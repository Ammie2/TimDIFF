(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param5739 = ((^((!(8'h9d)) ? {(8'had)} : (^~(8'ha2)))) + ((^(8'ha0)) ? ({(8'ha7)} - (~&(8'h9c))) : (~(~|(8'haa))))) )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h1651):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire4;
  input wire [(3'h4):(1'h0)] wire3;
  input wire [(2'h2):(1'h0)] wire2;
  input wire signed [(3'h4):(1'h0)] wire1;
  input wire signed [(4'he):(1'h0)] wire0;
  wire signed [(4'hd):(1'h0)] wire5737;
  wire [(3'h5):(1'h0)] wire553;
  wire [(3'h7):(1'h0)] wire552;
  reg signed [(4'hc):(1'h0)] reg551 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg550 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg549 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg548 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg547 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar546 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg545 = (1'h0);
  reg [(4'hc):(1'h0)] reg544 = (1'h0);
  reg [(3'h5):(1'h0)] forvar543 = (1'h0);
  reg [(2'h2):(1'h0)] reg542 = (1'h0);
  reg [(3'h7):(1'h0)] forvar541 = (1'h0);
  reg [(3'h6):(1'h0)] forvar540 = (1'h0);
  reg [(5'h10):(1'h0)] forvar539 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg538 = (1'h0);
  reg signed [(4'he):(1'h0)] reg537 = (1'h0);
  reg [(4'he):(1'h0)] forvar536 = (1'h0);
  reg signed [(4'he):(1'h0)] reg535 = (1'h0);
  reg [(5'h10):(1'h0)] reg534 = (1'h0);
  reg [(4'h8):(1'h0)] reg533 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg532 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg531 = (1'h0);
  reg [(4'ha):(1'h0)] forvar530 = (1'h0);
  reg [(4'h9):(1'h0)] reg528 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar527 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg529 = (1'h0);
  reg [(3'h5):(1'h0)] forvar528 = (1'h0);
  reg [(4'he):(1'h0)] reg527 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg526 = (1'h0);
  reg [(3'h5):(1'h0)] forvar525 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg520 = (1'h0);
  reg [(2'h3):(1'h0)] reg524 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg523 = (1'h0);
  reg [(3'h5):(1'h0)] reg522 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg521 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar520 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg519 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg518 = (1'h0);
  reg [(2'h2):(1'h0)] reg517 = (1'h0);
  reg [(4'h8):(1'h0)] reg516 = (1'h0);
  reg [(4'he):(1'h0)] forvar515 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar514 = (1'h0);
  reg [(4'ha):(1'h0)] forvar511 = (1'h0);
  reg [(4'h9):(1'h0)] reg510 = (1'h0);
  reg [(4'hf):(1'h0)] reg514 = (1'h0);
  reg [(3'h6):(1'h0)] reg513 = (1'h0);
  reg [(4'h8):(1'h0)] reg512 = (1'h0);
  reg [(2'h2):(1'h0)] reg511 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar510 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar509 = (1'h0);
  reg [(4'h8):(1'h0)] reg508 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar507 = (1'h0);
  reg [(4'h9):(1'h0)] reg506 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg505 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar504 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar503 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg502 = (1'h0);
  reg [(4'h9):(1'h0)] reg501 = (1'h0);
  reg [(3'h6):(1'h0)] forvar500 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg499 = (1'h0);
  reg [(4'he):(1'h0)] forvar498 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg496 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg495 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg494 = (1'h0);
  reg signed [(4'he):(1'h0)] reg493 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg492 = (1'h0);
  reg [(3'h4):(1'h0)] forvar491 = (1'h0);
  reg [(4'h8):(1'h0)] forvar490 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar489 = (1'h0);
  reg [(4'ha):(1'h0)] reg488 = (1'h0);
  reg [(5'h10):(1'h0)] reg487 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar486 = (1'h0);
  reg [(3'h6):(1'h0)] reg481 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg485 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg484 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg483 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar481 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg480 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg479 = (1'h0);
  reg [(4'hf):(1'h0)] reg478 = (1'h0);
  reg [(5'h10):(1'h0)] forvar476 = (1'h0);
  reg [(3'h4):(1'h0)] reg477 = (1'h0);
  reg [(4'hc):(1'h0)] reg476 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg475 = (1'h0);
  reg [(4'h9):(1'h0)] reg474 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg473 = (1'h0);
  reg [(3'h7):(1'h0)] reg472 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar471 = (1'h0);
  reg [(2'h2):(1'h0)] reg470 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg469 = (1'h0);
  reg [(4'h8):(1'h0)] reg468 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar466 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg467 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg466 = (1'h0);
  reg [(4'hf):(1'h0)] reg465 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg464 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar463 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg462 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg461 = (1'h0);
  reg [(4'ha):(1'h0)] reg460 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg459 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg458 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg457 = (1'h0);
  reg [(4'h9):(1'h0)] reg456 = (1'h0);
  reg [(4'h8):(1'h0)] reg455 = (1'h0);
  reg [(4'hd):(1'h0)] forvar454 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar453 = (1'h0);
  reg [(4'ha):(1'h0)] reg452 = (1'h0);
  reg [(3'h6):(1'h0)] reg451 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg450 = (1'h0);
  reg [(2'h2):(1'h0)] reg449 = (1'h0);
  reg [(4'he):(1'h0)] reg444 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar443 = (1'h0);
  reg [(4'h8):(1'h0)] reg448 = (1'h0);
  reg [(4'he):(1'h0)] reg447 = (1'h0);
  reg [(5'h10):(1'h0)] reg446 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg445 = (1'h0);
  reg [(3'h4):(1'h0)] forvar444 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg443 = (1'h0);
  reg [(4'hf):(1'h0)] reg442 = (1'h0);
  reg [(3'h4):(1'h0)] forvar441 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar428 = (1'h0);
  reg [(4'hc):(1'h0)] forvar427 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar424 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar415 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg418 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg414 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg413 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar410 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar405 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar399 = (1'h0);
  reg [(3'h6):(1'h0)] reg397 = (1'h0);
  reg [(3'h6):(1'h0)] reg393 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg392 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar391 = (1'h0);
  reg [(3'h5):(1'h0)] forvar430 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar429 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg425 = (1'h0);
  reg [(3'h4):(1'h0)] reg423 = (1'h0);
  reg [(4'hd):(1'h0)] forvar422 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar421 = (1'h0);
  reg [(4'hb):(1'h0)] forvar419 = (1'h0);
  reg [(3'h4):(1'h0)] reg417 = (1'h0);
  reg [(2'h2):(1'h0)] reg440 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar439 = (1'h0);
  reg [(3'h6):(1'h0)] reg438 = (1'h0);
  reg [(3'h4):(1'h0)] reg437 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg436 = (1'h0);
  reg [(3'h6):(1'h0)] reg435 = (1'h0);
  reg [(4'hc):(1'h0)] reg434 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg433 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg432 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg431 = (1'h0);
  reg [(5'h10):(1'h0)] reg430 = (1'h0);
  reg [(4'h8):(1'h0)] reg429 = (1'h0);
  reg [(2'h2):(1'h0)] reg428 = (1'h0);
  reg [(4'h8):(1'h0)] reg427 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar425 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg424 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar423 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg422 = (1'h0);
  reg [(4'hb):(1'h0)] reg421 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg420 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg419 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar418 = (1'h0);
  reg [(4'ha):(1'h0)] forvar417 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg415 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar414 = (1'h0);
  reg [(4'he):(1'h0)] forvar413 = (1'h0);
  reg [(2'h3):(1'h0)] forvar402 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg401 = (1'h0);
  reg [(3'h5):(1'h0)] reg412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg411 = (1'h0);
  reg [(5'h10):(1'h0)] reg410 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg408 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg407 = (1'h0);
  reg [(4'hb):(1'h0)] reg406 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg405 = (1'h0);
  reg [(4'he):(1'h0)] reg404 = (1'h0);
  reg [(4'h9):(1'h0)] reg403 = (1'h0);
  reg [(4'ha):(1'h0)] reg402 = (1'h0);
  reg [(3'h7):(1'h0)] forvar401 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg400 = (1'h0);
  reg [(3'h4):(1'h0)] reg399 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg398 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar397 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg395 = (1'h0);
  reg [(4'hd):(1'h0)] reg394 = (1'h0);
  reg [(4'h8):(1'h0)] forvar393 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar392 = (1'h0);
  reg [(4'hb):(1'h0)] reg391 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg390 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg389 = (1'h0);
  reg [(4'hf):(1'h0)] reg388 = (1'h0);
  reg [(4'he):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg386 = (1'h0);
  reg [(5'h10):(1'h0)] reg385 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg384 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg383 = (1'h0);
  reg [(2'h2):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg381 = (1'h0);
  reg [(3'h6):(1'h0)] forvar380 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg378 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg377 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar376 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg365 = (1'h0);
  reg [(3'h7):(1'h0)] reg375 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg374 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg373 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg372 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg371 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg370 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg368 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg367 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg366 = (1'h0);
  reg [(2'h3):(1'h0)] forvar365 = (1'h0);
  reg [(4'hd):(1'h0)] reg364 = (1'h0);
  reg [(2'h3):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg362 = (1'h0);
  reg [(4'ha):(1'h0)] reg361 = (1'h0);
  reg [(3'h6):(1'h0)] reg360 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg359 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar358 = (1'h0);
  reg [(4'h9):(1'h0)] reg357 = (1'h0);
  reg signed [(4'he):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar353 = (1'h0);
  reg [(3'h6):(1'h0)] reg341 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg351 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg350 = (1'h0);
  reg [(4'h8):(1'h0)] reg349 = (1'h0);
  reg [(4'hb):(1'h0)] reg348 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg347 = (1'h0);
  reg signed [(4'he):(1'h0)] reg346 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg345 = (1'h0);
  reg [(3'h7):(1'h0)] reg344 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg343 = (1'h0);
  reg [(3'h7):(1'h0)] reg342 = (1'h0);
  reg [(4'hd):(1'h0)] forvar341 = (1'h0);
  reg [(4'hc):(1'h0)] reg340 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg339 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg338 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg337 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg336 = (1'h0);
  reg [(2'h2):(1'h0)] forvar335 = (1'h0);
  reg [(3'h4):(1'h0)] reg334 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg333 = (1'h0);
  reg [(3'h6):(1'h0)] reg332 = (1'h0);
  reg [(3'h5):(1'h0)] reg331 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar330 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg329 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg328 = (1'h0);
  reg [(2'h2):(1'h0)] forvar327 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg326 = (1'h0);
  reg [(4'hf):(1'h0)] reg325 = (1'h0);
  reg [(3'h5):(1'h0)] reg324 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar323 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar322 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire321;
  wire signed [(4'he):(1'h0)] wire320;
  reg signed [(4'h9):(1'h0)] reg319 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg306 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg318 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar317 = (1'h0);
  reg [(4'hc):(1'h0)] reg316 = (1'h0);
  reg [(4'h9):(1'h0)] reg315 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg314 = (1'h0);
  reg [(4'hf):(1'h0)] reg313 = (1'h0);
  reg [(4'he):(1'h0)] reg312 = (1'h0);
  reg [(4'he):(1'h0)] reg311 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg310 = (1'h0);
  reg [(4'hf):(1'h0)] reg309 = (1'h0);
  reg signed [(4'he):(1'h0)] reg308 = (1'h0);
  reg [(2'h3):(1'h0)] reg307 = (1'h0);
  reg [(2'h2):(1'h0)] forvar306 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg301 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg305 = (1'h0);
  reg [(4'h9):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg303 = (1'h0);
  reg [(4'he):(1'h0)] reg302 = (1'h0);
  reg [(4'ha):(1'h0)] forvar301 = (1'h0);
  reg [(3'h6):(1'h0)] reg300 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar299 = (1'h0);
  reg [(3'h7):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg297 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar296 = (1'h0);
  reg [(4'hc):(1'h0)] reg295 = (1'h0);
  reg [(2'h3):(1'h0)] forvar294 = (1'h0);
  reg [(4'h9):(1'h0)] reg293 = (1'h0);
  reg signed [(4'he):(1'h0)] reg292 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg291 = (1'h0);
  reg [(2'h3):(1'h0)] forvar290 = (1'h0);
  reg signed [(4'he):(1'h0)] reg289 = (1'h0);
  reg signed [(4'he):(1'h0)] reg288 = (1'h0);
  reg [(3'h4):(1'h0)] reg287 = (1'h0);
  reg [(4'hb):(1'h0)] reg286 = (1'h0);
  reg [(3'h4):(1'h0)] forvar285 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar284 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg284 = (1'h0);
  reg [(3'h5):(1'h0)] reg283 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar280 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar275 = (1'h0);
  reg [(3'h4):(1'h0)] reg269 = (1'h0);
  reg [(3'h5):(1'h0)] reg268 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar267 = (1'h0);
  reg [(3'h5):(1'h0)] forvar262 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg282 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg281 = (1'h0);
  reg [(3'h6):(1'h0)] reg280 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg279 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg278 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg277 = (1'h0);
  reg signed [(4'he):(1'h0)] reg276 = (1'h0);
  reg [(3'h7):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg274 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg272 = (1'h0);
  reg signed [(4'he):(1'h0)] reg271 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg270 = (1'h0);
  reg [(4'hb):(1'h0)] forvar269 = (1'h0);
  reg [(4'ha):(1'h0)] forvar268 = (1'h0);
  reg [(5'h10):(1'h0)] reg267 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg263 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg265 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg264 = (1'h0);
  reg [(4'hc):(1'h0)] forvar263 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg261 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar260 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg259 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg258 = (1'h0);
  reg [(4'he):(1'h0)] reg257 = (1'h0);
  reg [(4'hd):(1'h0)] reg256 = (1'h0);
  reg [(3'h4):(1'h0)] forvar255 = (1'h0);
  reg [(3'h6):(1'h0)] forvar254 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg250 = (1'h0);
  reg [(4'h8):(1'h0)] reg244 = (1'h0);
  reg [(2'h2):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg245 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg254 = (1'h0);
  reg [(4'hf):(1'h0)] reg253 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar250 = (1'h0);
  reg [(4'hb):(1'h0)] reg249 = (1'h0);
  reg [(2'h3):(1'h0)] forvar248 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg247 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg246 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar245 = (1'h0);
  reg [(4'hb):(1'h0)] forvar244 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar243 = (1'h0);
  wire signed [(4'he):(1'h0)] wire242;
  wire [(4'hd):(1'h0)] wire241;
  reg signed [(4'h8):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg238 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg237 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg236 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg235 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg234 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar233 = (1'h0);
  reg [(2'h2):(1'h0)] forvar232 = (1'h0);
  reg [(3'h4):(1'h0)] reg231 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg230 = (1'h0);
  reg signed [(4'he):(1'h0)] reg229 = (1'h0);
  reg [(4'hf):(1'h0)] reg228 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg227 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg226 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg225 = (1'h0);
  reg [(5'h10):(1'h0)] forvar224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg223 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg222 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg220 = (1'h0);
  reg [(4'he):(1'h0)] forvar218 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg216 = (1'h0);
  reg [(3'h5):(1'h0)] forvar214 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar220 = (1'h0);
  reg [(4'hf):(1'h0)] reg219 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg217 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar216 = (1'h0);
  reg [(2'h3):(1'h0)] reg211 = (1'h0);
  reg [(3'h5):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg214 = (1'h0);
  reg [(2'h3):(1'h0)] reg213 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg212 = (1'h0);
  reg [(3'h5):(1'h0)] forvar211 = (1'h0);
  reg [(4'h8):(1'h0)] reg210 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg206 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg201 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg198 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar197 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar194 = (1'h0);
  reg [(4'ha):(1'h0)] forvar190 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg193 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar185 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar184 = (1'h0);
  reg [(5'h10):(1'h0)] reg183 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg179 = (1'h0);
  reg [(4'hf):(1'h0)] reg178 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg209 = (1'h0);
  reg [(2'h2):(1'h0)] reg208 = (1'h0);
  reg [(3'h5):(1'h0)] reg207 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar206 = (1'h0);
  reg [(4'hf):(1'h0)] reg205 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg204 = (1'h0);
  reg [(3'h5):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg202 = (1'h0);
  reg [(5'h10):(1'h0)] forvar201 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg199 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar198 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg196 = (1'h0);
  reg [(4'h8):(1'h0)] reg195 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg194 = (1'h0);
  reg [(2'h3):(1'h0)] forvar193 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg192 = (1'h0);
  reg signed [(4'he):(1'h0)] reg191 = (1'h0);
  reg [(4'hf):(1'h0)] forvar188 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg186 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg189 = (1'h0);
  reg [(3'h5):(1'h0)] reg188 = (1'h0);
  reg [(4'hc):(1'h0)] reg187 = (1'h0);
  reg [(4'hb):(1'h0)] forvar186 = (1'h0);
  reg [(4'h8):(1'h0)] reg185 = (1'h0);
  reg [(4'hc):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar183 = (1'h0);
  reg [(3'h7):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg181 = (1'h0);
  reg [(4'h9):(1'h0)] reg180 = (1'h0);
  reg [(4'hb):(1'h0)] forvar179 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar178 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg176 = (1'h0);
  reg [(4'hf):(1'h0)] reg175 = (1'h0);
  reg [(4'h9):(1'h0)] forvar174 = (1'h0);
  reg [(4'hc):(1'h0)] reg173 = (1'h0);
  reg [(3'h7):(1'h0)] reg172 = (1'h0);
  reg [(3'h6):(1'h0)] reg171 = (1'h0);
  reg [(4'hd):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar168 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg167 = (1'h0);
  reg [(4'hd):(1'h0)] reg166 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar165 = (1'h0);
  reg [(4'h9):(1'h0)] reg164 = (1'h0);
  reg [(4'hd):(1'h0)] reg163 = (1'h0);
  reg [(4'hb):(1'h0)] reg162 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg161 = (1'h0);
  reg [(4'he):(1'h0)] forvar160 = (1'h0);
  reg [(3'h5):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg159 = (1'h0);
  reg [(4'hb):(1'h0)] reg158 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar157 = (1'h0);
  reg [(3'h6):(1'h0)] reg156 = (1'h0);
  reg [(4'hf):(1'h0)] forvar155 = (1'h0);
  reg [(5'h10):(1'h0)] forvar154 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar153 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg152 = (1'h0);
  reg [(4'hd):(1'h0)] reg151 = (1'h0);
  reg [(3'h4):(1'h0)] reg150 = (1'h0);
  reg [(4'hf):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar147 = (1'h0);
  reg [(4'hb):(1'h0)] reg146 = (1'h0);
  reg [(4'hd):(1'h0)] reg145 = (1'h0);
  reg [(3'h5):(1'h0)] reg144 = (1'h0);
  reg [(3'h5):(1'h0)] reg143 = (1'h0);
  reg [(4'ha):(1'h0)] reg142 = (1'h0);
  reg [(2'h2):(1'h0)] reg141 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar140 = (1'h0);
  reg [(3'h6):(1'h0)] reg139 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg138 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg137 = (1'h0);
  reg [(4'hc):(1'h0)] reg136 = (1'h0);
  reg [(2'h3):(1'h0)] reg135 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar133 = (1'h0);
  reg [(4'hc):(1'h0)] reg132 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar131 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg130 = (1'h0);
  reg [(2'h3):(1'h0)] forvar129 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg128 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg127 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg126 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar125 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg124 = (1'h0);
  reg [(3'h5):(1'h0)] reg123 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg122 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg121 = (1'h0);
  reg [(4'he):(1'h0)] forvar120 = (1'h0);
  reg [(4'h8):(1'h0)] forvar119 = (1'h0);
  reg [(3'h4):(1'h0)] reg118 = (1'h0);
  reg [(4'ha):(1'h0)] reg117 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg115 = (1'h0);
  reg [(4'hf):(1'h0)] forvar114 = (1'h0);
  reg [(3'h4):(1'h0)] forvar113 = (1'h0);
  reg [(2'h3):(1'h0)] reg112 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar110 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg108 = (1'h0);
  reg [(4'hd):(1'h0)] reg107 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg106 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg104 = (1'h0);
  reg [(3'h5):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar102 = (1'h0);
  reg [(4'ha):(1'h0)] reg101 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg99 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg94 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg98 = (1'h0);
  reg [(5'h10):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg96 = (1'h0);
  reg [(4'hb):(1'h0)] reg95 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar94 = (1'h0);
  reg [(4'hc):(1'h0)] reg93 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar92 = (1'h0);
  reg [(5'h10):(1'h0)] reg91 = (1'h0);
  reg [(2'h2):(1'h0)] forvar79 = (1'h0);
  reg [(4'hb):(1'h0)] reg90 = (1'h0);
  reg [(4'h9):(1'h0)] forvar74 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar70 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg69 = (1'h0);
  reg [(4'hc):(1'h0)] reg89 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg88 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg87 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar86 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg85 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg84 = (1'h0);
  reg [(4'ha):(1'h0)] reg83 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg82 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg76 = (1'h0);
  reg [(4'h9):(1'h0)] forvar75 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg81 = (1'h0);
  reg [(4'hf):(1'h0)] reg80 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg79 = (1'h0);
  reg [(3'h6):(1'h0)] reg78 = (1'h0);
  reg [(4'he):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar76 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg75 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg74 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg73 = (1'h0);
  reg [(4'hf):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar69 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg68 = (1'h0);
  reg [(4'ha):(1'h0)] forvar67 = (1'h0);
  reg [(4'hd):(1'h0)] reg66 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar64 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg61 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar59 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar56 = (1'h0);
  reg [(3'h6):(1'h0)] reg55 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg53 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar52 = (1'h0);
  reg [(4'hd):(1'h0)] reg50 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar45 = (1'h0);
  reg [(4'he):(1'h0)] forvar37 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar36 = (1'h0);
  reg [(4'hc):(1'h0)] reg64 = (1'h0);
  reg [(4'hf):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg62 = (1'h0);
  reg [(3'h6):(1'h0)] forvar61 = (1'h0);
  reg [(4'hd):(1'h0)] reg60 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg58 = (1'h0);
  reg [(4'hd):(1'h0)] reg57 = (1'h0);
  reg [(3'h6):(1'h0)] reg56 = (1'h0);
  reg [(4'ha):(1'h0)] forvar55 = (1'h0);
  reg [(5'h10):(1'h0)] reg54 = (1'h0);
  reg [(4'hd):(1'h0)] forvar53 = (1'h0);
  reg [(3'h6):(1'h0)] reg52 = (1'h0);
  reg [(4'ha):(1'h0)] reg51 = (1'h0);
  reg [(4'h8):(1'h0)] forvar50 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg49 = (1'h0);
  reg [(3'h6):(1'h0)] forvar48 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg43 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar40 = (1'h0);
  reg [(4'h8):(1'h0)] reg39 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg47 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg46 = (1'h0);
  reg signed [(4'he):(1'h0)] reg45 = (1'h0);
  reg [(3'h7):(1'h0)] reg44 = (1'h0);
  reg [(4'ha):(1'h0)] forvar43 = (1'h0);
  reg [(4'h9):(1'h0)] reg42 = (1'h0);
  reg [(3'h5):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg40 = (1'h0);
  reg [(3'h5):(1'h0)] forvar39 = (1'h0);
  reg [(4'hc):(1'h0)] reg38 = (1'h0);
  reg [(4'ha):(1'h0)] reg37 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar11 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7 = (1'h0);
  reg [(3'h6):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg33 = (1'h0);
  reg [(3'h4):(1'h0)] reg32 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg31 = (1'h0);
  reg [(4'h9):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg27 = (1'h0);
  reg [(3'h5):(1'h0)] reg26 = (1'h0);
  reg [(4'hd):(1'h0)] reg25 = (1'h0);
  reg [(4'hf):(1'h0)] reg24 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg23 = (1'h0);
  reg [(3'h5):(1'h0)] reg22 = (1'h0);
  reg [(3'h5):(1'h0)] forvar21 = (1'h0);
  reg [(4'hb):(1'h0)] forvar20 = (1'h0);
  reg [(4'he):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg18 = (1'h0);
  reg [(3'h7):(1'h0)] reg17 = (1'h0);
  reg [(4'hb):(1'h0)] reg16 = (1'h0);
  reg [(3'h5):(1'h0)] reg15 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg13 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg12 = (1'h0);
  reg [(4'hc):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg10 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg9 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar8 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6 = (1'h0);
  wire [(2'h2):(1'h0)] wire5;
  assign y = {wire5737,
                 wire553,
                 wire552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 forvar546,
                 reg545,
                 reg544,
                 forvar543,
                 reg542,
                 forvar541,
                 forvar540,
                 forvar539,
                 reg538,
                 reg537,
                 forvar536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg531,
                 forvar530,
                 reg528,
                 forvar527,
                 reg529,
                 forvar528,
                 reg527,
                 reg526,
                 forvar525,
                 reg520,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 forvar520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 forvar515,
                 forvar514,
                 forvar511,
                 reg510,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 forvar510,
                 forvar509,
                 reg508,
                 forvar507,
                 reg506,
                 reg505,
                 forvar504,
                 forvar503,
                 reg502,
                 reg501,
                 forvar500,
                 reg499,
                 forvar498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 forvar491,
                 forvar490,
                 forvar489,
                 reg488,
                 reg487,
                 forvar486,
                 reg481,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 forvar481,
                 reg480,
                 reg479,
                 reg478,
                 forvar476,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 forvar471,
                 reg470,
                 reg469,
                 reg468,
                 forvar466,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 forvar463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 forvar454,
                 forvar453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg444,
                 forvar443,
                 reg448,
                 reg447,
                 reg446,
                 reg445,
                 forvar444,
                 reg443,
                 reg442,
                 forvar441,
                 forvar428,
                 forvar427,
                 forvar424,
                 forvar415,
                 reg418,
                 reg414,
                 reg413,
                 forvar410,
                 forvar405,
                 forvar399,
                 reg397,
                 reg393,
                 reg392,
                 forvar391,
                 forvar430,
                 forvar429,
                 reg425,
                 reg423,
                 forvar422,
                 forvar421,
                 forvar419,
                 reg417,
                 reg440,
                 forvar439,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 forvar425,
                 reg424,
                 forvar423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 forvar418,
                 forvar417,
                 reg416,
                 reg415,
                 forvar414,
                 forvar413,
                 forvar402,
                 reg401,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 forvar401,
                 reg400,
                 reg399,
                 reg398,
                 forvar397,
                 reg396,
                 reg395,
                 reg394,
                 forvar393,
                 forvar392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 forvar380,
                 reg379,
                 reg378,
                 reg377,
                 forvar376,
                 reg365,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 forvar365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 forvar358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 forvar353,
                 reg341,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg342,
                 forvar341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 forvar335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 forvar330,
                 reg329,
                 reg328,
                 forvar327,
                 reg326,
                 reg325,
                 reg324,
                 forvar323,
                 forvar322,
                 wire321,
                 wire320,
                 reg319,
                 reg306,
                 reg318,
                 forvar317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 forvar306,
                 reg301,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 forvar301,
                 reg300,
                 forvar299,
                 reg298,
                 reg297,
                 forvar296,
                 reg295,
                 forvar294,
                 reg293,
                 reg292,
                 reg291,
                 forvar290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 forvar285,
                 forvar284,
                 reg284,
                 reg283,
                 forvar280,
                 forvar275,
                 reg269,
                 reg268,
                 forvar267,
                 forvar262,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 forvar269,
                 forvar268,
                 reg267,
                 reg266,
                 reg263,
                 reg265,
                 reg264,
                 forvar263,
                 reg262,
                 reg261,
                 forvar260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 forvar255,
                 forvar254,
                 reg250,
                 reg244,
                 reg248,
                 reg245,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 forvar250,
                 reg249,
                 forvar248,
                 reg247,
                 reg246,
                 forvar245,
                 forvar244,
                 forvar243,
                 wire242,
                 wire241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 forvar233,
                 forvar232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 forvar224,
                 reg223,
                 reg222,
                 reg220,
                 forvar218,
                 reg216,
                 forvar214,
                 reg221,
                 forvar220,
                 reg219,
                 reg218,
                 reg217,
                 forvar216,
                 reg211,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 forvar211,
                 reg210,
                 reg206,
                 reg201,
                 reg198,
                 forvar197,
                 forvar194,
                 forvar190,
                 reg193,
                 forvar185,
                 forvar184,
                 reg183,
                 reg179,
                 reg178,
                 reg209,
                 reg208,
                 reg207,
                 forvar206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 forvar201,
                 reg200,
                 reg199,
                 forvar198,
                 reg197,
                 reg196,
                 reg195,
                 reg194,
                 forvar193,
                 reg192,
                 reg191,
                 forvar188,
                 reg186,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 forvar186,
                 reg185,
                 reg184,
                 forvar183,
                 reg182,
                 reg181,
                 reg180,
                 forvar179,
                 forvar178,
                 reg177,
                 reg176,
                 reg175,
                 forvar174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 forvar168,
                 reg167,
                 reg166,
                 forvar165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 forvar160,
                 reg157,
                 reg159,
                 reg158,
                 forvar157,
                 reg156,
                 forvar155,
                 forvar154,
                 forvar153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 forvar147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 forvar140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 forvar133,
                 reg132,
                 forvar131,
                 reg130,
                 forvar129,
                 reg128,
                 reg127,
                 reg126,
                 forvar125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 forvar120,
                 forvar119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 forvar114,
                 forvar113,
                 reg112,
                 reg111,
                 forvar110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 forvar102,
                 reg101,
                 reg100,
                 reg99,
                 reg94,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 forvar94,
                 reg93,
                 forvar92,
                 reg91,
                 forvar79,
                 reg90,
                 forvar74,
                 forvar70,
                 reg69,
                 reg89,
                 reg88,
                 reg87,
                 forvar86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg76,
                 forvar75,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 forvar76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 forvar69,
                 reg68,
                 forvar67,
                 reg66,
                 reg65,
                 forvar64,
                 reg61,
                 forvar59,
                 forvar56,
                 reg55,
                 reg53,
                 forvar52,
                 reg50,
                 forvar45,
                 forvar37,
                 forvar36,
                 reg64,
                 reg63,
                 reg62,
                 forvar61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 forvar55,
                 reg54,
                 forvar53,
                 reg52,
                 reg51,
                 forvar50,
                 reg49,
                 forvar48,
                 reg43,
                 forvar40,
                 reg39,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 forvar43,
                 reg42,
                 reg41,
                 reg40,
                 forvar39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 forvar11,
                 reg7,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 forvar21,
                 forvar20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 forvar8,
                 forvar7,
                 forvar6,
                 wire5,
                 (1'h0)};
  assign wire5 = (^(($signed(wire4) ?
                     $signed((8'hb1)) : wire1[(3'h4):(1'h1)]) || $signed($signed(wire4))));
  always
    @(posedge clk) begin
      for (forvar6 = (1'h0); (forvar6 < (1'h1)); forvar6 = (forvar6 + (1'h1)))
        begin
          if ($unsigned(($unsigned($unsigned(wire0)) && (8'hb4))))
            begin
              for (forvar7 = (1'h0); (forvar7 < (2'h3)); forvar7 = (forvar7 + (1'h1)))
                begin
                  for (forvar8 = (1'h0); (forvar8 < (2'h2)); forvar8 = (forvar8 + (1'h1)))
                    begin
                      reg9 <= ((forvar7 ? wire1 : forvar8) ^~ wire3);
                      reg10 <= ($unsigned($signed((wire0 == forvar6))) <<< ((~^wire0[(4'hd):(2'h3)]) + wire2));
                      reg11 <= {(wire3[(2'h2):(1'h0)] ~^ ((wire3 >> wire0) < $unsigned((8'ha8))))};
                    end
                  if (({reg10[(1'h1):(1'h1)]} ~^ $signed((forvar8 + {wire1}))))
                    begin
                      reg12 <= $unsigned((reg10 ?
                          $signed(((8'h9d) ? wire3 : reg9)) : wire5));
                      reg13 <= $signed($signed(reg9[(4'hb):(4'ha)]));
                    end
                  else
                    begin
                      reg12 <= reg13[(1'h0):(1'h0)];
                      reg13 <= $signed(($unsigned({reg12}) & (8'hab)));
                      reg14 <= reg9[(4'hd):(4'hd)];
                      reg15 <= wire1;
                    end
                  if ((~|wire1))
                    begin
                      reg16 <= $unsigned(reg9[(1'h0):(1'h0)]);
                      reg17 <= ((((^~(8'h9c)) | (wire1 ? reg9 : forvar7)) ?
                          (wire3 ?
                              reg13[(2'h3):(2'h2)] : forvar7) : wire1) >= (+{wire5}));
                      reg18 <= ($unsigned((|(^~reg9))) ?
                          (~^((reg9 > (8'hb8)) || $signed(reg10))) : {reg15[(3'h4):(3'h4)]});
                      reg19 <= reg18;
                    end
                  else
                    begin
                      reg16 <= $signed((~^((8'ha2) ?
                          $unsigned(reg12) : reg18)));
                      reg17 <= ((wire3 ?
                          (!$signed((8'h9e))) : ((~|wire2) >= wire2)) ^ (({forvar7} >>> (|reg14)) ~^ $signed(((8'hb1) <= forvar8))));
                      reg18 <= (8'h9e);
                    end
                end
              for (forvar20 = (1'h0); (forvar20 < (2'h3)); forvar20 = (forvar20 + (1'h1)))
                begin
                  for (forvar21 = (1'h0); (forvar21 < (2'h3)); forvar21 = (forvar21 + (1'h1)))
                    begin
                      reg22 <= (!$unsigned({{reg15}}));
                    end
                  if (reg22[(2'h3):(2'h3)])
                    begin
                      reg23 <= {reg17};
                      reg24 <= {(~|(+{reg16}))};
                    end
                  else
                    begin
                      reg23 <= reg18[(2'h2):(1'h0)];
                      reg24 <= $unsigned(($unsigned($unsigned(wire4)) ?
                          (((8'h9d) ? reg19 : (8'hb2)) ?
                              wire0 : $signed(forvar7)) : reg16[(2'h3):(2'h3)]));
                      reg25 <= ((($unsigned(forvar21) != (^~wire0)) << (reg15 ?
                          (reg22 * wire3) : (wire3 ^ wire4))) >>> ((^~$unsigned(wire1)) ?
                          $signed((8'hb0)) : {(forvar21 ? reg14 : (8'hb4))}));
                      reg26 <= (^wire1);
                    end
                  if ((wire0[(4'he):(3'h5)] ^ ((8'hb3) >= $signed(wire0))))
                    begin
                      reg27 <= forvar21;
                      reg28 <= reg16;
                    end
                  else
                    begin
                      reg27 <= (reg15[(3'h5):(3'h4)] ?
                          {(|(|reg10))} : (($unsigned((8'ha9)) ?
                                  (+reg23) : forvar20[(4'h9):(3'h4)]) ?
                              (8'hb6) : ($unsigned((8'h9d)) < $signed(wire3))));
                      reg28 <= {$unsigned(((wire5 & wire2) > (|reg11)))};
                      reg29 <= wire0[(4'ha):(3'h5)];
                      reg30 <= $unsigned(forvar21[(2'h3):(1'h0)]);
                    end
                  if ($signed($unsigned((reg18[(1'h1):(1'h0)] || reg24[(4'hf):(4'hd)]))))
                    begin
                      reg31 <= ($unsigned({(-reg25)}) >>> (8'ha1));
                      reg32 <= reg10[(4'ha):(1'h0)];
                      reg33 <= reg32[(1'h1):(1'h0)];
                      reg34 <= (($signed($unsigned(reg32)) ?
                          ((reg24 ? reg33 : wire5) ?
                              wire3 : (|forvar7)) : ($unsigned(reg15) ?
                              reg11 : {reg16})) < (+reg28[(5'h10):(2'h2)]));
                    end
                  else
                    begin
                      reg31 <= (((!reg10[(4'h9):(2'h3)]) == {(forvar8 ?
                              reg32 : reg12)}) ~^ $signed(({reg29} ?
                          $unsigned(reg16) : ((8'ha5) ? (8'h9e) : forvar20))));
                      reg32 <= (8'hb5);
                    end
                end
            end
          else
            begin
              if ($signed($signed($unsigned(wire3))))
                begin
                  reg7 <= $unsigned(wire1);
                end
              else
                begin
                  reg7 <= {(^~(8'hab))};
                  for (forvar8 = (1'h0); (forvar8 < (1'h0)); forvar8 = (forvar8 + (1'h1)))
                    begin
                      reg9 <= (^~($signed((reg16 ?
                          (8'hb1) : (8'hb5))) + (|(8'ha4))));
                      reg10 <= wire4;
                    end
                  for (forvar11 = (1'h0); (forvar11 < (1'h1)); forvar11 = (forvar11 + (1'h1)))
                    begin
                      reg12 <= (reg16[(1'h0):(1'h0)] ?
                          $unsigned($signed(forvar20)) : $signed(wire0[(4'ha):(3'h6)]));
                      reg13 <= ($unsigned((!forvar21[(3'h5):(2'h3)])) > {wire0[(4'ha):(3'h7)]});
                    end
                end
            end
          reg35 <= ($signed((((8'hb5) > reg17) && (reg13 ? reg11 : reg16))) ?
              (~&reg26[(3'h4):(2'h2)]) : forvar6);
          if (forvar11)
            begin
              reg36 <= ($signed(forvar11) - ({$unsigned(reg34)} ?
                  {$signed(reg31)} : $signed(((8'ha9) ? wire2 : reg18))));
              if ((~|($signed($unsigned(forvar7)) ?
                  (~&$unsigned(wire3)) : ((reg31 && (8'hb9)) ^~ reg18[(2'h2):(1'h0)]))))
                begin
                  if ({{reg32}})
                    begin
                      reg37 <= (&forvar11[(3'h6):(1'h0)]);
                      reg38 <= reg10;
                    end
                  else
                    begin
                      reg37 <= {$unsigned((&reg34[(1'h1):(1'h1)]))};
                      reg38 <= ({reg36} ?
                          {reg27[(4'hd):(4'hd)]} : $signed($signed((8'ha4))));
                    end
                  for (forvar39 = (1'h0); (forvar39 < (2'h2)); forvar39 = (forvar39 + (1'h1)))
                    begin
                      reg40 <= ($signed(reg18) ?
                          wire1[(2'h3):(1'h1)] : ((forvar6 ?
                                  $unsigned(reg12) : (forvar11 ?
                                      reg10 : reg32)) ?
                              $unsigned($signed(forvar6)) : (((8'hb8) == reg37) ?
                                  (^reg9) : reg18[(1'h0):(1'h0)])));
                      reg41 <= (wire5 ?
                          ((^~((8'hab) ?
                              reg30 : (8'haf))) ^~ (!$unsigned(reg40))) : $unsigned((-reg12)));
                      reg42 <= (^$unsigned($unsigned((^~reg7))));
                    end
                  for (forvar43 = (1'h0); (forvar43 < (1'h1)); forvar43 = (forvar43 + (1'h1)))
                    begin
                      reg44 <= ($signed(({forvar6} * reg27)) ?
                          reg27 : reg40[(1'h1):(1'h1)]);
                      reg45 <= ((8'h9e) | ($signed($signed(reg15)) < (~&(|wire5))));
                      reg46 <= reg18;
                      reg47 <= {(((reg45 ? reg33 : reg46) ? reg28 : (8'haf)) ?
                              (^(reg24 ?
                                  (8'ha4) : reg10)) : ((reg37 > reg25) << (wire5 > (8'haa))))};
                    end
                end
              else
                begin
                  if (({forvar39} < $unsigned((8'ha0))))
                    begin
                      reg37 <= (~$signed(((reg25 ? (8'hae) : reg31) ?
                          (^(8'hac)) : $unsigned((8'ha0)))));
                      reg38 <= forvar8[(3'h6):(1'h0)];
                      reg39 <= (!$unsigned($signed((reg9 > forvar39))));
                    end
                  else
                    begin
                      reg37 <= $signed(reg31[(3'h6):(3'h6)]);
                      reg38 <= $unsigned((reg13[(2'h2):(2'h2)] - (~reg12)));
                    end
                  for (forvar40 = (1'h0); (forvar40 < (1'h1)); forvar40 = (forvar40 + (1'h1)))
                    begin
                      reg41 <= $signed(reg23);
                      reg42 <= ((reg39[(2'h2):(1'h0)] ^~ ({forvar20} ?
                          (8'hba) : {reg14})) | reg31);
                    end
                  if (({$unsigned(reg35[(1'h1):(1'h1)])} <= ($unsigned($signed(reg32)) < $unsigned((reg9 ?
                      reg23 : reg13)))))
                    begin
                      reg43 <= $signed(({(~^reg9)} ?
                          $signed((^~(8'hb0))) : $signed(((8'hb0) ?
                              reg45 : (8'hb3)))));
                      reg44 <= $unsigned($unsigned(reg44[(1'h1):(1'h1)]));
                      reg45 <= $signed(($unsigned($signed((8'hac))) ?
                          reg43[(1'h0):(1'h0)] : $unsigned($signed(reg27))));
                    end
                  else
                    begin
                      reg43 <= ((~$unsigned({reg15})) ?
                          (^$signed(reg24)) : ((((8'haa) + reg15) ?
                                  reg19 : reg11[(3'h5):(2'h3)]) ?
                              reg17[(2'h3):(2'h3)] : (((8'ha9) >= reg35) << reg11[(2'h2):(2'h2)])));
                    end
                end
              for (forvar48 = (1'h0); (forvar48 < (1'h0)); forvar48 = (forvar48 + (1'h1)))
                begin
                  if (($signed($signed((!reg24))) ?
                      reg38[(1'h1):(1'h1)] : ($unsigned((reg38 ?
                              forvar7 : reg18)) ?
                          reg40[(1'h1):(1'h0)] : forvar7)))
                    begin
                      reg49 <= (8'haf);
                    end
                  else
                    begin
                      reg49 <= $unsigned((~&(reg32 >> $signed(reg15))));
                    end
                  for (forvar50 = (1'h0); (forvar50 < (1'h0)); forvar50 = (forvar50 + (1'h1)))
                    begin
                      reg51 <= (8'haf);
                      reg52 <= (wire4 ? $unsigned((+(~|forvar20))) : reg11);
                    end
                end
              for (forvar53 = (1'h0); (forvar53 < (1'h1)); forvar53 = (forvar53 + (1'h1)))
                begin
                  reg54 <= (~reg51[(3'h4):(1'h0)]);
                  for (forvar55 = (1'h0); (forvar55 < (2'h2)); forvar55 = (forvar55 + (1'h1)))
                    begin
                      reg56 <= $unsigned($signed(((-wire3) ?
                          (8'h9d) : (reg28 ? reg45 : reg52))));
                    end
                  if (reg49)
                    begin
                      reg57 <= ($signed(reg24) ?
                          {forvar7} : (({reg24} && (reg16 - reg23)) ^ (reg35 && reg15)));
                      reg58 <= $signed((reg52 ^~ (-((8'ha9) ? reg22 : reg57))));
                      reg59 <= (reg49 ?
                          forvar11 : ({forvar8[(1'h0):(1'h0)]} ?
                              (forvar20[(3'h4):(2'h3)] ?
                                  (|(8'hae)) : (^(8'hab))) : (&(8'h9e))));
                    end
                  else
                    begin
                      reg57 <= (((-(~|(8'haf))) && ($signed(forvar7) ?
                              (8'ha1) : {reg18})) ?
                          {reg34} : $signed((wire4 >> $unsigned((8'haa)))));
                      reg58 <= (($unsigned(reg46[(2'h3):(2'h3)]) - wire4[(3'h6):(2'h3)]) ?
                          (~{(forvar39 ?
                                  forvar50 : (8'ha8))}) : $signed((8'ha4)));
                      reg59 <= {$unsigned((forvar43[(4'h8):(1'h1)] ?
                              reg18 : reg51))};
                      reg60 <= ((8'h9d) == reg32[(2'h2):(1'h1)]);
                    end
                  for (forvar61 = (1'h0); (forvar61 < (2'h2)); forvar61 = (forvar61 + (1'h1)))
                    begin
                      reg62 <= reg36;
                      reg63 <= $signed({reg34[(2'h2):(1'h0)]});
                      reg64 <= reg39;
                    end
                end
            end
          else
            begin
              for (forvar36 = (1'h0); (forvar36 < (1'h1)); forvar36 = (forvar36 + (1'h1)))
                begin
                  for (forvar37 = (1'h0); (forvar37 < (1'h1)); forvar37 = (forvar37 + (1'h1)))
                    begin
                      reg38 <= (8'ha4);
                      reg39 <= (+(-(^(~|reg59))));
                      reg40 <= $unsigned((~^reg22[(2'h3):(2'h2)]));
                      reg41 <= (^~$signed(({reg25} ?
                          {reg54} : reg13[(3'h5):(3'h5)])));
                    end
                  if ($unsigned((forvar8 ?
                      ($unsigned(reg35) ?
                          (~^reg11) : reg35[(3'h4):(3'h4)]) : ((~&reg27) <= $signed(forvar40)))))
                    begin
                      reg42 <= (reg28 ?
                          ((-$signed((8'hb9))) + $unsigned((reg24 < reg31))) : reg51[(2'h2):(1'h1)]);
                      reg43 <= ($signed((|{reg63})) ^~ reg11[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg42 <= reg57;
                    end
                end
              reg44 <= $signed(($unsigned($signed(reg7)) ?
                  wire4[(3'h4):(2'h2)] : reg51[(1'h0):(1'h0)]));
              if (reg60)
                begin
                  for (forvar45 = (1'h0); (forvar45 < (2'h3)); forvar45 = (forvar45 + (1'h1)))
                    begin
                      reg46 <= forvar50;
                    end
                  reg47 <= (~^(((reg30 ? reg41 : (8'ha3)) ?
                      {(8'haf)} : $unsigned(forvar7)) << reg42));
                  for (forvar48 = (1'h0); (forvar48 < (2'h3)); forvar48 = (forvar48 + (1'h1)))
                    begin
                      reg49 <= {$signed(reg22)};
                      reg50 <= forvar7[(4'hb):(2'h2)];
                      reg51 <= $signed((+$unsigned(reg33)));
                    end
                  for (forvar52 = (1'h0); (forvar52 < (2'h2)); forvar52 = (forvar52 + (1'h1)))
                    begin
                      reg53 <= $unsigned((^~$unsigned((reg35 ~^ reg49))));
                      reg54 <= $signed(reg43);
                    end
                end
              else
                begin
                  for (forvar45 = (1'h0); (forvar45 < (1'h1)); forvar45 = (forvar45 + (1'h1)))
                    begin
                      reg46 <= ((8'hae) != $signed((reg64[(4'h9):(4'h9)] ?
                          forvar11 : forvar52)));
                      reg47 <= ((~|(~^reg47)) > reg33);
                    end
                  for (forvar48 = (1'h0); (forvar48 < (2'h3)); forvar48 = (forvar48 + (1'h1)))
                    begin
                      reg49 <= $signed(reg38);
                      reg50 <= reg44;
                      reg51 <= (8'had);
                    end
                  for (forvar52 = (1'h0); (forvar52 < (2'h2)); forvar52 = (forvar52 + (1'h1)))
                    begin
                      reg53 <= reg45[(4'h8):(3'h5)];
                      reg54 <= reg58[(1'h0):(1'h0)];
                      reg55 <= (~^(reg45 >>> $signed(forvar53)));
                    end
                end
              if (($signed((|(wire4 == reg60))) << forvar21))
                begin
                  for (forvar56 = (1'h0); (forvar56 < (1'h0)); forvar56 = (forvar56 + (1'h1)))
                    begin
                      reg57 <= wire1;
                      reg58 <= ((({reg41} ?
                                  (reg33 ? reg25 : (8'hb4)) : (|reg7)) ?
                              $unsigned(reg19) : {(reg50 == forvar8)}) ?
                          $unsigned(($unsigned(forvar43) == (reg10 ?
                              reg37 : (8'h9e)))) : (((reg36 ~^ reg30) ?
                              {reg19} : ((8'ha0) >>> reg7)) ^ $unsigned($unsigned((8'hba)))));
                      reg59 <= reg13;
                      reg60 <= ($signed((~^$signed((8'ha7)))) ?
                          {(reg31[(3'h4):(2'h3)] >> reg46)} : (({reg44} - $unsigned(reg13)) ?
                              $signed((^~(8'hb9))) : reg7[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  if (reg28)
                    begin
                      reg56 <= (^forvar20[(4'h9):(1'h0)]);
                      reg57 <= (|forvar7);
                    end
                  else
                    begin
                      reg56 <= $signed($signed((+forvar56[(2'h3):(1'h0)])));
                      reg57 <= forvar45;
                      reg58 <= (((~&$unsigned(forvar6)) ^~ forvar45[(1'h1):(1'h1)]) ?
                          reg49[(3'h6):(1'h0)] : reg47);
                    end
                  for (forvar59 = (1'h0); (forvar59 < (2'h3)); forvar59 = (forvar59 + (1'h1)))
                    begin
                      reg60 <= (~^forvar36[(1'h1):(1'h1)]);
                      reg61 <= (8'hb4);
                      reg62 <= (8'hba);
                      reg63 <= $unsigned(({(^~(8'hac))} ?
                          $signed($unsigned((8'ha6))) : (&(reg46 + forvar53))));
                    end
                  for (forvar64 = (1'h0); (forvar64 < (1'h1)); forvar64 = (forvar64 + (1'h1)))
                    begin
                      reg65 <= ($unsigned((~^wire4)) ?
                          {({reg54} && forvar56[(3'h5):(3'h5)])} : (~|reg26));
                    end
                end
            end
        end
      reg66 <= (8'hab);
      for (forvar67 = (1'h0); (forvar67 < (1'h0)); forvar67 = (forvar67 + (1'h1)))
        begin
          reg68 <= reg10;
          if (forvar11[(3'h5):(2'h3)])
            begin
              for (forvar69 = (1'h0); (forvar69 < (2'h2)); forvar69 = (forvar69 + (1'h1)))
                begin
                  if ($unsigned($unsigned(reg10[(4'hd):(4'hc)])))
                    begin
                      reg70 <= $unsigned(reg56);
                      reg71 <= forvar39;
                      reg72 <= forvar36;
                      reg73 <= reg31[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg70 <= ($signed(reg46) ?
                          (($signed(reg60) ? (reg44 - reg35) : $signed(wire1)) ?
                              reg31[(2'h3):(2'h2)] : (&reg65)) : forvar40);
                      reg71 <= ($signed(((^reg22) == (|reg52))) ?
                          ($signed((reg7 ? reg25 : forvar56)) ?
                              (8'hb6) : (forvar40[(4'h9):(2'h2)] ?
                                  $signed((8'hb3)) : (reg11 ^~ reg61))) : ($unsigned($signed(reg31)) ?
                              reg33 : {$signed((8'ha9))}));
                      reg72 <= $signed($signed(($unsigned(reg13) ?
                          (forvar48 ^ reg19) : reg53)));
                    end
                  reg74 <= $signed(reg49);
                end
              if ($unsigned(({$signed((8'had))} >> reg11)))
                begin
                  reg75 <= $unsigned(({reg38} ?
                      ((reg63 ^~ reg65) ?
                          reg40 : reg12[(1'h0):(1'h0)]) : (reg51[(3'h4):(1'h0)] ?
                          (|forvar53) : (~&reg38))));
                  for (forvar76 = (1'h0); (forvar76 < (1'h1)); forvar76 = (forvar76 + (1'h1)))
                    begin
                      reg77 <= reg49[(1'h1):(1'h1)];
                      reg78 <= $signed((^~({reg28} ?
                          $unsigned(forvar40) : $signed(reg18))));
                      reg79 <= (~|reg41);
                      reg80 <= ((+(-$signed(reg73))) ?
                          {reg70} : $unsigned(((reg40 ?
                              reg23 : wire4) ~^ reg57)));
                    end
                  reg81 <= $unsigned({((8'haf) ? reg77 : (~|forvar50))});
                end
              else
                begin
                  for (forvar75 = (1'h0); (forvar75 < (1'h1)); forvar75 = (forvar75 + (1'h1)))
                    begin
                      reg76 <= (8'hb1);
                      reg77 <= (reg40[(2'h3):(2'h2)] << (8'hac));
                      reg78 <= (($signed(reg30[(4'h9):(1'h0)]) ?
                          $unsigned((forvar43 <= reg56)) : ($unsigned(forvar53) >>> $unsigned(reg66))) << $unsigned($signed((reg59 ?
                          forvar56 : forvar64))));
                      reg79 <= ((~^$signed($unsigned(reg52))) * $unsigned(((reg26 & reg17) | $signed((8'h9f)))));
                    end
                  if (((reg33[(4'hc):(1'h0)] > reg55) ?
                      (8'ha1) : wire2[(1'h0):(1'h0)]))
                    begin
                      reg80 <= reg57[(4'hd):(3'h7)];
                      reg81 <= ($unsigned(reg14) ^ ($unsigned({(8'h9f)}) << ($signed(forvar48) + wire1)));
                    end
                  else
                    begin
                      reg80 <= {reg70[(1'h0):(1'h0)]};
                      reg81 <= forvar52[(3'h4):(2'h2)];
                    end
                  if ($unsigned($signed(($unsigned(reg14) ?
                      $signed(reg27) : reg55[(2'h2):(1'h1)]))))
                    begin
                      reg82 <= (&$signed(forvar48));
                    end
                  else
                    begin
                      reg82 <= ((8'ha8) ?
                          $signed(($unsigned(reg60) ?
                              reg57 : $unsigned(reg42))) : reg42[(3'h5):(2'h3)]);
                      reg83 <= (8'ha3);
                      reg84 <= $signed($signed($signed(reg11)));
                      reg85 <= wire4[(5'h10):(4'h9)];
                    end
                end
              for (forvar86 = (1'h0); (forvar86 < (1'h0)); forvar86 = (forvar86 + (1'h1)))
                begin
                  if ($unsigned({((reg28 ? (8'hba) : reg53) ?
                          forvar39 : $unsigned((8'hb7)))}))
                    begin
                      reg87 <= ((8'hb0) >> (((forvar43 <= (8'h9e)) && {reg17}) ?
                          (reg65 ?
                              ((8'hab) ?
                                  reg36 : reg26) : forvar53) : reg54[(4'h9):(3'h5)]));
                    end
                  else
                    begin
                      reg87 <= reg12[(3'h5):(1'h1)];
                      reg88 <= $signed(({$signed(reg73)} && reg72[(4'ha):(1'h0)]));
                      reg89 <= reg60;
                    end
                end
            end
          else
            begin
              if ($unsigned(((~&$unsigned(reg22)) ?
                  (forvar37 ?
                      (reg61 + reg74) : $signed(forvar56)) : (reg74[(4'ha):(3'h6)] ?
                      $unsigned(forvar75) : forvar52[(4'h8):(3'h6)]))))
                begin
                  reg69 <= (^~reg18);
                  for (forvar70 = (1'h0); (forvar70 < (2'h2)); forvar70 = (forvar70 + (1'h1)))
                    begin
                      reg71 <= $unsigned(forvar8[(1'h0):(1'h0)]);
                      reg72 <= forvar40;
                      reg73 <= reg70;
                    end
                  for (forvar74 = (1'h0); (forvar74 < (2'h3)); forvar74 = (forvar74 + (1'h1)))
                    begin
                      reg75 <= $unsigned(reg70);
                      reg76 <= ($unsigned(reg9[(1'h0):(1'h0)]) ?
                          (~&(~&$signed(reg12))) : $unsigned($signed($unsigned(reg77))));
                      reg77 <= ((((reg11 == reg83) ?
                          (-reg49) : reg17) != (reg71[(3'h7):(3'h7)] >>> (~(8'hba)))) && forvar67[(3'h5):(1'h0)]);
                      reg78 <= $signed($signed($signed($unsigned(reg43))));
                    end
                end
              else
                begin
                  reg69 <= $signed($signed($unsigned(((8'hb0) >= reg18))));
                end
              if ($unsigned(((^reg23) ?
                  (reg40[(3'h4):(3'h4)] >>> (~^forvar6)) : (~(8'hb9)))))
                begin
                  if (((8'hab) ?
                      $unsigned($signed((+reg89))) : $unsigned((|$unsigned(reg17)))))
                    begin
                      reg79 <= (($signed((forvar67 && (8'ha3))) ?
                          reg35[(3'h6):(1'h0)] : reg58[(1'h1):(1'h0)]) < $unsigned(reg50));
                      reg80 <= $unsigned(reg13[(1'h1):(1'h0)]);
                      reg81 <= {$signed($unsigned((reg61 | reg71)))};
                      reg82 <= (!$signed({{reg7}}));
                    end
                  else
                    begin
                      reg79 <= ((~|reg85[(3'h4):(1'h0)]) * {{{forvar11}}});
                      reg80 <= ((~reg89) >>> ({(reg71 < reg16)} ?
                          reg85 : (~&$unsigned(reg76))));
                      reg81 <= $signed($unsigned((+((8'hb0) ? wire5 : reg70))));
                      reg82 <= $signed($signed(reg33[(1'h1):(1'h1)]));
                    end
                  if ({reg62[(3'h4):(2'h2)]})
                    begin
                      reg83 <= (reg23[(4'hb):(3'h4)] ?
                          (reg31 * forvar45) : {($signed(reg75) ?
                                  forvar74[(4'h9):(3'h4)] : $signed(reg76))});
                      reg84 <= (~(($signed(reg14) | forvar37) ?
                          {$signed(reg68)} : (8'ha1)));
                    end
                  else
                    begin
                      reg83 <= {$unsigned(((|reg32) ~^ (reg37 <= (8'hac))))};
                      reg84 <= $unsigned((~|$unsigned(forvar6)));
                      reg85 <= (((8'h9e) ?
                          reg23 : ((reg70 >> (8'hb6)) ?
                              {(8'hae)} : $signed(reg84))) ^ {{(&forvar86)}});
                    end
                  for (forvar86 = (1'h0); (forvar86 < (2'h3)); forvar86 = (forvar86 + (1'h1)))
                    begin
                      reg87 <= (+($signed($unsigned(reg63)) ?
                          $signed(reg23) : reg59[(2'h2):(1'h0)]));
                      reg88 <= $signed($signed((^wire5)));
                      reg89 <= $signed(reg52);
                      reg90 <= reg85;
                    end
                end
              else
                begin
                  for (forvar79 = (1'h0); (forvar79 < (1'h0)); forvar79 = (forvar79 + (1'h1)))
                    begin
                      reg80 <= $unsigned(forvar21[(2'h3):(1'h0)]);
                    end
                  if (reg23)
                    begin
                      reg81 <= $unsigned(reg30[(4'h9):(3'h5)]);
                    end
                  else
                    begin
                      reg81 <= ((forvar55 <= ((forvar76 ? reg44 : forvar21) ?
                              reg9 : $unsigned(forvar8))) ?
                          (~|(forvar75[(1'h0):(1'h0)] || (forvar7 ?
                              reg71 : reg78))) : (~^(^~$signed(forvar37))));
                      reg82 <= reg78[(2'h3):(1'h0)];
                    end
                end
              reg91 <= {({$signed(reg46)} && ((reg30 ? reg75 : reg19) ?
                      forvar43 : (forvar8 ? reg80 : reg17)))};
            end
          if ((|reg57[(1'h1):(1'h0)]))
            begin
              for (forvar92 = (1'h0); (forvar92 < (2'h2)); forvar92 = (forvar92 + (1'h1)))
                begin
                  reg93 <= ((^$signed((forvar7 << wire1))) < reg76[(4'h9):(1'h1)]);
                  for (forvar94 = (1'h0); (forvar94 < (1'h1)); forvar94 = (forvar94 + (1'h1)))
                    begin
                      reg95 <= (reg27 > reg69[(4'h8):(3'h7)]);
                      reg96 <= $signed((forvar52 ?
                          $unsigned($unsigned((8'hb0))) : reg56[(3'h6):(3'h6)]));
                    end
                  reg97 <= reg16[(4'hb):(1'h1)];
                end
              reg98 <= {wire2[(1'h1):(1'h0)]};
            end
          else
            begin
              for (forvar92 = (1'h0); (forvar92 < (2'h3)); forvar92 = (forvar92 + (1'h1)))
                begin
                  if (forvar74[(4'h9):(2'h3)])
                    begin
                      reg93 <= (-reg77[(3'h7):(2'h3)]);
                      reg94 <= {(8'ha3)};
                    end
                  else
                    begin
                      reg93 <= reg98;
                      reg94 <= reg79[(3'h4):(3'h4)];
                    end
                  if (reg45[(3'h7):(3'h4)])
                    begin
                      reg95 <= (reg23 > $signed($unsigned(reg41[(2'h3):(1'h1)])));
                      reg96 <= (~{$signed(reg18)});
                      reg97 <= reg41;
                      reg98 <= forvar86;
                    end
                  else
                    begin
                      reg95 <= $signed(reg69[(4'h8):(2'h3)]);
                    end
                  if (forvar69[(1'h0):(1'h0)])
                    begin
                      reg99 <= $unsigned(reg96);
                      reg100 <= $signed(({(reg69 ?
                              reg89 : reg95)} < reg72[(4'ha):(2'h2)]));
                      reg101 <= $unsigned((^~reg75[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg99 <= (^~(8'hb9));
                      reg100 <= (reg16[(2'h2):(1'h1)] ?
                          ((~(reg33 ? reg10 : (8'hb4))) ?
                              $unsigned((!reg39)) : $unsigned((forvar6 & forvar48))) : $signed(reg18));
                      reg101 <= (-(($signed(reg64) >>> (8'hba)) ^ reg68[(3'h7):(2'h3)]));
                    end
                end
              for (forvar102 = (1'h0); (forvar102 < (1'h1)); forvar102 = (forvar102 + (1'h1)))
                begin
                  if ((reg85[(4'ha):(2'h3)] <= (8'haf)))
                    begin
                      reg103 <= forvar94[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg103 <= (^(reg61[(1'h0):(1'h0)] && (^reg24)));
                      reg104 <= $signed(({$unsigned(reg58)} ?
                          {$unsigned(reg41)} : {forvar6[(1'h1):(1'h1)]}));
                      reg105 <= $signed((|reg99));
                    end
                  if ($unsigned($unsigned(forvar59[(1'h0):(1'h0)])))
                    begin
                      reg106 <= reg50;
                    end
                  else
                    begin
                      reg106 <= (reg55[(3'h6):(2'h2)] >>> reg23[(4'hc):(2'h2)]);
                      reg107 <= reg12[(4'h8):(2'h3)];
                      reg108 <= (^~reg33);
                    end
                  reg109 <= reg74;
                  for (forvar110 = (1'h0); (forvar110 < (2'h3)); forvar110 = (forvar110 + (1'h1)))
                    begin
                      reg111 <= $signed((!($signed(forvar110) ^ $unsigned(forvar39))));
                      reg112 <= ((~((reg33 ? reg71 : reg57) ?
                              (+reg73) : (-(8'ha8)))) ?
                          reg99[(4'h9):(2'h2)] : reg88[(3'h4):(1'h0)]);
                    end
                end
              for (forvar113 = (1'h0); (forvar113 < (1'h0)); forvar113 = (forvar113 + (1'h1)))
                begin
                  for (forvar114 = (1'h0); (forvar114 < (2'h3)); forvar114 = (forvar114 + (1'h1)))
                    begin
                      reg115 <= reg103;
                      reg116 <= ((8'hb8) ?
                          $unsigned($unsigned($signed(reg50))) : (8'ha6));
                      reg117 <= (~^(forvar102 ? $unsigned({(8'hb9)}) : reg13));
                    end
                  reg118 <= (^~(({(8'ha4)} & reg73) ?
                      reg84[(4'h9):(2'h2)] : forvar6));
                end
            end
          for (forvar119 = (1'h0); (forvar119 < (1'h0)); forvar119 = (forvar119 + (1'h1)))
            begin
              for (forvar120 = (1'h0); (forvar120 < (2'h2)); forvar120 = (forvar120 + (1'h1)))
                begin
                  if ((forvar11[(3'h6):(1'h0)] > ($unsigned(reg16) == $signed(reg31))))
                    begin
                      reg121 <= ((&$unsigned({reg9})) || $signed(((&reg47) ?
                          (forvar74 * reg39) : (forvar20 || reg84))));
                      reg122 <= reg41[(3'h5):(2'h3)];
                      reg123 <= (reg81 ?
                          (+(reg27[(4'h8):(3'h6)] ?
                              reg96 : $unsigned((8'ha9)))) : (reg63 ?
                              $unsigned((~forvar21)) : ({reg117} - {reg62})));
                      reg124 <= $signed(((!(~^reg76)) ?
                          ({reg99} ?
                              {forvar94} : (~|reg122)) : (forvar37[(4'h9):(3'h5)] ?
                              (8'ha9) : $signed((8'hb2)))));
                    end
                  else
                    begin
                      reg121 <= $unsigned((((forvar86 || forvar61) << $unsigned(reg53)) ?
                          $signed($signed(reg112)) : reg12[(2'h3):(1'h0)]));
                    end
                  for (forvar125 = (1'h0); (forvar125 < (1'h0)); forvar125 = (forvar125 + (1'h1)))
                    begin
                      reg126 <= (~|reg89);
                      reg127 <= ($signed({reg78[(2'h2):(2'h2)]}) ?
                          forvar102 : reg52);
                    end
                  if ({$signed($unsigned((!reg98)))})
                    begin
                      reg128 <= forvar69;
                    end
                  else
                    begin
                      reg128 <= reg69[(3'h7):(3'h4)];
                    end
                  for (forvar129 = (1'h0); (forvar129 < (1'h1)); forvar129 = (forvar129 + (1'h1)))
                    begin
                      reg130 <= ($unsigned(($signed(reg14) + reg44[(3'h5):(1'h0)])) ?
                          $unsigned(((forvar7 ?
                              reg46 : reg87) <= reg126[(3'h6):(3'h4)])) : ((-$unsigned(reg108)) ?
                              (reg95[(4'hb):(1'h1)] ?
                                  $signed(forvar69) : reg56) : $unsigned((8'hb4))));
                    end
                end
              for (forvar131 = (1'h0); (forvar131 < (1'h1)); forvar131 = (forvar131 + (1'h1)))
                begin
                  reg132 <= $unsigned({reg115});
                  for (forvar133 = (1'h0); (forvar133 < (2'h2)); forvar133 = (forvar133 + (1'h1)))
                    begin
                      reg134 <= (&(~|((forvar125 >> reg85) | reg55[(1'h0):(1'h0)])));
                      reg135 <= (reg71 ?
                          (($signed(reg121) && (reg93 ? reg115 : reg35)) ?
                              reg101 : ((forvar11 ^~ (8'hb4)) ?
                                  $signed(reg25) : reg29)) : {(reg80 * $signed(reg39))});
                      reg136 <= $unsigned((&((&reg94) ^~ $unsigned(reg29))));
                      reg137 <= (reg108 * {$unsigned($signed(reg107))});
                    end
                  if (reg62)
                    begin
                      reg138 <= reg69[(1'h1):(1'h1)];
                      reg139 <= $unsigned((reg59 | $unsigned($signed(reg34))));
                    end
                  else
                    begin
                      reg138 <= $signed(($unsigned((wire4 - reg37)) ?
                          reg33[(3'h7):(1'h1)] : (|(forvar92 >= forvar53))));
                      reg139 <= (^~({reg52} ^ $signed((~^(8'haf)))));
                    end
                  for (forvar140 = (1'h0); (forvar140 < (1'h1)); forvar140 = (forvar140 + (1'h1)))
                    begin
                      reg141 <= $unsigned(forvar37[(2'h2):(2'h2)]);
                      reg142 <= ((reg96 ?
                              reg101[(1'h0):(1'h0)] : (((8'ha7) | (8'hb9)) ?
                                  reg141[(1'h0):(1'h0)] : $unsigned((8'h9c)))) ?
                          forvar11 : (~$signed(reg45)));
                      reg143 <= ((8'ha6) ?
                          ($signed((^~reg106)) ?
                              (^(reg107 != reg83)) : forvar125[(2'h2):(1'h1)]) : (~^reg51[(4'ha):(3'h5)]));
                      reg144 <= forvar50[(3'h4):(1'h1)];
                    end
                end
              if ((&$unsigned(reg144[(3'h5):(3'h4)])))
                begin
                  reg145 <= reg104;
                end
              else
                begin
                  reg145 <= reg126;
                  reg146 <= $unsigned($unsigned(forvar53[(4'hc):(3'h5)]));
                  for (forvar147 = (1'h0); (forvar147 < (1'h0)); forvar147 = (forvar147 + (1'h1)))
                    begin
                      reg148 <= ((reg122 >> {$signed(reg42)}) ?
                          {(|reg74)} : reg138);
                      reg149 <= reg33;
                      reg150 <= ((forvar11 <= ($unsigned(forvar125) << forvar52[(2'h3):(2'h3)])) ^ $unsigned(($signed(reg89) ?
                          (reg9 ? reg27 : reg124) : $signed(reg87))));
                      reg151 <= (8'ha6);
                    end
                end
              reg152 <= $signed(forvar53);
            end
        end
      for (forvar153 = (1'h0); (forvar153 < (2'h3)); forvar153 = (forvar153 + (1'h1)))
        begin
          if (((8'hb0) == (reg66[(1'h0):(1'h0)] ?
              reg100[(2'h3):(1'h0)] : (^~(8'hb3)))))
            begin
              for (forvar154 = (1'h0); (forvar154 < (2'h3)); forvar154 = (forvar154 + (1'h1)))
                begin
                  for (forvar155 = (1'h0); (forvar155 < (2'h3)); forvar155 = (forvar155 + (1'h1)))
                    begin
                      reg156 <= forvar36;
                    end
                  for (forvar157 = (1'h0); (forvar157 < (1'h1)); forvar157 = (forvar157 + (1'h1)))
                    begin
                      reg158 <= reg41;
                    end
                  reg159 <= (~^(forvar59 ?
                      $signed(reg15[(2'h3):(2'h3)]) : (((8'hb7) ?
                          reg90 : wire5) + $unsigned(reg31))));
                end
            end
          else
            begin
              for (forvar154 = (1'h0); (forvar154 < (2'h3)); forvar154 = (forvar154 + (1'h1)))
                begin
                  for (forvar155 = (1'h0); (forvar155 < (1'h0)); forvar155 = (forvar155 + (1'h1)))
                    begin
                      reg156 <= $unsigned(($unsigned({(8'hba)}) ?
                          {$unsigned(forvar70)} : $unsigned((~reg148))));
                      reg157 <= forvar154[(4'hc):(2'h3)];
                      reg158 <= (~|(($unsigned(reg74) && $unsigned((8'hb3))) == ((wire4 <<< (8'ha1)) ?
                          (|(8'hb5)) : reg123[(3'h4):(1'h0)])));
                      reg159 <= (~^($unsigned(forvar45) != {reg55[(2'h2):(2'h2)]}));
                    end
                  for (forvar160 = (1'h0); (forvar160 < (2'h2)); forvar160 = (forvar160 + (1'h1)))
                    begin
                      reg161 <= (!$unsigned(($signed(reg72) ?
                          (reg25 ? reg33 : reg141) : (!reg58))));
                      reg162 <= (forvar119 ? forvar48 : reg99);
                      reg163 <= $signed(reg9);
                      reg164 <= ($unsigned($signed((8'ha4))) > ($unsigned((reg45 ?
                          (8'hb5) : reg63)) == (-{(8'hb7)})));
                    end
                  for (forvar165 = (1'h0); (forvar165 < (2'h2)); forvar165 = (forvar165 + (1'h1)))
                    begin
                      reg166 <= $unsigned((~|((reg89 || reg22) - (!reg34))));
                      reg167 <= $unsigned(({$unsigned(reg52)} ?
                          reg27[(4'h9):(2'h3)] : (~^(wire3 ?
                              forvar92 : (8'hb8)))));
                    end
                  for (forvar168 = (1'h0); (forvar168 < (1'h1)); forvar168 = (forvar168 + (1'h1)))
                    begin
                      reg169 <= $signed(((~|(reg23 || (8'haa))) ?
                          forvar64[(4'h9):(4'h9)] : $signed((reg31 ?
                              reg106 : (8'haa)))));
                      reg170 <= (($unsigned($signed((8'hb2))) ?
                              ((reg128 >>> reg149) ^ $signed(reg72)) : ((forvar39 ?
                                  (8'ha7) : (8'had)) >= {forvar131})) ?
                          {(8'haa)} : reg107);
                      reg171 <= reg52[(3'h4):(1'h1)];
                      reg172 <= reg24;
                    end
                end
              reg173 <= ((8'hb4) | (forvar8 ?
                  $signed((~&reg79)) : forvar39[(3'h4):(1'h0)]));
              for (forvar174 = (1'h0); (forvar174 < (1'h0)); forvar174 = (forvar174 + (1'h1)))
                begin
                  if ((-(reg127 ?
                      ((+reg65) * $unsigned((8'ha1))) : (-$signed(reg171)))))
                    begin
                      reg175 <= (~reg56);
                      reg176 <= reg72[(3'h7):(3'h7)];
                      reg177 <= (forvar165 ?
                          (reg175 ^ ({reg60} != $unsigned(reg115))) : ($signed(forvar64) <<< ($signed((8'ha1)) <<< reg9)));
                    end
                  else
                    begin
                      reg175 <= reg148[(4'ha):(4'ha)];
                      reg176 <= (((wire0[(1'h0):(1'h0)] >= {forvar92}) ?
                          ((reg130 ?
                              reg66 : reg97) >>> (reg65 | reg148)) : {(reg18 ?
                                  reg115 : reg36)}) <<< $unsigned({(forvar119 == reg111)}));
                      reg177 <= {reg97[(1'h1):(1'h1)]};
                    end
                end
            end
          if ($signed((^((8'hb1) ? $signed(reg50) : $unsigned((8'ha9))))))
            begin
              for (forvar178 = (1'h0); (forvar178 < (2'h3)); forvar178 = (forvar178 + (1'h1)))
                begin
                  for (forvar179 = (1'h0); (forvar179 < (2'h2)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= $unsigned(reg93);
                      reg181 <= (!reg51[(3'h4):(3'h4)]);
                    end
                  reg182 <= (-forvar174[(1'h1):(1'h0)]);
                end
              if ($signed((^forvar48[(1'h1):(1'h1)])))
                begin
                  for (forvar183 = (1'h0); (forvar183 < (1'h1)); forvar183 = (forvar183 + (1'h1)))
                    begin
                      reg184 <= ((reg57[(3'h7):(3'h7)] ?
                          $signed(reg45) : $signed($unsigned(reg169))) ^ {{reg173[(3'h4):(2'h3)]}});
                      reg185 <= forvar140[(1'h0):(1'h0)];
                    end
                  for (forvar186 = (1'h0); (forvar186 < (1'h1)); forvar186 = (forvar186 + (1'h1)))
                    begin
                      reg187 <= ((|reg182[(3'h5):(3'h5)]) ?
                          (^reg181[(1'h0):(1'h0)]) : (!reg19[(4'hd):(3'h4)]));
                      reg188 <= ((!reg152) ^ ((+(reg118 ? reg143 : forvar165)) ?
                          (-reg187[(4'h8):(3'h7)]) : (reg24 ?
                              (reg27 == reg143) : (forvar168 | reg44))));
                      reg189 <= (^(8'ha6));
                      reg190 <= (+$unsigned(({forvar45} >>> $unsigned(reg144))));
                    end
                end
              else
                begin
                  for (forvar183 = (1'h0); (forvar183 < (1'h0)); forvar183 = (forvar183 + (1'h1)))
                    begin
                      reg184 <= (~&($signed(reg23[(4'h9):(1'h1)]) | reg115));
                      reg185 <= (($signed((-reg59)) ?
                              (~|(reg64 ? forvar8 : reg76)) : (8'hb6)) ?
                          $unsigned({forvar56[(1'h0):(1'h0)]}) : $signed(reg148));
                      reg186 <= (($signed((reg108 - reg158)) < $signed((reg158 ?
                              reg31 : reg50))) ?
                          $signed((8'hb5)) : ($signed($unsigned(forvar155)) ?
                              {(reg18 <= forvar133)} : reg136[(4'hb):(3'h5)]));
                    end
                  reg187 <= reg54;
                  for (forvar188 = (1'h0); (forvar188 < (1'h0)); forvar188 = (forvar188 + (1'h1)))
                    begin
                      reg189 <= ((reg157 ?
                              reg103[(3'h4):(2'h3)] : $signed({reg71})) ?
                          $signed($signed((reg95 + reg73))) : forvar113[(1'h1):(1'h1)]);
                      reg190 <= ((forvar40[(4'h9):(1'h0)] << {$unsigned(forvar7)}) ^ $unsigned(reg111));
                      reg191 <= {$signed((^~(+forvar53)))};
                      reg192 <= (((~&reg139) ?
                          ((reg33 ? reg189 : forvar155) ?
                              (forvar6 || forvar43) : ((8'ha9) >= reg17)) : {$signed((8'hb2))}) || $signed(reg29));
                    end
                  for (forvar193 = (1'h0); (forvar193 < (1'h0)); forvar193 = (forvar193 + (1'h1)))
                    begin
                      reg194 <= forvar61[(2'h2):(1'h0)];
                      reg195 <= $unsigned(($unsigned((reg136 >= reg33)) ?
                          {(~&forvar113)} : reg116[(1'h0):(1'h0)]));
                      reg196 <= forvar155;
                      reg197 <= reg72[(4'he):(4'h8)];
                    end
                end
              for (forvar198 = (1'h0); (forvar198 < (2'h2)); forvar198 = (forvar198 + (1'h1)))
                begin
                  reg199 <= $signed(reg181);
                  reg200 <= (+forvar174[(2'h2):(1'h1)]);
                  for (forvar201 = (1'h0); (forvar201 < (2'h2)); forvar201 = (forvar201 + (1'h1)))
                    begin
                      reg202 <= ({{$signed(reg127)}} ?
                          reg40[(2'h3):(1'h0)] : $signed(reg181[(4'ha):(3'h4)]));
                      reg203 <= $signed(reg103);
                      reg204 <= ($unsigned((&(~&reg203))) >= reg82);
                      reg205 <= $signed((8'ha9));
                    end
                end
              for (forvar206 = (1'h0); (forvar206 < (1'h1)); forvar206 = (forvar206 + (1'h1)))
                begin
                  reg207 <= reg99;
                  reg208 <= (reg141[(2'h2):(2'h2)] ?
                      (~&$unsigned(reg89)) : (reg40 <<< $unsigned($unsigned(reg176))));
                  reg209 <= $unsigned({(((8'ha2) | (8'hac)) ?
                          (forvar188 & reg51) : $unsigned((8'ha4)))});
                end
            end
          else
            begin
              if ($unsigned((^~(^$unsigned(reg116)))))
                begin
                  if ($unsigned((reg16 ^~ (~&(reg182 ? forvar125 : reg73)))))
                    begin
                      reg178 <= ({((reg203 ? reg91 : reg22) > reg167)} ?
                          $signed((forvar20[(3'h5):(3'h4)] ?
                              $signed(reg11) : reg170)) : reg97[(4'h9):(4'h8)]);
                    end
                  else
                    begin
                      reg178 <= (|(({reg40} ?
                              reg151 : (reg74 ? forvar56 : forvar201)) ?
                          (~&$signed((8'haf))) : ($signed((8'h9c)) == (^forvar69))));
                    end
                  if ($unsigned((|reg30)))
                    begin
                      reg179 <= $signed((reg107 * reg77[(3'h4):(2'h3)]));
                      reg180 <= ($signed($unsigned((reg202 ?
                          reg97 : reg172))) ~^ reg65);
                    end
                  else
                    begin
                      reg179 <= reg187[(4'hb):(3'h4)];
                      reg180 <= $signed(((^(reg181 && forvar125)) | (~|$signed(reg99))));
                    end
                  if (reg132[(3'h5):(3'h4)])
                    begin
                      reg181 <= {(reg122 << ((~&reg112) < (^reg68)))};
                      reg182 <= (reg98 >= forvar168[(1'h0):(1'h0)]);
                      reg183 <= ($signed(((reg90 != (8'hac)) ?
                              (forvar53 >= reg163) : $unsigned(reg112))) ?
                          {((forvar157 ?
                                  forvar64 : reg54) ^ reg192)} : {$unsigned((^reg203))});
                    end
                  else
                    begin
                      reg181 <= (~^reg77[(2'h2):(2'h2)]);
                      reg182 <= forvar154;
                    end
                end
              else
                begin
                  reg178 <= reg123[(1'h1):(1'h1)];
                  for (forvar179 = (1'h0); (forvar179 < (1'h1)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= $signed($unsigned((8'ha9)));
                      reg181 <= $unsigned(($unsigned(((8'hb6) * reg149)) ?
                          $unsigned((reg76 < (8'h9f))) : (|reg151[(3'h5):(3'h5)])));
                      reg182 <= ($unsigned(reg143) & reg47[(2'h2):(2'h2)]);
                    end
                  reg183 <= ($unsigned(((reg151 ? forvar69 : reg175) ?
                          (reg149 ? forvar110 : (8'hb0)) : reg163)) ?
                      (wire3 ~^ $unsigned(reg204[(3'h4):(1'h0)])) : (((reg72 ?
                              (8'h9f) : forvar94) ?
                          (^~reg192) : (8'hb0)) + ((~^(8'h9e)) < $unsigned(reg63))));
                end
              for (forvar184 = (1'h0); (forvar184 < (2'h3)); forvar184 = (forvar184 + (1'h1)))
                begin
                  for (forvar185 = (1'h0); (forvar185 < (1'h0)); forvar185 = (forvar185 + (1'h1)))
                    begin
                      reg186 <= reg69[(4'hf):(2'h2)];
                      reg187 <= forvar70;
                      reg188 <= $unsigned((((~^reg76) - (reg134 ?
                              wire4 : reg51)) ?
                          (^(forvar92 ?
                              reg203 : forvar6)) : (&$signed(reg171))));
                    end
                  reg189 <= reg209;
                end
              if (reg72)
                begin
                  if (({reg33[(3'h7):(1'h0)]} ?
                      reg156[(2'h2):(1'h1)] : $signed({((8'had) ?
                              forvar120 : reg132)})))
                    begin
                      reg190 <= (reg7 ? reg122 : (!forvar110));
                      reg191 <= forvar40;
                      reg192 <= ((~&($unsigned(reg23) <= $unsigned(reg138))) ?
                          (($signed(reg207) < (reg138 ? reg55 : reg182)) ?
                              reg75 : {forvar61}) : {$unsigned(forvar59)});
                      reg193 <= (reg82[(2'h2):(1'h1)] ?
                          reg98[(2'h3):(2'h3)] : reg179);
                    end
                  else
                    begin
                      reg190 <= (&forvar40[(3'h6):(3'h4)]);
                      reg191 <= reg190[(2'h2):(1'h0)];
                    end
                  if (({reg98} <<< $signed(reg65)))
                    begin
                      reg194 <= $unsigned(wire0);
                      reg195 <= reg170;
                    end
                  else
                    begin
                      reg194 <= forvar64[(4'hf):(2'h2)];
                      reg195 <= $unsigned(reg190[(1'h1):(1'h0)]);
                      reg196 <= reg79[(3'h7):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar190 = (1'h0); (forvar190 < (2'h2)); forvar190 = (forvar190 + (1'h1)))
                    begin
                      reg191 <= $signed((~^(reg146[(3'h7):(3'h6)] ?
                          reg25[(4'ha):(1'h0)] : (forvar69 ? reg16 : reg204))));
                      reg192 <= ({reg115} ?
                          $unsigned(forvar55[(3'h4):(1'h0)]) : $unsigned(($signed(forvar198) ?
                              $unsigned(reg41) : (reg175 <= forvar56))));
                      reg193 <= $unsigned($unsigned(reg37));
                    end
                  for (forvar194 = (1'h0); (forvar194 < (1'h1)); forvar194 = (forvar194 + (1'h1)))
                    begin
                      reg195 <= (reg87 >= (!$unsigned((forvar59 ?
                          (8'hb7) : reg32))));
                      reg196 <= ({((reg87 ~^ wire5) ^ $unsigned((8'ha6)))} <<< $signed($unsigned((reg185 ?
                          reg68 : (8'hac)))));
                    end
                end
              for (forvar197 = (1'h0); (forvar197 < (2'h3)); forvar197 = (forvar197 + (1'h1)))
                begin
                  if ((~^$signed((^(^forvar75)))))
                    begin
                      reg198 <= reg18[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg198 <= $unsigned(reg41);
                      reg199 <= $unsigned({reg100[(3'h4):(3'h4)]});
                      reg200 <= $signed($signed($signed({forvar64})));
                    end
                  if ($signed($unsigned(((reg95 == reg12) ?
                      (-reg204) : forvar20))))
                    begin
                      reg201 <= $signed(($unsigned(reg22[(2'h2):(1'h0)]) <<< forvar197[(1'h1):(1'h0)]));
                      reg202 <= reg31[(2'h2):(2'h2)];
                      reg203 <= ($unsigned((forvar64[(1'h1):(1'h0)] < (8'ha3))) != reg106);
                      reg204 <= (&((reg44[(3'h7):(2'h2)] <<< reg59) << ((^~reg194) ?
                          $signed(forvar113) : $unsigned(forvar70))));
                    end
                  else
                    begin
                      reg201 <= ((^(+$unsigned((8'ha7)))) ?
                          reg85 : ({(reg53 < forvar11)} + (~^$unsigned(forvar56))));
                      reg202 <= (|((forvar193 <= (~^reg179)) <= ((+forvar178) ?
                          reg197 : forvar74[(3'h7):(3'h5)])));
                      reg203 <= $unsigned($signed(reg195));
                      reg204 <= reg37;
                    end
                  if ({$unsigned((((8'haa) - (8'hb9)) >= (reg78 ?
                          (8'ha7) : forvar125)))})
                    begin
                      reg205 <= $unsigned((~&(reg171[(2'h3):(2'h3)] <= (reg128 ?
                          forvar190 : (8'ha2)))));
                    end
                  else
                    begin
                      reg205 <= forvar125[(3'h7):(1'h0)];
                      reg206 <= reg204;
                    end
                  if (($unsigned((forvar86 - {forvar125})) ?
                      $unsigned(reg127) : reg141[(1'h1):(1'h1)]))
                    begin
                      reg207 <= reg31[(2'h2):(2'h2)];
                      reg208 <= ($unsigned(reg198) ?
                          forvar56 : (~^(!$unsigned(reg181))));
                      reg209 <= forvar86[(3'h4):(2'h3)];
                      reg210 <= ((~$unsigned($signed(reg32))) ?
                          reg152[(3'h7):(3'h7)] : reg44[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg207 <= forvar69;
                      reg208 <= $signed({reg33});
                      reg209 <= reg161[(2'h2):(1'h1)];
                    end
                end
            end
          if ({reg182[(3'h5):(2'h2)]})
            begin
              if (reg74)
                begin
                  for (forvar211 = (1'h0); (forvar211 < (1'h1)); forvar211 = (forvar211 + (1'h1)))
                    begin
                      reg212 <= reg203;
                      reg213 <= reg17[(1'h0):(1'h0)];
                    end
                  if (reg109)
                    begin
                      reg214 <= $signed((reg141 || ((|reg127) ~^ (~^(8'hb2)))));
                    end
                  else
                    begin
                      reg214 <= {(^{(&reg54)})};
                      reg215 <= reg12[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  reg211 <= {reg150[(1'h1):(1'h1)]};
                end
              for (forvar216 = (1'h0); (forvar216 < (1'h1)); forvar216 = (forvar216 + (1'h1)))
                begin
                  if ($signed(reg164[(3'h6):(3'h6)]))
                    begin
                      reg217 <= ($unsigned($unsigned($signed(forvar193))) ?
                          $unsigned($signed(reg54[(4'hc):(3'h4)])) : $unsigned(($unsigned(reg127) ?
                              forvar179 : forvar52)));
                      reg218 <= reg157;
                      reg219 <= ((-reg122[(1'h0):(1'h0)]) << ($unsigned({reg98}) << $signed((8'ha3))));
                    end
                  else
                    begin
                      reg217 <= {(($signed(reg184) + {reg57}) ?
                              (reg198 ~^ (^~reg186)) : (~^(reg135 <<< reg105)))};
                      reg218 <= reg192[(3'h6):(3'h6)];
                    end
                  for (forvar220 = (1'h0); (forvar220 < (2'h3)); forvar220 = (forvar220 + (1'h1)))
                    begin
                      reg221 <= forvar92[(3'h6):(3'h4)];
                    end
                end
            end
          else
            begin
              for (forvar211 = (1'h0); (forvar211 < (2'h3)); forvar211 = (forvar211 + (1'h1)))
                begin
                  if (forvar39)
                    begin
                      reg212 <= (~|(~^((reg85 ~^ forvar198) ?
                          $signed((8'ha1)) : (forvar40 ? reg52 : reg169))));
                      reg213 <= (8'h9e);
                    end
                  else
                    begin
                      reg212 <= $unsigned((-reg206[(1'h1):(1'h0)]));
                      reg213 <= $signed(reg88);
                    end
                  for (forvar214 = (1'h0); (forvar214 < (1'h0)); forvar214 = (forvar214 + (1'h1)))
                    begin
                      reg215 <= (~&(~&$signed((^~reg103))));
                      reg216 <= {reg80};
                      reg217 <= forvar174;
                    end
                end
              if (reg50[(1'h1):(1'h1)])
                begin
                  reg218 <= (~&(~$signed(((8'hac) ? reg75 : reg126))));
                end
              else
                begin
                  for (forvar218 = (1'h0); (forvar218 < (1'h1)); forvar218 = (forvar218 + (1'h1)))
                    begin
                      reg219 <= (8'hb5);
                    end
                  if (reg214)
                    begin
                      reg220 <= ((~&forvar102[(1'h1):(1'h1)]) ?
                          (8'hb1) : ({(^reg94)} == (reg122 ^ reg136)));
                      reg221 <= $unsigned(reg189);
                      reg222 <= ((($signed(forvar201) ?
                          forvar40[(4'hd):(4'hd)] : reg11) && {$unsigned(reg204)}) | $unsigned(reg176));
                      reg223 <= (reg81 ?
                          (reg148[(4'hc):(4'h8)] + reg162[(3'h7):(3'h4)]) : ($unsigned((&reg96)) ?
                              ((forvar45 | forvar179) ?
                                  ((8'ha2) ?
                                      (8'ha9) : reg222) : (reg51 != (8'hb7))) : forvar185));
                    end
                  else
                    begin
                      reg220 <= $unsigned($signed((reg106 >= {reg211})));
                      reg221 <= ($signed(reg163) ^~ $signed((reg109 ?
                          (+reg76) : (^reg152))));
                    end
                end
              for (forvar224 = (1'h0); (forvar224 < (2'h2)); forvar224 = (forvar224 + (1'h1)))
                begin
                  reg225 <= (^((&forvar92) ^~ reg183[(3'h5):(1'h0)]));
                  if ($unsigned((reg132[(4'ha):(4'ha)] ?
                      $unsigned(reg176[(1'h0):(1'h0)]) : (8'haf))))
                    begin
                      reg226 <= reg126;
                      reg227 <= reg218[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg226 <= {reg91};
                    end
                  reg228 <= forvar67;
                  if (reg22)
                    begin
                      reg229 <= $unsigned(reg135);
                      reg230 <= reg156;
                    end
                  else
                    begin
                      reg229 <= {$signed(((forvar50 ? reg192 : (8'hac)) ?
                              {reg118} : $unsigned(reg191)))};
                      reg230 <= (reg38[(4'hc):(4'ha)] ?
                          $unsigned(forvar125[(3'h5):(2'h3)]) : ($unsigned(((8'hba) | reg141)) | reg136));
                      reg231 <= {($unsigned(reg60) ?
                              (~^$unsigned(reg94)) : (^~reg116))};
                    end
                end
              for (forvar232 = (1'h0); (forvar232 < (1'h0)); forvar232 = (forvar232 + (1'h1)))
                begin
                  for (forvar233 = (1'h0); (forvar233 < (1'h0)); forvar233 = (forvar233 + (1'h1)))
                    begin
                      reg234 <= (^~$unsigned((~(~^reg49))));
                      reg235 <= $signed(forvar147);
                      reg236 <= reg132;
                    end
                  if (($unsigned(($unsigned(reg19) & reg60)) - $unsigned({$unsigned(reg204)})))
                    begin
                      reg237 <= reg123;
                      reg238 <= reg230[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg237 <= reg199[(2'h2):(1'h1)];
                      reg238 <= (&$unsigned((reg75 >>> $signed(reg64))));
                      reg239 <= forvar67[(1'h0):(1'h0)];
                      reg240 <= forvar69;
                    end
                end
            end
        end
    end
  assign wire241 = (8'ha5);
  assign wire242 = $unsigned(((reg126[(3'h5):(1'h0)] && {reg44}) > (8'hb9)));
  always
    @(posedge clk) begin
      if ((($unsigned((reg42 && (8'ha2))) * reg35[(2'h2):(1'h1)]) ?
          $unsigned(wire242) : (reg23 ?
              ((forvar6 ? forvar232 : reg77) ?
                  reg187 : (^reg195)) : {reg99[(4'h9):(1'h1)]})))
        begin
          for (forvar243 = (1'h0); (forvar243 < (1'h0)); forvar243 = (forvar243 + (1'h1)))
            begin
              for (forvar244 = (1'h0); (forvar244 < (2'h2)); forvar244 = (forvar244 + (1'h1)))
                begin
                  for (forvar245 = (1'h0); (forvar245 < (2'h2)); forvar245 = (forvar245 + (1'h1)))
                    begin
                      reg246 <= forvar165;
                    end
                  reg247 <= ($unsigned((8'ha9)) ?
                      {$signed($unsigned(wire2))} : reg202[(1'h1):(1'h1)]);
                  for (forvar248 = (1'h0); (forvar248 < (1'h1)); forvar248 = (forvar248 + (1'h1)))
                    begin
                      reg249 <= forvar11[(3'h6):(3'h5)];
                    end
                  for (forvar250 = (1'h0); (forvar250 < (2'h3)); forvar250 = (forvar250 + (1'h1)))
                    begin
                      reg251 <= ((~|$unsigned((-forvar178))) && wire5);
                      reg252 <= reg137;
                      reg253 <= $signed({$unsigned((^reg76))});
                      reg254 <= reg116;
                    end
                end
            end
        end
      else
        begin
          for (forvar243 = (1'h0); (forvar243 < (2'h2)); forvar243 = (forvar243 + (1'h1)))
            begin
              if ($unsigned((&$unsigned((reg183 + (8'ha3))))))
                begin
                  for (forvar244 = (1'h0); (forvar244 < (2'h3)); forvar244 = (forvar244 + (1'h1)))
                    begin
                      reg245 <= ($signed(reg33[(1'h1):(1'h1)]) - {reg17[(3'h6):(2'h2)]});
                    end
                  if ($signed(forvar155))
                    begin
                      reg246 <= reg31;
                      reg247 <= (8'ha5);
                      reg248 <= (~|reg238);
                      reg249 <= $unsigned(($signed(forvar220) - ((+reg78) ?
                          (~&reg175) : (reg218 ? reg229 : forvar133))));
                    end
                  else
                    begin
                      reg246 <= (^$unsigned($signed($unsigned(reg164))));
                      reg247 <= (|$unsigned(((~&reg97) ?
                          {forvar79} : (forvar74 ? (8'hb0) : (8'haa)))));
                      reg248 <= $unsigned((~&($unsigned(reg30) ?
                          $signed((8'hb4)) : (+reg10))));
                      reg249 <= ((&($signed(reg228) ?
                              reg202[(3'h4):(2'h2)] : {reg77})) ?
                          {(((8'hb9) && forvar45) ?
                                  (reg122 ?
                                      (8'ha8) : reg190) : reg18[(3'h4):(3'h4)])} : reg195[(1'h0):(1'h0)]);
                    end
                  for (forvar250 = (1'h0); (forvar250 < (1'h0)); forvar250 = (forvar250 + (1'h1)))
                    begin
                      reg251 <= (&(^$signed((reg230 ~^ reg180))));
                      reg252 <= $unsigned((reg137 - (forvar198 >= forvar133)));
                      reg253 <= $signed((((reg235 - wire241) << {forvar198}) ?
                          $signed(reg204) : $unsigned($signed((8'hb3)))));
                    end
                end
              else
                begin
                  if ((reg7[(3'h5):(3'h4)] ?
                      (({forvar188} ? $signed(reg9) : $unsigned(forvar220)) ?
                          forvar69[(3'h4):(3'h4)] : (reg145[(3'h6):(1'h1)] <= reg58)) : $signed($signed(reg247))))
                    begin
                      reg244 <= reg226;
                      reg245 <= $signed($unsigned(($signed((8'ha3)) ?
                          reg42 : $signed(reg148))));
                      reg246 <= $unsigned(($signed($unsigned(forvar129)) && (forvar140[(2'h2):(1'h1)] ?
                          wire2[(1'h1):(1'h1)] : $signed(forvar36))));
                    end
                  else
                    begin
                      reg244 <= $unsigned({$signed((^forvar125))});
                      reg245 <= ($unsigned(forvar94[(2'h3):(2'h3)]) > ((~&(forvar248 ?
                          reg61 : (8'ha6))) & (~forvar43)));
                    end
                  if ((reg83[(1'h0):(1'h0)] ?
                      (reg121 ?
                          $unsigned((8'hb4)) : $unsigned(reg185[(3'h4):(1'h0)])) : $unsigned((^(reg247 ?
                          reg123 : (8'h9f))))))
                    begin
                      reg247 <= (&reg186);
                      reg248 <= {$unsigned(((wire242 & reg35) ?
                              $unsigned(forvar183) : {reg171}))};
                      reg249 <= reg195;
                      reg250 <= (~(forvar183[(4'h8):(3'h4)] ?
                          reg77[(3'h5):(3'h5)] : forvar131[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg247 <= reg88;
                    end
                end
              for (forvar254 = (1'h0); (forvar254 < (1'h0)); forvar254 = (forvar254 + (1'h1)))
                begin
                  for (forvar255 = (1'h0); (forvar255 < (1'h1)); forvar255 = (forvar255 + (1'h1)))
                    begin
                      reg256 <= reg36;
                      reg257 <= (((~(forvar79 ? wire4 : reg152)) > (~((8'haa) ?
                              reg100 : reg28))) ?
                          (forvar211 ?
                              reg167[(2'h2):(2'h2)] : (|(|(8'hb4)))) : ((forvar21 != (~|(8'hac))) ?
                              $unsigned((forvar188 << (8'hb9))) : ($signed(reg40) < forvar79[(1'h0):(1'h0)])));
                      reg258 <= ((($signed(reg203) <= $signed((8'had))) ~^ (reg207[(1'h0):(1'h0)] ?
                              reg45 : (~reg10))) ?
                          $unsigned(($unsigned(reg144) ?
                              forvar86[(3'h7):(2'h2)] : $signed(reg229))) : $signed(($signed(forvar211) & $unsigned(reg42))));
                      reg259 <= (reg225 ~^ (8'hb4));
                    end
                  for (forvar260 = (1'h0); (forvar260 < (2'h2)); forvar260 = (forvar260 + (1'h1)))
                    begin
                      reg261 <= $unsigned($signed({$unsigned((8'ha4))}));
                    end
                end
            end
          if ({$unsigned(forvar59)})
            begin
              if (reg12[(3'h5):(1'h0)])
                begin
                  reg262 <= ((((8'hb4) ?
                      reg136[(4'ha):(3'h7)] : $unsigned(reg57)) ^ $signed($unsigned(reg24))) >> ((&reg208) ?
                      $unsigned({forvar125}) : (-(^reg209))));
                  for (forvar263 = (1'h0); (forvar263 < (2'h2)); forvar263 = (forvar263 + (1'h1)))
                    begin
                      reg264 <= {$signed(((reg247 + reg96) ?
                              (reg66 ? reg180 : (8'h9f)) : (reg69 & reg15)))};
                    end
                  if (forvar185)
                    begin
                      reg265 <= (|((~&(+(8'hb8))) ^~ $unsigned(reg91[(3'h5):(1'h1)])));
                    end
                  else
                    begin
                      reg265 <= (forvar244[(4'hb):(3'h6)] ?
                          reg261[(1'h0):(1'h0)] : {reg161[(3'h4):(1'h0)]});
                    end
                end
              else
                begin
                  if (((forvar40[(4'hb):(3'h7)] ?
                      ((&reg64) ?
                          reg115 : reg157) : $signed((8'h9c))) || reg158))
                    begin
                      reg262 <= $unsigned(($unsigned(reg192) ?
                          (-(reg88 >> reg60)) : reg37));
                      reg263 <= ((~reg27[(3'h5):(3'h4)]) + (forvar211[(1'h1):(1'h1)] ?
                          reg244[(1'h0):(1'h0)] : $signed($unsigned(reg208))));
                    end
                  else
                    begin
                      reg262 <= reg89[(1'h0):(1'h0)];
                      reg263 <= $unsigned(($unsigned($signed(reg157)) ?
                          (~|$unsigned(forvar102)) : reg45));
                      reg264 <= reg162;
                      reg265 <= $signed((~$signed((reg172 + forvar184))));
                    end
                  reg266 <= reg79[(2'h3):(2'h2)];
                  reg267 <= (~&(($unsigned(reg205) | reg36[(3'h7):(2'h2)]) == ({reg19} && (~|forvar197))));
                end
              for (forvar268 = (1'h0); (forvar268 < (1'h0)); forvar268 = (forvar268 + (1'h1)))
                begin
                  for (forvar269 = (1'h0); (forvar269 < (1'h0)); forvar269 = (forvar269 + (1'h1)))
                    begin
                      reg270 <= reg210;
                      reg271 <= wire1;
                      reg272 <= $unsigned($signed({reg75[(3'h6):(1'h0)]}));
                    end
                  if ($signed((reg252 >= forvar243[(2'h2):(1'h1)])))
                    begin
                      reg273 <= $signed((~^$signed((8'ha5))));
                      reg274 <= ($signed(($unsigned(reg261) ?
                              (reg231 ^~ reg58) : (^reg112))) ?
                          ($unsigned(forvar268) ~^ (+(|reg17))) : (((~reg217) | $signed(reg248)) ?
                              (-$unsigned(reg220)) : ($unsigned((8'h9e)) ?
                                  reg239 : ((8'ha7) < reg158))));
                    end
                  else
                    begin
                      reg273 <= ((+$unsigned((reg245 >= (8'ha9)))) << ((&(|reg183)) < reg150));
                      reg274 <= {($unsigned((!reg175)) ?
                              ($signed(reg198) ?
                                  $signed(reg116) : {reg162}) : $signed(reg73))};
                      reg275 <= {(^(!(~^reg173)))};
                    end
                end
              if (((((^reg91) ?
                  (~|(8'h9e)) : (reg135 | wire241)) - $unsigned(((8'haf) == (8'ha9)))) * ($signed((^~reg230)) > reg136[(4'hb):(1'h0)])))
                begin
                  if ($unsigned((((~^reg183) ^ (^~forvar178)) ?
                      (^reg151) : (~&(reg22 ? forvar220 : forvar155)))))
                    begin
                      reg276 <= (8'hb2);
                      reg277 <= {$unsigned(($unsigned((8'haf)) ?
                              reg36[(3'h7):(3'h5)] : reg41[(2'h3):(1'h0)]))};
                      reg278 <= $unsigned({{reg18[(2'h3):(2'h3)]}});
                      reg279 <= (~|$unsigned($signed((forvar69 ?
                          reg12 : reg208))));
                    end
                  else
                    begin
                      reg276 <= (reg208[(1'h1):(1'h1)] && ($signed((8'hb5)) ?
                          ($unsigned(wire241) >> {reg151}) : {forvar157}));
                    end
                end
              else
                begin
                  if (($unsigned(reg262[(3'h6):(2'h2)]) ?
                      reg58 : (-$signed(reg274[(1'h0):(1'h0)]))))
                    begin
                      reg276 <= (|$signed(((reg231 ?
                          reg30 : (8'hb0)) | $signed(reg271))));
                      reg277 <= (~&((reg193[(2'h2):(1'h0)] & $signed(reg259)) | ((reg107 ?
                              reg195 : forvar129) ?
                          $unsigned(forvar61) : reg9)));
                      reg278 <= wire3[(1'h1):(1'h0)];
                      reg279 <= (~{forvar154});
                    end
                  else
                    begin
                      reg276 <= {(|(~&forvar255))};
                      reg277 <= $unsigned(reg263);
                    end
                  if ($signed(reg85[(3'h7):(1'h1)]))
                    begin
                      reg280 <= $unsigned(((8'hb9) & $signed($unsigned(reg35))));
                    end
                  else
                    begin
                      reg280 <= $signed(forvar232);
                      reg281 <= {(($unsigned((8'hb7)) <<< (forvar248 ?
                                  (8'hab) : (8'hb8))) ?
                              forvar119[(4'h8):(1'h1)] : forvar147[(4'he):(1'h0)])};
                    end
                end
              reg282 <= ($unsigned(reg211[(2'h3):(1'h0)]) ?
                  (^~$unsigned(reg36[(4'h8):(3'h6)])) : forvar64);
            end
          else
            begin
              if (forvar7[(4'ha):(1'h1)])
                begin
                  for (forvar262 = (1'h0); (forvar262 < (2'h2)); forvar262 = (forvar262 + (1'h1)))
                    begin
                      reg263 <= reg205;
                      reg264 <= $signed($unsigned($unsigned((reg7 + forvar244))));
                      reg265 <= reg263;
                    end
                end
              else
                begin
                  for (forvar262 = (1'h0); (forvar262 < (1'h0)); forvar262 = (forvar262 + (1'h1)))
                    begin
                      reg263 <= $signed($unsigned(reg196[(4'ha):(3'h4)]));
                      reg264 <= (^~(reg246[(3'h5):(2'h3)] ?
                          ($signed(reg77) >>> reg85) : forvar61));
                    end
                end
              reg266 <= $signed(reg206[(1'h1):(1'h1)]);
              if ($unsigned(forvar6[(4'he):(3'h6)]))
                begin
                  for (forvar267 = (1'h0); (forvar267 < (2'h2)); forvar267 = (forvar267 + (1'h1)))
                    begin
                      reg268 <= ($signed(((forvar198 >>> reg103) ?
                              reg214 : (+(8'ha6)))) ?
                          forvar147[(1'h0):(1'h0)] : $signed(((~|forvar211) ?
                              (&reg279) : (!reg9))));
                      reg269 <= (wire2 && (forvar262 && ((|reg116) ?
                          $unsigned(forvar45) : $unsigned(reg178))));
                      reg270 <= $unsigned($unsigned((!((8'ha9) ~^ reg142))));
                    end
                  if ($unsigned(({reg268} ?
                      (forvar48 ?
                          (reg61 ^~ forvar40) : reg78) : (reg49[(2'h2):(2'h2)] ?
                          $signed(reg211) : (forvar21 ? reg69 : forvar174)))))
                    begin
                      reg271 <= $signed(($unsigned($unsigned((8'ha0))) ?
                          ({forvar254} ^ forvar194) : ({(8'ha8)} >>> ((8'hb6) << reg12))));
                      reg272 <= ({forvar50} ?
                          (forvar129[(1'h0):(1'h0)] ^~ $unsigned(reg171[(2'h2):(2'h2)])) : {(reg202[(4'he):(2'h2)] ?
                                  $unsigned(reg55) : reg237[(2'h3):(1'h0)])});
                      reg273 <= $unsigned((|$unsigned((&reg207))));
                      reg274 <= (|(~&reg182[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg271 <= ((forvar147 >>> $signed($signed((8'hb3)))) >> (reg237[(2'h3):(1'h0)] ?
                          ((&reg43) >= $signed(forvar206)) : $unsigned(reg9[(4'hd):(3'h6)])));
                      reg272 <= ({((8'ha0) ?
                              {reg82} : (8'ha2))} != ($signed((~&reg235)) ?
                          reg11 : {(reg91 ? forvar198 : reg211)}));
                      reg273 <= reg272;
                      reg274 <= (($unsigned($signed(reg172)) - ($unsigned(forvar255) ?
                          $signed(reg228) : $signed(forvar178))) + (((~|(8'ha8)) == $unsigned(reg206)) > $unsigned((reg151 ?
                          reg59 : reg231))));
                    end
                  for (forvar275 = (1'h0); (forvar275 < (2'h2)); forvar275 = (forvar275 + (1'h1)))
                    begin
                      reg276 <= (!(((reg185 >> reg149) << $signed(reg22)) ?
                          $signed({forvar268}) : $unsigned($signed(reg227))));
                      reg277 <= (^(($signed(reg226) ?
                          (forvar255 ?
                              forvar39 : reg229) : $signed(reg227)) & $signed((+reg123))));
                      reg278 <= reg36;
                      reg279 <= $unsigned($signed((+forvar254)));
                    end
                  for (forvar280 = (1'h0); (forvar280 < (2'h2)); forvar280 = (forvar280 + (1'h1)))
                    begin
                      reg281 <= $signed(reg10[(3'h4):(1'h0)]);
                    end
                end
              else
                begin
                  reg267 <= (reg97[(4'hf):(3'h7)] - (^($signed(reg138) * (reg280 ?
                      reg36 : reg141))));
                end
              reg282 <= $signed($signed($unsigned(((8'ha5) << reg184))));
            end
        end
      reg283 <= (8'hb9);
      if (reg100)
        begin
          reg284 <= forvar52[(1'h0):(1'h0)];
        end
      else
        begin
          for (forvar284 = (1'h0); (forvar284 < (2'h3)); forvar284 = (forvar284 + (1'h1)))
            begin
              if ($unsigned((8'hb8)))
                begin
                  for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
                    begin
                      reg286 <= ($signed((|(reg65 > reg253))) ?
                          ($unsigned($unsigned(reg43)) ?
                              $signed(reg95[(3'h7):(3'h7)]) : ((~|reg280) < {reg150})) : reg211[(2'h3):(1'h0)]);
                      reg287 <= $unsigned($signed(forvar183[(4'h9):(1'h1)]));
                      reg288 <= {{(~^(!reg30))}};
                      reg289 <= $signed({{(!reg134)}});
                    end
                  for (forvar290 = (1'h0); (forvar290 < (1'h1)); forvar290 = (forvar290 + (1'h1)))
                    begin
                      reg291 <= (reg218 <= reg211);
                      reg292 <= reg73;
                      reg293 <= $unsigned(($unsigned($unsigned(reg276)) != $signed(reg228[(4'h8):(3'h7)])));
                    end
                  for (forvar294 = (1'h0); (forvar294 < (2'h2)); forvar294 = (forvar294 + (1'h1)))
                    begin
                      reg295 <= $signed(reg38);
                    end
                  for (forvar296 = (1'h0); (forvar296 < (1'h1)); forvar296 = (forvar296 + (1'h1)))
                    begin
                      reg297 <= reg93;
                      reg298 <= ($signed(((reg132 ? (8'hb9) : reg75) ?
                          $unsigned(forvar179) : $signed(wire241))) <= reg107);
                    end
                end
              else
                begin
                  for (forvar285 = (1'h0); (forvar285 < (1'h1)); forvar285 = (forvar285 + (1'h1)))
                    begin
                      reg286 <= ($signed($unsigned($unsigned(reg213))) != ((wire3[(1'h1):(1'h1)] + (reg291 ?
                          reg13 : forvar186)) < reg13));
                      reg287 <= ($unsigned(($unsigned((8'had)) ?
                              {reg25} : (reg264 != forvar285))) ?
                          (8'haf) : (^(((8'hb3) == reg272) != (reg263 <<< forvar185))));
                      reg288 <= (|$signed((reg193[(1'h1):(1'h1)] ?
                          (forvar233 ^ (8'hb6)) : ((8'hb5) ?
                              reg143 : (8'h9c)))));
                    end
                end
            end
          if ((^~{forvar8}))
            begin
              if ($unsigned({$unsigned(forvar250)}))
                begin
                  for (forvar299 = (1'h0); (forvar299 < (2'h3)); forvar299 = (forvar299 + (1'h1)))
                    begin
                      reg300 <= (8'hb4);
                    end
                  for (forvar301 = (1'h0); (forvar301 < (1'h0)); forvar301 = (forvar301 + (1'h1)))
                    begin
                      reg302 <= ($unsigned(forvar250[(2'h2):(1'h0)]) ~^ (($signed(reg170) ?
                          $unsigned((8'hb3)) : $signed(forvar86)) == $signed((reg234 >= forvar211))));
                      reg303 <= reg63[(4'hc):(2'h3)];
                      reg304 <= $signed((((~^forvar110) >> reg121) ?
                          {$unsigned(reg295)} : ((reg226 ? forvar245 : reg24) ?
                              (forvar133 + forvar179) : $signed(reg191))));
                      reg305 <= (reg251 ?
                          reg80[(4'h8):(3'h4)] : $signed(forvar262[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar299 = (1'h0); (forvar299 < (2'h2)); forvar299 = (forvar299 + (1'h1)))
                    begin
                      reg300 <= (8'ha1);
                      reg301 <= forvar43;
                      reg302 <= (^~reg29);
                      reg303 <= forvar36[(1'h0):(1'h0)];
                    end
                end
              if ((forvar254 ?
                  $unsigned(({forvar263} << reg280[(1'h1):(1'h0)])) : (!((reg121 ?
                      reg105 : forvar94) ^ reg231))))
                begin
                  for (forvar306 = (1'h0); (forvar306 < (1'h0)); forvar306 = (forvar306 + (1'h1)))
                    begin
                      reg307 <= $unsigned($signed(({reg43} ?
                          $unsigned(reg185) : (+reg281))));
                      reg308 <= ((+forvar113[(2'h3):(1'h0)]) > ((reg162 || {forvar59}) ?
                          reg293 : reg213[(1'h1):(1'h0)]));
                      reg309 <= (($signed((^~reg7)) ?
                              {{forvar214}} : $unsigned((^~(8'ha2)))) ?
                          {$signed((-reg186))} : reg280);
                    end
                  if (reg40[(1'h0):(1'h0)])
                    begin
                      reg310 <= (($unsigned({forvar45}) ~^ reg123[(2'h2):(2'h2)]) > (&$unsigned((&reg164))));
                      reg311 <= reg104[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg310 <= reg281;
                      reg311 <= ((-reg28[(3'h7):(3'h7)]) ^~ (8'hb0));
                      reg312 <= ({((~|reg226) > ((8'hb4) <= forvar45))} && (8'ha8));
                    end
                  if (reg192)
                    begin
                      reg313 <= (reg214[(4'ha):(3'h7)] ?
                          ((forvar74 && $unsigned((8'h9f))) < reg46[(4'hb):(2'h3)]) : ((((8'ha7) ?
                                      reg275 : reg29) ?
                                  $signed(forvar125) : reg170[(3'h5):(2'h2)]) ?
                              wire241[(3'h5):(1'h1)] : reg161));
                      reg314 <= (~^forvar39[(3'h4):(2'h3)]);
                      reg315 <= reg218[(2'h3):(1'h1)];
                      reg316 <= $unsigned(reg101[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg313 <= $signed(($signed((^(8'hb0))) ?
                          (^(8'hb9)) : $unsigned((!reg66))));
                      reg314 <= ((^~((reg123 ~^ reg28) && {reg53})) | $signed(((~&forvar178) + (^~reg201))));
                    end
                  for (forvar317 = (1'h0); (forvar317 < (1'h0)); forvar317 = (forvar317 + (1'h1)))
                    begin
                      reg318 <= ({($signed((8'had)) > (8'haf))} ?
                          $signed((reg313 == reg272[(1'h1):(1'h0)])) : $unsigned((~|$signed((8'ha8)))));
                    end
                end
              else
                begin
                  if (reg14)
                    begin
                      reg306 <= $unsigned(reg16);
                      reg307 <= $signed(reg170);
                      reg308 <= ((!((reg82 ^~ reg289) ?
                          ((8'ha7) ? reg35 : reg107) : (reg163 ?
                              reg146 : (8'h9e)))) ~^ $unsigned($signed((!reg78))));
                      reg309 <= ((&$signed((reg161 - reg77))) <= (~$signed({reg194})));
                    end
                  else
                    begin
                      reg306 <= reg167;
                      reg307 <= $unsigned($signed((reg167[(2'h3):(1'h1)] ?
                          ((8'ha6) ? reg237 : (8'hb5)) : $signed((8'hb7)))));
                    end
                  reg310 <= forvar129[(1'h0):(1'h0)];
                end
              reg319 <= $unsigned(({$unsigned(reg166)} ?
                  reg183 : $unsigned($unsigned(reg250))));
            end
          else
            begin
              for (forvar299 = (1'h0); (forvar299 < (2'h2)); forvar299 = (forvar299 + (1'h1)))
                begin
                  if (reg79)
                    begin
                      reg300 <= ((~^$unsigned($signed(reg148))) ?
                          ((+reg43) ?
                              ((~|reg138) ?
                                  reg98 : reg306) : {reg85}) : (~(((8'ha4) & reg196) ?
                              reg171 : (forvar56 | reg40))));
                      reg301 <= (($signed((~&reg257)) && $signed($unsigned(reg66))) - reg36[(2'h3):(2'h2)]);
                      reg302 <= forvar69;
                      reg303 <= $unsigned((reg23 != ($signed(reg14) <<< (reg71 ?
                          forvar301 : forvar6))));
                    end
                  else
                    begin
                      reg300 <= $unsigned($unsigned((~&(reg245 * reg215))));
                    end
                end
            end
        end
    end
  assign wire320 = (reg152 ?
                       $signed(((reg26 + (8'hb9)) == reg279)) : $signed($signed((8'haa))));
  assign wire321 = $signed(($unsigned($signed((8'hb9))) ?
                       ((~&forvar61) ^~ (reg272 ?
                           reg301 : reg286)) : $unsigned(forvar201[(3'h7):(1'h0)])));
  always
    @(posedge clk) begin
      for (forvar322 = (1'h0); (forvar322 < (1'h1)); forvar322 = (forvar322 + (1'h1)))
        begin
          for (forvar323 = (1'h0); (forvar323 < (1'h0)); forvar323 = (forvar323 + (1'h1)))
            begin
              if (($unsigned($signed((|forvar11))) ?
                  (~^forvar110) : $unsigned(((+reg230) ?
                      {forvar245} : (reg187 ? reg82 : (8'hac))))))
                begin
                  if ((!(reg203[(3'h5):(3'h4)] ?
                      ((+reg64) || (reg278 ?
                          forvar11 : reg180)) : reg15[(1'h1):(1'h0)])))
                    begin
                      reg324 <= reg41[(3'h5):(1'h1)];
                      reg325 <= (!$unsigned($unsigned($signed(reg267))));
                      reg326 <= reg96;
                    end
                  else
                    begin
                      reg324 <= (!(8'ha6));
                      reg325 <= ((reg79 ?
                              $signed($unsigned(reg64)) : $unsigned(((8'ha9) & (8'hac)))) ?
                          ($signed(((8'h9f) && reg266)) ?
                              $unsigned((forvar301 ?
                                  forvar255 : forvar61)) : ($signed((8'ha6)) ?
                                  $unsigned(forvar39) : ((8'had) <= reg206))) : ((((8'hb3) ?
                                      reg123 : forvar248) ?
                                  $signed(forvar294) : $signed(reg25)) ?
                              $signed((~|reg272)) : reg148));
                    end
                  for (forvar327 = (1'h0); (forvar327 < (2'h3)); forvar327 = (forvar327 + (1'h1)))
                    begin
                      reg328 <= $signed(reg256[(4'hb):(1'h0)]);
                      reg329 <= $unsigned(((~reg10[(1'h0):(1'h0)]) | $unsigned({reg45})));
                    end
                  for (forvar330 = (1'h0); (forvar330 < (1'h0)); forvar330 = (forvar330 + (1'h1)))
                    begin
                      reg331 <= ($unsigned(($signed((8'ha3)) ?
                          ((8'h9c) >= reg311) : $unsigned(reg196))) << (+$signed((forvar157 ?
                          reg14 : forvar11))));
                      reg332 <= ((~|reg157) ~^ forvar75);
                      reg333 <= reg249[(2'h3):(1'h1)];
                      reg334 <= (~|($unsigned((reg150 && (8'h9c))) == $unsigned((!forvar255))));
                    end
                end
              else
                begin
                  if (($unsigned($unsigned(reg94[(1'h0):(1'h0)])) >>> reg200))
                    begin
                      reg324 <= ($signed($unsigned(forvar6)) ?
                          $signed((((8'h9e) ~^ reg237) ~^ reg161[(2'h2):(2'h2)])) : reg49);
                      reg325 <= $unsigned($unsigned($unsigned($signed((8'hb3)))));
                      reg326 <= forvar119;
                    end
                  else
                    begin
                      reg324 <= $signed({((!reg58) ? {reg62} : reg238)});
                      reg325 <= reg121[(1'h1):(1'h1)];
                    end
                  for (forvar327 = (1'h0); (forvar327 < (2'h3)); forvar327 = (forvar327 + (1'h1)))
                    begin
                      reg328 <= (-{forvar255});
                      reg329 <= $unsigned($unsigned((reg115 ?
                          reg104 : ((8'h9c) - reg220))));
                    end
                  for (forvar330 = (1'h0); (forvar330 < (1'h0)); forvar330 = (forvar330 + (1'h1)))
                    begin
                      reg331 <= (($unsigned((reg167 ?
                          reg302 : reg47)) - (reg169[(3'h4):(2'h3)] ?
                          (~&reg272) : $unsigned(reg167))) - (reg50[(3'h4):(2'h3)] != reg176[(2'h2):(1'h1)]));
                      reg332 <= reg107;
                      reg333 <= ((!reg200[(1'h0):(1'h0)]) <<< (-(8'hae)));
                      reg334 <= (~^(((reg236 < reg88) ?
                              (^reg109) : (forvar125 ? reg12 : (8'ha0))) ?
                          forvar174[(3'h4):(1'h0)] : {$unsigned(forvar102)}));
                    end
                  for (forvar335 = (1'h0); (forvar335 < (1'h1)); forvar335 = (forvar335 + (1'h1)))
                    begin
                      reg336 <= (((reg208 <= forvar36[(2'h2):(1'h0)]) ?
                              $signed(reg64) : $unsigned($signed(forvar21))) ?
                          reg33 : $signed((8'ha5)));
                      reg337 <= reg231;
                      reg338 <= ($signed(((!forvar243) ?
                              forvar11[(2'h2):(1'h0)] : $signed((8'hb2)))) ?
                          (~^(wire241 ?
                              (forvar50 ~^ forvar194) : $signed((8'hb5)))) : (forvar190[(4'ha):(3'h6)] ~^ $unsigned((~forvar154))));
                      reg339 <= (&reg74[(3'h4):(1'h0)]);
                    end
                end
              if ((-(reg82 > ($unsigned(reg37) >>> forvar190[(4'h8):(2'h3)]))))
                begin
                  reg340 <= $signed(($unsigned((~|reg286)) ?
                      $unsigned($unsigned(reg205)) : forvar218));
                  for (forvar341 = (1'h0); (forvar341 < (1'h0)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= reg304;
                      reg343 <= (($unsigned((reg258 ?
                              forvar267 : (8'haa))) ^~ forvar269) ?
                          (&$unsigned(forvar206[(1'h1):(1'h1)])) : $unsigned($signed((~^reg223))));
                      reg344 <= (~^((-(~|reg103)) ?
                          {(forvar220 ?
                                  reg266 : reg288)} : ($signed(reg23) >= (forvar64 ?
                              (8'hb8) : (8'ha3)))));
                    end
                  if ({(+(wire3[(1'h1):(1'h0)] - {reg229}))})
                    begin
                      reg345 <= (~&(!(~&reg23)));
                      reg346 <= {forvar214[(3'h4):(3'h4)]};
                      reg347 <= (reg75 ^~ (((reg179 > reg244) || $unsigned(reg301)) >>> (reg244[(1'h1):(1'h0)] ?
                          (reg45 ? reg37 : reg304) : {reg198})));
                      reg348 <= ({$signed($signed(forvar232))} ?
                          reg46 : reg144);
                    end
                  else
                    begin
                      reg345 <= $unsigned(reg40[(3'h4):(2'h3)]);
                      reg346 <= reg122[(1'h0):(1'h0)];
                      reg347 <= ((reg312 || $unsigned((forvar190 ?
                              reg115 : reg103))) ?
                          {($signed((8'hb8)) && (reg279 ?
                                  reg261 : reg213))} : (|reg107[(4'h9):(4'h9)]));
                      reg348 <= ($unsigned(($signed(forvar155) ?
                          (reg107 ?
                              reg200 : forvar36) : reg109)) <<< (!$unsigned({reg74})));
                    end
                  if ((&(($unsigned(forvar322) ?
                      (~forvar285) : $unsigned(forvar50)) != $signed($unsigned(reg221)))))
                    begin
                      reg349 <= {$signed((8'ha9))};
                      reg350 <= $signed((~^forvar232));
                    end
                  else
                    begin
                      reg349 <= {$signed(reg214[(2'h3):(1'h1)])};
                      reg350 <= $signed($signed($unsigned($signed(reg127))));
                      reg351 <= (reg194[(4'hb):(2'h2)] - (((forvar131 <<< forvar254) ?
                          (reg88 ?
                              reg329 : reg158) : (reg262 << reg38)) <= $unsigned((&reg44))));
                      reg352 <= reg76[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  reg340 <= reg249[(3'h4):(2'h3)];
                  reg341 <= ($signed(reg87) ~^ ((|reg142) ?
                      ((|forvar56) >>> (forvar214 << forvar280)) : $unsigned((&forvar317))));
                  if (reg10)
                    begin
                      reg342 <= $unsigned((~|$unsigned((8'ha5))));
                      reg343 <= reg137;
                      reg344 <= ($signed(forvar114[(3'h7):(1'h0)]) * {reg152});
                    end
                  else
                    begin
                      reg342 <= $unsigned(((forvar6[(4'hc):(4'hc)] ?
                              reg275 : $unsigned((8'hb2))) ?
                          {(~&reg151)} : {$signed((8'hb1))}));
                      reg343 <= $unsigned(({reg214[(4'h9):(3'h5)]} ?
                          $unsigned(reg127) : forvar323));
                      reg344 <= (-{$signed((~|reg55))});
                      reg345 <= ($unsigned($signed((reg185 ?
                          reg23 : forvar254))) * reg259[(3'h6):(3'h6)]);
                    end
                end
              for (forvar353 = (1'h0); (forvar353 < (2'h2)); forvar353 = (forvar353 + (1'h1)))
                begin
                  if (reg276)
                    begin
                      reg354 <= reg222[(3'h4):(1'h0)];
                      reg355 <= ($unsigned(reg169) ?
                          $signed($signed(reg266[(2'h2):(1'h0)])) : forvar11);
                      reg356 <= ($unsigned($unsigned($signed(reg202))) ?
                          $unsigned(forvar120) : $unsigned(forvar214[(3'h4):(1'h1)]));
                      reg357 <= $unsigned((forvar157[(1'h1):(1'h0)] ?
                          ((forvar330 ? (8'hb7) : (8'hb0)) << (forvar6 ?
                              reg199 : forvar206)) : reg354));
                    end
                  else
                    begin
                      reg354 <= ($unsigned($signed(reg106[(4'h8):(4'h8)])) ?
                          forvar74 : {$unsigned($unsigned(reg157))});
                      reg355 <= ($unsigned((~&$unsigned(reg34))) ?
                          $signed(reg252) : reg105[(1'h0):(1'h0)]);
                      reg356 <= ((forvar160 ?
                              $unsigned(reg305) : ($unsigned(reg88) ?
                                  (~|reg338) : (|(8'ha5)))) ?
                          (reg73 > (~&forvar317)) : reg298);
                      reg357 <= $signed(forvar55);
                    end
                  for (forvar358 = (1'h0); (forvar358 < (2'h3)); forvar358 = (forvar358 + (1'h1)))
                    begin
                      reg359 <= $unsigned((+({reg111} ?
                          $signed((8'hb8)) : ((8'ha3) ? (8'hb9) : reg280))));
                      reg360 <= forvar232[(1'h0):(1'h0)];
                    end
                  if ($signed($unsigned(reg357)))
                    begin
                      reg361 <= forvar322;
                      reg362 <= (&forvar233);
                      reg363 <= $unsigned((reg98 ?
                          ($signed(reg145) == $unsigned(forvar21)) : ({reg238} ?
                              $unsigned((8'h9c)) : (reg284 >> (8'hb3)))));
                    end
                  else
                    begin
                      reg361 <= (&$signed($unsigned((reg334 ?
                          reg258 : reg359))));
                      reg362 <= ($signed(wire321[(4'h9):(4'h8)]) ?
                          (!reg211) : ($unsigned({reg117}) ?
                              $unsigned({reg203}) : ((reg221 ?
                                  (8'ha7) : reg170) >> reg218[(1'h1):(1'h0)])));
                    end
                  reg364 <= $unsigned(reg264);
                end
              if ($signed(reg52[(3'h5):(3'h5)]))
                begin
                  for (forvar365 = (1'h0); (forvar365 < (1'h1)); forvar365 = (forvar365 + (1'h1)))
                    begin
                      reg366 <= reg157[(3'h5):(3'h4)];
                      reg367 <= reg82[(1'h0):(1'h0)];
                    end
                  reg368 <= (8'hb8);
                  if ($unsigned(((&{reg319}) ?
                      $unsigned((8'hae)) : reg54[(3'h5):(2'h3)])))
                    begin
                      reg369 <= $signed($unsigned($signed($unsigned(reg227))));
                      reg370 <= (~|{forvar280[(2'h2):(1'h1)]});
                      reg371 <= reg225;
                    end
                  else
                    begin
                      reg369 <= $unsigned(($unsigned((reg308 | reg81)) ?
                          reg171 : reg200[(2'h2):(2'h2)]));
                      reg370 <= (^~(($signed(reg223) << (reg340 ?
                          (8'hb9) : reg16)) ^ reg11));
                    end
                  if ($unsigned(((^(^~reg199)) - reg126[(4'ha):(3'h7)])))
                    begin
                      reg372 <= (8'ha4);
                    end
                  else
                    begin
                      reg372 <= (|reg135);
                      reg373 <= $unsigned(reg47[(1'h0):(1'h0)]);
                      reg374 <= $signed((reg136 ?
                          $unsigned((~|(8'hba))) : forvar280));
                      reg375 <= (($unsigned(reg304[(3'h7):(1'h0)]) <<< reg202) ^ wire241);
                    end
                end
              else
                begin
                  if (({(8'hb6)} ?
                      $signed(($unsigned((8'ha7)) ?
                          (forvar201 <= (8'ha8)) : (^~reg166))) : reg304))
                    begin
                      reg365 <= ($signed((~^(reg248 <= reg159))) ?
                          forvar102 : (($unsigned(reg246) & (reg370 ?
                                  reg139 : reg112)) ?
                              (8'hb2) : (forvar75 ?
                                  forvar52 : $signed(reg186))));
                      reg366 <= wire3[(2'h2):(1'h0)];
                      reg367 <= reg94[(4'ha):(1'h1)];
                      reg368 <= {reg263[(1'h1):(1'h1)]};
                    end
                  else
                    begin
                      reg365 <= $signed($unsigned((!(forvar183 ?
                          (8'h9f) : reg275))));
                      reg366 <= forvar323[(4'hb):(3'h7)];
                      reg367 <= reg19;
                      reg368 <= $unsigned((reg161 <= reg363[(1'h1):(1'h1)]));
                    end
                  if (wire241)
                    begin
                      reg369 <= (forvar285 <<< (^(reg16 ?
                          (&reg304) : (!reg283))));
                    end
                  else
                    begin
                      reg369 <= reg372;
                      reg370 <= $unsigned({($unsigned(reg187) * (!reg117))});
                    end
                end
            end
          for (forvar376 = (1'h0); (forvar376 < (2'h2)); forvar376 = (forvar376 + (1'h1)))
            begin
              if ($signed({($signed(reg36) <<< reg10[(3'h5):(3'h4)])}))
                begin
                  reg377 <= (^~(($signed(forvar61) != (reg31 | reg205)) == (forvar206 & {reg173})));
                end
              else
                begin
                  if ((^(reg10[(3'h4):(1'h1)] & ((forvar262 ?
                      reg88 : reg209) ^~ (reg91 <= reg91)))))
                    begin
                      reg377 <= forvar183[(3'h7):(2'h2)];
                    end
                  else
                    begin
                      reg377 <= (~|$signed((((8'hb4) > reg348) == ((8'hae) ?
                          reg259 : reg194))));
                      reg378 <= $signed(reg35);
                    end
                  reg379 <= $signed($unsigned(reg341[(2'h3):(1'h1)]));
                  for (forvar380 = (1'h0); (forvar380 < (1'h1)); forvar380 = (forvar380 + (1'h1)))
                    begin
                      reg381 <= (({reg52} ?
                          (~(wire2 ? reg108 : reg202)) : ((8'ha0) ?
                              (8'h9e) : (|reg169))) ^~ forvar260[(3'h6):(1'h0)]);
                      reg382 <= reg306;
                    end
                end
              if (reg269)
                begin
                  reg383 <= (~((~(forvar254 ?
                      reg9 : reg25)) <= reg329[(3'h7):(3'h6)]));
                  reg384 <= ((&forvar36[(1'h0):(1'h0)]) != reg206);
                  if ((&reg378[(2'h3):(1'h1)]))
                    begin
                      reg385 <= forvar184;
                    end
                  else
                    begin
                      reg385 <= $signed({forvar37});
                      reg386 <= {$signed($unsigned(reg328))};
                      reg387 <= $unsigned(reg218[(2'h3):(2'h2)]);
                      reg388 <= ($signed(forvar67[(1'h0):(1'h0)]) ?
                          {(((8'h9c) ? forvar133 : reg383) ?
                                  $unsigned((8'hba)) : reg291[(3'h4):(2'h3)])} : ({$unsigned(reg66)} ?
                              $unsigned(reg104) : $unsigned((reg386 ?
                                  reg311 : reg254))));
                    end
                end
              else
                begin
                  if (((&reg288[(4'h8):(2'h3)]) ?
                      reg374[(1'h1):(1'h1)] : (~&$unsigned(reg78[(3'h5):(1'h0)]))))
                    begin
                      reg383 <= forvar157;
                      reg384 <= (|(&reg368[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg383 <= (~&reg34);
                      reg384 <= $unsigned((((forvar197 ? reg193 : reg145) ?
                              forvar185 : (&forvar94)) ?
                          (|reg152[(2'h3):(1'h1)]) : ((~reg193) ?
                              (reg313 ? reg59 : reg192) : ((8'h9d) ?
                                  reg230 : reg88))));
                      reg385 <= ((~^(reg238[(2'h3):(2'h2)] ?
                              (forvar232 | reg298) : reg316)) ?
                          reg267 : (|$signed(((8'hab) >> (8'ha8)))));
                    end
                  reg386 <= $signed(reg164[(3'h5):(2'h3)]);
                end
            end
          reg389 <= (reg90 << $unsigned($unsigned($signed(reg185))));
          reg390 <= reg370;
        end
      if ({$signed((reg256[(3'h4):(2'h2)] ?
              (reg202 ? wire4 : reg246) : (reg203 ? (8'hb7) : (8'ha6))))})
        begin
          reg391 <= reg221[(1'h0):(1'h0)];
          for (forvar392 = (1'h0); (forvar392 < (2'h3)); forvar392 = (forvar392 + (1'h1)))
            begin
              for (forvar393 = (1'h0); (forvar393 < (2'h2)); forvar393 = (forvar393 + (1'h1)))
                begin
                  if (reg250)
                    begin
                      reg394 <= reg313[(4'h8):(2'h3)];
                      reg395 <= reg336[(2'h2):(1'h1)];
                      reg396 <= $unsigned(reg17);
                    end
                  else
                    begin
                      reg394 <= reg196[(1'h0):(1'h0)];
                    end
                end
              if (forvar59)
                begin
                  for (forvar397 = (1'h0); (forvar397 < (1'h1)); forvar397 = (forvar397 + (1'h1)))
                    begin
                      reg398 <= $unsigned($signed({$unsigned(reg292)}));
                      reg399 <= (8'ha8);
                      reg400 <= $unsigned((($signed(reg139) ?
                              (reg72 < reg284) : $signed((8'hac))) ?
                          (^~reg69) : ((~reg82) ?
                              $signed(reg227) : $signed(reg267))));
                    end
                  for (forvar401 = (1'h0); (forvar401 < (2'h3)); forvar401 = (forvar401 + (1'h1)))
                    begin
                      reg402 <= $unsigned($signed(forvar21[(1'h0):(1'h0)]));
                      reg403 <= reg318[(1'h0):(1'h0)];
                      reg404 <= reg307;
                    end
                  if (reg387[(3'h6):(1'h0)])
                    begin
                      reg405 <= {(~|$signed(reg166[(4'h8):(3'h7)]))};
                    end
                  else
                    begin
                      reg405 <= reg25;
                      reg406 <= $unsigned($signed((~&reg22[(1'h1):(1'h0)])));
                      reg407 <= (reg280[(3'h6):(1'h0)] <= (^$signed((^(8'ha2)))));
                      reg408 <= reg79;
                    end
                  if ({reg202[(2'h2):(1'h1)]})
                    begin
                      reg409 <= $signed({reg404});
                      reg410 <= (((reg58[(1'h1):(1'h0)] ?
                              (^~forvar323) : (reg240 ? forvar6 : reg132)) ?
                          ((reg274 ? (8'hae) : (8'haf)) ?
                              (&(8'haf)) : reg186[(3'h7):(3'h5)]) : ((reg239 ?
                                  forvar376 : reg342) ?
                              (8'hb9) : $unsigned(reg408))) >> ($unsigned($signed(forvar76)) ?
                          $unsigned(reg177[(2'h2):(2'h2)]) : (wire2 ?
                              (reg258 ?
                                  reg293 : reg104) : reg356[(1'h1):(1'h0)])));
                      reg411 <= reg116;
                      reg412 <= forvar155;
                    end
                  else
                    begin
                      reg409 <= reg248[(2'h2):(2'h2)];
                      reg410 <= $signed($signed($unsigned(reg254)));
                    end
                end
              else
                begin
                  for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
                    begin
                      reg398 <= {reg170[(3'h5):(1'h1)]};
                      reg399 <= (~^reg385[(4'hf):(3'h4)]);
                      reg400 <= forvar267;
                      reg401 <= {$unsigned(reg16[(2'h3):(2'h3)])};
                    end
                  for (forvar402 = (1'h0); (forvar402 < (1'h0)); forvar402 = (forvar402 + (1'h1)))
                    begin
                      reg403 <= ($unsigned((+(reg267 ? reg192 : reg411))) ?
                          (~|reg379[(3'h6):(2'h2)]) : forvar275);
                    end
                end
              for (forvar413 = (1'h0); (forvar413 < (1'h0)); forvar413 = (forvar413 + (1'h1)))
                begin
                  for (forvar414 = (1'h0); (forvar414 < (2'h2)); forvar414 = (forvar414 + (1'h1)))
                    begin
                      reg415 <= $unsigned((reg161 >> $unsigned($unsigned((8'haa)))));
                      reg416 <= ((&$unsigned(forvar79[(2'h2):(1'h1)])) ?
                          (+(8'hb8)) : (reg45 ~^ ((&forvar244) ?
                              {reg213} : (forvar414 && reg246))));
                    end
                end
            end
          if ({reg18[(3'h5):(2'h2)]})
            begin
              for (forvar417 = (1'h0); (forvar417 < (2'h3)); forvar417 = (forvar417 + (1'h1)))
                begin
                  for (forvar418 = (1'h0); (forvar418 < (1'h0)); forvar418 = (forvar418 + (1'h1)))
                    begin
                      reg419 <= $signed($unsigned(reg308));
                      reg420 <= $unsigned($unsigned(reg23[(1'h0):(1'h0)]));
                    end
                  reg421 <= $unsigned($unsigned((reg249 ?
                      reg79 : $signed(reg401))));
                end
              if (((^$signed({forvar43})) ^~ $unsigned(((reg169 == reg30) * $unsigned(reg17)))))
                begin
                  reg422 <= ($unsigned(((reg412 && reg302) || $signed(forvar7))) <= $unsigned((reg304[(2'h3):(2'h3)] ?
                      reg109 : (reg107 ? (8'hb3) : reg360))));
                end
              else
                begin
                  reg422 <= {$unsigned(forvar248)};
                  for (forvar423 = (1'h0); (forvar423 < (2'h3)); forvar423 = (forvar423 + (1'h1)))
                    begin
                      reg424 <= forvar110;
                    end
                  for (forvar425 = (1'h0); (forvar425 < (1'h0)); forvar425 = (forvar425 + (1'h1)))
                    begin
                      reg426 <= $signed($unsigned(forvar299));
                      reg427 <= $unsigned(reg371);
                      reg428 <= (({reg411} ?
                              $unsigned($unsigned(reg345)) : (^reg333)) ?
                          $unsigned(reg329[(4'h8):(4'h8)]) : $signed($unsigned((-reg382))));
                      reg429 <= ((reg111[(1'h0):(1'h0)] * reg314) >> $signed($unsigned((reg310 && (8'hb9)))));
                    end
                  if ($signed($signed((reg47[(2'h2):(2'h2)] * (~|reg313)))))
                    begin
                      reg430 <= reg277[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg430 <= ($signed(((|reg283) && reg211[(1'h0):(1'h0)])) ^ (8'hba));
                      reg431 <= $unsigned(reg117[(3'h5):(3'h4)]);
                      reg432 <= reg409[(3'h7):(2'h2)];
                      reg433 <= $unsigned(reg199[(3'h4):(1'h1)]);
                    end
                end
              if (reg94)
                begin
                  reg434 <= {(($signed(reg223) & (^~(8'hab))) ?
                          (reg314[(2'h2):(1'h1)] + $unsigned(reg9)) : ($unsigned(reg141) ?
                              (reg76 ? (8'hac) : reg90) : {reg399}))};
                end
              else
                begin
                  if ((~&($signed($unsigned(forvar21)) ?
                      $unsigned($signed(reg210)) : forvar414[(4'h8):(1'h1)])))
                    begin
                      reg434 <= $unsigned($signed($signed(reg7)));
                      reg435 <= {reg292[(4'hc):(1'h1)]};
                    end
                  else
                    begin
                      reg434 <= reg276[(4'he):(1'h1)];
                    end
                  if (reg49)
                    begin
                      reg436 <= reg138;
                      reg437 <= {($unsigned((^reg263)) && $unsigned(forvar92[(1'h0):(1'h0)]))};
                    end
                  else
                    begin
                      reg436 <= (((+$signed(forvar201)) ?
                          $signed((^~(8'ha9))) : ($unsigned(reg43) ?
                              reg69 : {forvar284})) ^~ reg188[(2'h3):(2'h2)]);
                    end
                  reg438 <= reg389;
                end
              for (forvar439 = (1'h0); (forvar439 < (2'h3)); forvar439 = (forvar439 + (1'h1)))
                begin
                  reg440 <= $unsigned((reg237 ?
                      forvar39 : ((&reg100) ?
                          (^forvar244) : (forvar299 ? reg405 : reg37))));
                end
            end
          else
            begin
              reg417 <= {$unsigned({(~|forvar260)})};
              for (forvar418 = (1'h0); (forvar418 < (1'h1)); forvar418 = (forvar418 + (1'h1)))
                begin
                  for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
                    begin
                      reg420 <= (&reg361);
                    end
                end
              for (forvar421 = (1'h0); (forvar421 < (2'h2)); forvar421 = (forvar421 + (1'h1)))
                begin
                  for (forvar422 = (1'h0); (forvar422 < (1'h0)); forvar422 = (forvar422 + (1'h1)))
                    begin
                      reg423 <= reg421[(1'h0):(1'h0)];
                      reg424 <= reg284[(1'h0):(1'h0)];
                    end
                  if ((-((~|((8'ha1) ? (8'hb2) : reg204)) < {reg25})))
                    begin
                      reg425 <= $signed(({(reg107 >= reg223)} ?
                          {(reg65 ? (8'hae) : reg254)} : (~|(~|reg25))));
                      reg426 <= ((reg212 ?
                              $signed(reg245[(2'h3):(2'h3)]) : $unsigned((reg97 ?
                                  reg277 : (8'hb3)))) ?
                          ((~|(reg309 ?
                              forvar102 : (8'ha4))) & {$unsigned(reg117)}) : (forvar275 ?
                              $signed(reg139) : ($unsigned(forvar439) ?
                                  forvar129 : ((8'ha4) + reg108))));
                    end
                  else
                    begin
                      reg425 <= $signed(reg430);
                      reg426 <= $signed($signed(reg387));
                      reg427 <= $signed((reg28[(2'h2):(2'h2)] ^~ $unsigned(reg404)));
                      reg428 <= reg24;
                    end
                end
              for (forvar429 = (1'h0); (forvar429 < (2'h2)); forvar429 = (forvar429 + (1'h1)))
                begin
                  for (forvar430 = (1'h0); (forvar430 < (2'h3)); forvar430 = (forvar430 + (1'h1)))
                    begin
                      reg431 <= (+reg162[(3'h6):(2'h2)]);
                      reg432 <= reg301[(3'h5):(2'h2)];
                      reg433 <= (((~$signed(reg423)) ?
                          forvar186[(1'h1):(1'h1)] : (reg172[(3'h7):(3'h5)] ?
                              $signed(reg40) : reg263[(1'h1):(1'h0)])) ^ $signed((reg411[(3'h4):(1'h1)] != $unsigned((8'h9c)))));
                    end
                  reg434 <= $signed($signed($unsigned((8'hb5))));
                end
            end
        end
      else
        begin
          for (forvar391 = (1'h0); (forvar391 < (2'h2)); forvar391 = (forvar391 + (1'h1)))
            begin
              if ({(~^$signed($signed(reg337)))})
                begin
                  reg392 <= ($signed(forvar323[(3'h6):(2'h2)]) << $signed(reg286));
                  if ({reg19[(1'h0):(1'h0)]})
                    begin
                      reg393 <= $signed($unsigned(((~^reg123) ?
                          (reg284 ? forvar147 : reg95) : {(8'hb4)})));
                      reg394 <= reg146;
                      reg395 <= reg419[(3'h6):(3'h6)];
                    end
                  else
                    begin
                      reg393 <= $unsigned(($signed({reg344}) ?
                          $signed(reg148) : ((forvar418 - reg430) >>> (^~reg313))));
                      reg394 <= (forvar36[(2'h2):(1'h1)] ?
                          $signed($unsigned($unsigned(forvar358))) : (forvar11[(2'h3):(2'h3)] ?
                              $signed({reg324}) : (reg28 && $unsigned(reg58))));
                      reg395 <= reg251[(2'h2):(1'h0)];
                      reg396 <= {((((8'haf) ^ reg196) + forvar275[(3'h4):(2'h3)]) ?
                              forvar20 : reg185)};
                    end
                end
              else
                begin
                  reg392 <= (-$signed((forvar285 | (reg403 ?
                      (8'hb8) : reg247))));
                  for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
                    begin
                      reg394 <= ((8'hab) | (reg262 + reg32[(2'h3):(1'h1)]));
                    end
                  if ({$signed(((+(8'h9c)) ? reg117 : wire242[(1'h1):(1'h0)]))})
                    begin
                      reg395 <= (^~reg204);
                      reg396 <= $unsigned((8'ha1));
                      reg397 <= (({$signed(reg122)} >> ((^~wire242) ?
                              reg398 : (-forvar74))) ?
                          $signed($unsigned((forvar285 ?
                              forvar197 : reg148))) : reg191);
                    end
                  else
                    begin
                      reg395 <= forvar341;
                    end
                  reg398 <= reg171[(3'h5):(1'h0)];
                end
              for (forvar399 = (1'h0); (forvar399 < (1'h0)); forvar399 = (forvar399 + (1'h1)))
                begin
                  if ($unsigned(reg261[(2'h2):(2'h2)]))
                    begin
                      reg400 <= $unsigned(({reg162} ^ (^$signed(reg130))));
                      reg401 <= $unsigned((8'hab));
                      reg402 <= reg318;
                      reg403 <= $unsigned((~&$unsigned((wire0 && reg278))));
                    end
                  else
                    begin
                      reg400 <= $signed((-$signed(reg164)));
                      reg401 <= (($signed({(8'ha2)}) > $signed($signed(reg211))) & reg46);
                      reg402 <= ((8'hb4) ?
                          (reg311 <<< (~^(reg261 ?
                              reg180 : (8'hae)))) : {{(|forvar301)}});
                      reg403 <= reg70;
                    end
                end
              reg404 <= {(reg350[(1'h1):(1'h1)] ?
                      ((~|forvar330) ? forvar79 : reg42) : $unsigned((reg273 ?
                          forvar376 : reg229)))};
              for (forvar405 = (1'h0); (forvar405 < (1'h1)); forvar405 = (forvar405 + (1'h1)))
                begin
                  if ({forvar11})
                    begin
                      reg406 <= $unsigned($unsigned((reg393 ~^ reg356[(3'h7):(3'h6)])));
                      reg407 <= (|forvar56[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg406 <= {{reg144[(2'h3):(1'h0)]}};
                      reg407 <= reg415[(4'h9):(2'h2)];
                      reg408 <= $unsigned(((wire242[(4'h9):(4'h9)] ?
                          forvar110[(2'h3):(2'h3)] : reg105[(1'h0):(1'h0)]) && forvar131));
                      reg409 <= reg57[(3'h5):(3'h4)];
                    end
                end
            end
          for (forvar410 = (1'h0); (forvar410 < (2'h2)); forvar410 = (forvar410 + (1'h1)))
            begin
              reg411 <= reg313[(1'h1):(1'h1)];
              if ({$signed((|$unsigned(forvar301)))})
                begin
                  if ({reg93})
                    begin
                      reg412 <= (~^reg10[(3'h4):(1'h1)]);
                      reg413 <= $unsigned(($unsigned({forvar147}) + $unsigned(forvar160[(4'h9):(3'h6)])));
                    end
                  else
                    begin
                      reg412 <= ({(8'ha5)} * reg42[(3'h4):(3'h4)]);
                    end
                  if ((^{$unsigned(reg164)}))
                    begin
                      reg414 <= ($signed(((forvar306 ? (8'ha1) : reg372) ?
                          reg393[(3'h6):(1'h0)] : $signed(reg266))) ^~ $unsigned(forvar11));
                    end
                  else
                    begin
                      reg414 <= ($unsigned(({reg49} <<< forvar86)) ?
                          ((reg230[(4'h8):(2'h3)] ?
                                  forvar45 : forvar391[(1'h1):(1'h1)]) ?
                              reg407[(4'h9):(1'h0)] : (+$signed(reg301))) : ((|(forvar267 << reg145)) ?
                              reg248[(1'h1):(1'h0)] : $unsigned($signed(wire2))));
                      reg415 <= (reg270 <= reg236);
                      reg416 <= $unsigned((+$unsigned($signed(reg188))));
                      reg417 <= $signed((((reg433 ^~ reg254) * (&reg280)) ?
                          forvar327[(2'h2):(2'h2)] : reg314[(3'h7):(3'h7)]));
                    end
                  if ($unsigned((|$signed($signed(reg273)))))
                    begin
                      reg418 <= (reg316[(1'h1):(1'h1)] && (reg249[(3'h4):(1'h0)] ?
                          (~|$unsigned((8'hb5))) : (~|$unsigned(reg173))));
                      reg419 <= (($signed($signed(reg319)) <<< $unsigned(((8'ha4) ?
                              forvar402 : reg146))) ?
                          (!($signed(forvar190) * reg328[(3'h5):(2'h2)])) : reg68[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg418 <= ((({(8'hb1)} ?
                          reg28 : {reg138}) && (~reg145)) < reg245);
                      reg419 <= ($signed((reg96 == $signed(forvar153))) - $signed(reg410[(4'h8):(3'h6)]));
                      reg420 <= reg284;
                    end
                  for (forvar421 = (1'h0); (forvar421 < (1'h0)); forvar421 = (forvar421 + (1'h1)))
                    begin
                      reg422 <= {reg137};
                      reg423 <= $unsigned((~^($signed(reg234) <= {(8'ha5)})));
                    end
                end
              else
                begin
                  reg412 <= reg370[(3'h5):(1'h1)];
                  for (forvar413 = (1'h0); (forvar413 < (2'h2)); forvar413 = (forvar413 + (1'h1)))
                    begin
                      reg414 <= reg139;
                    end
                  for (forvar415 = (1'h0); (forvar415 < (1'h0)); forvar415 = (forvar415 + (1'h1)))
                    begin
                      reg416 <= (($signed($unsigned(reg101)) ?
                          ((reg34 < reg79) ?
                              (8'had) : (~|forvar168)) : {(forvar397 < reg409)}) < {($unsigned(reg329) ?
                              $signed(reg228) : (reg53 >> forvar296))});
                      reg417 <= $signed(reg220);
                      reg418 <= ({$unsigned((reg413 == reg272))} ^~ (^~reg91));
                    end
                  for (forvar419 = (1'h0); (forvar419 < (1'h0)); forvar419 = (forvar419 + (1'h1)))
                    begin
                      reg420 <= (($signed((~|reg400)) * reg415) ?
                          (((~reg426) > {reg379}) ?
                              $unsigned((reg99 >>> reg7)) : ($signed((8'hb9)) ?
                                  (~|reg203) : $signed(reg217))) : (((reg24 ^~ forvar193) && (+forvar263)) & {(forvar243 >= reg281)}));
                      reg421 <= reg126;
                      reg422 <= (reg35[(3'h4):(1'h0)] << $signed(((8'h9e) ?
                          (reg430 >>> reg336) : {forvar120})));
                    end
                end
            end
          for (forvar424 = (1'h0); (forvar424 < (2'h2)); forvar424 = (forvar424 + (1'h1)))
            begin
              reg425 <= (8'ha3);
              reg426 <= $unsigned((forvar184 ? (~|(8'h9f)) : {reg83}));
              for (forvar427 = (1'h0); (forvar427 < (1'h0)); forvar427 = (forvar427 + (1'h1)))
                begin
                  for (forvar428 = (1'h0); (forvar428 < (1'h1)); forvar428 = (forvar428 + (1'h1)))
                    begin
                      reg429 <= reg247;
                      reg430 <= reg252[(3'h4):(1'h0)];
                      reg431 <= (|{(8'ha3)});
                      reg432 <= (8'ha0);
                    end
                end
            end
        end
      for (forvar441 = (1'h0); (forvar441 < (1'h0)); forvar441 = (forvar441 + (1'h1)))
        begin
          reg442 <= (8'haf);
          if ($signed((!(!$signed(reg244)))))
            begin
              if (($signed(reg206[(1'h1):(1'h0)]) ~^ $signed((|{forvar153}))))
                begin
                  reg443 <= $signed((&((reg204 ?
                      wire242 : forvar185) - $signed(reg149))));
                  for (forvar444 = (1'h0); (forvar444 < (1'h1)); forvar444 = (forvar444 + (1'h1)))
                    begin
                      reg445 <= $signed(forvar186);
                      reg446 <= {forvar401};
                      reg447 <= ((~^$unsigned((~&reg135))) ?
                          (8'haf) : (reg253 ^~ reg45));
                      reg448 <= reg391[(3'h6):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar443 = (1'h0); (forvar443 < (1'h0)); forvar443 = (forvar443 + (1'h1)))
                    begin
                      reg444 <= $unsigned({{$signed(reg209)}});
                      reg445 <= $unsigned($unsigned(reg220[(3'h4):(2'h2)]));
                      reg446 <= (reg360[(3'h4):(3'h4)] ?
                          reg105 : (^$unsigned(forvar190)));
                      reg447 <= $unsigned($signed((-$unsigned((8'had)))));
                    end
                  reg448 <= reg431;
                  if ($signed((|((reg375 ?
                      forvar418 : forvar160) <<< ((8'hb0) * reg281)))))
                    begin
                      reg449 <= ((reg412[(1'h0):(1'h0)] ?
                              (((8'hab) - reg17) != {reg366}) : $signed({(8'ha2)})) ?
                          (-(~^((8'hb4) >>> reg72))) : $signed(wire242));
                      reg450 <= $unsigned({forvar365});
                      reg451 <= (reg187[(4'h9):(3'h4)] <<< $unsigned(forvar299[(4'h8):(1'h0)]));
                    end
                  else
                    begin
                      reg449 <= reg222[(4'h9):(3'h6)];
                      reg450 <= reg422;
                      reg451 <= (reg306[(2'h3):(1'h1)] * ((8'ha6) ?
                          $unsigned(reg264[(3'h5):(3'h4)]) : (|forvar417)));
                    end
                end
            end
          else
            begin
              if ((reg50 ?
                  $unsigned(forvar36) : ((reg373[(2'h3):(2'h2)] & (reg447 ?
                          reg53 : reg275)) ?
                      (8'hb3) : forvar439[(4'h8):(3'h5)])))
                begin
                  for (forvar443 = (1'h0); (forvar443 < (1'h1)); forvar443 = (forvar443 + (1'h1)))
                    begin
                      reg444 <= (~^$signed(reg305));
                      reg445 <= {($unsigned({(8'ha1)}) ~^ reg449)};
                      reg446 <= (~|((8'hba) ?
                          reg184[(3'h6):(3'h4)] : ($unsigned((8'h9e)) <= {forvar133})));
                      reg447 <= $signed(reg264);
                    end
                  if ($unsigned(((forvar52[(3'h4):(1'h1)] ?
                      (reg101 << reg62) : $signed(reg201)) < reg145)))
                    begin
                      reg448 <= ((-reg126) ~^ $unsigned($signed((reg222 ?
                          reg89 : reg136))));
                      reg449 <= $signed({(~|(reg70 ~^ reg279))});
                      reg450 <= (^reg329);
                    end
                  else
                    begin
                      reg448 <= (~&(reg418 << $unsigned((reg146 + reg156))));
                    end
                  reg451 <= (reg389[(1'h1):(1'h1)] ?
                      $unsigned(reg108[(4'h8):(3'h5)]) : reg311[(4'h9):(3'h6)]);
                end
              else
                begin
                  for (forvar443 = (1'h0); (forvar443 < (1'h1)); forvar443 = (forvar443 + (1'h1)))
                    begin
                      reg444 <= $unsigned({(~&{reg283})});
                    end
                end
              reg452 <= {(+(~&(forvar335 ~^ forvar322)))};
              for (forvar453 = (1'h0); (forvar453 < (1'h0)); forvar453 = (forvar453 + (1'h1)))
                begin
                  for (forvar454 = (1'h0); (forvar454 < (1'h1)); forvar454 = (forvar454 + (1'h1)))
                    begin
                      reg455 <= (&reg77);
                      reg456 <= $signed(reg173[(4'ha):(1'h0)]);
                      reg457 <= $signed({$signed(reg413)});
                      reg458 <= (^$unsigned((-(~^reg134))));
                    end
                  if (reg172)
                    begin
                      reg459 <= $unsigned(((~|{(8'h9d)}) ^~ $unsigned(wire2[(1'h0):(1'h0)])));
                      reg460 <= (forvar317 <= reg282[(1'h0):(1'h0)]);
                      reg461 <= (~&$signed($signed($signed((8'hb3)))));
                      reg462 <= ((reg149[(4'h9):(3'h4)] <= $unsigned($signed(reg340))) <<< $unsigned(reg148[(3'h4):(1'h1)]));
                    end
                  else
                    begin
                      reg459 <= (~|$signed($signed((forvar69 ?
                          forvar55 : (8'hb4)))));
                      reg460 <= (~(|((reg14 <= reg186) ?
                          {(8'hb4)} : $unsigned((8'ha9)))));
                    end
                end
              if ($unsigned($unsigned(((^reg213) < $signed(forvar376)))))
                begin
                  for (forvar463 = (1'h0); (forvar463 < (1'h0)); forvar463 = (forvar463 + (1'h1)))
                    begin
                      reg464 <= reg49;
                      reg465 <= (8'hae);
                      reg466 <= ((+$signed(reg444[(3'h7):(1'h1)])) ?
                          (reg103[(3'h4):(1'h0)] ?
                              ($signed(forvar198) ?
                                  ((8'ha1) ? (8'hb9) : reg292) : (forvar198 ?
                                      forvar418 : (8'hba))) : {$unsigned(reg65)}) : (-reg307[(1'h0):(1'h0)]));
                      reg467 <= $signed($unsigned(reg195));
                    end
                end
              else
                begin
                  for (forvar463 = (1'h0); (forvar463 < (1'h1)); forvar463 = (forvar463 + (1'h1)))
                    begin
                      reg464 <= $unsigned(reg96[(3'h5):(3'h4)]);
                      reg465 <= ($signed((^reg18)) ^ reg457);
                    end
                  for (forvar466 = (1'h0); (forvar466 < (2'h2)); forvar466 = (forvar466 + (1'h1)))
                    begin
                      reg467 <= $unsigned({((^~reg267) + (reg252 != forvar37))});
                      reg468 <= (reg364 | reg444[(4'hb):(3'h6)]);
                      reg469 <= (8'haa);
                      reg470 <= reg280;
                    end
                  for (forvar471 = (1'h0); (forvar471 < (2'h2)); forvar471 = (forvar471 + (1'h1)))
                    begin
                      reg472 <= (($signed({reg338}) ~^ $unsigned((8'had))) ?
                          reg405[(3'h4):(3'h4)] : (reg83[(2'h2):(1'h1)] == $signed(forvar102)));
                      reg473 <= (((forvar179 != $unsigned(reg395)) ?
                          forvar299 : (~|$signed(reg367))) <= $unsigned($unsigned(reg256)));
                    end
                  if (reg385[(5'h10):(4'hf)])
                    begin
                      reg474 <= ((($signed(forvar341) >>> (forvar184 ?
                          reg270 : (8'ha0))) >>> reg30[(1'h1):(1'h1)]) ^~ (!((forvar119 > reg150) ?
                          forvar114[(3'h6):(3'h6)] : reg287[(2'h3):(1'h1)])));
                      reg475 <= forvar405;
                    end
                  else
                    begin
                      reg474 <= $signed($unsigned($signed(reg104)));
                    end
                end
            end
          if ({{((forvar188 ? reg458 : reg121) ?
                      (reg178 ? reg399 : forvar365) : $signed(reg63))}})
            begin
              reg476 <= forvar353;
              reg477 <= ((&reg158) ?
                  (forvar290 || $unsigned((forvar322 ?
                      reg179 : reg187))) : ((8'hba) ?
                      ((reg24 && reg462) ?
                          ((8'ha2) > (8'h9d)) : (reg35 == reg148)) : (-$unsigned(forvar294))));
            end
          else
            begin
              if ($signed($unsigned(((~^reg198) ?
                  $unsigned(reg109) : (reg73 | reg10)))))
                begin
                  if (reg98[(3'h6):(2'h2)])
                    begin
                      reg476 <= $signed(forvar113);
                      reg477 <= reg430[(5'h10):(4'h8)];
                    end
                  else
                    begin
                      reg476 <= reg350;
                      reg477 <= (~|(+{(&reg356)}));
                    end
                end
              else
                begin
                  for (forvar476 = (1'h0); (forvar476 < (1'h0)); forvar476 = (forvar476 + (1'h1)))
                    begin
                      reg477 <= {forvar280[(1'h1):(1'h1)]};
                      reg478 <= reg214[(4'ha):(4'h9)];
                    end
                  if ({((reg383 ?
                          $signed(reg245) : (reg57 ?
                              forvar454 : reg97)) > {{reg135}})})
                    begin
                      reg479 <= $signed($unsigned($unsigned((reg475 < reg116))));
                    end
                  else
                    begin
                      reg479 <= (|{(^~(~|reg269))});
                      reg480 <= $unsigned($signed($signed(forvar296)));
                    end
                end
              if (reg189[(1'h1):(1'h1)])
                begin
                  for (forvar481 = (1'h0); (forvar481 < (2'h2)); forvar481 = (forvar481 + (1'h1)))
                    begin
                      reg482 <= $unsigned(((~|$signed(reg218)) == ($signed((8'ha5)) ?
                          reg297[(4'h8):(4'h8)] : {reg370})));
                      reg483 <= $signed($unsigned(reg375[(1'h1):(1'h1)]));
                      reg484 <= (+$signed((8'hb3)));
                    end
                  reg485 <= ($unsigned(((forvar301 ?
                          reg56 : (8'hb0)) <<< reg416[(2'h3):(2'h3)])) ?
                      (forvar267 ?
                          reg287 : $unsigned(reg422)) : $signed((~|(forvar439 ?
                          reg389 : reg135))));
                end
              else
                begin
                  reg481 <= (|(^$signed((~^reg377))));
                end
              for (forvar486 = (1'h0); (forvar486 < (2'h2)); forvar486 = (forvar486 + (1'h1)))
                begin
                  reg487 <= $signed({$signed((forvar244 ^ (8'hb1)))});
                end
              reg488 <= $signed((((reg76 | (8'ha7)) & ((8'ha9) ?
                  reg341 : forvar418)) || $signed((8'hb2))));
            end
          for (forvar489 = (1'h0); (forvar489 < (1'h0)); forvar489 = (forvar489 + (1'h1)))
            begin
              for (forvar490 = (1'h0); (forvar490 < (1'h0)); forvar490 = (forvar490 + (1'h1)))
                begin
                  for (forvar491 = (1'h0); (forvar491 < (1'h1)); forvar491 = (forvar491 + (1'h1)))
                    begin
                      reg492 <= $signed($signed(reg275));
                      reg493 <= $signed(forvar423[(4'hb):(4'ha)]);
                      reg494 <= reg446;
                      reg495 <= (&(+reg384));
                    end
                  reg496 <= reg276;
                  reg497 <= (|(^$signed((~&forvar79))));
                end
              for (forvar498 = (1'h0); (forvar498 < (1'h0)); forvar498 = (forvar498 + (1'h1)))
                begin
                  reg499 <= reg220[(3'h4):(2'h3)];
                  for (forvar500 = (1'h0); (forvar500 < (1'h1)); forvar500 = (forvar500 + (1'h1)))
                    begin
                      reg501 <= reg17[(3'h7):(3'h4)];
                    end
                end
              reg502 <= $signed((($unsigned((8'h9c)) ? forvar185 : reg341) ?
                  reg157 : reg53[(2'h3):(2'h3)]));
              for (forvar503 = (1'h0); (forvar503 < (1'h0)); forvar503 = (forvar503 + (1'h1)))
                begin
                  for (forvar504 = (1'h0); (forvar504 < (2'h3)); forvar504 = (forvar504 + (1'h1)))
                    begin
                      reg505 <= reg368;
                      reg506 <= (8'ha6);
                    end
                  for (forvar507 = (1'h0); (forvar507 < (1'h0)); forvar507 = (forvar507 + (1'h1)))
                    begin
                      reg508 <= wire321[(2'h3):(1'h0)];
                    end
                end
            end
        end
      for (forvar509 = (1'h0); (forvar509 < (1'h0)); forvar509 = (forvar509 + (1'h1)))
        begin
          if (reg396[(4'h9):(2'h2)])
            begin
              if ((~^(($unsigned(forvar301) <= $signed(reg423)) && $unsigned($unsigned(reg12)))))
                begin
                  for (forvar510 = (1'h0); (forvar510 < (2'h3)); forvar510 = (forvar510 + (1'h1)))
                    begin
                      reg511 <= (reg87[(1'h0):(1'h0)] ?
                          $signed($unsigned($unsigned(reg145))) : forvar413);
                      reg512 <= reg499;
                      reg513 <= reg173[(1'h1):(1'h0)];
                    end
                  reg514 <= (~&(~&(&(-forvar401))));
                end
              else
                begin
                  if (({($unsigned((8'ha2)) ? {reg472} : reg442)} ?
                      $signed($unsigned($unsigned((8'hb1)))) : $signed(reg208[(2'h2):(2'h2)])))
                    begin
                      reg510 <= (~&($unsigned($signed((8'haa))) ?
                          $unsigned($signed(reg115)) : reg385));
                      reg511 <= {$unsigned((reg495[(3'h4):(1'h1)] ?
                              reg406 : reg95[(4'hb):(4'h9)]))};
                      reg512 <= (~&forvar61);
                      reg513 <= reg470[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg510 <= ($signed((((8'hb6) ?
                              reg28 : (8'ha7)) + $signed(forvar110))) ?
                          $signed({{reg159}}) : {forvar290});
                    end
                end
            end
          else
            begin
              reg510 <= forvar194[(4'hb):(4'h9)];
              for (forvar511 = (1'h0); (forvar511 < (2'h3)); forvar511 = (forvar511 + (1'h1)))
                begin
                  reg512 <= $signed(reg482);
                  reg513 <= {({$unsigned(reg16)} >>> ($unsigned(reg35) ?
                          (8'ha8) : {forvar507}))};
                end
              for (forvar514 = (1'h0); (forvar514 < (2'h3)); forvar514 = (forvar514 + (1'h1)))
                begin
                  for (forvar515 = (1'h0); (forvar515 < (2'h3)); forvar515 = (forvar515 + (1'h1)))
                    begin
                      reg516 <= ((+reg354[(3'h6):(3'h4)]) + $signed(($unsigned(forvar232) ?
                          (~(8'ha2)) : (&(8'hab)))));
                      reg517 <= $signed((+forvar424));
                      reg518 <= $signed({forvar69[(4'h9):(4'h8)]});
                    end
                  reg519 <= $signed((8'ha5));
                end
              if ((reg116 <= (!{$signed(forvar510)})))
                begin
                  for (forvar520 = (1'h0); (forvar520 < (2'h2)); forvar520 = (forvar520 + (1'h1)))
                    begin
                      reg521 <= $signed((+(|(reg408 <= reg417))));
                      reg522 <= ((forvar418 ?
                              reg66[(1'h0):(1'h0)] : (reg445 <<< (reg343 ?
                                  reg41 : reg37))) ?
                          $unsigned(reg211[(2'h3):(2'h2)]) : $signed({reg302}));
                      reg523 <= (!(reg280[(2'h2):(2'h2)] ^~ reg43[(2'h2):(1'h0)]));
                    end
                  reg524 <= (forvar131 ?
                      $signed(((reg151 || reg50) ^~ ((8'ha6) ~^ forvar481))) : $signed($signed((reg191 ?
                          reg178 : reg252))));
                end
              else
                begin
                  if ((reg488 <= reg480[(1'h0):(1'h0)]))
                    begin
                      reg520 <= (reg171[(3'h6):(3'h6)] ?
                          reg481 : forvar119[(3'h4):(1'h1)]);
                      reg521 <= reg222;
                      reg522 <= $signed(((~reg55[(2'h2):(1'h0)]) ?
                          (+((8'ha5) ? reg434 : reg511)) : {(8'hae)}));
                      reg523 <= $signed(reg210);
                    end
                  else
                    begin
                      reg520 <= $signed(($signed((8'ha6)) - (~^forvar503)));
                      reg521 <= $signed(($signed($signed(reg388)) ?
                          reg482[(3'h4):(3'h4)] : reg440[(2'h2):(1'h1)]));
                      reg522 <= (~($signed($signed(reg211)) ?
                          $signed(reg253) : ($signed((8'ha7)) ?
                              ((8'haf) ? (8'hb3) : reg146) : {reg319})));
                    end
                  reg524 <= {((&(reg13 ?
                          reg340 : reg485)) == $unsigned(reg47))};
                end
            end
          for (forvar525 = (1'h0); (forvar525 < (1'h0)); forvar525 = (forvar525 + (1'h1)))
            begin
              reg526 <= (8'ha9);
              if (reg213[(1'h0):(1'h0)])
                begin
                  reg527 <= (+(((reg111 != reg37) >> {reg526}) ?
                      $signed(forvar376[(2'h2):(1'h0)]) : $unsigned((reg118 != forvar40))));
                  for (forvar528 = (1'h0); (forvar528 < (1'h0)); forvar528 = (forvar528 + (1'h1)))
                    begin
                      reg529 <= forvar401;
                    end
                end
              else
                begin
                  for (forvar527 = (1'h0); (forvar527 < (1'h1)); forvar527 = (forvar527 + (1'h1)))
                    begin
                      reg528 <= $unsigned((reg348[(3'h7):(2'h3)] <<< $unsigned($signed(forvar20))));
                      reg529 <= forvar48[(1'h1):(1'h0)];
                    end
                  for (forvar530 = (1'h0); (forvar530 < (1'h0)); forvar530 = (forvar530 + (1'h1)))
                    begin
                      reg531 <= reg450;
                      reg532 <= $signed($signed(forvar190));
                      reg533 <= reg415[(3'h6):(1'h1)];
                    end
                  if ($unsigned((8'h9e)))
                    begin
                      reg534 <= {$unsigned(forvar79[(1'h1):(1'h0)])};
                    end
                  else
                    begin
                      reg534 <= (($signed({forvar491}) ?
                          $signed($unsigned(forvar43)) : {(8'h9d)}) << {reg257[(2'h2):(1'h0)]});
                      reg535 <= (((-(+forvar463)) ?
                              ($signed(reg481) ?
                                  ((8'hb3) ?
                                      (8'ha4) : forvar422) : $signed((8'hb9))) : $unsigned($unsigned(wire3))) ?
                          $unsigned((8'ha6)) : (^~$signed(reg339[(3'h4):(1'h0)])));
                    end
                  for (forvar536 = (1'h0); (forvar536 < (2'h2)); forvar536 = (forvar536 + (1'h1)))
                    begin
                      reg537 <= (($unsigned((forvar466 ?
                              (8'hba) : reg274)) != reg136) ?
                          $signed(reg389[(2'h3):(1'h1)]) : reg214[(2'h2):(1'h0)]);
                      reg538 <= $unsigned(forvar341);
                    end
                end
            end
          for (forvar539 = (1'h0); (forvar539 < (2'h2)); forvar539 = (forvar539 + (1'h1)))
            begin
              for (forvar540 = (1'h0); (forvar540 < (1'h1)); forvar540 = (forvar540 + (1'h1)))
                begin
                  for (forvar541 = (1'h0); (forvar541 < (1'h1)); forvar541 = (forvar541 + (1'h1)))
                    begin
                      reg542 <= ($signed(((8'ha5) ~^ reg438)) ?
                          (((&reg141) & forvar6[(4'ha):(4'h9)]) || reg166) : $signed(reg273[(2'h3):(1'h1)]));
                    end
                  for (forvar543 = (1'h0); (forvar543 < (2'h2)); forvar543 = (forvar543 + (1'h1)))
                    begin
                      reg544 <= reg14[(1'h1):(1'h0)];
                      reg545 <= forvar285[(3'h4):(2'h2)];
                    end
                  for (forvar546 = (1'h0); (forvar546 < (1'h0)); forvar546 = (forvar546 + (1'h1)))
                    begin
                      reg547 <= (((reg170 || (|reg483)) <= (reg103 ?
                              reg402[(1'h1):(1'h1)] : reg394[(2'h2):(1'h0)])) ?
                          (8'ha6) : (($signed(reg473) >> reg283) ?
                              (reg244[(1'h1):(1'h1)] ?
                                  (&forvar254) : (reg483 ?
                                      reg94 : (8'ha6))) : (reg87[(4'ha):(3'h7)] != forvar70)));
                      reg548 <= (forvar184 ?
                          $unsigned(($unsigned(reg36) + reg488)) : reg144);
                      reg549 <= $signed({(~&reg32[(3'h4):(2'h3)])});
                      reg550 <= ($unsigned((&(reg529 >>> reg431))) ?
                          ($unsigned((reg9 && reg531)) + ((reg38 ~^ (8'hb0)) >>> $signed(forvar206))) : ($signed($signed((8'ha7))) ?
                              (reg381 >= forvar536) : {reg472}));
                    end
                end
              reg551 <= (~(&$unsigned($signed(reg175))));
            end
        end
    end
  assign wire552 = (~^($signed($signed((8'ha2))) == $signed(reg467)));
  assign wire553 = ($unsigned((reg510 && (forvar263 ? forvar294 : forvar52))) ?
                       (($signed(forvar540) <= (reg263 - reg459)) ?
                           ({reg173} && (8'hb1)) : (+reg179)) : (8'h9d));
  module554 modinst5738 (.wire556(reg549), .y(wire5737), .wire555(reg357), .wire558(reg66), .wire557(reg435), .clk(clk));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module554
#(parameter param5736 = ({(-{(8'ha1)})} >> ((8'ha1) - ((8'haa) < (!(8'ha4))))))
(y, clk, wire558, wire557, wire556, wire555);
  output wire [(32'h1e01):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire558;
  input wire signed [(3'h6):(1'h0)] wire557;
  input wire [(2'h3):(1'h0)] wire556;
  input wire signed [(4'h9):(1'h0)] wire555;
  reg [(3'h7):(1'h0)] reg5735 = (1'h0);
  reg [(4'h9):(1'h0)] reg5734 = (1'h0);
  reg [(3'h4):(1'h0)] reg5733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5732 = (1'h0);
  reg [(4'ha):(1'h0)] reg5731 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5730 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5729 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5725 = (1'h0);
  reg [(4'he):(1'h0)] reg5722 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5717 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5713 = (1'h0);
  reg [(5'h10):(1'h0)] reg5712 = (1'h0);
  reg [(4'he):(1'h0)] forvar5702 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5698 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5694 = (1'h0);
  reg [(4'h9):(1'h0)] reg5693 = (1'h0);
  reg [(3'h4):(1'h0)] reg5707 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5705 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5703 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5701 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5697 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5692 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5688 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5686 = (1'h0);
  reg [(5'h10):(1'h0)] reg5682 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5679 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5678 = (1'h0);
  reg [(3'h4):(1'h0)] reg5677 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5670 = (1'h0);
  reg [(4'hd):(1'h0)] reg5669 = (1'h0);
  reg [(3'h4):(1'h0)] reg5730 = (1'h0);
  reg [(3'h4):(1'h0)] reg5729 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5728 = (1'h0);
  reg [(4'hb):(1'h0)] reg5727 = (1'h0);
  reg [(4'he):(1'h0)] reg5726 = (1'h0);
  reg [(2'h2):(1'h0)] reg5725 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5724 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5723 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5722 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5721 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5720 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5719 = (1'h0);
  reg [(3'h6):(1'h0)] reg5718 = (1'h0);
  reg [(5'h10):(1'h0)] reg5715 = (1'h0);
  reg [(4'h9):(1'h0)] reg5717 = (1'h0);
  reg [(4'hb):(1'h0)] reg5716 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5715 = (1'h0);
  reg [(4'h9):(1'h0)] reg5714 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5713 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5712 = (1'h0);
  reg [(5'h10):(1'h0)] reg5711 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5710 = (1'h0);
  reg [(4'h8):(1'h0)] reg5709 = (1'h0);
  reg [(2'h3):(1'h0)] reg5708 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5707 = (1'h0);
  reg [(3'h6):(1'h0)] reg5706 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5705 = (1'h0);
  reg [(4'h8):(1'h0)] reg5704 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5703 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5702 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5701 = (1'h0);
  reg [(4'hc):(1'h0)] reg5700 = (1'h0);
  reg [(5'h10):(1'h0)] reg5699 = (1'h0);
  reg [(3'h4):(1'h0)] reg5698 = (1'h0);
  reg [(3'h6):(1'h0)] reg5697 = (1'h0);
  reg [(4'hb):(1'h0)] reg5696 = (1'h0);
  reg [(3'h4):(1'h0)] reg5695 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5694 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5693 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5692 = (1'h0);
  reg [(5'h10):(1'h0)] reg5691 = (1'h0);
  reg [(4'hd):(1'h0)] reg5690 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5689 = (1'h0);
  reg [(4'h9):(1'h0)] reg5688 = (1'h0);
  reg [(4'h9):(1'h0)] reg5687 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5686 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5685 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5684 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5683 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5682 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5681 = (1'h0);
  reg [(4'he):(1'h0)] reg5680 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5679 = (1'h0);
  reg [(4'hd):(1'h0)] reg5678 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5677 = (1'h0);
  reg [(4'h8):(1'h0)] reg5676 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5675 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5674 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5673 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5672 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5671 = (1'h0);
  reg [(4'h8):(1'h0)] reg5670 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5669 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5668 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5667 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5660 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5666 = (1'h0);
  reg [(3'h4):(1'h0)] reg5665 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5664 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5663 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5662 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5661 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5660 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5659 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5654 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5649 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5658 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5657 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5656 = (1'h0);
  reg [(2'h2):(1'h0)] reg5655 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5654 = (1'h0);
  reg [(4'hb):(1'h0)] reg5653 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5650 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5652 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5651 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5650 = (1'h0);
  reg [(4'h8):(1'h0)] reg5649 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5648 = (1'h0);
  wire [(4'hd):(1'h0)] wire5647;
  reg signed [(2'h2):(1'h0)] reg5646 = (1'h0);
  reg [(4'hb):(1'h0)] reg5645 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5644 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5643 = (1'h0);
  reg [(4'hc):(1'h0)] reg5642 = (1'h0);
  reg [(3'h7):(1'h0)] reg5641 = (1'h0);
  reg [(3'h4):(1'h0)] reg5640 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5639 = (1'h0);
  reg [(3'h4):(1'h0)] reg5638 = (1'h0);
  reg [(3'h6):(1'h0)] reg5637 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5636 = (1'h0);
  reg [(4'hf):(1'h0)] reg5635 = (1'h0);
  reg [(4'he):(1'h0)] reg5634 = (1'h0);
  reg [(4'hb):(1'h0)] reg5633 = (1'h0);
  reg [(4'hf):(1'h0)] reg5632 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5630 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5631 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5630 = (1'h0);
  reg [(2'h3):(1'h0)] reg5629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5628 = (1'h0);
  reg [(4'ha):(1'h0)] reg5627 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5626 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5625 = (1'h0);
  reg [(4'hc):(1'h0)] reg5624 = (1'h0);
  reg [(2'h3):(1'h0)] reg5623 = (1'h0);
  reg [(3'h5):(1'h0)] reg5622 = (1'h0);
  reg [(4'ha):(1'h0)] reg5621 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5620 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5617 = (1'h0);
  reg [(4'hf):(1'h0)] reg5615 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5612 = (1'h0);
  reg [(3'h7):(1'h0)] reg5620 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5619 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5618 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5617 = (1'h0);
  reg [(4'hb):(1'h0)] reg5616 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5615 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5614 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5613 = (1'h0);
  reg [(4'ha):(1'h0)] reg5612 = (1'h0);
  reg [(4'hc):(1'h0)] reg5611 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5610 = (1'h0);
  reg [(4'h8):(1'h0)] reg5609 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5608 = (1'h0);
  reg [(3'h7):(1'h0)] reg5607 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5606 = (1'h0);
  reg [(2'h3):(1'h0)] reg5605 = (1'h0);
  reg [(3'h5):(1'h0)] reg5604 = (1'h0);
  reg [(4'hf):(1'h0)] reg5603 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5602 = (1'h0);
  reg [(4'he):(1'h0)] forvar5601 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5600 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5591 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5588 = (1'h0);
  reg [(4'h9):(1'h0)] reg5586 = (1'h0);
  reg [(5'h10):(1'h0)] reg5599 = (1'h0);
  reg [(3'h4):(1'h0)] reg5598 = (1'h0);
  reg [(4'hc):(1'h0)] reg5597 = (1'h0);
  reg [(4'hc):(1'h0)] reg5596 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5595 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5594 = (1'h0);
  reg [(4'hd):(1'h0)] reg5593 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5592 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5591 = (1'h0);
  reg [(4'h9):(1'h0)] reg5590 = (1'h0);
  reg [(4'h8):(1'h0)] reg5589 = (1'h0);
  reg [(5'h10):(1'h0)] reg5588 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5587 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5586 = (1'h0);
  reg [(4'ha):(1'h0)] reg5585 = (1'h0);
  reg [(5'h10):(1'h0)] reg5584 = (1'h0);
  reg [(4'he):(1'h0)] forvar5583 = (1'h0);
  reg [(4'h9):(1'h0)] reg5581 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5579 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5582 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5581 = (1'h0);
  reg [(5'h10):(1'h0)] reg5580 = (1'h0);
  reg [(4'he):(1'h0)] forvar5579 = (1'h0);
  reg [(5'h10):(1'h0)] reg5578 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5577 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5576 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5575 = (1'h0);
  reg [(4'hd):(1'h0)] reg5574 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5573 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5572 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5571 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5570 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5569 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5568 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5567 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5564 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5557 = (1'h0);
  reg [(4'h9):(1'h0)] reg5561 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5559 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5566 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5565 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5564 = (1'h0);
  reg [(2'h2):(1'h0)] reg5563 = (1'h0);
  reg [(4'ha):(1'h0)] reg5562 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5561 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5560 = (1'h0);
  reg [(4'ha):(1'h0)] reg5559 = (1'h0);
  reg [(4'hb):(1'h0)] reg5558 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5557 = (1'h0);
  reg [(4'ha):(1'h0)] reg5556 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5555 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5554 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5553 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5552 = (1'h0);
  reg [(4'hd):(1'h0)] reg5551 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5550 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5549 = (1'h0);
  reg [(5'h10):(1'h0)] reg5548 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5547 = (1'h0);
  reg [(5'h10):(1'h0)] reg5546 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5545 = (1'h0);
  reg [(3'h6):(1'h0)] reg5544 = (1'h0);
  reg [(2'h3):(1'h0)] reg5543 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5542 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5541 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5540 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5539 = (1'h0);
  reg [(5'h10):(1'h0)] reg5538 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5537 = (1'h0);
  reg [(5'h10):(1'h0)] reg5536 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5535 = (1'h0);
  reg [(3'h7):(1'h0)] reg5534 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5533 = (1'h0);
  reg [(4'h8):(1'h0)] reg5533 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5532 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire5531;
  wire [(3'h4):(1'h0)] wire5530;
  wire signed [(4'h9):(1'h0)] wire5529;
  wire signed [(3'h6):(1'h0)] wire5528;
  wire signed [(3'h4):(1'h0)] wire5527;
  wire [(4'hc):(1'h0)] wire5526;
  wire signed [(4'hd):(1'h0)] wire5524;
  wire [(5'h10):(1'h0)] wire1020;
  reg signed [(4'hd):(1'h0)] forvar961 = (1'h0);
  reg [(4'hb):(1'h0)] reg969 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar963 = (1'h0);
  reg [(2'h3):(1'h0)] reg962 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg956 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar955 = (1'h0);
  reg [(2'h3):(1'h0)] reg954 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg952 = (1'h0);
  reg [(4'hf):(1'h0)] reg1019 = (1'h0);
  reg [(4'ha):(1'h0)] reg1018 = (1'h0);
  reg [(4'hd):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1016 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1015 = (1'h0);
  reg [(4'h9):(1'h0)] reg1014 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1013 = (1'h0);
  reg [(4'h8):(1'h0)] reg1012 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1011 = (1'h0);
  reg [(4'hb):(1'h0)] reg1010 = (1'h0);
  reg [(2'h2):(1'h0)] reg1009 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1008 = (1'h0);
  reg [(4'hd):(1'h0)] reg1007 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1006 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1005 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1004 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1003 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1002 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1001 = (1'h0);
  reg [(4'h8):(1'h0)] reg1000 = (1'h0);
  reg [(2'h2):(1'h0)] reg999 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar998 = (1'h0);
  reg [(5'h10):(1'h0)] forvar997 = (1'h0);
  reg [(3'h6):(1'h0)] forvar996 = (1'h0);
  reg [(3'h4):(1'h0)] reg995 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg994 = (1'h0);
  reg [(4'hd):(1'h0)] reg993 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg992 = (1'h0);
  reg [(4'he):(1'h0)] forvar991 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg990 = (1'h0);
  reg [(5'h10):(1'h0)] reg989 = (1'h0);
  reg [(4'ha):(1'h0)] reg988 = (1'h0);
  reg [(4'he):(1'h0)] forvar987 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg986 = (1'h0);
  reg [(4'hb):(1'h0)] reg985 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg984 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar980 = (1'h0);
  reg [(3'h5):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg982 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg981 = (1'h0);
  reg [(4'hc):(1'h0)] reg980 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg975 = (1'h0);
  reg [(5'h10):(1'h0)] reg971 = (1'h0);
  reg [(2'h2):(1'h0)] reg979 = (1'h0);
  reg [(2'h2):(1'h0)] reg978 = (1'h0);
  reg [(5'h10):(1'h0)] reg977 = (1'h0);
  reg [(4'hb):(1'h0)] reg976 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar975 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg974 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg973 = (1'h0);
  reg [(3'h5):(1'h0)] reg972 = (1'h0);
  reg [(4'hd):(1'h0)] forvar971 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg970 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar969 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg968 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg967 = (1'h0);
  reg [(3'h6):(1'h0)] reg966 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar965 = (1'h0);
  reg [(3'h7):(1'h0)] reg964 = (1'h0);
  reg [(4'h9):(1'h0)] reg963 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar962 = (1'h0);
  reg [(3'h5):(1'h0)] reg961 = (1'h0);
  reg [(3'h4):(1'h0)] forvar960 = (1'h0);
  reg [(4'he):(1'h0)] reg960 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg959 = (1'h0);
  reg [(4'hf):(1'h0)] reg958 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg957 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar956 = (1'h0);
  reg [(4'hc):(1'h0)] reg955 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar954 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar953 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar952 = (1'h0);
  reg [(4'he):(1'h0)] forvar900 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar931 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg926 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg925 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar924 = (1'h0);
  reg [(4'ha):(1'h0)] reg922 = (1'h0);
  reg [(2'h2):(1'h0)] reg920 = (1'h0);
  reg [(2'h3):(1'h0)] forvar919 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg918 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg917 = (1'h0);
  reg [(4'h9):(1'h0)] reg907 = (1'h0);
  reg [(4'he):(1'h0)] reg906 = (1'h0);
  reg [(2'h3):(1'h0)] forvar902 = (1'h0);
  reg [(4'hc):(1'h0)] forvar892 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar885 = (1'h0);
  reg [(4'hd):(1'h0)] reg951 = (1'h0);
  reg [(3'h7):(1'h0)] reg942 = (1'h0);
  reg [(3'h5):(1'h0)] reg950 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg949 = (1'h0);
  reg [(4'h9):(1'h0)] reg948 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg947 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg946 = (1'h0);
  reg [(4'hf):(1'h0)] forvar945 = (1'h0);
  reg [(3'h5):(1'h0)] reg944 = (1'h0);
  reg [(4'hc):(1'h0)] reg943 = (1'h0);
  reg [(4'h9):(1'h0)] forvar942 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg941 = (1'h0);
  reg [(4'hb):(1'h0)] reg940 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg939 = (1'h0);
  reg [(4'h9):(1'h0)] reg938 = (1'h0);
  reg [(3'h4):(1'h0)] reg937 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg936 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg935 = (1'h0);
  reg [(4'hb):(1'h0)] reg934 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg933 = (1'h0);
  reg [(4'hf):(1'h0)] reg932 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg931 = (1'h0);
  reg [(5'h10):(1'h0)] reg930 = (1'h0);
  reg [(5'h10):(1'h0)] reg929 = (1'h0);
  reg [(4'h8):(1'h0)] reg928 = (1'h0);
  reg [(3'h7):(1'h0)] forvar927 = (1'h0);
  reg [(4'h9):(1'h0)] forvar926 = (1'h0);
  reg [(3'h5):(1'h0)] forvar925 = (1'h0);
  reg [(4'ha):(1'h0)] reg924 = (1'h0);
  reg [(3'h4):(1'h0)] reg923 = (1'h0);
  reg [(2'h3):(1'h0)] forvar922 = (1'h0);
  reg [(3'h5):(1'h0)] reg921 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar920 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg919 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar918 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar917 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg915 = (1'h0);
  reg [(2'h2):(1'h0)] reg914 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg913 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg912 = (1'h0);
  reg [(3'h7):(1'h0)] forvar911 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg910 = (1'h0);
  reg [(4'he):(1'h0)] reg909 = (1'h0);
  reg [(3'h6):(1'h0)] reg908 = (1'h0);
  reg [(4'h9):(1'h0)] forvar907 = (1'h0);
  reg [(2'h3):(1'h0)] forvar906 = (1'h0);
  reg [(3'h7):(1'h0)] reg901 = (1'h0);
  reg [(3'h4):(1'h0)] forvar899 = (1'h0);
  reg [(2'h3):(1'h0)] forvar897 = (1'h0);
  reg [(4'h8):(1'h0)] reg905 = (1'h0);
  reg [(4'h9):(1'h0)] reg904 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg903 = (1'h0);
  reg [(3'h5):(1'h0)] reg902 = (1'h0);
  reg [(3'h7):(1'h0)] forvar901 = (1'h0);
  reg [(2'h2):(1'h0)] forvar895 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg894 = (1'h0);
  reg [(2'h2):(1'h0)] forvar893 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg889 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg888 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar887 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg886 = (1'h0);
  reg [(3'h6):(1'h0)] forvar884 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg900 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg899 = (1'h0);
  reg [(4'h9):(1'h0)] reg898 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg897 = (1'h0);
  reg [(4'hf):(1'h0)] reg896 = (1'h0);
  reg [(4'hd):(1'h0)] reg895 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar894 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg893 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg892 = (1'h0);
  reg [(3'h5):(1'h0)] reg891 = (1'h0);
  reg [(3'h7):(1'h0)] reg890 = (1'h0);
  reg [(4'hb):(1'h0)] forvar889 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar888 = (1'h0);
  reg [(4'h8):(1'h0)] reg887 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar886 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg885 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg884 = (1'h0);
  reg [(4'ha):(1'h0)] forvar883 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg882 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar881 = (1'h0);
  reg [(3'h6):(1'h0)] reg880 = (1'h0);
  reg [(2'h3):(1'h0)] reg879 = (1'h0);
  reg [(4'h8):(1'h0)] reg878 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg877 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg876 = (1'h0);
  reg signed [(4'he):(1'h0)] reg875 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg874 = (1'h0);
  reg [(3'h7):(1'h0)] reg872 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar871 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar870 = (1'h0);
  reg [(3'h7):(1'h0)] reg867 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar866 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar865 = (1'h0);
  reg [(2'h2):(1'h0)] forvar862 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar858 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg851 = (1'h0);
  reg signed [(4'he):(1'h0)] reg863 = (1'h0);
  reg [(4'h9):(1'h0)] forvar861 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg859 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg873 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar872 = (1'h0);
  reg [(4'he):(1'h0)] reg871 = (1'h0);
  reg [(4'hd):(1'h0)] reg870 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg869 = (1'h0);
  reg signed [(4'he):(1'h0)] reg868 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar867 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg866 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg865 = (1'h0);
  reg [(4'hb):(1'h0)] reg864 = (1'h0);
  reg [(4'h9):(1'h0)] forvar863 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg862 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg861 = (1'h0);
  reg [(3'h7):(1'h0)] reg860 = (1'h0);
  reg [(4'hb):(1'h0)] forvar859 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar853 = (1'h0);
  reg [(4'he):(1'h0)] reg858 = (1'h0);
  reg [(4'hc):(1'h0)] reg857 = (1'h0);
  reg [(2'h3):(1'h0)] reg856 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg855 = (1'h0);
  reg [(2'h2):(1'h0)] reg854 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg853 = (1'h0);
  reg [(5'h10):(1'h0)] reg852 = (1'h0);
  reg [(3'h6):(1'h0)] forvar851 = (1'h0);
  reg [(4'hb):(1'h0)] forvar843 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar836 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar834 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar831 = (1'h0);
  reg [(4'he):(1'h0)] reg832 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg829 = (1'h0);
  reg [(4'ha):(1'h0)] reg828 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg844 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar840 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg850 = (1'h0);
  reg signed [(4'he):(1'h0)] reg849 = (1'h0);
  reg [(2'h2):(1'h0)] reg848 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg847 = (1'h0);
  reg [(4'hd):(1'h0)] reg846 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg845 = (1'h0);
  reg [(3'h7):(1'h0)] forvar844 = (1'h0);
  reg [(2'h2):(1'h0)] reg843 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg842 = (1'h0);
  reg [(3'h4):(1'h0)] reg841 = (1'h0);
  reg [(3'h7):(1'h0)] reg840 = (1'h0);
  reg [(3'h4):(1'h0)] reg839 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg838 = (1'h0);
  reg [(4'he):(1'h0)] reg837 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg836 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg835 = (1'h0);
  reg [(3'h7):(1'h0)] reg834 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg833 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar832 = (1'h0);
  reg [(4'ha):(1'h0)] reg831 = (1'h0);
  reg [(4'hd):(1'h0)] reg830 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar829 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar828 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg827 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg826 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg825 = (1'h0);
  reg [(4'ha):(1'h0)] forvar824 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg823 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg822 = (1'h0);
  reg [(4'hc):(1'h0)] reg821 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg820 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar819 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg818 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg817 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg816 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg815 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar814 = (1'h0);
  reg [(4'hc):(1'h0)] reg813 = (1'h0);
  reg [(4'hf):(1'h0)] reg812 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar811 = (1'h0);
  reg [(4'hb):(1'h0)] reg810 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg809 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg808 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg807 = (1'h0);
  reg [(2'h2):(1'h0)] forvar806 = (1'h0);
  reg [(3'h7):(1'h0)] reg806 = (1'h0);
  reg [(2'h2):(1'h0)] reg805 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg804 = (1'h0);
  reg [(4'ha):(1'h0)] reg803 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg802 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg801 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg800 = (1'h0);
  reg [(4'h9):(1'h0)] reg799 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar798 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg797 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg796 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg795 = (1'h0);
  reg [(4'hf):(1'h0)] reg794 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg793 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg792 = (1'h0);
  reg [(3'h7):(1'h0)] reg791 = (1'h0);
  reg [(4'hd):(1'h0)] forvar790 = (1'h0);
  reg [(3'h4):(1'h0)] reg789 = (1'h0);
  reg [(4'ha):(1'h0)] reg788 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar787 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg786 = (1'h0);
  reg [(4'hc):(1'h0)] reg785 = (1'h0);
  reg [(4'hb):(1'h0)] forvar784 = (1'h0);
  reg [(4'h8):(1'h0)] forvar783 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg782 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg781 = (1'h0);
  reg [(3'h6):(1'h0)] reg780 = (1'h0);
  reg [(4'hb):(1'h0)] reg779 = (1'h0);
  reg [(4'h8):(1'h0)] forvar778 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg777 = (1'h0);
  reg [(4'h9):(1'h0)] reg776 = (1'h0);
  reg [(4'hb):(1'h0)] forvar775 = (1'h0);
  reg [(3'h6):(1'h0)] reg774 = (1'h0);
  reg [(2'h3):(1'h0)] forvar771 = (1'h0);
  reg [(4'hb):(1'h0)] reg773 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg772 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg771 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar770 = (1'h0);
  reg [(4'hc):(1'h0)] forvar746 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg748 = (1'h0);
  reg [(4'hb):(1'h0)] forvar742 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg741 = (1'h0);
  reg [(3'h7):(1'h0)] reg769 = (1'h0);
  reg [(4'hb):(1'h0)] forvar768 = (1'h0);
  reg [(3'h6):(1'h0)] reg767 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg766 = (1'h0);
  reg [(4'h9):(1'h0)] reg765 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg764 = (1'h0);
  reg [(4'hc):(1'h0)] forvar763 = (1'h0);
  reg [(4'he):(1'h0)] reg761 = (1'h0);
  reg [(4'he):(1'h0)] forvar759 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg756 = (1'h0);
  reg [(4'hc):(1'h0)] reg763 = (1'h0);
  reg [(4'hf):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar761 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg760 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg759 = (1'h0);
  reg [(4'hb):(1'h0)] reg758 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg757 = (1'h0);
  reg [(3'h4):(1'h0)] forvar756 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg755 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg754 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg753 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg752 = (1'h0);
  reg [(4'hd):(1'h0)] reg751 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg750 = (1'h0);
  reg [(3'h6):(1'h0)] reg749 = (1'h0);
  reg [(4'hc):(1'h0)] forvar748 = (1'h0);
  reg [(3'h7):(1'h0)] reg747 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg746 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar745 = (1'h0);
  reg [(4'h9):(1'h0)] reg745 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg744 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg743 = (1'h0);
  reg [(3'h6):(1'h0)] reg742 = (1'h0);
  reg [(5'h10):(1'h0)] forvar741 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg740 = (1'h0);
  reg [(2'h2):(1'h0)] reg739 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg738 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar737 = (1'h0);
  reg [(4'hc):(1'h0)] reg736 = (1'h0);
  reg [(3'h7):(1'h0)] reg735 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg734 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar733 = (1'h0);
  reg [(4'hd):(1'h0)] forvar731 = (1'h0);
  reg [(3'h6):(1'h0)] reg732 = (1'h0);
  reg [(4'hb):(1'h0)] reg731 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar730 = (1'h0);
  reg [(4'he):(1'h0)] reg729 = (1'h0);
  reg [(5'h10):(1'h0)] reg728 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg727 = (1'h0);
  reg [(4'hb):(1'h0)] reg726 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg725 = (1'h0);
  reg [(4'h9):(1'h0)] reg724 = (1'h0);
  reg signed [(4'he):(1'h0)] reg723 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar722 = (1'h0);
  reg [(4'he):(1'h0)] reg721 = (1'h0);
  reg [(2'h3):(1'h0)] reg720 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg719 = (1'h0);
  reg [(3'h6):(1'h0)] reg718 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg717 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg716 = (1'h0);
  reg [(3'h7):(1'h0)] reg715 = (1'h0);
  reg [(3'h5):(1'h0)] reg714 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar713 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg712 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar711 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg710 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg709 = (1'h0);
  reg [(2'h3):(1'h0)] reg708 = (1'h0);
  reg [(3'h7):(1'h0)] forvar707 = (1'h0);
  reg [(5'h10):(1'h0)] reg704 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar702 = (1'h0);
  reg [(3'h5):(1'h0)] forvar700 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg707 = (1'h0);
  reg [(5'h10):(1'h0)] reg706 = (1'h0);
  reg [(4'hc):(1'h0)] reg705 = (1'h0);
  reg [(4'ha):(1'h0)] forvar704 = (1'h0);
  reg [(4'he):(1'h0)] reg703 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg702 = (1'h0);
  reg [(4'hd):(1'h0)] reg701 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg700 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar699 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar695 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar693 = (1'h0);
  reg [(4'hb):(1'h0)] forvar689 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar688 = (1'h0);
  reg [(3'h5):(1'h0)] reg698 = (1'h0);
  reg [(4'h8):(1'h0)] forvar697 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg696 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg695 = (1'h0);
  reg signed [(4'he):(1'h0)] reg694 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg693 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg692 = (1'h0);
  reg [(3'h4):(1'h0)] reg691 = (1'h0);
  reg [(3'h6):(1'h0)] forvar687 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg689 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg688 = (1'h0);
  reg [(4'hb):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg686 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg685 = (1'h0);
  reg [(4'ha):(1'h0)] reg684 = (1'h0);
  reg [(4'hb):(1'h0)] reg683 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar682 = (1'h0);
  reg [(4'hd):(1'h0)] forvar681 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg680 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar676 = (1'h0);
  reg [(3'h4):(1'h0)] reg674 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar671 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar650 = (1'h0);
  reg [(3'h6):(1'h0)] forvar648 = (1'h0);
  reg [(4'hf):(1'h0)] forvar644 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg669 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg664 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar661 = (1'h0);
  reg signed [(4'he):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar656 = (1'h0);
  reg [(3'h7):(1'h0)] reg655 = (1'h0);
  reg [(5'h10):(1'h0)] forvar652 = (1'h0);
  reg [(2'h3):(1'h0)] forvar649 = (1'h0);
  reg [(4'hb):(1'h0)] reg647 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg660 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg679 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg678 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg677 = (1'h0);
  reg [(3'h7):(1'h0)] reg676 = (1'h0);
  reg [(3'h7):(1'h0)] reg675 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar674 = (1'h0);
  reg [(3'h6):(1'h0)] reg673 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg672 = (1'h0);
  reg [(4'hd):(1'h0)] reg671 = (1'h0);
  reg [(3'h6):(1'h0)] reg670 = (1'h0);
  reg [(3'h6):(1'h0)] forvar669 = (1'h0);
  reg [(3'h6):(1'h0)] forvar668 = (1'h0);
  reg [(5'h10):(1'h0)] reg667 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg666 = (1'h0);
  reg [(4'hd):(1'h0)] reg665 = (1'h0);
  reg [(2'h2):(1'h0)] forvar664 = (1'h0);
  reg [(4'he):(1'h0)] reg663 = (1'h0);
  reg signed [(4'he):(1'h0)] reg662 = (1'h0);
  reg [(4'h9):(1'h0)] reg661 = (1'h0);
  reg [(3'h7):(1'h0)] forvar660 = (1'h0);
  reg [(4'ha):(1'h0)] forvar659 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg658 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg657 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg656 = (1'h0);
  reg [(3'h6):(1'h0)] forvar655 = (1'h0);
  reg [(2'h3):(1'h0)] reg654 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg653 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg652 = (1'h0);
  reg [(4'he):(1'h0)] reg651 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg650 = (1'h0);
  reg [(4'hb):(1'h0)] reg649 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg648 = (1'h0);
  reg [(4'hf):(1'h0)] forvar647 = (1'h0);
  reg [(4'h9):(1'h0)] reg646 = (1'h0);
  reg [(4'hb):(1'h0)] reg645 = (1'h0);
  reg [(4'h8):(1'h0)] reg644 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar643 = (1'h0);
  reg [(4'ha):(1'h0)] reg643 = (1'h0);
  reg [(4'ha):(1'h0)] reg642 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar641 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar640 = (1'h0);
  reg [(4'he):(1'h0)] reg639 = (1'h0);
  reg [(2'h3):(1'h0)] forvar638 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg637 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg636 = (1'h0);
  reg [(3'h7):(1'h0)] reg635 = (1'h0);
  reg [(4'h8):(1'h0)] reg634 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar633 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg632 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar631 = (1'h0);
  reg [(4'hf):(1'h0)] forvar630 = (1'h0);
  reg [(3'h6):(1'h0)] forvar629 = (1'h0);
  reg signed [(4'he):(1'h0)] reg628 = (1'h0);
  reg [(4'ha):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar626 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg625 = (1'h0);
  reg [(4'ha):(1'h0)] reg624 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg623 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg622 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar621 = (1'h0);
  reg [(4'hd):(1'h0)] forvar620 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg619 = (1'h0);
  reg [(2'h2):(1'h0)] reg618 = (1'h0);
  reg [(3'h4):(1'h0)] reg617 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg616 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar615 = (1'h0);
  reg [(4'he):(1'h0)] reg614 = (1'h0);
  reg [(4'h9):(1'h0)] reg613 = (1'h0);
  reg [(4'hc):(1'h0)] reg612 = (1'h0);
  reg [(4'h8):(1'h0)] forvar608 = (1'h0);
  reg [(4'hf):(1'h0)] reg611 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg610 = (1'h0);
  reg [(3'h7):(1'h0)] reg609 = (1'h0);
  reg [(4'ha):(1'h0)] reg608 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar607 = (1'h0);
  reg [(2'h3):(1'h0)] forvar602 = (1'h0);
  reg [(3'h7):(1'h0)] reg601 = (1'h0);
  reg [(4'ha):(1'h0)] reg606 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg605 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg604 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg603 = (1'h0);
  reg [(3'h7):(1'h0)] reg602 = (1'h0);
  reg [(4'he):(1'h0)] forvar601 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar600 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg599 = (1'h0);
  reg [(4'h8):(1'h0)] reg598 = (1'h0);
  reg [(4'h8):(1'h0)] reg597 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg592 = (1'h0);
  reg [(3'h5):(1'h0)] reg591 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg596 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar595 = (1'h0);
  reg [(4'hc):(1'h0)] reg594 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg593 = (1'h0);
  reg [(4'ha):(1'h0)] forvar592 = (1'h0);
  reg [(4'ha):(1'h0)] forvar591 = (1'h0);
  reg [(3'h4):(1'h0)] reg590 = (1'h0);
  reg [(4'h8):(1'h0)] forvar589 = (1'h0);
  reg [(4'he):(1'h0)] forvar588 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg587 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg586 = (1'h0);
  reg signed [(4'he):(1'h0)] reg585 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar584 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg583 = (1'h0);
  reg [(4'hd):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg581 = (1'h0);
  reg [(4'ha):(1'h0)] reg580 = (1'h0);
  reg [(5'h10):(1'h0)] forvar579 = (1'h0);
  reg [(4'h8):(1'h0)] reg578 = (1'h0);
  reg [(3'h5):(1'h0)] reg577 = (1'h0);
  reg [(4'ha):(1'h0)] forvar575 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar571 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg573 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar570 = (1'h0);
  reg [(3'h7):(1'h0)] reg576 = (1'h0);
  reg [(3'h6):(1'h0)] reg575 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg574 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar573 = (1'h0);
  reg [(4'ha):(1'h0)] reg567 = (1'h0);
  reg [(3'h6):(1'h0)] reg572 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg571 = (1'h0);
  reg [(4'he):(1'h0)] reg570 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg569 = (1'h0);
  reg [(4'h8):(1'h0)] reg568 = (1'h0);
  reg [(2'h2):(1'h0)] forvar567 = (1'h0);
  reg [(4'he):(1'h0)] reg566 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg565 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar564 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg563 = (1'h0);
  reg [(4'ha):(1'h0)] forvar562 = (1'h0);
  wire [(4'he):(1'h0)] wire561;
  wire signed [(3'h6):(1'h0)] wire560;
  wire signed [(4'h9):(1'h0)] wire559;
  assign y = {reg5735,
                 reg5734,
                 reg5733,
                 reg5732,
                 reg5731,
                 forvar5730,
                 forvar5729,
                 forvar5725,
                 reg5722,
                 forvar5717,
                 forvar5713,
                 reg5712,
                 forvar5702,
                 forvar5698,
                 forvar5694,
                 reg5693,
                 reg5707,
                 reg5705,
                 reg5703,
                 forvar5701,
                 forvar5697,
                 forvar5692,
                 forvar5688,
                 forvar5686,
                 reg5682,
                 forvar5679,
                 forvar5678,
                 reg5677,
                 forvar5670,
                 reg5669,
                 reg5730,
                 reg5729,
                 reg5728,
                 reg5727,
                 reg5726,
                 reg5725,
                 reg5724,
                 reg5723,
                 forvar5722,
                 reg5721,
                 reg5720,
                 reg5719,
                 reg5718,
                 reg5715,
                 reg5717,
                 reg5716,
                 forvar5715,
                 reg5714,
                 reg5713,
                 forvar5712,
                 reg5711,
                 reg5710,
                 reg5709,
                 reg5708,
                 forvar5707,
                 reg5706,
                 forvar5705,
                 reg5704,
                 forvar5703,
                 reg5702,
                 reg5701,
                 reg5700,
                 reg5699,
                 reg5698,
                 reg5697,
                 reg5696,
                 reg5695,
                 reg5694,
                 forvar5693,
                 reg5692,
                 reg5691,
                 reg5690,
                 reg5689,
                 reg5688,
                 reg5687,
                 reg5686,
                 reg5685,
                 forvar5684,
                 reg5683,
                 forvar5682,
                 reg5681,
                 reg5680,
                 reg5679,
                 reg5678,
                 forvar5677,
                 reg5676,
                 reg5675,
                 reg5674,
                 reg5673,
                 reg5672,
                 reg5671,
                 reg5670,
                 forvar5669,
                 forvar5668,
                 reg5667,
                 forvar5660,
                 reg5666,
                 reg5665,
                 reg5664,
                 reg5663,
                 reg5662,
                 reg5661,
                 reg5660,
                 reg5659,
                 reg5654,
                 forvar5649,
                 reg5658,
                 reg5657,
                 reg5656,
                 reg5655,
                 forvar5654,
                 reg5653,
                 forvar5650,
                 reg5652,
                 reg5651,
                 reg5650,
                 reg5649,
                 forvar5648,
                 wire5647,
                 reg5646,
                 reg5645,
                 forvar5644,
                 reg5643,
                 reg5642,
                 reg5641,
                 reg5640,
                 reg5639,
                 reg5638,
                 reg5637,
                 reg5636,
                 reg5635,
                 reg5634,
                 reg5633,
                 reg5632,
                 forvar5630,
                 reg5631,
                 reg5630,
                 reg5629,
                 reg5628,
                 reg5627,
                 reg5626,
                 forvar5625,
                 reg5624,
                 reg5623,
                 reg5622,
                 reg5621,
                 forvar5620,
                 forvar5617,
                 reg5615,
                 forvar5612,
                 reg5620,
                 reg5619,
                 reg5618,
                 reg5617,
                 reg5616,
                 forvar5615,
                 reg5614,
                 reg5613,
                 reg5612,
                 reg5611,
                 forvar5610,
                 reg5609,
                 reg5608,
                 reg5607,
                 forvar5606,
                 reg5605,
                 reg5604,
                 reg5603,
                 reg5602,
                 forvar5601,
                 forvar5600,
                 reg5591,
                 forvar5588,
                 reg5586,
                 reg5599,
                 reg5598,
                 reg5597,
                 reg5596,
                 reg5595,
                 reg5594,
                 reg5593,
                 reg5592,
                 forvar5591,
                 reg5590,
                 reg5589,
                 reg5588,
                 reg5587,
                 forvar5586,
                 reg5585,
                 reg5584,
                 forvar5583,
                 reg5581,
                 reg5579,
                 reg5582,
                 forvar5581,
                 reg5580,
                 forvar5579,
                 reg5578,
                 forvar5577,
                 reg5576,
                 reg5575,
                 reg5574,
                 reg5573,
                 forvar5572,
                 reg5571,
                 reg5570,
                 forvar5569,
                 reg5568,
                 reg5567,
                 forvar5564,
                 reg5557,
                 reg5561,
                 forvar5559,
                 reg5566,
                 reg5565,
                 reg5564,
                 reg5563,
                 reg5562,
                 forvar5561,
                 reg5560,
                 reg5559,
                 reg5558,
                 forvar5557,
                 reg5556,
                 forvar5555,
                 reg5554,
                 forvar5553,
                 reg5552,
                 reg5551,
                 forvar5550,
                 reg5549,
                 reg5548,
                 reg5547,
                 reg5546,
                 reg5545,
                 reg5544,
                 reg5543,
                 reg5542,
                 forvar5541,
                 forvar5540,
                 reg5539,
                 reg5538,
                 reg5537,
                 reg5536,
                 reg5535,
                 reg5534,
                 forvar5533,
                 reg5533,
                 forvar5532,
                 wire5531,
                 wire5530,
                 wire5529,
                 wire5528,
                 wire5527,
                 wire5526,
                 wire5524,
                 wire1020,
                 forvar961,
                 reg969,
                 forvar963,
                 reg962,
                 reg956,
                 forvar955,
                 reg954,
                 reg952,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 forvar1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1008,
                 reg1007,
                 reg1006,
                 forvar1005,
                 reg1004,
                 forvar1003,
                 forvar1002,
                 reg1001,
                 reg1000,
                 reg999,
                 forvar998,
                 forvar997,
                 forvar996,
                 reg995,
                 reg994,
                 reg993,
                 reg992,
                 forvar991,
                 reg990,
                 reg989,
                 reg988,
                 forvar987,
                 reg986,
                 reg985,
                 reg984,
                 forvar980,
                 reg983,
                 reg982,
                 reg981,
                 reg980,
                 reg975,
                 reg971,
                 reg979,
                 reg978,
                 reg977,
                 reg976,
                 forvar975,
                 reg974,
                 reg973,
                 reg972,
                 forvar971,
                 reg970,
                 forvar969,
                 reg968,
                 reg967,
                 reg966,
                 forvar965,
                 reg964,
                 reg963,
                 forvar962,
                 reg961,
                 forvar960,
                 reg960,
                 reg959,
                 reg958,
                 reg957,
                 forvar956,
                 reg955,
                 forvar954,
                 forvar953,
                 forvar952,
                 forvar900,
                 forvar931,
                 reg926,
                 reg925,
                 forvar924,
                 reg922,
                 reg920,
                 forvar919,
                 reg918,
                 reg917,
                 reg907,
                 reg906,
                 forvar902,
                 forvar892,
                 forvar885,
                 reg951,
                 reg942,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 forvar945,
                 reg944,
                 reg943,
                 forvar942,
                 reg941,
                 reg940,
                 reg939,
                 reg938,
                 reg937,
                 reg936,
                 reg935,
                 reg934,
                 reg933,
                 reg932,
                 reg931,
                 reg930,
                 reg929,
                 reg928,
                 forvar927,
                 forvar926,
                 forvar925,
                 reg924,
                 reg923,
                 forvar922,
                 reg921,
                 forvar920,
                 reg919,
                 forvar918,
                 forvar917,
                 reg916,
                 reg915,
                 reg914,
                 reg913,
                 reg912,
                 forvar911,
                 reg910,
                 reg909,
                 reg908,
                 forvar907,
                 forvar906,
                 reg901,
                 forvar899,
                 forvar897,
                 reg905,
                 reg904,
                 reg903,
                 reg902,
                 forvar901,
                 forvar895,
                 reg894,
                 forvar893,
                 reg889,
                 reg888,
                 forvar887,
                 reg886,
                 forvar884,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 forvar894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 forvar889,
                 forvar888,
                 reg887,
                 forvar886,
                 reg885,
                 reg884,
                 forvar883,
                 reg882,
                 forvar881,
                 reg880,
                 reg879,
                 reg878,
                 reg877,
                 reg876,
                 reg875,
                 reg874,
                 reg872,
                 forvar871,
                 forvar870,
                 reg867,
                 forvar866,
                 forvar865,
                 forvar862,
                 forvar858,
                 reg851,
                 reg863,
                 forvar861,
                 reg859,
                 reg873,
                 forvar872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 forvar867,
                 reg866,
                 reg865,
                 reg864,
                 forvar863,
                 reg862,
                 reg861,
                 reg860,
                 forvar859,
                 forvar853,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 reg853,
                 reg852,
                 forvar851,
                 forvar843,
                 forvar836,
                 forvar834,
                 forvar831,
                 reg832,
                 reg829,
                 reg828,
                 reg844,
                 forvar840,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 reg845,
                 forvar844,
                 reg843,
                 reg842,
                 reg841,
                 reg840,
                 reg839,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 reg834,
                 reg833,
                 forvar832,
                 reg831,
                 reg830,
                 forvar829,
                 forvar828,
                 reg827,
                 reg826,
                 reg825,
                 forvar824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 forvar819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 forvar814,
                 reg813,
                 reg812,
                 forvar811,
                 reg810,
                 reg809,
                 reg808,
                 reg807,
                 forvar806,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 reg801,
                 reg800,
                 reg799,
                 forvar798,
                 reg797,
                 reg796,
                 reg795,
                 reg794,
                 reg793,
                 reg792,
                 reg791,
                 forvar790,
                 reg789,
                 reg788,
                 forvar787,
                 reg786,
                 reg785,
                 forvar784,
                 forvar783,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 forvar778,
                 reg777,
                 reg776,
                 forvar775,
                 reg774,
                 forvar771,
                 reg773,
                 reg772,
                 reg771,
                 forvar770,
                 forvar746,
                 reg748,
                 forvar742,
                 reg741,
                 reg769,
                 forvar768,
                 reg767,
                 reg766,
                 reg765,
                 reg764,
                 forvar763,
                 reg761,
                 forvar759,
                 reg756,
                 reg763,
                 reg762,
                 forvar761,
                 reg760,
                 reg759,
                 reg758,
                 reg757,
                 forvar756,
                 reg755,
                 reg754,
                 reg753,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 forvar748,
                 reg747,
                 reg746,
                 forvar745,
                 reg745,
                 reg744,
                 reg743,
                 reg742,
                 forvar741,
                 reg740,
                 reg739,
                 reg738,
                 forvar737,
                 reg736,
                 reg735,
                 reg734,
                 forvar733,
                 forvar731,
                 reg732,
                 reg731,
                 forvar730,
                 reg729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 reg723,
                 forvar722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 forvar713,
                 reg712,
                 forvar711,
                 reg710,
                 reg709,
                 reg708,
                 forvar707,
                 reg704,
                 forvar702,
                 forvar700,
                 reg707,
                 reg706,
                 reg705,
                 forvar704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 forvar699,
                 forvar695,
                 forvar693,
                 forvar689,
                 forvar688,
                 reg698,
                 forvar697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 forvar687,
                 reg690,
                 reg689,
                 reg688,
                 reg687,
                 reg686,
                 reg685,
                 reg684,
                 reg683,
                 forvar682,
                 forvar681,
                 reg680,
                 forvar676,
                 reg674,
                 forvar671,
                 forvar650,
                 forvar648,
                 forvar644,
                 reg669,
                 reg664,
                 forvar661,
                 reg659,
                 forvar656,
                 reg655,
                 forvar652,
                 forvar649,
                 reg647,
                 reg668,
                 reg660,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 reg675,
                 forvar674,
                 reg673,
                 reg672,
                 reg671,
                 reg670,
                 forvar669,
                 forvar668,
                 reg667,
                 reg666,
                 reg665,
                 forvar664,
                 reg663,
                 reg662,
                 reg661,
                 forvar660,
                 forvar659,
                 reg658,
                 reg657,
                 reg656,
                 forvar655,
                 reg654,
                 reg653,
                 reg652,
                 reg651,
                 reg650,
                 reg649,
                 reg648,
                 forvar647,
                 reg646,
                 reg645,
                 reg644,
                 forvar643,
                 reg643,
                 reg642,
                 forvar641,
                 forvar640,
                 reg639,
                 forvar638,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 forvar633,
                 reg632,
                 forvar631,
                 forvar630,
                 forvar629,
                 reg628,
                 reg627,
                 forvar626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 forvar621,
                 forvar620,
                 reg619,
                 reg618,
                 reg617,
                 reg616,
                 forvar615,
                 reg614,
                 reg613,
                 reg612,
                 forvar608,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 forvar607,
                 forvar602,
                 reg601,
                 reg606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 forvar601,
                 forvar600,
                 reg599,
                 reg598,
                 reg597,
                 reg592,
                 reg591,
                 reg596,
                 forvar595,
                 reg594,
                 reg593,
                 forvar592,
                 forvar591,
                 reg590,
                 forvar589,
                 forvar588,
                 reg587,
                 reg586,
                 reg585,
                 forvar584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 forvar579,
                 reg578,
                 reg577,
                 forvar575,
                 forvar571,
                 reg573,
                 forvar570,
                 reg576,
                 reg575,
                 reg574,
                 forvar573,
                 reg567,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 forvar567,
                 reg566,
                 reg565,
                 forvar564,
                 reg563,
                 forvar562,
                 wire561,
                 wire560,
                 wire559,
                 (1'h0)};
  assign wire559 = (~^$signed(($signed(wire555) != $signed(wire556))));
  assign wire560 = (((wire559[(1'h0):(1'h0)] == $signed(wire559)) ?
                       (8'h9d) : ({wire557} ~^ ((8'h9c) != wire557))) ~^ (wire557 & (^$unsigned(wire559))));
  assign wire561 = wire555[(3'h5):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar562 = (1'h0); (forvar562 < (2'h3)); forvar562 = (forvar562 + (1'h1)))
        begin
          reg563 <= $signed(wire557[(1'h0):(1'h0)]);
          if ($unsigned(wire558[(3'h5):(3'h4)]))
            begin
              if ($signed((~&$signed((^wire558)))))
                begin
                  for (forvar564 = (1'h0); (forvar564 < (2'h3)); forvar564 = (forvar564 + (1'h1)))
                    begin
                      reg565 <= ($signed((^~wire558)) ^ forvar564[(1'h1):(1'h0)]);
                      reg566 <= (^~(($unsigned(wire557) > (wire559 - wire558)) ?
                          wire558[(3'h7):(3'h6)] : (8'ha7)));
                    end
                  for (forvar567 = (1'h0); (forvar567 < (2'h2)); forvar567 = (forvar567 + (1'h1)))
                    begin
                      reg568 <= (({(~^wire555)} >>> $unsigned({(8'ha5)})) ?
                          wire556[(2'h2):(1'h1)] : (({forvar562} ?
                                  (wire561 ^ forvar564) : wire558) ?
                              {$unsigned(wire558)} : {(wire557 ?
                                      forvar564 : wire559)}));
                      reg569 <= $unsigned(forvar567[(2'h2):(1'h1)]);
                      reg570 <= reg563[(3'h6):(1'h1)];
                      reg571 <= (({(wire560 && wire558)} ?
                          wire556 : {{(8'hb5)}}) ^~ (wire557[(1'h0):(1'h0)] ?
                          $unsigned({reg570}) : $signed((8'haf))));
                    end
                  reg572 <= (-$unsigned(reg570[(4'h9):(1'h0)]));
                end
              else
                begin
                  for (forvar564 = (1'h0); (forvar564 < (2'h2)); forvar564 = (forvar564 + (1'h1)))
                    begin
                      reg565 <= wire556;
                      reg566 <= (reg563 < {$signed((wire560 ^ wire555))});
                      reg567 <= ((reg566[(4'h9):(2'h2)] == $unsigned((reg570 != reg563))) ?
                          ((&wire555) ^ $unsigned((~(8'ha2)))) : ((wire561[(3'h7):(1'h1)] ?
                                  (reg570 || (8'ha7)) : (reg563 ?
                                      reg572 : (8'h9e))) ?
                              wire556 : {$signed(wire560)}));
                      reg568 <= (($unsigned(forvar564[(3'h4):(1'h0)]) ?
                              {(~&forvar562)} : $unsigned((reg565 ?
                                  wire561 : (8'h9f)))) ?
                          ((!(&reg570)) * ($unsigned(forvar564) << $signed(reg565))) : (reg569[(2'h2):(1'h1)] ?
                              (((8'ha3) < wire561) ?
                                  $signed(reg570) : (reg571 >>> wire555)) : $unsigned((forvar562 ^~ reg570))));
                    end
                end
              for (forvar573 = (1'h0); (forvar573 < (2'h2)); forvar573 = (forvar573 + (1'h1)))
                begin
                  if ($unsigned((!$unsigned((reg571 ^ wire559)))))
                    begin
                      reg574 <= reg569[(3'h5):(1'h0)];
                      reg575 <= forvar562[(3'h4):(3'h4)];
                      reg576 <= reg574;
                    end
                  else
                    begin
                      reg574 <= (^(^{$signed((8'h9d))}));
                      reg575 <= ($unsigned(((wire560 ?
                              (8'ha1) : wire558) << {wire555})) ?
                          $signed(wire558) : (((8'h9d) ?
                                  $unsigned((8'hab)) : ((8'haf) ?
                                      wire559 : reg575)) ?
                              forvar573[(4'hb):(4'h9)] : $unsigned($unsigned((8'had)))));
                      reg576 <= (((&reg576) ?
                              (!forvar564[(2'h2):(1'h0)]) : (^forvar567)) ?
                          ({$signed((8'hb3))} || forvar573[(2'h2):(2'h2)]) : $signed(wire556));
                    end
                end
            end
          else
            begin
              for (forvar564 = (1'h0); (forvar564 < (2'h3)); forvar564 = (forvar564 + (1'h1)))
                begin
                  if ({($unsigned($unsigned(wire561)) == ($unsigned(forvar567) ?
                          $unsigned((8'h9d)) : reg576))})
                    begin
                      reg565 <= reg565[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg565 <= $signed((8'h9e));
                      reg566 <= $unsigned((8'hab));
                      reg567 <= $unsigned(((8'ha3) ?
                          (+(forvar564 ? reg565 : reg571)) : (~|reg572)));
                      reg568 <= (-(((8'h9e) ?
                          $signed(reg569) : wire558[(4'hc):(1'h1)]) == {{reg570}}));
                    end
                end
              if ((~&($unsigned((reg576 <= reg574)) ^~ ({reg568} ?
                  reg567[(2'h2):(1'h1)] : reg566[(4'h9):(3'h6)]))))
                begin
                  reg569 <= {wire559[(3'h5):(1'h0)]};
                  for (forvar570 = (1'h0); (forvar570 < (2'h2)); forvar570 = (forvar570 + (1'h1)))
                    begin
                      reg571 <= $unsigned($signed(((^~wire561) ?
                          ((8'haa) ? reg566 : wire558) : forvar573)));
                      reg572 <= (~&{reg572[(3'h4):(2'h3)]});
                      reg573 <= wire561[(4'ha):(3'h6)];
                      reg574 <= (!(reg566 ?
                          $signed({reg568}) : $unsigned(reg565)));
                    end
                  reg575 <= (~&reg574[(3'h4):(1'h1)]);
                end
              else
                begin
                  if ($signed(forvar567[(2'h2):(2'h2)]))
                    begin
                      reg569 <= forvar573;
                      reg570 <= ((|(reg566 < (8'hb0))) <= $signed($unsigned(reg573)));
                    end
                  else
                    begin
                      reg569 <= ((-reg571[(3'h4):(2'h3)]) < ($unsigned((reg569 & reg563)) ?
                          (^~$signed(reg566)) : reg573[(2'h2):(1'h0)]));
                    end
                  for (forvar571 = (1'h0); (forvar571 < (1'h0)); forvar571 = (forvar571 + (1'h1)))
                    begin
                      reg572 <= $signed((&{$signed(forvar571)}));
                      reg573 <= ($unsigned($unsigned((+wire556))) << ((~|wire560) != {(forvar571 ?
                              reg563 : (8'ha7))}));
                      reg574 <= wire558;
                    end
                  for (forvar575 = (1'h0); (forvar575 < (2'h3)); forvar575 = (forvar575 + (1'h1)))
                    begin
                      reg576 <= wire559;
                      reg577 <= $unsigned(((~&reg567[(3'h4):(2'h3)]) ?
                          wire560 : $unsigned($unsigned((8'ha0)))));
                      reg578 <= (forvar570 ?
                          {((wire557 + forvar567) < (~&wire559))} : (|$signed((wire560 ?
                              wire557 : wire557))));
                    end
                end
              for (forvar579 = (1'h0); (forvar579 < (1'h1)); forvar579 = (forvar579 + (1'h1)))
                begin
                  if ((~|((~|forvar562[(4'h9):(3'h4)]) ?
                      $unsigned((reg568 == wire555)) : $signed((reg563 >= (8'h9d))))))
                    begin
                      reg580 <= reg569;
                      reg581 <= ($unsigned($signed((8'haa))) | (|(~^(~&reg573))));
                    end
                  else
                    begin
                      reg580 <= {({(wire561 >= (8'ha9))} ?
                              (-(forvar575 ?
                                  reg565 : reg568)) : $signed((forvar564 || (8'hb7))))};
                      reg581 <= (reg580[(2'h3):(1'h0)] ?
                          (~$signed(wire555)) : wire559[(2'h3):(1'h1)]);
                      reg582 <= ((((reg569 * reg563) < (wire560 ~^ reg576)) ?
                          (~^(reg580 << wire557)) : reg577) ~^ $unsigned(wire560[(3'h6):(1'h1)]));
                    end
                  reg583 <= ((8'hb6) < reg572);
                  for (forvar584 = (1'h0); (forvar584 < (2'h2)); forvar584 = (forvar584 + (1'h1)))
                    begin
                      reg585 <= forvar570[(3'h4):(1'h0)];
                      reg586 <= reg572[(2'h2):(1'h0)];
                      reg587 <= (^~{(~&(reg570 * (8'ha3)))});
                    end
                end
            end
        end
      for (forvar588 = (1'h0); (forvar588 < (2'h3)); forvar588 = (forvar588 + (1'h1)))
        begin
          for (forvar589 = (1'h0); (forvar589 < (1'h0)); forvar589 = (forvar589 + (1'h1)))
            begin
              reg590 <= reg566[(3'h6):(2'h3)];
            end
          if (((~^reg581) ?
              reg581 : $signed(($unsigned(forvar579) && (reg563 <<< reg573)))))
            begin
              for (forvar591 = (1'h0); (forvar591 < (1'h0)); forvar591 = (forvar591 + (1'h1)))
                begin
                  for (forvar592 = (1'h0); (forvar592 < (1'h1)); forvar592 = (forvar592 + (1'h1)))
                    begin
                      reg593 <= $unsigned(reg582);
                      reg594 <= {($signed($unsigned(wire558)) <= {(^reg567)})};
                    end
                  for (forvar595 = (1'h0); (forvar595 < (2'h2)); forvar595 = (forvar595 + (1'h1)))
                    begin
                      reg596 <= forvar584;
                    end
                end
            end
          else
            begin
              if (wire558)
                begin
                  if ({wire555})
                    begin
                      reg591 <= (($signed((8'hba)) - reg568) - forvar595);
                      reg592 <= $signed($signed(($unsigned(wire559) ^~ (forvar571 ?
                          reg567 : forvar579))));
                      reg593 <= $signed((^(+reg566[(4'he):(4'hd)])));
                      reg594 <= $unsigned($unsigned((^~reg586[(3'h5):(2'h3)])));
                    end
                  else
                    begin
                      reg591 <= reg580[(3'h7):(3'h4)];
                      reg592 <= forvar570;
                    end
                end
              else
                begin
                  for (forvar591 = (1'h0); (forvar591 < (2'h3)); forvar591 = (forvar591 + (1'h1)))
                    begin
                      reg592 <= (~|$signed((~|reg580)));
                      reg593 <= reg582;
                      reg594 <= (~|{((reg567 ^~ reg569) ?
                              $signed(forvar573) : (wire557 ?
                                  reg578 : wire557))});
                    end
                  for (forvar595 = (1'h0); (forvar595 < (2'h2)); forvar595 = (forvar595 + (1'h1)))
                    begin
                      reg596 <= reg567;
                      reg597 <= $signed({reg596[(1'h1):(1'h0)]});
                    end
                  reg598 <= ((~|(+$signed(reg576))) ^ (^~(8'hb5)));
                  reg599 <= $unsigned((forvar591 ?
                      forvar591 : $signed($signed(reg580))));
                end
            end
        end
      for (forvar600 = (1'h0); (forvar600 < (2'h2)); forvar600 = (forvar600 + (1'h1)))
        begin
          if (wire557[(1'h0):(1'h0)])
            begin
              if ((wire561[(3'h7):(2'h2)] <<< ($unsigned($unsigned(reg577)) ?
                  ({reg583} ? $unsigned(forvar588) : forvar592) : {(forvar584 ?
                          forvar571 : reg575)})))
                begin
                  for (forvar601 = (1'h0); (forvar601 < (1'h1)); forvar601 = (forvar601 + (1'h1)))
                    begin
                      reg602 <= reg599;
                      reg603 <= (($unsigned((-reg599)) ?
                              ((forvar575 | reg583) > (~|wire560)) : ($signed(reg602) != (&reg566))) ?
                          {(~(reg573 != forvar567))} : $signed(((reg582 ?
                              forvar592 : (8'ha6)) <<< reg567[(3'h4):(2'h2)])));
                      reg604 <= (wire555[(3'h5):(2'h3)] && (reg571[(4'h8):(3'h4)] ?
                          reg573 : forvar589[(3'h4):(3'h4)]));
                      reg605 <= $signed($signed((reg587[(4'ha):(3'h7)] ~^ forvar575)));
                    end
                  reg606 <= (wire558 || (^~reg587));
                end
              else
                begin
                  reg601 <= reg572[(2'h2):(2'h2)];
                  for (forvar602 = (1'h0); (forvar602 < (2'h3)); forvar602 = (forvar602 + (1'h1)))
                    begin
                      reg603 <= ((forvar584[(4'h8):(1'h1)] << (8'hb1)) ?
                          (~forvar579[(4'h8):(2'h2)]) : $unsigned($unsigned((reg585 ^ (8'hb3)))));
                    end
                end
              for (forvar607 = (1'h0); (forvar607 < (1'h0)); forvar607 = (forvar607 + (1'h1)))
                begin
                  if (((~&wire560[(1'h1):(1'h0)]) ?
                      $signed(forvar595[(2'h3):(1'h0)]) : (~($unsigned(reg585) ?
                          (&(8'haa)) : (forvar567 < forvar564)))))
                    begin
                      reg608 <= $signed((($signed(forvar571) ?
                          $signed(reg572) : (reg598 ^~ (8'hb3))) - wire557[(3'h5):(1'h1)]));
                      reg609 <= wire555[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg608 <= ((reg563[(3'h6):(2'h3)] >>> (&(forvar600 ?
                          forvar588 : reg603))) >>> {$signed(reg576[(2'h3):(2'h3)])});
                      reg609 <= (reg605[(4'h8):(4'h8)] == reg578[(1'h1):(1'h0)]);
                      reg610 <= (8'haa);
                      reg611 <= reg582;
                    end
                end
            end
          else
            begin
              for (forvar601 = (1'h0); (forvar601 < (1'h0)); forvar601 = (forvar601 + (1'h1)))
                begin
                  for (forvar602 = (1'h0); (forvar602 < (1'h0)); forvar602 = (forvar602 + (1'h1)))
                    begin
                      reg603 <= ($unsigned(reg601[(3'h5):(3'h5)]) ?
                          $signed($signed((reg593 ?
                              (8'ha2) : reg585))) : (|($signed((8'ha9)) | (reg578 ?
                              reg606 : forvar570))));
                      reg604 <= (+reg576[(3'h4):(3'h4)]);
                      reg605 <= $unsigned((reg603 ?
                          reg605[(3'h4):(1'h0)] : (((8'hb9) == reg610) << (reg581 << reg611))));
                      reg606 <= {{reg596}};
                    end
                end
              for (forvar607 = (1'h0); (forvar607 < (1'h1)); forvar607 = (forvar607 + (1'h1)))
                begin
                  for (forvar608 = (1'h0); (forvar608 < (2'h2)); forvar608 = (forvar608 + (1'h1)))
                    begin
                      reg609 <= {$signed(wire561[(4'he):(1'h0)])};
                      reg610 <= (reg592 ?
                          $unsigned(reg572) : $unsigned((&forvar600)));
                      reg611 <= (((forvar570[(1'h0):(1'h0)] + (8'h9e)) * forvar571[(3'h6):(3'h4)]) ?
                          (8'ha9) : {($unsigned(forvar600) ?
                                  (reg609 - reg586) : (forvar570 < forvar571))});
                    end
                  if ((reg575[(3'h4):(3'h4)] >>> (forvar589 ?
                      $signed($unsigned(forvar571)) : ((+forvar589) <= wire556))))
                    begin
                      reg612 <= $unsigned(reg603[(2'h2):(1'h1)]);
                      reg613 <= reg605;
                      reg614 <= forvar588[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg612 <= reg585;
                      reg613 <= reg591[(2'h3):(1'h1)];
                    end
                  for (forvar615 = (1'h0); (forvar615 < (2'h3)); forvar615 = (forvar615 + (1'h1)))
                    begin
                      reg616 <= $signed((forvar571[(3'h6):(2'h3)] < ({(8'ha6)} ?
                          forvar573[(4'h8):(2'h3)] : {reg574})));
                      reg617 <= {(^forvar608[(4'h8):(3'h4)])};
                      reg618 <= $unsigned($signed($signed(((8'ha2) ~^ reg613))));
                      reg619 <= (($signed($signed(forvar584)) != ((forvar575 >> reg585) ?
                              reg580 : (reg597 ? forvar615 : reg601))) ?
                          $signed($signed(reg618[(2'h2):(2'h2)])) : $signed($signed((reg582 ?
                              forvar564 : reg609))));
                    end
                end
            end
          for (forvar620 = (1'h0); (forvar620 < (1'h0)); forvar620 = (forvar620 + (1'h1)))
            begin
              for (forvar621 = (1'h0); (forvar621 < (2'h2)); forvar621 = (forvar621 + (1'h1)))
                begin
                  if ((8'ha1))
                    begin
                      reg622 <= (reg572 < reg601[(1'h1):(1'h1)]);
                      reg623 <= ($signed(reg573[(1'h0):(1'h0)]) | (+({reg596} ?
                          $signed(forvar607) : {(8'ha6)})));
                      reg624 <= ($signed(($unsigned(forvar564) * reg592)) || {$signed(((8'h9d) ?
                              reg565 : forvar584))});
                      reg625 <= reg592[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg622 <= wire556;
                    end
                  for (forvar626 = (1'h0); (forvar626 < (1'h1)); forvar626 = (forvar626 + (1'h1)))
                    begin
                      reg627 <= (^~$unsigned($unsigned((reg570 ?
                          reg617 : reg604))));
                      reg628 <= (($unsigned($unsigned(reg612)) ?
                              $signed(reg616) : ($unsigned((8'hb7)) & {reg604})) ?
                          $signed(reg592[(3'h4):(2'h3)]) : (((reg618 >>> wire561) >>> (reg587 ?
                              reg614 : reg567)) > $unsigned($unsigned(reg585))));
                    end
                end
            end
          for (forvar629 = (1'h0); (forvar629 < (1'h1)); forvar629 = (forvar629 + (1'h1)))
            begin
              for (forvar630 = (1'h0); (forvar630 < (2'h2)); forvar630 = (forvar630 + (1'h1)))
                begin
                  for (forvar631 = (1'h0); (forvar631 < (1'h1)); forvar631 = (forvar631 + (1'h1)))
                    begin
                      reg632 <= reg609[(3'h5):(2'h3)];
                    end
                  for (forvar633 = (1'h0); (forvar633 < (1'h1)); forvar633 = (forvar633 + (1'h1)))
                    begin
                      reg634 <= {($unsigned(forvar571[(4'hc):(2'h2)]) ?
                              forvar570 : {(~^reg586)})};
                      reg635 <= $signed($unsigned((wire556[(1'h0):(1'h0)] << {forvar600})));
                      reg636 <= reg598[(3'h4):(2'h2)];
                      reg637 <= {reg591};
                    end
                end
              for (forvar638 = (1'h0); (forvar638 < (2'h2)); forvar638 = (forvar638 + (1'h1)))
                begin
                  reg639 <= ($unsigned($signed($unsigned(reg576))) - $unsigned((^reg571[(3'h7):(3'h7)])));
                end
              for (forvar640 = (1'h0); (forvar640 < (2'h3)); forvar640 = (forvar640 + (1'h1)))
                begin
                  for (forvar641 = (1'h0); (forvar641 < (1'h0)); forvar641 = (forvar641 + (1'h1)))
                    begin
                      reg642 <= ($unsigned(reg606[(1'h1):(1'h1)]) << ($unsigned(((8'hba) ?
                          reg634 : wire559)) | (^~(reg567 ?
                          reg592 : (8'haa)))));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned({((&reg578) ? (^(8'ha1)) : $unsigned(forvar600))}))
        begin
          if ($signed(($signed(reg593) ?
              (!reg635[(3'h7):(2'h3)]) : forvar573[(4'h8):(3'h4)])))
            begin
              reg643 <= reg636;
            end
          else
            begin
              for (forvar643 = (1'h0); (forvar643 < (2'h2)); forvar643 = (forvar643 + (1'h1)))
                begin
                  if (((~&(~&{forvar615})) ^ {($unsigned(forvar579) ?
                          (~|forvar564) : (reg604 & forvar608))}))
                    begin
                      reg644 <= reg566[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg644 <= reg594[(3'h7):(1'h1)];
                      reg645 <= ((~$unsigned((forvar641 ?
                          forvar584 : reg616))) * $unsigned(forvar608));
                      reg646 <= ($signed($signed((wire559 ?
                              (8'hb5) : forvar640))) ?
                          reg623[(2'h3):(1'h0)] : (8'hb1));
                    end
                  for (forvar647 = (1'h0); (forvar647 < (2'h2)); forvar647 = (forvar647 + (1'h1)))
                    begin
                      reg648 <= {reg604};
                      reg649 <= $unsigned(reg625);
                      reg650 <= {(~&wire558)};
                      reg651 <= (8'h9e);
                    end
                  if (reg634)
                    begin
                      reg652 <= ((((reg599 ? reg593 : (8'haa)) ?
                                  (~&forvar584) : (~|reg582)) ?
                              (!reg611[(3'h4):(1'h0)]) : reg635[(2'h3):(1'h0)]) ?
                          (~^forvar564[(1'h0):(1'h0)]) : ({(forvar591 >> (8'ha3))} < ($signed(reg581) ?
                              (-reg563) : (reg639 <<< reg586))));
                    end
                  else
                    begin
                      reg652 <= ((|((~|reg577) | (forvar575 || forvar567))) == reg593[(1'h1):(1'h1)]);
                      reg653 <= reg590[(3'h4):(2'h3)];
                      reg654 <= ({((!reg596) ?
                                  (reg623 | reg605) : $signed(reg582))} ?
                          wire558[(4'hd):(3'h5)] : (8'hb4));
                    end
                  for (forvar655 = (1'h0); (forvar655 < (1'h0)); forvar655 = (forvar655 + (1'h1)))
                    begin
                      reg656 <= forvar562;
                      reg657 <= (+((reg645[(1'h0):(1'h0)] & (wire559 * (8'hb5))) & ((|wire560) > (reg587 ?
                          (8'hb9) : forvar621))));
                      reg658 <= {($signed((reg653 != (8'hb8))) > (((8'ha2) <= reg650) >>> reg649))};
                    end
                end
            end
          if ((($signed(reg585[(1'h1):(1'h0)]) || $unsigned($unsigned(reg628))) ?
              forvar615[(3'h6):(3'h5)] : (~|(reg573[(1'h1):(1'h1)] != (wire558 ?
                  forvar630 : (8'ha7))))))
            begin
              for (forvar659 = (1'h0); (forvar659 < (1'h0)); forvar659 = (forvar659 + (1'h1)))
                begin
                  for (forvar660 = (1'h0); (forvar660 < (2'h2)); forvar660 = (forvar660 + (1'h1)))
                    begin
                      reg661 <= (reg653[(1'h0):(1'h0)] >= ((~((8'h9c) && forvar584)) << (&forvar579)));
                      reg662 <= (((~|reg618) || forvar620) ?
                          reg648 : (~^{(reg627 ? (8'hb9) : (8'haa))}));
                      reg663 <= (8'hae);
                    end
                  for (forvar664 = (1'h0); (forvar664 < (2'h2)); forvar664 = (forvar664 + (1'h1)))
                    begin
                      reg665 <= reg653[(1'h0):(1'h0)];
                      reg666 <= {($signed(((8'hac) ?
                              forvar573 : reg628)) <<< {(reg613 ?
                                  reg661 : reg576)})};
                    end
                end
              reg667 <= $unsigned(forvar600);
              for (forvar668 = (1'h0); (forvar668 < (2'h2)); forvar668 = (forvar668 + (1'h1)))
                begin
                  for (forvar669 = (1'h0); (forvar669 < (2'h3)); forvar669 = (forvar669 + (1'h1)))
                    begin
                      reg670 <= reg642;
                      reg671 <= ((reg565[(1'h1):(1'h0)] << (wire557 * (~&(8'hb1)))) ?
                          ((forvar588 ?
                                  (reg657 ^ reg616) : reg657[(3'h4):(2'h2)]) ?
                              reg586 : (^{reg663})) : (~^((forvar621 ~^ (8'hae)) << (&reg606))));
                      reg672 <= $signed(reg637);
                      reg673 <= forvar601;
                    end
                  for (forvar674 = (1'h0); (forvar674 < (1'h1)); forvar674 = (forvar674 + (1'h1)))
                    begin
                      reg675 <= (!$signed({$signed(reg567)}));
                      reg676 <= {reg575};
                      reg677 <= ($unsigned({(^~reg565)}) ?
                          reg587 : wire559[(3'h7):(3'h6)]);
                    end
                end
              if ($signed(wire555))
                begin
                  reg678 <= reg598[(3'h4):(3'h4)];
                end
              else
                begin
                  reg678 <= reg653[(2'h3):(2'h2)];
                  if (forvar608[(1'h0):(1'h0)])
                    begin
                      reg679 <= (+$unsigned({forvar595}));
                    end
                  else
                    begin
                      reg679 <= ((forvar674 & $signed((reg673 || reg677))) ?
                          (($signed(reg605) ?
                                  (reg614 & reg597) : (forvar602 == reg623)) ?
                              $signed($unsigned(reg574)) : forvar655[(2'h2):(2'h2)]) : $unsigned((^$unsigned(reg635))));
                    end
                end
            end
          else
            begin
              for (forvar659 = (1'h0); (forvar659 < (2'h3)); forvar659 = (forvar659 + (1'h1)))
                begin
                  if (reg613)
                    begin
                      reg660 <= $signed((&$signed((reg565 & reg597))));
                    end
                  else
                    begin
                      reg660 <= $signed(reg654[(1'h0):(1'h0)]);
                      reg661 <= reg614[(1'h1):(1'h1)];
                      reg662 <= (|reg605);
                    end
                end
              reg663 <= (($unsigned(reg572[(1'h0):(1'h0)]) ?
                      $unsigned(reg672) : forvar659) ?
                  $signed(((+forvar591) ?
                      $unsigned(reg619) : reg586)) : (^~{{reg591}}));
              for (forvar664 = (1'h0); (forvar664 < (2'h3)); forvar664 = (forvar664 + (1'h1)))
                begin
                  if (reg678)
                    begin
                      reg665 <= forvar607;
                      reg666 <= forvar641;
                      reg667 <= $unsigned(reg578[(1'h1):(1'h0)]);
                      reg668 <= reg594[(3'h7):(3'h6)];
                    end
                  else
                    begin
                      reg665 <= (reg679 ? $signed($signed((^reg573))) : reg634);
                      reg666 <= (~&$signed($unsigned(reg628[(3'h6):(2'h3)])));
                    end
                end
            end
        end
      else
        begin
          if ({reg644[(1'h0):(1'h0)]})
            begin
              for (forvar643 = (1'h0); (forvar643 < (1'h1)); forvar643 = (forvar643 + (1'h1)))
                begin
                  if ((($signed($signed(reg651)) ?
                      ($unsigned(reg651) ?
                          (forvar660 ?
                              forvar647 : reg602) : reg662[(2'h2):(1'h1)]) : reg663) <= forvar591))
                    begin
                      reg644 <= (($signed((-reg616)) || ((reg617 & reg627) ?
                          (reg671 ^~ reg617) : (reg627 || forvar631))) && ($unsigned((&forvar631)) || $unsigned($unsigned(reg645))));
                      reg645 <= (forvar630[(3'h7):(3'h5)] <<< reg625);
                    end
                  else
                    begin
                      reg644 <= (forvar570 ?
                          {reg585[(4'hc):(4'hb)]} : ((((8'ha7) ?
                                  forvar638 : (8'haa)) ~^ (reg566 != (8'h9f))) ?
                              wire560 : reg653));
                      reg645 <= (+{$signed({reg643})});
                    end
                  if ((&(!(~&(forvar660 ? reg602 : reg667)))))
                    begin
                      reg646 <= reg658[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg646 <= $unsigned(reg583);
                      reg647 <= (~&$unsigned((&reg592[(1'h1):(1'h1)])));
                      reg648 <= (~&({reg671[(4'hd):(3'h4)]} ?
                          $signed(reg660) : (wire557[(2'h3):(1'h1)] ?
                              (~&(8'h9c)) : {reg627})));
                    end
                  for (forvar649 = (1'h0); (forvar649 < (1'h1)); forvar649 = (forvar649 + (1'h1)))
                    begin
                      reg650 <= ($signed(forvar584) | ({(reg609 ?
                                  forvar643 : (8'hb9))} ?
                          $unsigned((reg642 ?
                              forvar570 : forvar592)) : {(reg606 > forvar564)}));
                      reg651 <= reg652;
                    end
                end
              if ($unsigned($signed(reg608[(1'h0):(1'h0)])))
                begin
                  for (forvar652 = (1'h0); (forvar652 < (2'h3)); forvar652 = (forvar652 + (1'h1)))
                    begin
                      reg653 <= ($signed(reg606[(4'h9):(4'h9)]) == ((^~$unsigned(forvar595)) + ((~&reg569) ^~ reg677[(1'h0):(1'h0)])));
                    end
                  if ($unsigned((reg634[(2'h3):(1'h0)] ?
                      reg591[(3'h5):(1'h1)] : $signed(reg599))))
                    begin
                      reg654 <= (reg643[(3'h6):(1'h0)] ^ reg660);
                      reg655 <= (|(!$unsigned($unsigned(forvar570))));
                      reg656 <= (8'ha5);
                      reg657 <= (($signed((reg637 != wire555)) & (reg602[(1'h0):(1'h0)] ^~ (reg585 != reg678))) ?
                          forvar567[(2'h2):(1'h1)] : ($signed(reg576) ?
                              (((8'h9c) & reg666) >= (forvar600 ?
                                  forvar600 : forvar607)) : (|$unsigned(reg650))));
                    end
                  else
                    begin
                      reg654 <= $unsigned(($signed($unsigned(reg671)) ?
                          ({reg665} < $unsigned(forvar571)) : reg657[(2'h3):(2'h3)]));
                      reg655 <= $unsigned(reg617);
                      reg656 <= (!reg647);
                      reg657 <= reg563[(3'h4):(2'h3)];
                    end
                end
              else
                begin
                  if (((|$signed((8'hb0))) ? {(~&(-reg602))} : reg665))
                    begin
                      reg652 <= (~&(~&forvar664));
                      reg653 <= reg663;
                      reg654 <= (^~reg653[(3'h6):(3'h5)]);
                      reg655 <= $signed(($signed(reg570[(3'h6):(3'h4)]) == ($signed((8'h9c)) <= $unsigned((8'hb1)))));
                    end
                  else
                    begin
                      reg652 <= $unsigned((^{(forvar640 <<< reg627)}));
                      reg653 <= $unsigned(forvar664);
                    end
                  for (forvar656 = (1'h0); (forvar656 < (2'h2)); forvar656 = (forvar656 + (1'h1)))
                    begin
                      reg657 <= wire558;
                      reg658 <= forvar674[(2'h3):(2'h3)];
                      reg659 <= (|({(reg655 ~^ reg585)} ?
                          {reg604[(2'h2):(2'h2)]} : reg643));
                      reg660 <= (~^($signed($signed(reg606)) ?
                          forvar607[(3'h5):(1'h0)] : reg642));
                    end
                  for (forvar661 = (1'h0); (forvar661 < (2'h2)); forvar661 = (forvar661 + (1'h1)))
                    begin
                      reg662 <= ((wire556 ?
                              $signed(reg679[(4'h8):(3'h5)]) : reg573) ?
                          {$unsigned(forvar669)} : ((~|(~|forvar655)) ?
                              $signed($unsigned(forvar607)) : $signed($unsigned(reg659))));
                      reg663 <= $signed($unsigned($signed($unsigned(reg678))));
                      reg664 <= ($signed(reg572[(1'h1):(1'h1)]) >> $signed(($unsigned(forvar564) >>> reg672)));
                      reg665 <= $signed({$signed(reg612)});
                    end
                  if (((~^$signed(((8'ha1) - reg659))) & (^~reg643)))
                    begin
                      reg666 <= (-reg578);
                      reg667 <= {$unsigned((^~{reg671}))};
                    end
                  else
                    begin
                      reg666 <= reg624;
                      reg667 <= forvar601;
                      reg668 <= reg598;
                      reg669 <= (-(!$signed((reg671 >>> reg663))));
                    end
                end
              reg670 <= reg604;
            end
          else
            begin
              for (forvar643 = (1'h0); (forvar643 < (2'h2)); forvar643 = (forvar643 + (1'h1)))
                begin
                  for (forvar644 = (1'h0); (forvar644 < (1'h0)); forvar644 = (forvar644 + (1'h1)))
                    begin
                      reg645 <= ($unsigned($signed(forvar584)) ?
                          {forvar647[(4'he):(3'h6)]} : {(((8'had) << reg649) ?
                                  (reg663 ?
                                      (8'hba) : reg654) : reg676[(1'h0):(1'h0)])});
                      reg646 <= reg666[(3'h7):(3'h7)];
                      reg647 <= forvar661[(1'h0):(1'h0)];
                    end
                end
              if ($unsigned((-reg567[(2'h2):(1'h1)])))
                begin
                  for (forvar648 = (1'h0); (forvar648 < (1'h1)); forvar648 = (forvar648 + (1'h1)))
                    begin
                      reg649 <= ((~|reg596) < {((8'hb4) ?
                              forvar629[(3'h4):(3'h4)] : {(8'hb6)})});
                    end
                  for (forvar650 = (1'h0); (forvar650 < (1'h0)); forvar650 = (forvar650 + (1'h1)))
                    begin
                      reg651 <= reg657[(2'h2):(1'h0)];
                      reg652 <= reg668[(3'h5):(3'h4)];
                      reg653 <= ((8'ha7) ?
                          reg571 : $unsigned(({reg632} ?
                              (forvar588 ?
                                  reg671 : (8'ha9)) : $signed(forvar571))));
                      reg654 <= reg646[(3'h7):(2'h2)];
                    end
                  for (forvar655 = (1'h0); (forvar655 < (1'h1)); forvar655 = (forvar655 + (1'h1)))
                    begin
                      reg656 <= $signed((reg658 ?
                          $unsigned((~&reg608)) : (!$unsigned(reg676))));
                      reg657 <= $unsigned(forvar648);
                      reg658 <= reg676[(3'h7):(1'h0)];
                      reg659 <= (((|(wire557 <<< reg665)) <= ((reg670 ?
                              forvar629 : reg652) <= $signed((8'hb4)))) ?
                          reg639[(4'ha):(3'h5)] : reg665[(4'hd):(4'ha)]);
                    end
                  if (reg605)
                    begin
                      reg660 <= (^~((forvar567 ?
                          $signed(forvar626) : (reg567 ?
                              reg661 : (8'ha3))) + forvar615[(3'h4):(2'h3)]));
                      reg661 <= {$signed($unsigned($unsigned((8'hb7))))};
                      reg662 <= reg659;
                    end
                  else
                    begin
                      reg660 <= ($unsigned(((reg585 + forvar629) != (&forvar641))) ?
                          reg670[(3'h5):(3'h5)] : $signed(forvar652));
                      reg661 <= $signed((($unsigned(wire558) == (forvar661 ?
                          forvar664 : reg622)) && $signed($signed(forvar641))));
                      reg662 <= $unsigned($unsigned(reg656[(4'ha):(3'h6)]));
                      reg663 <= ($unsigned($unsigned((reg592 ~^ (8'h9d)))) ?
                          (reg671[(2'h3):(1'h0)] ?
                              $signed($signed(reg669)) : {{forvar661}}) : $signed(($unsigned(reg569) || (|reg585))));
                    end
                end
              else
                begin
                  reg648 <= $unsigned(forvar592);
                end
              if (reg567)
                begin
                  if ($signed(forvar631[(4'ha):(4'h9)]))
                    begin
                      reg664 <= {($signed((^~(8'h9e))) ?
                              $unsigned($unsigned(reg661)) : reg610[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg664 <= (^~(forvar579 | $unsigned((reg625 * reg571))));
                      reg665 <= $signed($unsigned((-$unsigned(forvar608))));
                    end
                  reg666 <= forvar641[(2'h2):(2'h2)];
                end
              else
                begin
                  if ($signed(($unsigned($unsigned(reg628)) || {{wire557}})))
                    begin
                      reg664 <= reg578[(3'h6):(3'h6)];
                      reg665 <= (wire558 * {$unsigned((~|reg666))});
                      reg666 <= (($unsigned(forvar620[(1'h0):(1'h0)]) ?
                          $unsigned(reg652) : $unsigned((reg613 ?
                              forvar584 : forvar630))) && (^(forvar650 ?
                          reg592[(2'h2):(1'h0)] : {reg656})));
                      reg667 <= (-$unsigned(($unsigned((8'h9d)) && $unsigned(forvar640))));
                    end
                  else
                    begin
                      reg664 <= (8'hb4);
                    end
                  for (forvar668 = (1'h0); (forvar668 < (2'h2)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg669 <= reg610;
                      reg670 <= (reg567[(2'h2):(1'h0)] ?
                          (((reg643 ?
                                  forvar668 : (8'hab)) != $unsigned(reg661)) ?
                              $unsigned((!reg570)) : wire561[(4'hb):(3'h4)]) : $signed((^(~|(8'hb5)))));
                    end
                  for (forvar671 = (1'h0); (forvar671 < (2'h2)); forvar671 = (forvar671 + (1'h1)))
                    begin
                      reg672 <= reg636[(2'h2):(1'h0)];
                      reg673 <= reg670;
                      reg674 <= (({$signed((8'hb6))} >= (|reg645[(3'h7):(2'h2)])) && {((forvar671 ?
                              reg675 : forvar626) ^ reg625)});
                      reg675 <= {$signed(reg601)};
                    end
                  for (forvar676 = (1'h0); (forvar676 < (1'h0)); forvar676 = (forvar676 + (1'h1)))
                    begin
                      reg677 <= {reg614[(2'h3):(2'h2)]};
                      reg678 <= $signed(reg614);
                      reg679 <= $signed(reg603[(2'h2):(1'h1)]);
                      reg680 <= (~(!($signed(reg590) ?
                          $signed(forvar649) : (reg667 ?
                              (8'had) : forvar562))));
                    end
                end
              for (forvar681 = (1'h0); (forvar681 < (2'h3)); forvar681 = (forvar681 + (1'h1)))
                begin
                  for (forvar682 = (1'h0); (forvar682 < (1'h0)); forvar682 = (forvar682 + (1'h1)))
                    begin
                      reg683 <= {$unsigned({reg667[(3'h4):(1'h0)]})};
                      reg684 <= (reg665 <= (forvar573[(2'h2):(1'h1)] ?
                          reg596[(4'ha):(3'h7)] : (~&(forvar629 ?
                              (8'ha6) : forvar671))));
                    end
                end
            end
          reg685 <= $signed(forvar602);
          reg686 <= ({((reg568 ? forvar567 : reg571) ?
                  (8'ha7) : {reg650})} <= reg669);
          if ($signed(forvar591))
            begin
              if (forvar656[(4'hc):(4'ha)])
                begin
                  if ((8'ha9))
                    begin
                      reg687 <= (forvar638 != reg658[(3'h7):(1'h0)]);
                      reg688 <= reg659[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg687 <= (forvar630 ?
                          (($unsigned(reg573) ?
                              (&wire556) : (^reg635)) - $unsigned($unsigned(reg599))) : reg665);
                      reg688 <= (reg590[(2'h3):(2'h2)] ^ forvar641);
                    end
                  if (((reg687[(1'h0):(1'h0)] ?
                      ((~&reg590) ~^ reg660[(2'h3):(1'h1)]) : $signed($signed(reg582))) * {((forvar570 ?
                          reg583 : reg656) == reg571[(4'hf):(4'h9)])}))
                    begin
                      reg689 <= (8'ha4);
                      reg690 <= $signed(reg657);
                    end
                  else
                    begin
                      reg689 <= reg598[(4'h8):(4'h8)];
                      reg690 <= $signed({$unsigned((reg645 ?
                              reg565 : (8'hb4)))});
                    end
                end
              else
                begin
                  for (forvar687 = (1'h0); (forvar687 < (1'h0)); forvar687 = (forvar687 + (1'h1)))
                    begin
                      reg688 <= $signed(reg617[(1'h0):(1'h0)]);
                      reg689 <= $unsigned(reg643[(4'ha):(2'h2)]);
                      reg690 <= reg602[(3'h7):(3'h6)];
                      reg691 <= ({(~$signed(reg674))} <<< forvar630);
                    end
                  reg692 <= (^~($signed(forvar671[(4'h8):(3'h6)]) - (-forvar633)));
                  reg693 <= ($unsigned(reg612[(3'h7):(3'h4)]) && (~|reg680[(4'ha):(3'h6)]));
                end
              if ($unsigned(reg592))
                begin
                  if (reg625[(1'h1):(1'h1)])
                    begin
                      reg694 <= (~(!$signed($unsigned(reg582))));
                      reg695 <= (((forvar649[(1'h0):(1'h0)] | $unsigned((8'haa))) ^ reg616[(3'h4):(2'h2)]) << (~|$unsigned((reg577 ?
                          (8'ha9) : reg661))));
                    end
                  else
                    begin
                      reg694 <= ($unsigned($signed((~&forvar668))) < (((8'h9e) ?
                          (reg605 ?
                              reg694 : reg692) : $unsigned(reg570)) == forvar589[(1'h0):(1'h0)]));
                      reg695 <= $signed((((reg646 ?
                          reg603 : reg647) && {reg568}) != reg580[(4'ha):(3'h6)]));
                    end
                end
              else
                begin
                  if (($signed($unsigned(reg597[(1'h1):(1'h0)])) ?
                      (+{(reg680 ?
                              forvar656 : forvar650)}) : reg670[(2'h2):(1'h1)]))
                    begin
                      reg694 <= ($signed($signed((reg650 << forvar641))) ?
                          $signed((forvar638[(2'h2):(2'h2)] >> (forvar649 || wire561))) : (-(forvar615[(1'h0):(1'h0)] * {forvar592})));
                      reg695 <= ((-reg570) << reg676);
                      reg696 <= (~(({(8'hb4)} ?
                          $signed(forvar607) : ((8'hb1) ?
                              reg667 : reg668)) * $unsigned((forvar575 ?
                          reg645 : forvar575))));
                    end
                  else
                    begin
                      reg694 <= reg616;
                    end
                  for (forvar697 = (1'h0); (forvar697 < (2'h3)); forvar697 = (forvar697 + (1'h1)))
                    begin
                      reg698 <= $unsigned((~(reg662[(3'h7):(1'h0)] != $signed(forvar595))));
                    end
                end
            end
          else
            begin
              reg687 <= {(8'ha4)};
              for (forvar688 = (1'h0); (forvar688 < (2'h2)); forvar688 = (forvar688 + (1'h1)))
                begin
                  for (forvar689 = (1'h0); (forvar689 < (1'h1)); forvar689 = (forvar689 + (1'h1)))
                    begin
                      reg690 <= ((-(~^(wire561 ? forvar676 : reg612))) ?
                          $signed($signed($unsigned((8'hb6)))) : $signed(((forvar588 == reg618) ?
                              reg582[(1'h1):(1'h1)] : $signed(reg650))));
                      reg691 <= forvar671;
                      reg692 <= forvar626;
                    end
                  for (forvar693 = (1'h0); (forvar693 < (2'h3)); forvar693 = (forvar693 + (1'h1)))
                    begin
                      reg694 <= ($unsigned(reg580[(2'h2):(2'h2)]) ?
                          ((reg597 < $signed((8'ha4))) <= reg648) : (reg602 ^~ (8'hab)));
                    end
                  for (forvar695 = (1'h0); (forvar695 < (2'h2)); forvar695 = (forvar695 + (1'h1)))
                    begin
                      reg696 <= ((~reg693) ?
                          $unsigned(((reg575 | reg659) - (reg592 ?
                              (8'hba) : reg690))) : ((-(&forvar601)) ?
                              (((8'hb7) || forvar643) ?
                                  (~&forvar676) : $unsigned(reg666)) : forvar573[(2'h3):(1'h1)]));
                    end
                end
            end
        end
      for (forvar699 = (1'h0); (forvar699 < (1'h0)); forvar699 = (forvar699 + (1'h1)))
        begin
          if ($unsigned(($signed(reg606[(4'h8):(1'h0)]) ?
              forvar575[(4'h8):(3'h4)] : $unsigned(reg652[(3'h4):(2'h3)]))))
            begin
              if ($unsigned((^~(|reg611))))
                begin
                  if ({(~&((reg611 << reg578) ?
                          (reg667 ? reg604 : forvar562) : (reg571 || reg614)))})
                    begin
                      reg700 <= {((((8'hb5) & reg692) ?
                              (reg645 ? forvar693 : reg685) : (forvar697 ?
                                  reg571 : reg563)) != $unsigned({reg611}))};
                      reg701 <= (^~reg672);
                      reg702 <= reg675[(3'h7):(3'h5)];
                      reg703 <= ($signed((^forvar682)) ?
                          $signed(forvar660) : reg693);
                    end
                  else
                    begin
                      reg700 <= (&($unsigned($signed(reg667)) ?
                          forvar669 : $unsigned((^~reg687))));
                      reg701 <= $unsigned(((|(8'hab)) <= ((~&reg700) ?
                          $unsigned(reg664) : reg587)));
                      reg702 <= {($signed((8'hb3)) ?
                              $unsigned((reg590 ?
                                  reg660 : wire556)) : reg689[(4'h9):(2'h2)])};
                      reg703 <= (-reg703[(4'ha):(3'h7)]);
                    end
                end
              else
                begin
                  if ($signed($unsigned(forvar674)))
                    begin
                      reg700 <= forvar649[(1'h0):(1'h0)];
                      reg701 <= $signed(reg694[(3'h6):(1'h1)]);
                      reg702 <= (~{forvar695});
                      reg703 <= {$signed(($signed(reg594) ?
                              forvar664[(2'h2):(1'h1)] : $unsigned(reg637)))};
                    end
                  else
                    begin
                      reg700 <= (($unsigned((reg690 ? reg605 : reg685)) ?
                              (~|(reg627 ?
                                  reg673 : wire560)) : $signed((reg632 ?
                                  reg698 : forvar671))) ?
                          {((forvar633 ? reg577 : (8'ha5)) ?
                                  {reg669} : reg671[(2'h3):(1'h0)])} : (~|{(8'hba)}));
                      reg701 <= $signed($signed(reg667));
                    end
                  for (forvar704 = (1'h0); (forvar704 < (2'h3)); forvar704 = (forvar704 + (1'h1)))
                    begin
                      reg705 <= reg634[(4'h8):(4'h8)];
                      reg706 <= ({((~(8'h9d)) <<< (reg571 << reg654))} ?
                          (+((8'hac) ?
                              (reg606 == reg596) : $unsigned(forvar704))) : reg613[(4'h8):(1'h0)]);
                      reg707 <= ($unsigned($signed((forvar629 ?
                          reg674 : reg601))) >>> {{forvar591[(3'h6):(1'h1)]}});
                    end
                end
            end
          else
            begin
              if ({(~($signed(reg667) ? reg692 : (8'ha3)))})
                begin
                  for (forvar700 = (1'h0); (forvar700 < (1'h0)); forvar700 = (forvar700 + (1'h1)))
                    begin
                      reg701 <= ((^~((reg669 ^~ reg634) >> $unsigned(reg671))) < (!{(reg625 - forvar631)}));
                    end
                  for (forvar702 = (1'h0); (forvar702 < (2'h2)); forvar702 = (forvar702 + (1'h1)))
                    begin
                      reg703 <= (~(|($signed(reg698) ?
                          $signed(forvar591) : (reg678 || reg583))));
                      reg704 <= $unsigned(forvar595);
                      reg705 <= $unsigned((reg690[(3'h7):(3'h7)] << $unsigned(reg691[(3'h4):(2'h3)])));
                    end
                  reg706 <= (^(!reg623[(3'h5):(3'h4)]));
                  for (forvar707 = (1'h0); (forvar707 < (2'h3)); forvar707 = (forvar707 + (1'h1)))
                    begin
                      reg708 <= forvar629;
                      reg709 <= $signed((reg596[(4'h9):(3'h7)] ?
                          $unsigned($signed((8'hac))) : $unsigned((^(8'ha2)))));
                      reg710 <= forvar638;
                    end
                end
              else
                begin
                  if ((-$signed({forvar588})))
                    begin
                      reg700 <= reg566;
                    end
                  else
                    begin
                      reg700 <= (^~(reg647 <= (~&(!reg689))));
                      reg701 <= (($signed((reg611 ? reg700 : reg661)) ?
                          ((reg645 ? (8'hba) : reg664) ?
                              $signed(forvar687) : ((8'hb6) ?
                                  reg672 : reg573)) : {(^reg587)}) ^ forvar660[(2'h3):(2'h3)]);
                      reg702 <= reg642;
                      reg703 <= (forvar592[(3'h4):(3'h4)] > reg565[(3'h7):(2'h2)]);
                    end
                  for (forvar704 = (1'h0); (forvar704 < (1'h1)); forvar704 = (forvar704 + (1'h1)))
                    begin
                      reg705 <= $signed($unsigned(((-forvar650) + (~^forvar608))));
                      reg706 <= ((|(reg656 + $unsigned((8'hab)))) ?
                          wire555 : ((reg670[(2'h2):(1'h1)] >= (8'had)) ?
                              $signed(forvar644[(4'h8):(3'h5)]) : reg690[(1'h1):(1'h1)]));
                      reg707 <= $signed($signed(wire555));
                    end
                  if ((~^$signed($signed(reg576[(1'h0):(1'h0)]))))
                    begin
                      reg708 <= $unsigned(forvar664);
                      reg709 <= ($signed((-reg651)) ?
                          $signed($unsigned(reg646)) : {((8'ha4) ?
                                  (~reg674) : forvar588)});
                      reg710 <= {(((~&reg582) ?
                                  $signed(forvar626) : $signed(reg575)) ?
                              $signed(((8'hba) ?
                                  reg571 : reg569)) : $signed((forvar589 ?
                                  forvar564 : reg686)))};
                    end
                  else
                    begin
                      reg708 <= ((~&reg657[(2'h3):(1'h1)]) ?
                          $unsigned($unsigned($unsigned((8'hb2)))) : reg594);
                      reg709 <= (({reg628} ?
                              reg677[(1'h0):(1'h0)] : (forvar607[(3'h4):(2'h2)] & forvar682[(3'h5):(1'h1)])) ?
                          ((+$signed(reg662)) ?
                              (^~(reg632 << reg705)) : $unsigned(reg693)) : (&(|reg683[(3'h4):(1'h0)])));
                      reg710 <= $signed(forvar579);
                    end
                  for (forvar711 = (1'h0); (forvar711 < (2'h2)); forvar711 = (forvar711 + (1'h1)))
                    begin
                      reg712 <= forvar573[(4'hd):(4'hb)];
                    end
                end
              for (forvar713 = (1'h0); (forvar713 < (2'h3)); forvar713 = (forvar713 + (1'h1)))
                begin
                  if ((({(!reg591)} ?
                          forvar655[(3'h4):(3'h4)] : (forvar711 ?
                              {forvar643} : (+forvar615))) ?
                      reg701[(4'ha):(3'h6)] : $unsigned((8'ha8))))
                    begin
                      reg714 <= $signed({forvar575[(3'h7):(1'h1)]});
                      reg715 <= reg582;
                      reg716 <= $signed((forvar584[(4'h8):(3'h4)] ^~ (reg674[(2'h3):(1'h0)] ?
                          $unsigned(forvar693) : (forvar700 == (8'hb0)))));
                    end
                  else
                    begin
                      reg714 <= ($unsigned((8'h9f)) > $signed({wire558}));
                      reg715 <= forvar695[(1'h0):(1'h0)];
                      reg716 <= $unsigned(forvar688);
                    end
                  if ($unsigned($signed(reg597)))
                    begin
                      reg717 <= (reg603[(1'h1):(1'h0)] ?
                          {forvar669[(2'h3):(2'h2)]} : forvar713[(1'h1):(1'h0)]);
                      reg718 <= reg673;
                    end
                  else
                    begin
                      reg717 <= forvar588;
                    end
                  if (forvar688)
                    begin
                      reg719 <= {($signed((reg576 ? reg654 : forvar567)) ?
                              reg712[(4'hf):(2'h3)] : ((!reg672) ?
                                  $unsigned(reg669) : reg597[(3'h4):(3'h4)]))};
                      reg720 <= (!($unsigned((~^reg676)) != $unsigned({reg714})));
                      reg721 <= ((~$signed((reg580 ?
                          reg583 : reg672))) || (forvar682 ?
                          (forvar589[(3'h4):(1'h1)] ~^ {reg696}) : ((reg680 ?
                              forvar674 : forvar643) && {(8'hab)})));
                    end
                  else
                    begin
                      reg719 <= reg627;
                      reg720 <= (reg617 ?
                          $unsigned(((reg662 ?
                              forvar600 : reg705) != ((8'hb8) >>> reg672))) : forvar567);
                      reg721 <= (^(-$signed(((8'hab) && reg656))));
                    end
                end
              for (forvar722 = (1'h0); (forvar722 < (2'h3)); forvar722 = (forvar722 + (1'h1)))
                begin
                  if ($signed((reg683[(4'h8):(2'h3)] ?
                      $signed($signed(forvar707)) : forvar664[(1'h1):(1'h0)])))
                    begin
                      reg723 <= (forvar695 | $unsigned($signed($signed(reg606))));
                    end
                  else
                    begin
                      reg723 <= $signed($unsigned((^$signed(forvar629))));
                      reg724 <= {(((forvar713 ?
                              (8'hb8) : reg649) && reg567) - (&forvar722[(2'h3):(2'h2)]))};
                      reg725 <= (|$signed($unsigned($unsigned(reg612))));
                      reg726 <= reg576[(3'h7):(3'h6)];
                    end
                  reg727 <= $signed(((&$signed(reg602)) ?
                      ((~|reg725) ^ reg632[(4'hf):(4'ha)]) : ((reg666 ^ reg602) ^~ (~^(8'h9f)))));
                  reg728 <= forvar707[(3'h4):(2'h3)];
                  reg729 <= $unsigned($signed((8'ha4)));
                end
            end
        end
      for (forvar730 = (1'h0); (forvar730 < (2'h3)); forvar730 = (forvar730 + (1'h1)))
        begin
          if ($signed({reg576}))
            begin
              reg731 <= (reg625 ~^ forvar630);
              reg732 <= ({(reg725[(1'h0):(1'h0)] ^~ forvar630[(3'h5):(1'h0)])} ?
                  $unsigned(((-reg672) && reg653)) : reg678[(3'h5):(3'h4)]);
            end
          else
            begin
              for (forvar731 = (1'h0); (forvar731 < (1'h1)); forvar731 = (forvar731 + (1'h1)))
                begin
                  reg732 <= (8'ha9);
                  for (forvar733 = (1'h0); (forvar733 < (2'h2)); forvar733 = (forvar733 + (1'h1)))
                    begin
                      reg734 <= reg574[(3'h4):(2'h3)];
                      reg735 <= ((reg639[(4'hb):(4'ha)] ?
                              reg646 : $signed(((8'h9d) ?
                                  forvar697 : wire560))) ?
                          (reg670 ?
                              $unsigned({reg671}) : (8'hb0)) : ({((8'hb9) != forvar629)} | reg676));
                      reg736 <= (forvar669[(2'h2):(2'h2)] == ($unsigned((forvar602 ?
                          reg569 : (8'ha5))) < ((&wire555) >> (reg734 ?
                          reg673 : reg691))));
                    end
                end
              for (forvar737 = (1'h0); (forvar737 < (2'h2)); forvar737 = (forvar737 + (1'h1)))
                begin
                  reg738 <= ($signed(reg694) ? (^~$signed(reg670)) : reg571);
                end
              reg739 <= (reg568 == $signed(((~|reg578) ?
                  $unsigned(reg706) : $signed(forvar704))));
              reg740 <= ($unsigned(($unsigned(wire558) == ((8'had) ?
                      forvar730 : forvar674))) ?
                  (forvar699 > (|((8'had) ? reg627 : reg637))) : (8'hb5));
            end
          if ($signed(((reg643 ? forvar647 : forvar676) ?
              $unsigned({(8'hb8)}) : (reg717[(3'h5):(1'h0)] || $signed(forvar584)))))
            begin
              if ({{{reg705}}})
                begin
                  for (forvar741 = (1'h0); (forvar741 < (2'h2)); forvar741 = (forvar741 + (1'h1)))
                    begin
                      reg742 <= $unsigned((|($signed((8'hb7)) ^ (&forvar730))));
                      reg743 <= (~&forvar562);
                      reg744 <= $signed(forvar722[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar741 = (1'h0); (forvar741 < (2'h2)); forvar741 = (forvar741 + (1'h1)))
                    begin
                      reg742 <= (((|(reg606 != reg663)) >= ($signed(forvar697) == reg657)) ?
                          reg642 : {forvar570});
                    end
                end
              if (reg565)
                begin
                  reg745 <= $unsigned(((forvar588 ^ reg574[(1'h1):(1'h0)]) & ($unsigned(reg637) * $signed(reg603))));
                end
              else
                begin
                  for (forvar745 = (1'h0); (forvar745 < (2'h3)); forvar745 = (forvar745 + (1'h1)))
                    begin
                      reg746 <= reg720;
                      reg747 <= $signed($unsigned((reg695 & ((8'h9d) ?
                          reg598 : forvar733))));
                    end
                  for (forvar748 = (1'h0); (forvar748 < (1'h0)); forvar748 = (forvar748 + (1'h1)))
                    begin
                      reg749 <= ($unsigned(((forvar660 ?
                              reg707 : reg673) >= $signed(forvar671))) ?
                          $unsigned(forvar588) : (~^forvar649[(1'h1):(1'h1)]));
                      reg750 <= (forvar697 <<< (+((~reg613) ^ $unsigned(reg650))));
                      reg751 <= $unsigned((((forvar630 && reg636) ?
                          (reg734 ?
                              reg627 : reg694) : (^~reg565)) != ($unsigned((8'h9f)) ?
                          (^~reg603) : $signed(reg578))));
                      reg752 <= ($unsigned(forvar626[(1'h0):(1'h0)]) < forvar573);
                    end
                  reg753 <= $unsigned(reg567);
                  reg754 <= ((($unsigned(reg663) ?
                          reg671 : $unsigned(reg598)) >>> reg593) ?
                      forvar702[(3'h5):(1'h1)] : $unsigned(($unsigned(reg752) ?
                          {reg614} : {reg691})));
                end
              if ((8'h9c))
                begin
                  reg755 <= reg571;
                  for (forvar756 = (1'h0); (forvar756 < (1'h1)); forvar756 = (forvar756 + (1'h1)))
                    begin
                      reg757 <= ($unsigned((&reg701)) ?
                          (~^((!reg750) && $unsigned(reg666))) : ($unsigned((8'hb1)) || reg742));
                      reg758 <= forvar699;
                      reg759 <= $signed(($signed($signed(reg746)) ?
                          (forvar722[(1'h1):(1'h1)] >= {forvar648}) : $unsigned($signed((8'hb6)))));
                      reg760 <= $signed(({(reg622 ? reg751 : forvar643)} ?
                          (~|(reg576 << reg571)) : ($unsigned(reg751) > $unsigned(reg735))));
                    end
                  for (forvar761 = (1'h0); (forvar761 < (1'h0)); forvar761 = (forvar761 + (1'h1)))
                    begin
                      reg762 <= (reg724 ?
                          (reg678 ?
                              $signed((forvar671 == forvar669)) : ((~^(8'h9c)) ?
                                  ((8'had) ?
                                      forvar702 : (8'ha8)) : (-forvar737))) : $signed(reg650));
                      reg763 <= (forvar620[(4'hb):(1'h1)] && {(reg698[(3'h4):(1'h1)] > reg685)});
                    end
                end
              else
                begin
                  if (($unsigned((~^{forvar660})) ?
                      (&($signed(reg669) < $signed(reg754))) : reg701))
                    begin
                      reg755 <= ({(^(&reg724))} - ((8'haf) ?
                          reg563 : ({forvar575} ? reg660 : $unsigned(reg634))));
                      reg756 <= ($unsigned((+(reg603 > forvar592))) <= forvar592);
                    end
                  else
                    begin
                      reg755 <= $unsigned((reg661 ?
                          (^~reg671[(4'hb):(3'h4)]) : {$unsigned((8'h9e))}));
                      reg756 <= reg692[(2'h2):(1'h1)];
                      reg757 <= {((^(+reg717)) ?
                              (8'ha4) : ({forvar584} ?
                                  reg569 : reg718[(2'h3):(1'h1)]))};
                      reg758 <= $unsigned((|(|reg586)));
                    end
                  for (forvar759 = (1'h0); (forvar759 < (1'h0)); forvar759 = (forvar759 + (1'h1)))
                    begin
                      reg760 <= reg593;
                      reg761 <= (|$unsigned((reg725[(1'h1):(1'h1)] ?
                          ((8'hb7) ? reg654 : forvar633) : {reg593})));
                      reg762 <= (~^$unsigned(reg677[(2'h2):(2'h2)]));
                    end
                  for (forvar763 = (1'h0); (forvar763 < (2'h2)); forvar763 = (forvar763 + (1'h1)))
                    begin
                      reg764 <= (8'hb6);
                      reg765 <= (((&(~|forvar722)) || ((!reg685) ?
                              reg738[(3'h4):(3'h4)] : $unsigned(reg727))) ?
                          reg718[(2'h3):(1'h1)] : $unsigned({(forvar571 ?
                                  forvar595 : (8'had))}));
                      reg766 <= (reg571 ? reg644 : (&wire560));
                      reg767 <= (~^(8'hb4));
                    end
                  for (forvar768 = (1'h0); (forvar768 < (2'h3)); forvar768 = (forvar768 + (1'h1)))
                    begin
                      reg769 <= reg616[(3'h5):(1'h1)];
                    end
                end
            end
          else
            begin
              reg741 <= (reg578[(1'h0):(1'h0)] ?
                  $signed({forvar638[(2'h3):(1'h0)]}) : (&{forvar655}));
              if (forvar761)
                begin
                  for (forvar742 = (1'h0); (forvar742 < (1'h0)); forvar742 = (forvar742 + (1'h1)))
                    begin
                      reg743 <= ((forvar601 ?
                          $unsigned((reg721 ?
                              reg613 : reg727)) : reg628[(4'hc):(4'h8)]) < (((+forvar745) ?
                              $signed(forvar600) : $signed(reg750)) ?
                          $unsigned((reg719 ?
                              reg597 : reg700)) : $unsigned({reg611})));
                      reg744 <= $unsigned((((forvar591 ?
                              reg724 : reg718) + {reg635}) ?
                          reg756 : reg611[(4'hf):(4'h9)]));
                      reg745 <= reg714[(3'h4):(1'h1)];
                      reg746 <= (-(~|reg758));
                    end
                  if (reg671[(4'hb):(4'h8)])
                    begin
                      reg747 <= ($signed((&(-reg565))) == ({reg708} - ($unsigned(reg675) ?
                          $signed(reg578) : forvar702)));
                      reg748 <= $unsigned((forvar638 ?
                          reg687[(1'h1):(1'h1)] : forvar648[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg747 <= (-(|(^forvar687)));
                      reg748 <= reg586[(1'h0):(1'h0)];
                      reg749 <= (~^$unsigned($signed(forvar763)));
                      reg750 <= forvar626[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if (($signed(reg706[(5'h10):(5'h10)]) ?
                      $signed((~|$unsigned(reg580))) : ((reg568[(2'h3):(2'h2)] ?
                              (~|(8'hb3)) : forvar733[(1'h1):(1'h1)]) ?
                          $unsigned((~forvar570)) : $unsigned(reg575[(3'h4):(2'h3)]))))
                    begin
                      reg742 <= (reg757[(4'hf):(4'hd)] ~^ reg565);
                      reg743 <= $signed((reg712 ?
                          forvar664 : (reg659 ?
                              (8'ha1) : reg742[(3'h5):(2'h3)])));
                      reg744 <= reg686[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg742 <= {$signed((-$unsigned(reg598)))};
                      reg743 <= reg676[(3'h6):(3'h5)];
                      reg744 <= reg680;
                      reg745 <= ((((reg617 ? reg753 : reg767) ?
                              (~reg643) : (^reg749)) ^~ (forvar668[(2'h2):(2'h2)] ?
                              {reg577} : $unsigned(reg757))) ?
                          (8'ha6) : ((~&(+forvar702)) * $unsigned((&(8'hb1)))));
                    end
                  for (forvar746 = (1'h0); (forvar746 < (1'h1)); forvar746 = (forvar746 + (1'h1)))
                    begin
                      reg747 <= reg619;
                      reg748 <= forvar697[(4'h8):(3'h4)];
                      reg749 <= (!$unsigned(((forvar695 ?
                          reg691 : wire556) > (!forvar756))));
                    end
                end
            end
          for (forvar770 = (1'h0); (forvar770 < (2'h2)); forvar770 = (forvar770 + (1'h1)))
            begin
              if ((reg758[(4'h9):(3'h7)] ?
                  $unsigned({(reg726 ? forvar731 : (8'ha4))}) : (8'h9e)))
                begin
                  if ({((^(|forvar589)) ?
                          (reg598 <<< $unsigned(reg676)) : $signed(forvar759[(4'he):(4'h8)]))})
                    begin
                      reg771 <= $signed({(~&((8'hb4) ~^ reg717))});
                      reg772 <= reg657;
                      reg773 <= $signed((forvar770[(1'h1):(1'h0)] <= $unsigned((8'h9f))));
                    end
                  else
                    begin
                      reg771 <= reg574;
                      reg772 <= $unsigned(reg606[(4'h9):(4'h9)]);
                      reg773 <= $signed($signed({(reg674 ?
                              forvar661 : reg680)}));
                    end
                end
              else
                begin
                  for (forvar771 = (1'h0); (forvar771 < (1'h0)); forvar771 = (forvar771 + (1'h1)))
                    begin
                      reg772 <= $unsigned((((reg602 ?
                          reg658 : reg662) | (forvar629 || reg767)) ^ $unsigned((|(8'haf)))));
                      reg773 <= $signed((~^$signed((~forvar745))));
                      reg774 <= ($signed((!$signed(reg710))) * (reg732 ?
                          {reg613} : $unsigned($unsigned(reg689))));
                    end
                  for (forvar775 = (1'h0); (forvar775 < (1'h1)); forvar775 = (forvar775 + (1'h1)))
                    begin
                      reg776 <= $unsigned((~&((^~reg650) ?
                          (reg570 ? reg694 : reg769) : (^~forvar671))));
                      reg777 <= ($signed(($signed(forvar745) ?
                          reg683[(1'h1):(1'h0)] : $signed(reg765))) <<< (+reg723[(3'h4):(2'h2)]));
                    end
                  for (forvar778 = (1'h0); (forvar778 < (2'h2)); forvar778 = (forvar778 + (1'h1)))
                    begin
                      reg779 <= (((&{reg648}) + $unsigned((reg577 && (8'hac)))) ^~ (((^~wire558) == (forvar741 ?
                          wire558 : forvar768)) << (reg661[(2'h2):(1'h1)] ?
                          {reg565} : reg632)));
                      reg780 <= (reg606[(4'h9):(1'h0)] ?
                          $signed(reg710[(3'h6):(3'h4)]) : reg678);
                      reg781 <= {(~^$signed($signed((8'ha9))))};
                      reg782 <= $signed({reg570[(3'h7):(3'h6)]});
                    end
                end
              for (forvar783 = (1'h0); (forvar783 < (2'h3)); forvar783 = (forvar783 + (1'h1)))
                begin
                  for (forvar784 = (1'h0); (forvar784 < (1'h1)); forvar784 = (forvar784 + (1'h1)))
                    begin
                      reg785 <= (|$signed(((reg565 ~^ reg581) > forvar681[(4'hc):(3'h6)])));
                      reg786 <= (($signed($unsigned(reg716)) ?
                              ((&(8'ha1)) ?
                                  (forvar783 < reg659) : forvar676[(2'h2):(2'h2)]) : (~&forvar571)) ?
                          $unsigned(reg602) : (forvar647[(2'h3):(1'h0)] ^~ reg734[(3'h5):(1'h1)]));
                    end
                  for (forvar787 = (1'h0); (forvar787 < (2'h2)); forvar787 = (forvar787 + (1'h1)))
                    begin
                      reg788 <= (reg779[(3'h4):(1'h0)] + ({reg780} - reg709[(4'hc):(3'h4)]));
                      reg789 <= (^~forvar652[(4'hb):(3'h6)]);
                    end
                  for (forvar790 = (1'h0); (forvar790 < (2'h3)); forvar790 = (forvar790 + (1'h1)))
                    begin
                      reg791 <= reg767[(3'h5):(2'h2)];
                      reg792 <= $unsigned($unsigned({(&(8'hb8))}));
                    end
                end
              if ((~|reg792))
                begin
                  reg793 <= reg616[(1'h1):(1'h1)];
                end
              else
                begin
                  reg793 <= (reg741[(2'h2):(2'h2)] ?
                      $unsigned(({(8'h9e)} ?
                          $signed(reg637) : (|forvar689))) : $unsigned($signed(reg702)));
                  if (($unsigned((8'h9f)) ?
                      $signed((reg573[(1'h1):(1'h0)] ?
                          (forvar737 ^~ reg758) : reg724[(4'h8):(3'h6)])) : (reg663[(4'ha):(2'h2)] != {{reg597}})))
                    begin
                      reg794 <= (reg703 && (8'haf));
                      reg795 <= (({reg570[(1'h1):(1'h1)]} ?
                          forvar626 : $unsigned(forvar745)) - $unsigned($signed((reg758 << forvar595))));
                      reg796 <= $signed(reg785);
                      reg797 <= ($unsigned({(reg577 ? reg710 : reg772)}) ?
                          reg767 : $signed(((|reg610) ?
                              (reg777 ^ (8'haa)) : (~reg744))));
                    end
                  else
                    begin
                      reg794 <= ($signed((~^(8'hb5))) ?
                          $signed((~^$signed(reg762))) : (((8'haf) << {forvar778}) ?
                              (~|reg728[(1'h1):(1'h1)]) : $signed({forvar668})));
                      reg795 <= {$signed((reg606[(4'h8):(1'h1)] ?
                              (reg686 ?
                                  reg661 : (8'h9e)) : reg695[(3'h7):(2'h2)]))};
                      reg796 <= (reg636[(3'h6):(3'h5)] ~^ $signed($signed(reg645[(2'h2):(1'h0)])));
                    end
                  for (forvar798 = (1'h0); (forvar798 < (1'h0)); forvar798 = (forvar798 + (1'h1)))
                    begin
                      reg799 <= $unsigned(reg779[(3'h6):(2'h2)]);
                      reg800 <= $unsigned($signed(((8'haa) ?
                          $unsigned((8'ha7)) : reg719[(1'h0):(1'h0)])));
                      reg801 <= (reg580[(3'h7):(2'h3)] * reg661[(1'h0):(1'h0)]);
                      reg802 <= {reg576[(3'h6):(2'h2)]};
                    end
                  if ($unsigned((({reg609} != reg612[(1'h1):(1'h1)]) ?
                      (!forvar644[(4'ha):(3'h4)]) : $unsigned({reg618}))))
                    begin
                      reg803 <= forvar770;
                      reg804 <= {(+(~(reg688 ^ (8'ha0))))};
                      reg805 <= (reg744[(3'h6):(2'h3)] ?
                          (((&forvar775) || ((8'hb3) || (8'h9c))) ?
                              (&(reg670 ?
                                  reg712 : (8'h9c))) : reg752[(4'h8):(3'h7)]) : reg747);
                    end
                  else
                    begin
                      reg803 <= {$unsigned($signed((reg721 > forvar630)))};
                      reg804 <= $signed({(8'haf)});
                      reg805 <= reg665;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(reg625[(4'h8):(3'h7)]))
        begin
          if ($unsigned(($unsigned(reg759[(1'h1):(1'h0)]) ?
              $signed((forvar775 ? (8'ha9) : (8'hb2))) : (^~(forvar644 ?
                  (8'h9d) : (8'ha3))))))
            begin
              if ((forvar650 ?
                  reg666[(3'h7):(2'h3)] : (($unsigned(reg684) * ((8'hba) ?
                          forvar784 : (8'ha6))) ?
                      ((forvar570 < forvar626) - reg735) : (~&reg574[(3'h4):(2'h2)]))))
                begin
                  reg806 <= ((!$unsigned((reg776 ?
                      reg575 : reg701))) ~^ $signed((reg692 ?
                      (wire557 ^~ reg580) : $signed(reg672))));
                end
              else
                begin
                  for (forvar806 = (1'h0); (forvar806 < (2'h3)); forvar806 = (forvar806 + (1'h1)))
                    begin
                      reg807 <= $signed($unsigned(forvar664));
                      reg808 <= reg674;
                      reg809 <= (&(~&forvar731));
                      reg810 <= forvar722[(2'h3):(1'h1)];
                    end
                  for (forvar811 = (1'h0); (forvar811 < (1'h1)); forvar811 = (forvar811 + (1'h1)))
                    begin
                      reg812 <= {reg732};
                    end
                  reg813 <= ($signed(forvar591) >> (+(^~$signed(reg678))));
                end
              for (forvar814 = (1'h0); (forvar814 < (2'h3)); forvar814 = (forvar814 + (1'h1)))
                begin
                  if ($unsigned(((!(reg723 ?
                      forvar660 : reg669)) ^ ((forvar652 <<< reg580) >> $signed(reg781)))))
                    begin
                      reg815 <= (~|forvar633[(1'h1):(1'h0)]);
                      reg816 <= (~&({$signed(reg767)} ?
                          ((reg634 * reg659) ?
                              (reg667 ?
                                  reg591 : reg668) : reg732) : (-(forvar608 ?
                              (8'hb6) : reg694))));
                    end
                  else
                    begin
                      reg815 <= forvar608;
                      reg816 <= $unsigned(($unsigned((-reg644)) ?
                          $signed(forvar652) : (reg704 >> $unsigned(reg639))));
                      reg817 <= $signed(reg610[(2'h3):(1'h1)]);
                      reg818 <= $unsigned(($unsigned((reg577 ^ (8'h9c))) ?
                          $unsigned(forvar601[(3'h6):(3'h5)]) : $signed($unsigned(forvar640))));
                    end
                  for (forvar819 = (1'h0); (forvar819 < (1'h1)); forvar819 = (forvar819 + (1'h1)))
                    begin
                      reg820 <= (^(((reg672 - (8'h9c)) == reg601) ~^ $signed((reg712 ?
                          (8'hac) : reg575))));
                      reg821 <= forvar575[(4'h9):(3'h6)];
                      reg822 <= {(((forvar783 ? forvar722 : forvar652) ?
                                  (forvar621 + reg690) : (8'ha1)) ?
                              reg805 : ((~reg750) ?
                                  (~&(8'h9d)) : (reg646 ^ forvar652)))};
                      reg823 <= reg606;
                    end
                end
              for (forvar824 = (1'h0); (forvar824 < (2'h3)); forvar824 = (forvar824 + (1'h1)))
                begin
                  reg825 <= reg669;
                  reg826 <= ((^($unsigned((8'ha3)) || {reg718})) || (^~$unsigned((-(8'ha1)))));
                end
            end
          else
            begin
              for (forvar806 = (1'h0); (forvar806 < (1'h0)); forvar806 = (forvar806 + (1'h1)))
                begin
                  reg807 <= {(!forvar775)};
                end
            end
        end
      else
        begin
          reg806 <= ($signed(reg720) <= $unsigned($unsigned(forvar768[(2'h3):(1'h1)])));
          reg807 <= ($unsigned((reg816 ?
              $unsigned(reg807) : reg651)) ^ reg786[(1'h1):(1'h0)]);
        end
      if ((^(8'ha7)))
        begin
          reg827 <= $signed((!reg647[(4'ha):(4'h8)]));
          if (reg616[(2'h2):(2'h2)])
            begin
              for (forvar828 = (1'h0); (forvar828 < (2'h2)); forvar828 = (forvar828 + (1'h1)))
                begin
                  for (forvar829 = (1'h0); (forvar829 < (2'h2)); forvar829 = (forvar829 + (1'h1)))
                    begin
                      reg830 <= $unsigned((8'hb7));
                    end
                  if ($unsigned(reg758))
                    begin
                      reg831 <= wire557[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg831 <= (($signed((reg648 & reg590)) ?
                              ($unsigned(forvar819) ?
                                  (~reg613) : (reg703 ?
                                      forvar731 : forvar811)) : $signed((^~reg747))) ?
                          (((reg587 ? reg608 : forvar656) ?
                              reg645[(3'h6):(3'h4)] : $unsigned(reg772)) & $unsigned((reg793 ?
                              reg635 : wire557))) : reg567);
                    end
                  for (forvar832 = (1'h0); (forvar832 < (2'h3)); forvar832 = (forvar832 + (1'h1)))
                    begin
                      reg833 <= (($unsigned(reg746[(1'h1):(1'h1)]) ?
                              ({forvar668} * (forvar763 <= reg618)) : reg701) ?
                          $unsigned(($signed(forvar798) < (~&reg735))) : forvar819[(2'h2):(1'h1)]);
                      reg834 <= (|reg774);
                    end
                  if ({({((8'hb9) ^~ reg634)} & (|(reg637 - (8'hba))))})
                    begin
                      reg835 <= $unsigned($unsigned({{forvar562}}));
                      reg836 <= forvar674;
                      reg837 <= reg599[(3'h5):(3'h5)];
                      reg838 <= reg687;
                    end
                  else
                    begin
                      reg835 <= $unsigned(reg628[(1'h0):(1'h0)]);
                      reg836 <= $unsigned(forvar615);
                    end
                end
              reg839 <= (^reg624[(3'h4):(1'h0)]);
              if (($unsigned((~^(!reg666))) - $signed((reg804[(4'h9):(3'h4)] ?
                  (forvar589 ? reg651 : reg765) : forvar659[(2'h3):(2'h3)]))))
                begin
                  if (reg701[(3'h5):(1'h0)])
                    begin
                      reg840 <= (8'h9c);
                      reg841 <= ($signed((-(^~(8'ha4)))) ?
                          ($signed(forvar713) <<< (~{reg753})) : (|((reg796 * reg813) - reg659)));
                      reg842 <= $signed($unsigned(reg774));
                      reg843 <= ({(~&reg728)} + reg754);
                    end
                  else
                    begin
                      reg840 <= {reg702[(1'h1):(1'h0)]};
                      reg841 <= $signed(reg614);
                    end
                  for (forvar844 = (1'h0); (forvar844 < (1'h1)); forvar844 = (forvar844 + (1'h1)))
                    begin
                      reg845 <= {{(reg732[(1'h0):(1'h0)] ^ (forvar745 << reg580))}};
                      reg846 <= $unsigned((($signed(reg791) >> ((8'hb8) ?
                          (8'hb4) : forvar746)) + ($unsigned(reg647) ?
                          reg635[(3'h5):(3'h4)] : reg764[(2'h3):(1'h1)])));
                      reg847 <= reg818[(1'h0):(1'h0)];
                    end
                  if ($signed({$signed(forvar564[(3'h6):(3'h4)])}))
                    begin
                      reg848 <= forvar713[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg848 <= (8'hae);
                      reg849 <= $unsigned($signed((8'ha5)));
                      reg850 <= ($signed({(~&reg709)}) ?
                          ((reg700 > (reg601 ? reg772 : reg571)) ?
                              $signed((reg612 <<< reg618)) : forvar731[(4'ha):(4'h9)]) : $signed(reg836));
                    end
                end
              else
                begin
                  for (forvar840 = (1'h0); (forvar840 < (1'h1)); forvar840 = (forvar840 + (1'h1)))
                    begin
                      reg841 <= (reg635 ?
                          ((!reg590) <= reg568[(3'h4):(2'h2)]) : (({forvar571} ?
                                  (reg715 <<< reg583) : reg781) ?
                              reg764[(4'hc):(1'h1)] : reg666));
                      reg842 <= ((~|wire557[(1'h0):(1'h0)]) ?
                          ((|(|(8'h9d))) > ($unsigned(reg680) ?
                              reg585 : (~(8'hb6)))) : (|(((8'ha2) || forvar631) ?
                              forvar730[(3'h6):(3'h6)] : reg797)));
                      reg843 <= $signed((^$unsigned((~&reg684))));
                      reg844 <= (&(($unsigned(reg831) ?
                          $unsigned(forvar650) : (^~forvar633)) <<< (^(reg706 ?
                          (8'ha1) : reg649))));
                    end
                  if ({wire559[(3'h5):(1'h1)]})
                    begin
                      reg845 <= (({$signed(reg706)} && $unsigned($unsigned(forvar575))) ?
                          (^(-(~^forvar664))) : (({reg661} ^~ (reg707 & reg769)) ?
                              $unsigned((~^forvar564)) : reg833));
                      reg846 <= {{(reg769[(2'h3):(1'h0)] ?
                                  (forvar828 * forvar756) : reg801)}};
                    end
                  else
                    begin
                      reg845 <= forvar592[(3'h6):(3'h6)];
                      reg846 <= reg645;
                      reg847 <= (reg820 < (8'hb4));
                    end
                end
            end
          else
            begin
              if (($unsigned(forvar806) ?
                  {reg568} : (($unsigned(reg650) ?
                      (^(8'hb9)) : (forvar704 ?
                          (8'ha3) : reg769)) | forvar629)))
                begin
                  if (({reg804} ?
                      $signed((^~((8'haf) <<< forvar770))) : reg759[(3'h5):(2'h2)]))
                    begin
                      reg828 <= reg751;
                      reg829 <= ($unsigned(reg845) ?
                          $signed(reg666[(2'h3):(1'h1)]) : $unsigned(($signed(reg797) ?
                              (reg804 + forvar819) : {(8'hb7)})));
                      reg830 <= (reg844[(3'h6):(3'h4)] ?
                          (~^(reg605 ? (reg625 && (8'hb2)) : reg751)) : reg642);
                    end
                  else
                    begin
                      reg828 <= (~$unsigned(reg780));
                      reg829 <= reg605;
                      reg830 <= $unsigned(reg788[(1'h0):(1'h0)]);
                      reg831 <= $signed(reg846[(2'h3):(2'h2)]);
                    end
                  reg832 <= reg590[(2'h3):(1'h1)];
                end
              else
                begin
                  for (forvar828 = (1'h0); (forvar828 < (1'h0)); forvar828 = (forvar828 + (1'h1)))
                    begin
                      reg829 <= ((((reg698 ?
                              reg649 : reg578) ^ $unsigned(reg816)) >= reg829[(4'hb):(3'h7)]) ?
                          reg777 : $signed((forvar702 ?
                              (reg651 + reg671) : (~^reg680))));
                    end
                  reg830 <= $signed(({$unsigned((8'ha1))} == $unsigned(reg752)));
                  for (forvar831 = (1'h0); (forvar831 < (2'h2)); forvar831 = (forvar831 + (1'h1)))
                    begin
                      reg832 <= $signed(forvar759[(4'hd):(1'h1)]);
                      reg833 <= (|{((~|forvar832) ~^ reg708[(2'h3):(2'h3)])});
                    end
                end
              for (forvar834 = (1'h0); (forvar834 < (2'h3)); forvar834 = (forvar834 + (1'h1)))
                begin
                  reg835 <= reg608;
                  for (forvar836 = (1'h0); (forvar836 < (2'h3)); forvar836 = (forvar836 + (1'h1)))
                    begin
                      reg837 <= $unsigned(reg738[(4'h9):(2'h3)]);
                      reg838 <= ($signed((&$unsigned(forvar643))) >>> reg723);
                    end
                  if (reg782[(1'h0):(1'h0)])
                    begin
                      reg839 <= ({$signed(reg764)} <= (forvar790 || (~&{(8'ha8)})));
                      reg840 <= (reg796 - (({forvar763} <<< ((8'hb7) >> reg692)) ?
                          $signed($signed(reg659)) : (+forvar704)));
                      reg841 <= (8'ha6);
                      reg842 <= $unsigned({(-reg837)});
                    end
                  else
                    begin
                      reg839 <= ($signed(($signed(reg654) >> reg748)) ?
                          reg803 : forvar697[(4'h8):(3'h5)]);
                    end
                end
              for (forvar843 = (1'h0); (forvar843 < (1'h1)); forvar843 = (forvar843 + (1'h1)))
                begin
                  for (forvar844 = (1'h0); (forvar844 < (2'h3)); forvar844 = (forvar844 + (1'h1)))
                    begin
                      reg845 <= reg729[(4'hd):(1'h1)];
                      reg846 <= {($unsigned($signed(reg714)) ^ reg731[(3'h5):(3'h4)])};
                    end
                  reg847 <= {(~&{reg706[(2'h3):(2'h2)]})};
                end
            end
          if (((+(!reg807[(3'h5):(3'h4)])) != reg646[(3'h7):(3'h7)]))
            begin
              if ({$signed(reg735)})
                begin
                  for (forvar851 = (1'h0); (forvar851 < (2'h3)); forvar851 = (forvar851 + (1'h1)))
                    begin
                      reg852 <= reg712;
                      reg853 <= ((~^reg572) ?
                          ($unsigned(reg846) < reg572[(2'h3):(2'h2)]) : ((^$signed(reg729)) << reg574));
                      reg854 <= forvar591[(3'h6):(3'h5)];
                    end
                  if ($unsigned($unsigned((&(8'ha9)))))
                    begin
                      reg855 <= {(!(+reg636))};
                      reg856 <= forvar602;
                      reg857 <= (8'hb0);
                      reg858 <= $signed((^$unsigned((forvar630 ?
                          (8'ha4) : reg702))));
                    end
                  else
                    begin
                      reg855 <= $signed($unsigned({(reg810 == reg727)}));
                      reg856 <= reg692;
                      reg857 <= (!(8'ha9));
                      reg858 <= (^~reg761[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar851 = (1'h0); (forvar851 < (2'h3)); forvar851 = (forvar851 + (1'h1)))
                    begin
                      reg852 <= $signed($unsigned($unsigned(reg718[(3'h6):(2'h3)])));
                    end
                  for (forvar853 = (1'h0); (forvar853 < (2'h2)); forvar853 = (forvar853 + (1'h1)))
                    begin
                      reg854 <= reg591[(2'h2):(1'h0)];
                      reg855 <= (((-(reg817 >= reg802)) >>> (|forvar600[(2'h3):(2'h3)])) <<< $unsigned($unsigned((-(8'hb9)))));
                      reg856 <= $signed(reg645);
                      reg857 <= $signed(({$unsigned(reg714)} ?
                          (~|forvar595) : $unsigned($signed(reg773))));
                    end
                  reg858 <= $unsigned(((8'hb5) ?
                      (~|$unsigned(reg832)) : reg718[(1'h1):(1'h0)]));
                end
              if ({$unsigned(((^forvar602) ? reg664[(3'h6):(2'h2)] : reg773))})
                begin
                  for (forvar859 = (1'h0); (forvar859 < (1'h1)); forvar859 = (forvar859 + (1'h1)))
                    begin
                      reg860 <= (reg628 | $unsigned(($unsigned(reg841) ?
                          $signed(forvar641) : $signed(reg812))));
                      reg861 <= (({reg843} ~^ ((reg714 >>> reg761) ?
                          {reg747} : (reg726 ?
                              reg602 : reg734))) == $signed(reg781));
                      reg862 <= (forvar787 ?
                          forvar775 : {forvar671[(4'h8):(1'h1)]});
                    end
                  for (forvar863 = (1'h0); (forvar863 < (1'h0)); forvar863 = (forvar863 + (1'h1)))
                    begin
                      reg864 <= reg763[(2'h3):(1'h1)];
                      reg865 <= $signed(reg772);
                      reg866 <= (+(^($signed(reg754) | $signed(reg683))));
                    end
                  for (forvar867 = (1'h0); (forvar867 < (1'h1)); forvar867 = (forvar867 + (1'h1)))
                    begin
                      reg868 <= (~^$signed($unsigned({reg583})));
                      reg869 <= forvar768;
                      reg870 <= $signed($signed((~^reg569[(1'h0):(1'h0)])));
                      reg871 <= (8'had);
                    end
                  for (forvar872 = (1'h0); (forvar872 < (2'h3)); forvar872 = (forvar872 + (1'h1)))
                    begin
                      reg873 <= reg624;
                    end
                end
              else
                begin
                  if ((8'ha2))
                    begin
                      reg859 <= $signed((reg603[(1'h0):(1'h0)] || $unsigned($unsigned(reg801))));
                      reg860 <= ((($unsigned(reg835) - (forvar584 - reg767)) - $unsigned(reg616)) || ($signed((reg623 > (8'h9f))) ?
                          reg796 : ((forvar638 * reg765) ?
                              reg674[(3'h4):(1'h0)] : {reg712})));
                    end
                  else
                    begin
                      reg859 <= ((($unsigned((8'hb4)) - $signed(forvar591)) ?
                              {reg569} : forvar629) ?
                          reg703[(4'ha):(2'h3)] : (reg846[(3'h4):(3'h4)] ?
                              {(~|forvar851)} : {reg771[(3'h5):(2'h2)]}));
                      reg860 <= $signed(reg614);
                    end
                  for (forvar861 = (1'h0); (forvar861 < (1'h1)); forvar861 = (forvar861 + (1'h1)))
                    begin
                      reg862 <= {forvar704};
                      reg863 <= {forvar693};
                      reg864 <= reg568;
                      reg865 <= (!$unsigned($unsigned({forvar828})));
                    end
                end
            end
          else
            begin
              if (($unsigned($unsigned(forvar640[(2'h3):(1'h1)])) ?
                  forvar584 : ($signed((^reg672)) ?
                      ({reg813} ?
                          reg625[(1'h0):(1'h0)] : (reg808 ?
                              reg763 : forvar650)) : reg792)))
                begin
                  reg851 <= ($signed($signed((~&reg821))) > ($signed($unsigned(forvar771)) + ($signed(reg856) + (~|reg716))));
                end
              else
                begin
                  for (forvar851 = (1'h0); (forvar851 < (2'h2)); forvar851 = (forvar851 + (1'h1)))
                    begin
                      reg852 <= $signed((forvar730 ?
                          reg602[(2'h2):(1'h1)] : $unsigned($signed((8'hab)))));
                    end
                  for (forvar853 = (1'h0); (forvar853 < (2'h2)); forvar853 = (forvar853 + (1'h1)))
                    begin
                      reg854 <= reg613;
                      reg855 <= (8'hb6);
                      reg856 <= reg785;
                      reg857 <= (reg742[(2'h3):(1'h1)] * $unsigned(reg613[(1'h0):(1'h0)]));
                    end
                  for (forvar858 = (1'h0); (forvar858 < (2'h2)); forvar858 = (forvar858 + (1'h1)))
                    begin
                      reg859 <= forvar851[(3'h6):(2'h2)];
                      reg860 <= $signed($unsigned(forvar595[(4'ha):(3'h4)]));
                    end
                end
              for (forvar861 = (1'h0); (forvar861 < (2'h3)); forvar861 = (forvar861 + (1'h1)))
                begin
                  for (forvar862 = (1'h0); (forvar862 < (2'h2)); forvar862 = (forvar862 + (1'h1)))
                    begin
                      reg863 <= ($signed($unsigned(reg785[(1'h1):(1'h0)])) ^~ $unsigned(($unsigned(reg652) ?
                          $signed(forvar649) : reg632[(4'h9):(2'h3)])));
                      reg864 <= (~&$unsigned(forvar669));
                    end
                end
              for (forvar865 = (1'h0); (forvar865 < (1'h1)); forvar865 = (forvar865 + (1'h1)))
                begin
                  for (forvar866 = (1'h0); (forvar866 < (1'h0)); forvar866 = (forvar866 + (1'h1)))
                    begin
                      reg867 <= (forvar733[(4'h9):(3'h6)] && (8'ha8));
                      reg868 <= reg573[(2'h2):(1'h0)];
                    end
                  reg869 <= ((|reg832) < (reg694 ?
                      $unsigned((|reg665)) : reg858));
                end
              for (forvar870 = (1'h0); (forvar870 < (2'h2)); forvar870 = (forvar870 + (1'h1)))
                begin
                  for (forvar871 = (1'h0); (forvar871 < (1'h1)); forvar871 = (forvar871 + (1'h1)))
                    begin
                      reg872 <= (~&(reg822 ? (8'hb0) : reg708[(1'h0):(1'h0)]));
                    end
                  if ((reg637[(3'h7):(1'h0)] ?
                      $unsigned(reg808[(2'h3):(2'h2)]) : (((~|reg808) ?
                          (~&(8'hba)) : $signed((8'ha9))) ^~ $signed({reg839}))))
                    begin
                      reg873 <= (forvar562 + reg757);
                      reg874 <= {reg870};
                      reg875 <= ($signed((^$unsigned(reg580))) | (reg741 > ((+forvar870) ^~ reg687[(4'ha):(2'h2)])));
                      reg876 <= forvar756[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg873 <= (!$signed($signed(forvar688)));
                      reg874 <= ($signed((~|reg705[(4'ha):(3'h4)])) && (~^((reg812 - reg702) ^ forvar746)));
                    end
                  if ((reg808[(1'h0):(1'h0)] ?
                      {$unsigned(reg734)} : reg586[(2'h2):(2'h2)]))
                    begin
                      reg877 <= forvar871;
                      reg878 <= $signed((!$unsigned($signed((8'hb7)))));
                    end
                  else
                    begin
                      reg877 <= (8'ha3);
                      reg878 <= forvar676;
                      reg879 <= forvar778;
                      reg880 <= {reg714[(2'h3):(2'h3)]};
                    end
                  for (forvar881 = (1'h0); (forvar881 < (1'h0)); forvar881 = (forvar881 + (1'h1)))
                    begin
                      reg882 <= reg761[(4'hd):(4'h8)];
                    end
                end
            end
        end
      else
        begin
          reg827 <= (8'ha0);
        end
      if ((&(^~reg776)))
        begin
          if ((+($signed((reg793 || reg786)) ?
              $signed(reg694[(2'h3):(2'h3)]) : (reg771[(2'h3):(2'h3)] << (reg797 - reg841)))))
            begin
              if ((~|({reg719} >> {(forvar770 ? forvar601 : reg856)})))
                begin
                  for (forvar883 = (1'h0); (forvar883 < (1'h1)); forvar883 = (forvar883 + (1'h1)))
                    begin
                      reg884 <= (reg760 ?
                          ({$signed(reg646)} ?
                              ($signed(reg810) ?
                                  $signed((8'hb3)) : {(8'haa)}) : ($signed(reg875) ?
                                  (8'ha8) : (reg863 * forvar644))) : (^forvar621));
                      reg885 <= $signed($signed(($unsigned(forvar761) ?
                          $signed(reg573) : (forvar649 && forvar853))));
                    end
                  for (forvar886 = (1'h0); (forvar886 < (1'h1)); forvar886 = (forvar886 + (1'h1)))
                    begin
                      reg887 <= reg797[(3'h4):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar883 = (1'h0); (forvar883 < (2'h2)); forvar883 = (forvar883 + (1'h1)))
                    begin
                      reg884 <= (($signed({reg648}) ?
                          (^forvar640[(4'hb):(4'h9)]) : (8'hb7)) >= ({$unsigned(reg745)} && $signed($signed((8'ha5)))));
                    end
                end
              for (forvar888 = (1'h0); (forvar888 < (2'h2)); forvar888 = (forvar888 + (1'h1)))
                begin
                  for (forvar889 = (1'h0); (forvar889 < (2'h3)); forvar889 = (forvar889 + (1'h1)))
                    begin
                      reg890 <= wire557;
                      reg891 <= (((!forvar564) ?
                          (8'hb1) : reg592[(3'h4):(1'h1)]) << (&reg827[(1'h0):(1'h0)]));
                      reg892 <= (reg808[(2'h2):(1'h0)] != (!(~|$unsigned(reg635))));
                      reg893 <= (reg603[(1'h0):(1'h0)] ? forvar671 : (+reg565));
                    end
                end
              for (forvar894 = (1'h0); (forvar894 < (1'h0)); forvar894 = (forvar894 + (1'h1)))
                begin
                  if ($unsigned({reg695[(2'h3):(2'h2)]}))
                    begin
                      reg895 <= reg612[(4'h8):(1'h0)];
                      reg896 <= $signed({(!{reg652})});
                      reg897 <= $unsigned($unsigned(forvar608[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg895 <= $signed($unsigned(reg792));
                      reg896 <= (reg726 || $unsigned((reg796 ?
                          (8'ha8) : (reg846 ? reg721 : (8'ha8)))));
                      reg897 <= {reg801};
                      reg898 <= (~|(reg785 - ($unsigned(reg795) ?
                          (8'ha8) : (|reg884))));
                    end
                  reg899 <= ($signed(((forvar652 ~^ forvar881) == forvar731)) > (8'ha3));
                  reg900 <= (8'hae);
                end
            end
          else
            begin
              for (forvar883 = (1'h0); (forvar883 < (1'h1)); forvar883 = (forvar883 + (1'h1)))
                begin
                  for (forvar884 = (1'h0); (forvar884 < (2'h2)); forvar884 = (forvar884 + (1'h1)))
                    begin
                      reg885 <= $unsigned({(~|forvar819)});
                      reg886 <= ((reg654[(2'h2):(2'h2)] ?
                          (^(!reg625)) : (|(~(8'hb7)))) >> ({$unsigned(reg801)} ?
                          $signed($unsigned((8'ha0))) : $signed($unsigned(reg782))));
                    end
                  for (forvar887 = (1'h0); (forvar887 < (2'h3)); forvar887 = (forvar887 + (1'h1)))
                    begin
                      reg888 <= $signed((8'hb8));
                      reg889 <= $signed(reg575[(3'h5):(1'h1)]);
                      reg890 <= $unsigned(reg669);
                      reg891 <= ((($unsigned((8'haf)) ?
                                  (8'hb5) : ((8'hac) | reg671)) ?
                              ((^~reg810) ?
                                  forvar859 : reg849[(3'h7):(3'h4)]) : $unsigned(reg666)) ?
                          $signed((&(-(8'h9e)))) : (8'ha5));
                    end
                  reg892 <= forvar870;
                end
              if (forvar626)
                begin
                  for (forvar893 = (1'h0); (forvar893 < (2'h2)); forvar893 = (forvar893 + (1'h1)))
                    begin
                      reg894 <= forvar671;
                    end
                  for (forvar895 = (1'h0); (forvar895 < (2'h3)); forvar895 = (forvar895 + (1'h1)))
                    begin
                      reg896 <= $signed(reg859[(3'h4):(1'h1)]);
                      reg897 <= (|$unsigned($signed(forvar674[(4'ha):(3'h5)])));
                    end
                  if (($signed($signed($signed((8'ha2)))) >= forvar629))
                    begin
                      reg898 <= forvar824;
                      reg899 <= reg825;
                      reg900 <= $signed($unsigned(($signed(reg838) && (reg601 ?
                          forvar742 : reg886))));
                    end
                  else
                    begin
                      reg898 <= (+reg834);
                      reg899 <= (^~$unsigned(((reg714 || reg888) ?
                          (|reg592) : (reg793 ? (8'hba) : reg842))));
                    end
                  for (forvar901 = (1'h0); (forvar901 < (1'h0)); forvar901 = (forvar901 + (1'h1)))
                    begin
                      reg902 <= reg850[(2'h3):(2'h3)];
                      reg903 <= {($unsigned((~|forvar689)) ?
                              ((^(8'hac)) | {forvar699}) : (^$signed(reg898)))};
                      reg904 <= $signed($signed(($unsigned(reg898) ?
                          reg815[(3'h6):(3'h4)] : $unsigned(forvar570))));
                      reg905 <= forvar778[(4'h8):(4'h8)];
                    end
                end
              else
                begin
                  reg893 <= forvar771[(1'h1):(1'h1)];
                  for (forvar894 = (1'h0); (forvar894 < (2'h3)); forvar894 = (forvar894 + (1'h1)))
                    begin
                      reg895 <= reg635;
                      reg896 <= {((wire555 <= reg738[(4'ha):(3'h7)]) <= (&forvar886[(3'h7):(3'h5)]))};
                    end
                  for (forvar897 = (1'h0); (forvar897 < (1'h0)); forvar897 = (forvar897 + (1'h1)))
                    begin
                      reg898 <= $signed({($unsigned(reg800) ?
                              $unsigned(reg869) : $signed((8'ha5)))});
                    end
                  for (forvar899 = (1'h0); (forvar899 < (1'h0)); forvar899 = (forvar899 + (1'h1)))
                    begin
                      reg900 <= $unsigned((forvar733[(1'h1):(1'h0)] ^ $unsigned($signed(reg862))));
                      reg901 <= (({forvar897[(2'h2):(2'h2)]} >> ($signed(reg720) || $unsigned(reg667))) ?
                          {forvar647[(4'hc):(4'h8)]} : $signed(reg812));
                      reg902 <= reg835;
                    end
                end
              for (forvar906 = (1'h0); (forvar906 < (1'h0)); forvar906 = (forvar906 + (1'h1)))
                begin
                  for (forvar907 = (1'h0); (forvar907 < (1'h0)); forvar907 = (forvar907 + (1'h1)))
                    begin
                      reg908 <= wire561;
                      reg909 <= forvar722;
                      reg910 <= (~(({reg690} ?
                              reg693[(1'h0):(1'h0)] : $signed(forvar676)) ?
                          (reg625[(4'hc):(4'ha)] ?
                              forvar591 : (&reg803)) : (!reg887)));
                    end
                  for (forvar911 = (1'h0); (forvar911 < (2'h3)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= ({(!reg575)} ?
                          reg647[(2'h3):(2'h2)] : ($unsigned(reg657[(3'h5):(2'h2)]) ?
                              $signed($unsigned(reg617)) : (((8'haf) ?
                                  (8'hab) : forvar607) * {forvar620})));
                      reg913 <= reg843;
                      reg914 <= ((^reg726) ?
                          (~^{$signed(forvar867)}) : {$signed($signed(reg813))});
                      reg915 <= $signed(reg577);
                    end
                end
            end
          reg916 <= {$unsigned(($signed(forvar745) ? reg755 : (&reg601)))};
          for (forvar917 = (1'h0); (forvar917 < (2'h2)); forvar917 = (forvar917 + (1'h1)))
            begin
              for (forvar918 = (1'h0); (forvar918 < (1'h1)); forvar918 = (forvar918 + (1'h1)))
                begin
                  reg919 <= (forvar746 ?
                      (~|(~^((8'hba) & reg863))) : $unsigned((~forvar615[(3'h7):(3'h7)])));
                  for (forvar920 = (1'h0); (forvar920 < (2'h3)); forvar920 = (forvar920 + (1'h1)))
                    begin
                      reg921 <= ((reg616 ?
                          {(reg793 - wire560)} : (~|(reg850 ^~ forvar918))) || $signed(reg875[(3'h4):(2'h2)]));
                    end
                  for (forvar922 = (1'h0); (forvar922 < (1'h1)); forvar922 = (forvar922 + (1'h1)))
                    begin
                      reg923 <= ($signed(forvar861) | reg894[(4'h9):(1'h1)]);
                      reg924 <= (reg660 ? {reg664} : reg634);
                    end
                end
            end
          for (forvar925 = (1'h0); (forvar925 < (1'h0)); forvar925 = (forvar925 + (1'h1)))
            begin
              for (forvar926 = (1'h0); (forvar926 < (1'h0)); forvar926 = (forvar926 + (1'h1)))
                begin
                  for (forvar927 = (1'h0); (forvar927 < (2'h3)); forvar927 = (forvar927 + (1'h1)))
                    begin
                      reg928 <= forvar661[(1'h1):(1'h0)];
                      reg929 <= forvar894[(2'h3):(1'h1)];
                      reg930 <= reg605;
                    end
                  if ((reg829[(3'h6):(3'h5)] ?
                      reg854[(2'h2):(2'h2)] : (+(~|(reg647 ?
                          forvar843 : forvar649)))))
                    begin
                      reg931 <= (+$signed($unsigned(reg719)));
                    end
                  else
                    begin
                      reg931 <= $signed(($signed((reg904 | reg850)) ?
                          reg614 : (reg793[(4'h9):(4'h9)] ?
                              forvar798[(4'ha):(4'h8)] : (forvar862 > reg854))));
                      reg932 <= reg757;
                      reg933 <= (&$unsigned((reg739[(2'h2):(1'h1)] ?
                          (+forvar922) : $signed(forvar763))));
                    end
                  if (reg596[(3'h4):(2'h3)])
                    begin
                      reg934 <= $unsigned((forvar722[(1'h1):(1'h1)] || ($signed(reg843) << $signed(reg897))));
                      reg935 <= ((^~reg842) ?
                          (~&((reg815 ? reg649 : (8'h9d)) ?
                              ((8'hb5) ?
                                  reg761 : reg724) : ((8'ha2) > forvar655))) : $signed(($unsigned(reg764) | $unsigned(forvar863))));
                      reg936 <= ($signed($signed((reg845 ?
                              (8'ha3) : forvar620))) ?
                          reg708[(2'h3):(2'h3)] : reg890);
                      reg937 <= ($signed($signed(forvar925[(2'h2):(1'h0)])) ?
                          $unsigned((reg900[(1'h1):(1'h1)] > $unsigned(reg757))) : $unsigned(reg695[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg934 <= $signed((^~(!reg785[(3'h4):(1'h1)])));
                      reg935 <= $signed(($signed((&forvar629)) ?
                          {{forvar595}} : $unsigned(((8'hb3) ?
                              reg721 : (8'hb0)))));
                      reg936 <= reg745[(3'h5):(3'h5)];
                    end
                  if ({(!($signed(reg876) ?
                          (forvar562 ? reg806 : reg669) : $signed(reg867)))})
                    begin
                      reg938 <= forvar660;
                      reg939 <= ((~|$signed($unsigned((8'hb9)))) && $unsigned((forvar595 && reg624[(4'h8):(3'h5)])));
                      reg940 <= $unsigned($signed($unsigned((reg874 ?
                          reg899 : reg684))));
                    end
                  else
                    begin
                      reg938 <= (($unsigned($unsigned(reg747)) ?
                          $unsigned(reg761) : (8'haf)) >> $unsigned($signed($signed(reg822))));
                      reg939 <= reg841[(3'h4):(1'h1)];
                    end
                end
              reg941 <= {reg581};
              if ($unsigned(reg636))
                begin
                  for (forvar942 = (1'h0); (forvar942 < (2'h2)); forvar942 = (forvar942 + (1'h1)))
                    begin
                      reg943 <= reg710[(1'h0):(1'h0)];
                      reg944 <= $unsigned(((^~{forvar759}) ?
                          (reg885 || $signed(forvar872)) : $signed($signed(forvar770))));
                    end
                  for (forvar945 = (1'h0); (forvar945 < (2'h2)); forvar945 = (forvar945 + (1'h1)))
                    begin
                      reg946 <= forvar600;
                      reg947 <= forvar851[(1'h1):(1'h1)];
                    end
                  if (wire560)
                    begin
                      reg948 <= (reg882[(3'h7):(2'h2)] != $unsigned(((reg884 ?
                              (8'h9e) : forvar834) ?
                          forvar872 : (reg841 ? reg714 : forvar756))));
                      reg949 <= (+$signed(reg844[(3'h4):(1'h1)]));
                      reg950 <= $signed($signed($signed({reg611})));
                    end
                  else
                    begin
                      reg948 <= $unsigned(forvar688);
                      reg949 <= (8'h9c);
                    end
                end
              else
                begin
                  reg942 <= (8'haf);
                end
              reg951 <= (|reg838);
            end
        end
      else
        begin
          for (forvar883 = (1'h0); (forvar883 < (1'h0)); forvar883 = (forvar883 + (1'h1)))
            begin
              for (forvar884 = (1'h0); (forvar884 < (1'h1)); forvar884 = (forvar884 + (1'h1)))
                begin
                  for (forvar885 = (1'h0); (forvar885 < (1'h1)); forvar885 = (forvar885 + (1'h1)))
                    begin
                      reg886 <= $unsigned($unsigned((reg847[(3'h5):(3'h4)] ?
                          reg839 : reg746)));
                    end
                  reg887 <= ((~forvar927) & (reg567[(2'h3):(2'h3)] + reg889));
                  if (forvar945)
                    begin
                      reg888 <= (~&reg900[(4'ha):(3'h7)]);
                      reg889 <= reg804;
                      reg890 <= (~|$signed(reg941[(4'h9):(3'h7)]));
                      reg891 <= reg943[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg888 <= ($unsigned((~&{forvar806})) == {forvar865});
                      reg889 <= forvar787;
                    end
                end
            end
          if ((({(reg714 < reg898)} && $signed($unsigned(forvar798))) ?
              reg766[(3'h5):(2'h3)] : (-(+(reg809 >= reg576)))))
            begin
              for (forvar892 = (1'h0); (forvar892 < (1'h1)); forvar892 = (forvar892 + (1'h1)))
                begin
                  for (forvar893 = (1'h0); (forvar893 < (1'h1)); forvar893 = (forvar893 + (1'h1)))
                    begin
                      reg894 <= ((8'h9d) ?
                          {reg765[(4'h9):(3'h5)]} : $unsigned(((reg704 ^~ reg618) != (!(8'ha6)))));
                      reg895 <= $signed(((forvar761 & forvar884) ?
                          reg571 : (reg946[(1'h1):(1'h1)] ?
                              $unsigned(reg809) : $signed((8'hba)))));
                      reg896 <= (reg897[(2'h3):(1'h1)] ?
                          $unsigned((^forvar742)) : (8'hb2));
                      reg897 <= reg850;
                    end
                  if ($unsigned((^reg716)))
                    begin
                      reg898 <= (reg655 == $signed({$signed(reg719)}));
                      reg899 <= reg901;
                      reg900 <= reg800;
                    end
                  else
                    begin
                      reg898 <= ($signed({{(8'ha9)}}) <<< reg680[(2'h3):(1'h1)]);
                      reg899 <= forvar589[(4'h8):(2'h2)];
                      reg900 <= (forvar853 - $unsigned(({(8'hba)} ?
                          $unsigned(reg700) : forvar867[(2'h3):(2'h3)])));
                    end
                end
              for (forvar901 = (1'h0); (forvar901 < (2'h2)); forvar901 = (forvar901 + (1'h1)))
                begin
                  for (forvar902 = (1'h0); (forvar902 < (2'h3)); forvar902 = (forvar902 + (1'h1)))
                    begin
                      reg903 <= (&($signed((-reg690)) & reg719));
                      reg904 <= $signed(reg762[(4'hb):(2'h3)]);
                      reg905 <= (reg884 ^ (-reg580));
                      reg906 <= reg891;
                    end
                  if ($signed(forvar649[(2'h3):(1'h0)]))
                    begin
                      reg907 <= (!$unsigned(($unsigned(reg732) ?
                          reg777[(1'h1):(1'h0)] : reg678[(2'h2):(1'h1)])));
                      reg908 <= (((!$signed(reg619)) ?
                          (8'hb7) : forvar832) <<< (reg590[(2'h2):(2'h2)] >> $unsigned((reg695 ?
                          reg693 : reg653))));
                      reg909 <= {(((forvar702 ? forvar660 : (8'hab)) ?
                                  $unsigned(reg788) : (8'ha4)) ?
                              $signed(((8'ha0) ^ reg816)) : {reg644})};
                      reg910 <= reg813[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg907 <= $unsigned($signed(((-(8'ha3)) >> ((8'ha3) ?
                          (8'ha7) : reg897))));
                      reg908 <= (~reg739[(1'h0):(1'h0)]);
                      reg909 <= (8'hab);
                    end
                  for (forvar911 = (1'h0); (forvar911 < (2'h3)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= (reg599 ? (8'ha8) : (~&reg720[(1'h1):(1'h1)]));
                      reg913 <= (~^((&forvar647) != ($unsigned(reg762) ?
                          $signed((8'hb4)) : (forvar756 ?
                              forvar819 : reg851))));
                      reg914 <= (!forvar733);
                    end
                  if (($unsigned($signed(reg674)) >= ((forvar669[(3'h5):(2'h2)] ?
                      reg762[(2'h2):(1'h0)] : $signed(reg786)) - forvar778)))
                    begin
                      reg915 <= (($signed($signed(reg870)) ?
                          ($signed(forvar901) ?
                              forvar759[(4'hc):(4'hb)] : reg941) : (^~(8'ha9))) && $unsigned($unsigned($signed(forvar562))));
                      reg916 <= (forvar668[(2'h3):(1'h0)] * (^~$signed($signed(forvar722))));
                    end
                  else
                    begin
                      reg915 <= (forvar652 < (~&(forvar790[(3'h4):(1'h1)] && (~^reg644))));
                      reg916 <= ($unsigned(reg565) >= (|{$signed(reg693)}));
                      reg917 <= reg702;
                      reg918 <= $signed((((reg712 && reg679) > reg644[(3'h4):(1'h1)]) > ((~|forvar687) ?
                          (forvar859 >= (8'ha6)) : $unsigned(reg718))));
                    end
                end
              if (reg939[(1'h1):(1'h1)])
                begin
                  for (forvar919 = (1'h0); (forvar919 < (1'h0)); forvar919 = (forvar919 + (1'h1)))
                    begin
                      reg920 <= (reg567[(2'h3):(1'h0)] ~^ forvar844);
                      reg921 <= $unsigned(reg944);
                      reg922 <= $unsigned((({reg863} ? reg827 : reg678) ?
                          {$unsigned(reg828)} : (8'ha6)));
                    end
                  reg923 <= (~&($unsigned($signed(reg567)) ?
                      reg622[(1'h0):(1'h0)] : $signed((&reg851))));
                  for (forvar924 = (1'h0); (forvar924 < (2'h3)); forvar924 = (forvar924 + (1'h1)))
                    begin
                      reg925 <= ((forvar722[(1'h1):(1'h0)] ?
                              ((+(8'ha5)) ?
                                  forvar871 : (reg872 ?
                                      forvar897 : (8'ha5))) : (~|$signed(reg895))) ?
                          (!reg888[(4'hc):(3'h5)]) : (|reg805[(1'h1):(1'h1)]));
                      reg926 <= ($unsigned($signed({reg668})) >= $unsigned(((reg779 && reg876) >= reg634[(4'h8):(2'h2)])));
                    end
                end
              else
                begin
                  if (reg712[(5'h10):(4'ha)])
                    begin
                      reg919 <= (($signed($unsigned(reg807)) ?
                              {$signed(reg855)} : (reg858[(2'h2):(1'h1)] > (reg650 ?
                                  reg923 : reg695))) ?
                          ($signed((reg698 ? reg580 : reg643)) ?
                              $signed({reg843}) : (~^reg807[(4'h9):(4'h9)])) : $signed($signed($unsigned(forvar564))));
                      reg920 <= $unsigned($unsigned(($signed(forvar562) <= $signed(forvar881))));
                      reg921 <= ((+forvar811) << ($signed(reg732) ?
                          reg845[(2'h3):(1'h0)] : ((reg930 ?
                                  forvar922 : reg830) ?
                              (-reg693) : (reg646 >> reg914))));
                      reg922 <= ($signed($unsigned((~&forvar620))) ?
                          reg624 : ($signed((reg735 || forvar844)) + (8'ha8)));
                    end
                  else
                    begin
                      reg919 <= (~|(|((|reg565) ~^ reg853[(2'h3):(1'h0)])));
                    end
                  if (reg602[(2'h2):(1'h1)])
                    begin
                      reg923 <= {(8'hb9)};
                    end
                  else
                    begin
                      reg923 <= forvar836;
                      reg924 <= (&(({reg886} ? $unsigned((8'ha1)) : {reg701}) ?
                          $unsigned(forvar664[(1'h0):(1'h0)]) : $unsigned($signed((8'ha1)))));
                      reg925 <= {(~^$unsigned($signed(reg947)))};
                      reg926 <= reg653;
                    end
                  for (forvar927 = (1'h0); (forvar927 < (1'h1)); forvar927 = (forvar927 + (1'h1)))
                    begin
                      reg928 <= (~$signed(forvar770[(2'h2):(2'h2)]));
                      reg929 <= {((forvar862[(2'h2):(2'h2)] ?
                                  (~|(8'ha7)) : $unsigned((8'h9e))) ?
                              $unsigned((reg849 ?
                                  reg717 : reg863)) : forvar814)};
                      reg930 <= reg873[(3'h4):(2'h2)];
                    end
                end
              if ((~^$unsigned(((reg752 <= forvar699) ?
                  (forvar659 ? reg781 : forvar783) : reg617))))
                begin
                  reg931 <= (+$unsigned((reg795[(3'h7):(1'h1)] && {reg922})));
                end
              else
                begin
                  for (forvar931 = (1'h0); (forvar931 < (2'h3)); forvar931 = (forvar931 + (1'h1)))
                    begin
                      reg932 <= (({(reg704 ?
                              forvar737 : reg632)} >> ($signed(reg676) ?
                          reg598[(3'h6):(2'h2)] : (^~reg707))) >> (forvar699 - forvar602[(1'h0):(1'h0)]));
                      reg933 <= forvar659;
                      reg934 <= (forvar620[(2'h3):(2'h2)] & reg948);
                      reg935 <= $unsigned(((forvar570[(4'ha):(3'h5)] ?
                              $unsigned(reg916) : (^~forvar629)) ?
                          forvar733 : $unsigned(forvar681[(3'h6):(3'h4)])));
                    end
                end
            end
          else
            begin
              if ({($signed(reg896) ?
                      ((&reg617) ?
                          (^~reg603) : $signed(forvar844)) : ($unsigned(reg609) - {forvar829}))})
                begin
                  reg892 <= reg923[(1'h1):(1'h1)];
                  for (forvar893 = (1'h0); (forvar893 < (2'h3)); forvar893 = (forvar893 + (1'h1)))
                    begin
                      reg894 <= reg757[(4'ha):(3'h7)];
                      reg895 <= reg779[(4'hb):(2'h3)];
                      reg896 <= $signed($signed(reg951));
                      reg897 <= forvar770;
                    end
                  if ((reg908[(1'h0):(1'h0)] ~^ reg935[(1'h1):(1'h0)]))
                    begin
                      reg898 <= (~|reg576);
                      reg899 <= $unsigned($signed(forvar589));
                      reg900 <= ({$unsigned($unsigned(reg593))} && ($signed((reg940 == forvar745)) ?
                          ((~reg669) + (reg635 <= forvar588)) : (reg578 && $signed(reg833))));
                    end
                  else
                    begin
                      reg898 <= ($unsigned({$unsigned((8'haa))}) <<< reg578[(3'h7):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar892 = (1'h0); (forvar892 < (1'h0)); forvar892 = (forvar892 + (1'h1)))
                    begin
                      reg893 <= forvar884;
                      reg894 <= reg727;
                      reg895 <= reg677[(1'h1):(1'h1)];
                    end
                  if ($unsigned(({reg916} ?
                      ((^reg941) ? ((8'hb7) ^ (8'hae)) : reg568) : (^~((8'hb6) ?
                          forvar853 : reg747)))))
                    begin
                      reg896 <= (8'hb6);
                      reg897 <= $signed(({reg899} ?
                          $signed((reg769 >> reg923)) : (^(reg684 <<< forvar831))));
                      reg898 <= ((~&($signed(wire558) ?
                              ((8'ha8) || (8'hb2)) : (&forvar894))) ?
                          reg706[(4'hc):(1'h1)] : $signed(reg592));
                      reg899 <= (+(8'hb4));
                    end
                  else
                    begin
                      reg896 <= (|(-$signed({reg743})));
                    end
                  for (forvar900 = (1'h0); (forvar900 < (1'h1)); forvar900 = (forvar900 + (1'h1)))
                    begin
                      reg901 <= {reg791[(3'h7):(3'h4)]};
                      reg902 <= $unsigned(forvar644[(4'hc):(3'h7)]);
                      reg903 <= ({reg719[(2'h3):(2'h3)]} <= reg891);
                      reg904 <= reg794;
                    end
                end
            end
          reg936 <= $signed((^((^~reg871) < reg852[(3'h6):(1'h0)])));
        end
      if (forvar644)
        begin
          for (forvar952 = (1'h0); (forvar952 < (1'h0)); forvar952 = (forvar952 + (1'h1)))
            begin
              for (forvar953 = (1'h0); (forvar953 < (2'h2)); forvar953 = (forvar953 + (1'h1)))
                begin
                  for (forvar954 = (1'h0); (forvar954 < (2'h3)); forvar954 = (forvar954 + (1'h1)))
                    begin
                      reg955 <= ({$unsigned($unsigned(forvar787))} * reg840[(1'h1):(1'h1)]);
                    end
                  for (forvar956 = (1'h0); (forvar956 < (2'h3)); forvar956 = (forvar956 + (1'h1)))
                    begin
                      reg957 <= $unsigned($signed(forvar655[(1'h0):(1'h0)]));
                      reg958 <= reg797[(1'h0):(1'h0)];
                    end
                end
              reg959 <= (reg891 ?
                  ((8'hab) ?
                      forvar668 : ((~&reg662) && (reg643 ?
                          forvar573 : forvar588))) : $unsigned(reg754));
              if ($signed(($unsigned($signed(reg665)) ?
                  {$unsigned((8'ha2))} : reg728[(3'h7):(3'h6)])))
                begin
                  reg960 <= (reg653[(3'h6):(3'h6)] ?
                      (+$unsigned(reg801[(4'ha):(4'h9)])) : {$signed($unsigned(reg709))});
                end
              else
                begin
                  for (forvar960 = (1'h0); (forvar960 < (1'h1)); forvar960 = (forvar960 + (1'h1)))
                    begin
                      reg961 <= {reg838};
                    end
                  for (forvar962 = (1'h0); (forvar962 < (2'h3)); forvar962 = (forvar962 + (1'h1)))
                    begin
                      reg963 <= $signed($unsigned(({(8'ha3)} ?
                          (8'hb3) : $unsigned((8'ha8)))));
                      reg964 <= (reg788[(2'h3):(2'h3)] >> (($signed(forvar707) && reg642[(4'h9):(3'h7)]) & reg661));
                    end
                  for (forvar965 = (1'h0); (forvar965 < (1'h0)); forvar965 = (forvar965 + (1'h1)))
                    begin
                      reg966 <= $unsigned($unsigned((+forvar806[(1'h1):(1'h1)])));
                      reg967 <= $signed(forvar814);
                    end
                end
              reg968 <= ((&reg909) ? forvar784 : reg912);
            end
          if ((~|($signed(reg943) * reg678[(1'h1):(1'h0)])))
            begin
              for (forvar969 = (1'h0); (forvar969 < (1'h0)); forvar969 = (forvar969 + (1'h1)))
                begin
                  reg970 <= (~^forvar892);
                  for (forvar971 = (1'h0); (forvar971 < (2'h2)); forvar971 = (forvar971 + (1'h1)))
                    begin
                      reg972 <= ($unsigned(($unsigned(reg708) ?
                              (+reg762) : (reg731 ? reg861 : reg591))) ?
                          forvar853[(3'h4):(1'h1)] : $signed(($signed(reg855) <= (reg742 ?
                              reg619 : forvar681))));
                      reg973 <= reg767;
                      reg974 <= ((&((~&(8'hb6)) ^~ (|forvar648))) ?
                          wire555 : (|$signed(reg890[(3'h4):(2'h2)])));
                    end
                  for (forvar975 = (1'h0); (forvar975 < (2'h3)); forvar975 = (forvar975 + (1'h1)))
                    begin
                      reg976 <= (reg874[(3'h5):(3'h5)] == (8'hb6));
                      reg977 <= $signed($unsigned(reg964[(1'h0):(1'h0)]));
                      reg978 <= ({reg833} ^ ({(reg878 | (8'ha7))} >> $unsigned({reg808})));
                      reg979 <= forvar853[(2'h2):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar969 = (1'h0); (forvar969 < (1'h1)); forvar969 = (forvar969 + (1'h1)))
                begin
                  reg970 <= (reg645[(3'h5):(2'h2)] + (&(~^(~^forvar962))));
                  reg971 <= {$unsigned({(+forvar659)})};
                end
              if (reg663[(4'ha):(2'h2)])
                begin
                  if ((reg780[(1'h0):(1'h0)] ?
                      ($signed((reg748 ?
                          forvar600 : (8'hb3))) ~^ $unsigned(reg928)) : (forvar922[(2'h2):(1'h1)] * $signed($signed((8'ha3))))))
                    begin
                      reg972 <= $unsigned(reg802[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg972 <= {reg941[(4'ha):(3'h7)]};
                      reg973 <= (~^(($unsigned(reg747) + (-reg802)) ^~ {(~|reg905)}));
                    end
                  if ((^forvar911[(3'h7):(3'h7)]))
                    begin
                      reg974 <= ($signed(((forvar895 && forvar895) ?
                              (8'ha4) : reg616)) ?
                          ((reg779 ^ (reg750 ? forvar778 : (8'haf))) ?
                              (reg566[(4'h8):(3'h5)] ?
                                  forvar659[(3'h5):(3'h4)] : ((8'hba) ?
                                      reg628 : forvar866)) : $unsigned(reg616[(4'h8):(3'h5)])) : ($signed($signed((8'ha6))) ?
                              (|(reg755 ?
                                  reg815 : reg793)) : forvar722[(2'h2):(2'h2)]));
                      reg975 <= $signed(($unsigned(reg593[(3'h4):(1'h1)]) ?
                          (|$unsigned(reg593)) : (forvar889[(1'h1):(1'h0)] && $signed(reg590))));
                      reg976 <= ((&(~(reg601 && reg828))) ?
                          $unsigned({(reg838 >> reg744)}) : $unsigned((~$signed((8'ha8)))));
                      reg977 <= (&forvar630);
                    end
                  else
                    begin
                      reg974 <= (reg759 < $unsigned(((reg850 ?
                          forvar571 : reg795) == (reg834 ?
                          reg816 : forvar840))));
                      reg975 <= ($unsigned((~^((8'hab) ? reg821 : forvar615))) ?
                          (reg763 ?
                              ((reg756 ?
                                  (8'haa) : reg796) + {(8'ha3)}) : ((reg769 >> forvar870) || $unsigned(reg671))) : $signed($unsigned($signed(forvar942))));
                      reg976 <= $signed($unsigned((~&$unsigned(reg871))));
                      reg977 <= $signed(((~{reg632}) & ($signed((8'ha2)) || reg747[(2'h3):(2'h3)])));
                    end
                  if ({forvar865[(2'h3):(1'h1)]})
                    begin
                      reg978 <= (reg698[(2'h2):(1'h1)] && (^$unsigned((^~reg571))));
                    end
                  else
                    begin
                      reg978 <= {$unsigned($signed({reg757}))};
                      reg979 <= $unsigned($unsigned({(!reg750)}));
                    end
                end
              else
                begin
                  reg972 <= (-($signed($signed(reg749)) <= reg688[(1'h0):(1'h0)]));
                end
              if (((^~(8'hb3)) - {$signed((8'hae))}))
                begin
                  if ({reg892})
                    begin
                      reg980 <= reg565;
                      reg981 <= (($signed(forvar615) >> ((!reg599) << reg794)) ?
                          (reg738[(4'ha):(2'h2)] <= $unsigned({forvar644})) : (~$signed(reg857[(3'h7):(1'h1)])));
                      reg982 <= {forvar836[(1'h0):(1'h0)]};
                      reg983 <= $unsigned($signed(((reg858 ?
                          reg715 : forvar656) << $unsigned(forvar595))));
                    end
                  else
                    begin
                      reg980 <= reg658[(2'h2):(1'h1)];
                      reg981 <= {(reg591[(3'h4):(3'h4)] ?
                              {reg591} : $signed(reg884[(1'h0):(1'h0)]))};
                    end
                end
              else
                begin
                  for (forvar980 = (1'h0); (forvar980 < (2'h3)); forvar980 = (forvar980 + (1'h1)))
                    begin
                      reg981 <= (forvar629[(3'h5):(1'h0)] <= ($unsigned((~&reg875)) ?
                          ($unsigned(reg567) ~^ forvar591) : forvar648[(3'h6):(1'h1)]));
                      reg982 <= $signed(($signed((!forvar562)) ~^ $signed(reg596)));
                      reg983 <= (~&(~&forvar870[(1'h1):(1'h0)]));
                    end
                  if ($signed($signed(((~|forvar962) >= $unsigned(forvar620)))))
                    begin
                      reg984 <= (forvar870 >= reg728);
                      reg985 <= {forvar861[(2'h2):(1'h1)]};
                      reg986 <= $signed($signed(reg734[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg984 <= reg897[(2'h2):(1'h0)];
                      reg985 <= (~^(!$signed({forvar900})));
                    end
                  for (forvar987 = (1'h0); (forvar987 < (2'h3)); forvar987 = (forvar987 + (1'h1)))
                    begin
                      reg988 <= $signed(forvar962[(3'h7):(2'h3)]);
                      reg989 <= ({{(~&reg928)}} ?
                          ((~(forvar704 ?
                              forvar840 : reg655)) == ($signed(forvar922) ?
                              (reg677 ?
                                  forvar926 : forvar828) : {forvar844})) : {(reg628[(4'ha):(2'h3)] ?
                                  forvar695 : reg802[(3'h4):(1'h1)])});
                      reg990 <= (!reg943);
                    end
                  for (forvar991 = (1'h0); (forvar991 < (2'h3)); forvar991 = (forvar991 + (1'h1)))
                    begin
                      reg992 <= $signed(((~&(reg716 ? forvar643 : (8'hb0))) ?
                          reg829 : ((+forvar713) == $signed((8'h9f)))));
                      reg993 <= $unsigned((({reg695} & (+forvar656)) ?
                          $unsigned(reg655[(3'h6):(2'h3)]) : (~{forvar676})));
                      reg994 <= reg873[(3'h4):(2'h3)];
                      reg995 <= {({reg760[(4'hc):(3'h4)]} + ((~reg929) ?
                              forvar571[(1'h1):(1'h0)] : $unsigned(reg863)))};
                    end
                end
            end
          for (forvar996 = (1'h0); (forvar996 < (1'h0)); forvar996 = (forvar996 + (1'h1)))
            begin
              for (forvar997 = (1'h0); (forvar997 < (2'h2)); forvar997 = (forvar997 + (1'h1)))
                begin
                  for (forvar998 = (1'h0); (forvar998 < (1'h0)); forvar998 = (forvar998 + (1'h1)))
                    begin
                      reg999 <= $unsigned(($signed((reg796 > reg898)) ?
                          $signed((forvar676 < reg603)) : reg590[(2'h3):(2'h2)]));
                      reg1000 <= ($unsigned(reg751[(3'h7):(1'h0)]) << (forvar621[(3'h7):(3'h6)] ?
                          $signed($signed(reg738)) : reg706[(3'h5):(3'h4)]));
                    end
                  reg1001 <= (reg743[(3'h7):(1'h0)] ?
                      (^((reg792 ?
                          reg834 : (8'ha6)) <= (^~forvar722))) : ((8'hac) || $signed({reg747})));
                end
              for (forvar1002 = (1'h0); (forvar1002 < (1'h1)); forvar1002 = (forvar1002 + (1'h1)))
                begin
                  for (forvar1003 = (1'h0); (forvar1003 < (2'h2)); forvar1003 = (forvar1003 + (1'h1)))
                    begin
                      reg1004 <= (reg801[(3'h4):(3'h4)] ?
                          reg785[(4'h8):(3'h6)] : $unsigned(((|forvar713) <= reg825[(3'h4):(2'h2)])));
                    end
                end
              for (forvar1005 = (1'h0); (forvar1005 < (2'h3)); forvar1005 = (forvar1005 + (1'h1)))
                begin
                  if ((~^$unsigned($unsigned($unsigned((8'hb1))))))
                    begin
                      reg1006 <= (^~($unsigned((reg904 | (8'ha6))) >= reg871[(4'hd):(1'h0)]));
                      reg1007 <= $unsigned($unsigned($signed((reg749 != reg890))));
                      reg1008 <= reg599;
                      reg1009 <= reg636[(3'h7):(2'h3)];
                    end
                  else
                    begin
                      reg1006 <= ($unsigned((^{reg803})) ^~ $unsigned(reg823[(3'h7):(3'h5)]));
                      reg1007 <= ($unsigned($signed((~&reg866))) ?
                          $unsigned($unsigned($unsigned(forvar844))) : $unsigned($signed((reg856 != reg856))));
                    end
                  if ((($signed((8'hb6)) ? reg982 : reg575[(3'h5):(1'h1)]) ?
                      reg568[(3'h7):(3'h5)] : (^reg929[(3'h4):(1'h0)])))
                    begin
                      reg1010 <= $signed(reg691);
                      reg1011 <= $unsigned((~|$unsigned((reg593 ?
                          reg568 : forvar655))));
                    end
                  else
                    begin
                      reg1010 <= (+(~|reg917[(4'ha):(2'h3)]));
                      reg1011 <= reg872[(3'h6):(2'h3)];
                      reg1012 <= reg601[(1'h0):(1'h0)];
                    end
                  for (forvar1013 = (1'h0); (forvar1013 < (2'h3)); forvar1013 = (forvar1013 + (1'h1)))
                    begin
                      reg1014 <= $signed($signed(((-reg642) ^~ (!(8'hba)))));
                      reg1015 <= (($unsigned($signed((8'ha4))) <= $signed((-reg892))) ?
                          reg693 : (reg958[(4'h8):(4'h8)] || (^~(reg806 ?
                              reg815 : reg772))));
                      reg1016 <= {{{forvar901}}};
                      reg1017 <= reg1007[(3'h5):(2'h3)];
                    end
                  reg1018 <= (~|(($signed(reg593) ?
                      (reg988 ~^ reg648) : reg864) > reg872));
                end
              reg1019 <= ((~^({reg940} ?
                  {reg951} : forvar871[(3'h5):(3'h5)])) ^~ reg940[(1'h1):(1'h1)]);
            end
        end
      else
        begin
          reg952 <= $signed({(!(forvar674 ? reg901 : reg569))});
          if (($signed(forvar761[(4'h9):(2'h2)]) ?
              {$signed(forvar631[(1'h0):(1'h0)])} : (^~$unsigned($unsigned(reg613)))))
            begin
              for (forvar953 = (1'h0); (forvar953 < (1'h1)); forvar953 = (forvar953 + (1'h1)))
                begin
                  reg954 <= $signed($signed(reg938[(1'h1):(1'h0)]));
                  for (forvar955 = (1'h0); (forvar955 < (1'h0)); forvar955 = (forvar955 + (1'h1)))
                    begin
                      reg956 <= (forvar925 >= ({(reg799 >= reg689)} <<< (reg995 << (|forvar668))));
                    end
                end
            end
          else
            begin
              for (forvar953 = (1'h0); (forvar953 < (2'h2)); forvar953 = (forvar953 + (1'h1)))
                begin
                  for (forvar954 = (1'h0); (forvar954 < (1'h0)); forvar954 = (forvar954 + (1'h1)))
                    begin
                      reg955 <= {({{reg567}} <= reg990[(3'h7):(2'h2)])};
                      reg956 <= $unsigned((((+forvar955) ?
                              (forvar608 ?
                                  (8'ha0) : reg903) : $unsigned((8'hb6))) ?
                          $signed($unsigned(forvar699)) : {$signed(reg586)}));
                      reg957 <= (reg926[(3'h4):(1'h0)] ?
                          ({forvar843[(3'h5):(2'h2)]} ?
                              {reg598} : ($unsigned(reg577) ?
                                  (~&(8'hb5)) : $unsigned(reg843))) : reg786);
                    end
                  if (($unsigned((8'ha3)) && reg955[(4'h8):(3'h5)]))
                    begin
                      reg958 <= (|reg980[(4'h9):(3'h7)]);
                      reg959 <= forvar669[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg958 <= reg619;
                    end
                end
              reg960 <= ((&((8'hba) || (!reg644))) <= {reg882});
              if ($signed((^~$signed(forvar900[(3'h7):(3'h6)]))))
                begin
                  if (reg698[(3'h5):(1'h1)])
                    begin
                      reg961 <= $unsigned(reg947[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg961 <= (&(8'h9d));
                      reg962 <= reg858[(4'h9):(4'h9)];
                    end
                  for (forvar963 = (1'h0); (forvar963 < (1'h0)); forvar963 = (forvar963 + (1'h1)))
                    begin
                      reg964 <= $signed(reg956[(4'h9):(3'h6)]);
                    end
                  for (forvar965 = (1'h0); (forvar965 < (2'h2)); forvar965 = (forvar965 + (1'h1)))
                    begin
                      reg966 <= (+$unsigned({(reg563 ? (8'h9e) : reg590)}));
                    end
                  if (((8'h9e) ?
                      $unsigned({reg802}) : forvar656[(5'h10):(4'hc)]))
                    begin
                      reg967 <= $signed(((8'ha2) ?
                          $signed((reg823 ? (8'hb3) : forvar600)) : ({(8'ha1)} ?
                              reg627 : (forvar798 ? forvar655 : reg740))));
                      reg968 <= $unsigned(($unsigned((8'hb3)) ?
                          (forvar960 << forvar756[(1'h1):(1'h1)]) : (!$signed(forvar901))));
                      reg969 <= reg1001;
                    end
                  else
                    begin
                      reg967 <= (forvar907[(4'h9):(4'h8)] ?
                          $signed(reg614[(1'h0):(1'h0)]) : (forvar649[(2'h3):(1'h0)] <<< $signed((reg852 * (8'ha0)))));
                      reg968 <= (reg916[(1'h0):(1'h0)] ?
                          $unsigned(($signed(reg587) & $signed(reg660))) : $signed(reg839));
                      reg969 <= reg567;
                      reg970 <= $signed((^$signed(forvar664)));
                    end
                end
              else
                begin
                  for (forvar961 = (1'h0); (forvar961 < (1'h1)); forvar961 = (forvar961 + (1'h1)))
                    begin
                      reg962 <= (~|$unsigned({$signed(reg895)}));
                    end
                  if (forvar664)
                    begin
                      reg963 <= ($unsigned(reg832[(4'hb):(4'ha)]) >>> forvar859[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg963 <= ((^~$signed((reg827 ?
                          forvar620 : reg692))) & ((8'hae) | (!(^~reg624))));
                    end
                end
            end
        end
    end
  assign wire1020 = (!$signed({(-reg788)}));
  module1021 modinst5525 (.clk(clk), .y(wire5524), .wire1025(reg796), .wire1024(reg820), .wire1023(reg929), .wire1022(forvar881));
  assign wire5526 = (!$unsigned($signed($signed(forvar702))));
  assign wire5527 = (~^$signed(((reg693 != forvar996) > $unsigned(reg744))));
  assign wire5528 = reg918[(4'hd):(2'h3)];
  assign wire5529 = forvar745[(3'h4):(1'h0)];
  assign wire5530 = ($signed((forvar866[(3'h5):(1'h0)] || $signed((8'ha6)))) ?
                        reg594 : forvar844[(3'h5):(1'h0)]);
  assign wire5531 = {((!(^reg862)) || forvar920)};
  always
    @(posedge clk) begin
      for (forvar5532 = (1'h0); (forvar5532 < (1'h0)); forvar5532 = (forvar5532 + (1'h1)))
        begin
          if ($unsigned(reg840))
            begin
              reg5533 <= $unsigned((^(~(reg1018 ? reg923 : reg867))));
            end
          else
            begin
              if (reg707[(2'h2):(1'h0)])
                begin
                  for (forvar5533 = (1'h0); (forvar5533 < (1'h1)); forvar5533 = (forvar5533 + (1'h1)))
                    begin
                      reg5534 <= $unsigned($unsigned($unsigned((&(8'hb1)))));
                    end
                end
              else
                begin
                  for (forvar5533 = (1'h0); (forvar5533 < (2'h3)); forvar5533 = (forvar5533 + (1'h1)))
                    begin
                      reg5534 <= forvar592[(1'h1):(1'h0)];
                      reg5535 <= (forvar641[(4'ha):(3'h4)] ?
                          {(~^$unsigned(reg946))} : $signed((forvar704 ?
                              (~^wire5531) : (reg740 << reg835))));
                    end
                  if ((|forvar695))
                    begin
                      reg5536 <= reg586;
                      reg5537 <= (+$signed((reg889[(2'h3):(1'h0)] - $signed(reg5533))));
                      reg5538 <= $signed($signed(reg660[(2'h3):(2'h2)]));
                      reg5539 <= ($signed(((~(8'h9c)) == (reg887 ?
                              reg1004 : forvar733))) ?
                          (&(forvar742[(3'h5):(2'h2)] ?
                              $unsigned(reg831) : {reg679})) : $signed(forvar759[(4'he):(4'hd)]));
                    end
                  else
                    begin
                      reg5536 <= forvar711;
                    end
                end
              for (forvar5540 = (1'h0); (forvar5540 < (2'h3)); forvar5540 = (forvar5540 + (1'h1)))
                begin
                  for (forvar5541 = (1'h0); (forvar5541 < (1'h1)); forvar5541 = (forvar5541 + (1'h1)))
                    begin
                      reg5542 <= (reg973[(2'h3):(2'h2)] >= $unsigned(($unsigned(reg597) << $signed(forvar676))));
                      reg5543 <= reg677;
                      reg5544 <= $unsigned($unsigned((reg937[(1'h1):(1'h1)] ?
                          (|reg756) : (reg780 ? reg837 : wire559))));
                    end
                  reg5545 <= ($signed($unsigned((reg759 | forvar741))) ?
                      (+reg896) : forvar5540);
                  if ((!reg873))
                    begin
                      reg5546 <= (reg877 != reg940);
                      reg5547 <= (((|{reg576}) ?
                          $signed(forvar811[(3'h4):(1'h1)]) : (reg833 - $unsigned(reg611))) > forvar584);
                      reg5548 <= reg956;
                      reg5549 <= $unsigned((((reg707 ? reg969 : forvar922) ?
                              reg692 : reg854[(1'h1):(1'h0)]) ?
                          forvar836 : (forvar831 ?
                              $signed(forvar741) : (reg985 >= reg650))));
                    end
                  else
                    begin
                      reg5546 <= (~&(~$unsigned((8'h9f))));
                    end
                  for (forvar5550 = (1'h0); (forvar5550 < (1'h1)); forvar5550 = (forvar5550 + (1'h1)))
                    begin
                      reg5551 <= ((^({reg914} || reg838[(4'hb):(1'h0)])) || (reg5533 >= forvar832));
                      reg5552 <= {({(-reg902)} ?
                              reg867[(3'h5):(1'h1)] : wire558)};
                    end
                end
              for (forvar5553 = (1'h0); (forvar5553 < (1'h1)); forvar5553 = (forvar5553 + (1'h1)))
                begin
                  reg5554 <= $signed(forvar962);
                end
            end
          for (forvar5555 = (1'h0); (forvar5555 < (2'h2)); forvar5555 = (forvar5555 + (1'h1)))
            begin
              reg5556 <= (&{{(wire560 ? reg658 : reg679)}});
            end
          if ((forvar906[(2'h3):(1'h0)] << $signed($unsigned(forvar745[(1'h1):(1'h0)]))))
            begin
              for (forvar5557 = (1'h0); (forvar5557 < (2'h3)); forvar5557 = (forvar5557 + (1'h1)))
                begin
                  if ($unsigned(reg596[(3'h7):(3'h4)]))
                    begin
                      reg5558 <= $signed({(8'hb3)});
                      reg5559 <= (reg862 ^~ $unsigned(((^(8'hb6)) ?
                          $signed(reg622) : reg645)));
                      reg5560 <= {{$unsigned((reg922 & forvar814))}};
                    end
                  else
                    begin
                      reg5558 <= reg704[(4'h8):(1'h0)];
                      reg5559 <= ((((8'ha2) != (reg967 && wire556)) != reg567[(1'h0):(1'h0)]) ?
                          (!(&reg728)) : $unsigned(wire558));
                    end
                  for (forvar5561 = (1'h0); (forvar5561 < (1'h1)); forvar5561 = (forvar5561 + (1'h1)))
                    begin
                      reg5562 <= forvar886[(3'h7):(3'h4)];
                      reg5563 <= ((!($signed(forvar952) | $signed((8'hab)))) > forvar955);
                    end
                  if ($unsigned(reg781[(2'h2):(2'h2)]))
                    begin
                      reg5564 <= ($signed((reg890[(3'h7):(3'h5)] ?
                          $signed(reg840) : $unsigned(reg900))) * ($signed({reg683}) ?
                          $signed((reg779 ?
                              reg769 : reg647)) : $unsigned($signed(forvar998))));
                      reg5565 <= {$signed(reg916)};
                    end
                  else
                    begin
                      reg5564 <= reg906;
                      reg5565 <= $signed(((!reg923[(3'h4):(1'h0)]) ?
                          ((-reg659) ?
                              $unsigned(reg985) : {reg725}) : (8'ha0)));
                      reg5566 <= $unsigned($unsigned($signed((reg598 ?
                          (8'ha9) : forvar759))));
                    end
                end
            end
          else
            begin
              if (reg614[(3'h7):(3'h4)])
                begin
                  for (forvar5557 = (1'h0); (forvar5557 < (1'h0)); forvar5557 = (forvar5557 + (1'h1)))
                    begin
                      reg5558 <= wire559[(3'h4):(1'h1)];
                    end
                  for (forvar5559 = (1'h0); (forvar5559 < (1'h0)); forvar5559 = (forvar5559 + (1'h1)))
                    begin
                      reg5560 <= (forvar600 ?
                          forvar579[(1'h0):(1'h0)] : forvar952[(1'h0):(1'h0)]);
                      reg5561 <= (&($signed({reg738}) ^ ($unsigned(reg827) && (reg988 > reg835))));
                      reg5562 <= $signed($signed(($signed(forvar889) ?
                          (wire557 ? forvar589 : (8'hb5)) : (&reg812))));
                    end
                  if (forvar866[(4'hc):(2'h3)])
                    begin
                      reg5563 <= $unsigned(reg769[(3'h7):(1'h0)]);
                      reg5564 <= ($unsigned((wire558 >= (reg813 == reg624))) > reg990[(3'h7):(2'h3)]);
                    end
                  else
                    begin
                      reg5563 <= $signed((forvar5541 ?
                          {(forvar737 || reg5559)} : (+$signed(forvar775))));
                      reg5564 <= ((~^(forvar707 ?
                              (~|reg874) : $unsigned(reg951))) ?
                          reg724 : ($unsigned((8'ha7)) ?
                              $unsigned(forvar1013[(1'h0):(1'h0)]) : (reg861 ?
                                  (8'ha0) : (-reg802))));
                      reg5565 <= forvar567[(2'h2):(2'h2)];
                      reg5566 <= {reg594};
                    end
                end
              else
                begin
                  if ((^~{(~|(forvar5555 < reg758))}))
                    begin
                      reg5557 <= reg856[(1'h0):(1'h0)];
                      reg5558 <= $signed(forvar843);
                      reg5559 <= $signed(forvar907[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg5557 <= $unsigned(forvar980);
                    end
                  if ((&reg705))
                    begin
                      reg5560 <= $unsigned(reg986[(3'h7):(3'h4)]);
                      reg5561 <= reg959;
                      reg5562 <= ({$unsigned($unsigned(reg563))} > (($unsigned(reg921) ?
                              reg983 : reg741[(2'h2):(1'h0)]) ?
                          ((reg950 ?
                              (8'hb7) : reg5547) << (forvar5553 * (8'hb3))) : (+{reg873})));
                      reg5563 <= $signed($unsigned($unsigned(reg796[(3'h7):(1'h0)])));
                    end
                  else
                    begin
                      reg5560 <= (~|($signed($signed(reg762)) ?
                          ($unsigned(wire555) + (reg5548 <= reg893)) : {$signed(reg816)}));
                      reg5561 <= (((~^reg898) - reg934[(1'h0):(1'h0)]) >> ((&$unsigned((8'ha9))) ?
                          reg710 : $unsigned((+reg992))));
                    end
                  for (forvar5564 = (1'h0); (forvar5564 < (2'h3)); forvar5564 = (forvar5564 + (1'h1)))
                    begin
                      reg5565 <= reg817[(4'h8):(3'h6)];
                      reg5566 <= (~&reg820[(2'h3):(1'h1)]);
                      reg5567 <= ((reg5561[(4'h8):(3'h5)] != ($unsigned(reg590) ~^ (8'hb2))) ?
                          (reg568 ?
                              {{forvar763}} : forvar626) : ({forvar889[(4'hb):(2'h2)]} << (-((8'hb8) < (8'ha1)))));
                      reg5568 <= {$unsigned((reg628 <<< $signed(forvar644)))};
                    end
                end
              for (forvar5569 = (1'h0); (forvar5569 < (2'h2)); forvar5569 = (forvar5569 + (1'h1)))
                begin
                  if (reg692)
                    begin
                      reg5570 <= (~$unsigned({(8'hb1)}));
                    end
                  else
                    begin
                      reg5570 <= $signed((forvar886[(1'h0):(1'h0)] - (^{reg700})));
                    end
                  reg5571 <= $signed(reg982[(3'h7):(2'h3)]);
                  for (forvar5572 = (1'h0); (forvar5572 < (2'h3)); forvar5572 = (forvar5572 + (1'h1)))
                    begin
                      reg5573 <= reg5565[(2'h2):(1'h1)];
                      reg5574 <= forvar630;
                      reg5575 <= reg673;
                    end
                end
              reg5576 <= reg5536;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar5577 = (1'h0); (forvar5577 < (1'h1)); forvar5577 = (forvar5577 + (1'h1)))
        begin
          if (reg648[(3'h5):(2'h2)])
            begin
              reg5578 <= $signed($signed((reg985 < reg932)));
            end
          else
            begin
              if ((&reg936[(2'h2):(1'h1)]))
                begin
                  reg5578 <= $signed($signed(($signed(forvar661) ?
                      $signed(reg838) : forvar689)));
                  for (forvar5579 = (1'h0); (forvar5579 < (1'h0)); forvar5579 = (forvar5579 + (1'h1)))
                    begin
                      reg5580 <= $unsigned(((8'hae) ?
                          $signed({reg659}) : (reg859[(3'h5):(3'h4)] ^ ((8'ha7) << forvar886))));
                    end
                  for (forvar5581 = (1'h0); (forvar5581 < (1'h1)); forvar5581 = (forvar5581 + (1'h1)))
                    begin
                      reg5582 <= (~(!reg1010));
                    end
                end
              else
                begin
                  reg5578 <= reg882[(4'ha):(2'h3)];
                  if ((($signed((reg931 ?
                      reg5547 : reg764)) - ($unsigned(reg843) ?
                      $signed(reg765) : (reg5561 < forvar730))) >>> ((reg958[(3'h4):(2'h3)] << forvar997) ?
                      ($unsigned(forvar969) && forvar919[(2'h3):(2'h3)]) : (((8'hac) * reg743) | {forvar924}))))
                    begin
                      reg5579 <= $signed(((-(forvar687 != reg627)) >= $signed(reg984)));
                      reg5580 <= reg975;
                      reg5581 <= (($signed((reg675 ? reg904 : reg818)) ?
                              $unsigned($signed(reg648)) : {(forvar631 * forvar798)}) ?
                          $signed(((^reg897) ?
                              $unsigned(reg938) : (~^reg719))) : $signed((+reg979[(1'h0):(1'h0)])));
                      reg5582 <= {($signed((reg5575 ?
                              reg847 : forvar731)) >= (8'ha7))};
                    end
                  else
                    begin
                      reg5579 <= forvar573[(4'hc):(4'hc)];
                    end
                  for (forvar5583 = (1'h0); (forvar5583 < (1'h1)); forvar5583 = (forvar5583 + (1'h1)))
                    begin
                      reg5584 <= ($unsigned((!$unsigned(forvar626))) ?
                          {reg896[(2'h3):(2'h3)]} : ((wire5529[(1'h0):(1'h0)] * $signed(reg896)) ?
                              reg959[(1'h1):(1'h0)] : $signed((!(8'hac)))));
                      reg5585 <= ((reg749 || $unsigned({reg632})) ?
                          {((reg698 ? forvar834 : wire558) ?
                                  (8'hac) : {forvar865})} : reg994[(3'h7):(3'h5)]);
                    end
                end
            end
          if (((!reg903) <<< {$unsigned(forvar649[(1'h0):(1'h0)])}))
            begin
              if ((!reg577[(2'h2):(1'h0)]))
                begin
                  for (forvar5586 = (1'h0); (forvar5586 < (2'h3)); forvar5586 = (forvar5586 + (1'h1)))
                    begin
                      reg5587 <= (^~($unsigned($unsigned(reg829)) ^~ $unsigned($unsigned(reg803))));
                      reg5588 <= reg567;
                      reg5589 <= ($signed($signed($signed(forvar907))) << (^~reg757));
                    end
                end
              else
                begin
                  for (forvar5586 = (1'h0); (forvar5586 < (1'h0)); forvar5586 = (forvar5586 + (1'h1)))
                    begin
                      reg5587 <= $unsigned((~|$unsigned($unsigned(forvar942))));
                      reg5588 <= $signed(reg946);
                      reg5589 <= forvar608[(3'h5):(3'h4)];
                      reg5590 <= ((((reg646 ? (8'hae) : reg736) ?
                              (+forvar700) : (+reg634)) ?
                          {(~^forvar927)} : (&$signed(reg614))) & (reg823 ?
                          $signed($signed(reg5533)) : reg563[(3'h6):(3'h6)]));
                    end
                end
              for (forvar5591 = (1'h0); (forvar5591 < (1'h1)); forvar5591 = (forvar5591 + (1'h1)))
                begin
                  if ($signed($signed(($unsigned(reg706) | $signed(forvar640)))))
                    begin
                      reg5592 <= $unsigned(((-reg989) <<< ((&reg822) ?
                          reg5564 : (^forvar926))));
                    end
                  else
                    begin
                      reg5592 <= forvar5581;
                      reg5593 <= (((forvar631[(2'h3):(1'h0)] - (~|reg5546)) >= ({reg715} >= $unsigned(reg720))) ?
                          $signed(reg800[(3'h4):(2'h2)]) : wire5531[(1'h0):(1'h0)]);
                      reg5594 <= $unsigned(($signed({reg645}) ?
                          ($unsigned(reg738) ?
                              {reg5576} : reg1008[(4'hb):(3'h4)]) : $signed((forvar671 ?
                              (8'hba) : (8'had)))));
                    end
                  reg5595 <= forvar895[(2'h2):(1'h0)];
                  if ((8'hb1))
                    begin
                      reg5596 <= (reg805[(2'h2):(1'h1)] ^ (8'had));
                      reg5597 <= {$signed(reg962[(2'h3):(2'h2)])};
                    end
                  else
                    begin
                      reg5596 <= $signed(($unsigned($signed(reg5582)) ?
                          {$signed((8'ha1))} : (forvar952 ?
                              reg5545[(4'ha):(3'h4)] : $unsigned(reg5562))));
                      reg5597 <= $unsigned(forvar644[(3'h6):(3'h6)]);
                      reg5598 <= {$signed($unsigned((-reg686)))};
                    end
                end
              reg5599 <= {forvar693[(1'h1):(1'h0)]};
            end
          else
            begin
              reg5586 <= forvar832[(1'h1):(1'h1)];
              reg5587 <= (reg928[(2'h3):(1'h0)] ?
                  $unsigned((forvar621[(2'h2):(2'h2)] ?
                      forvar832 : reg900)) : ((^~$signed(forvar897)) ?
                      reg760 : forvar858[(4'hd):(4'h9)]));
              for (forvar5588 = (1'h0); (forvar5588 < (1'h0)); forvar5588 = (forvar5588 + (1'h1)))
                begin
                  reg5589 <= $unsigned({reg939});
                  reg5590 <= $unsigned((reg896 ^ $unsigned((reg915 ?
                      (8'hb5) : forvar573))));
                  if (((reg919 <<< $unsigned(forvar629[(3'h6):(3'h4)])) ?
                      ((&(reg826 ~^ reg636)) ?
                          reg605[(1'h1):(1'h0)] : ((^reg671) ?
                              $signed(reg817) : $unsigned(reg975))) : (reg936[(4'h9):(1'h0)] ?
                          (((8'hb3) && reg663) <= (reg744 & reg602)) : {$unsigned(forvar814)})))
                    begin
                      reg5591 <= $unsigned({(((8'h9d) ?
                              forvar859 : reg729) * (~^reg594))});
                      reg5592 <= (+{reg921});
                      reg5593 <= (8'hb8);
                    end
                  else
                    begin
                      reg5591 <= reg719;
                      reg5592 <= $unsigned($signed({reg889}));
                      reg5593 <= ((^(reg5548[(4'hd):(4'h9)] ?
                              $signed(forvar756) : $signed(reg791))) ?
                          $signed($signed(forvar640[(4'h9):(3'h5)])) : $unsigned(reg944[(2'h3):(1'h1)]));
                      reg5594 <= {(^$unsigned(((8'haa) && forvar763)))};
                    end
                  reg5595 <= (~^reg908);
                end
            end
          for (forvar5600 = (1'h0); (forvar5600 < (1'h0)); forvar5600 = (forvar5600 + (1'h1)))
            begin
              for (forvar5601 = (1'h0); (forvar5601 < (2'h3)); forvar5601 = (forvar5601 + (1'h1)))
                begin
                  if (((~&($signed(reg943) ^ (~|reg576))) & $signed(forvar998[(1'h1):(1'h1)])))
                    begin
                      reg5602 <= $signed(forvar871);
                    end
                  else
                    begin
                      reg5602 <= (forvar660[(3'h7):(3'h4)] ?
                          (|$unsigned($unsigned(reg801))) : ($unsigned(reg961) + reg729));
                      reg5603 <= (forvar647[(4'he):(4'he)] ?
                          reg565[(1'h0):(1'h0)] : reg916);
                      reg5604 <= (((~forvar761[(4'hd):(3'h4)]) == $signed($unsigned(forvar911))) ?
                          {(|((8'hb0) ? forvar756 : reg756))} : (8'h9c));
                      reg5605 <= ($signed(reg578[(3'h7):(1'h1)]) ?
                          $unsigned(($signed(reg926) ?
                              reg764[(3'h6):(2'h3)] : forvar5555)) : reg856[(2'h2):(1'h1)]);
                    end
                  for (forvar5606 = (1'h0); (forvar5606 < (2'h2)); forvar5606 = (forvar5606 + (1'h1)))
                    begin
                      reg5607 <= (($signed({reg816}) ?
                          $unsigned((reg946 << forvar858)) : (8'ha2)) - $unsigned(forvar682));
                    end
                  if ($signed({((-reg856) ?
                          (reg876 ? forvar883 : reg879) : $unsigned(reg572))}))
                    begin
                      reg5608 <= reg794[(4'hd):(4'hd)];
                      reg5609 <= ((|{(forvar798 ? reg896 : (8'h9c))}) ?
                          $unsigned($unsigned(reg594[(4'h9):(4'h9)])) : (~forvar5601));
                    end
                  else
                    begin
                      reg5608 <= forvar942;
                      reg5609 <= $signed({$unsigned((-reg728))});
                    end
                end
            end
          for (forvar5610 = (1'h0); (forvar5610 < (2'h3)); forvar5610 = (forvar5610 + (1'h1)))
            begin
              if (forvar920)
                begin
                  if ((~|$unsigned(forvar641)))
                    begin
                      reg5611 <= $signed(($unsigned(reg5558) ?
                          reg774[(1'h1):(1'h0)] : reg5574[(2'h2):(1'h0)]));
                      reg5612 <= $signed({reg1000[(3'h7):(3'h7)]});
                      reg5613 <= $signed(forvar954[(3'h5):(3'h5)]);
                      reg5614 <= (($unsigned(((8'h9c) && reg665)) ?
                              reg5558[(4'h8):(1'h0)] : (8'hb4)) ?
                          reg647[(3'h4):(2'h2)] : reg750);
                    end
                  else
                    begin
                      reg5611 <= $signed({({reg974} ?
                              (forvar5583 ?
                                  reg5598 : reg706) : reg728[(1'h1):(1'h0)])});
                    end
                  for (forvar5615 = (1'h0); (forvar5615 < (1'h0)); forvar5615 = (forvar5615 + (1'h1)))
                    begin
                      reg5616 <= forvar689;
                      reg5617 <= ({$signed(reg980)} ?
                          reg895[(4'hb):(4'h8)] : (~&($signed(reg834) <<< $unsigned(reg646))));
                      reg5618 <= (+forvar722[(3'h4):(2'h2)]);
                      reg5619 <= (^$signed(($signed(reg5564) ?
                          (!forvar5606) : $unsigned(forvar853))));
                    end
                  reg5620 <= (forvar962[(1'h1):(1'h1)] - $unsigned(reg755));
                end
              else
                begin
                  reg5611 <= (forvar5583 ? $signed(reg834) : reg772);
                  for (forvar5612 = (1'h0); (forvar5612 < (2'h2)); forvar5612 = (forvar5612 + (1'h1)))
                    begin
                      reg5613 <= $unsigned(reg946[(3'h4):(2'h2)]);
                      reg5614 <= (~|($signed((reg864 >= reg942)) > forvar5553));
                      reg5615 <= $signed((~|({reg929} ? reg668 : reg954)));
                      reg5616 <= (~{reg613[(3'h5):(2'h2)]});
                    end
                  for (forvar5617 = (1'h0); (forvar5617 < (1'h1)); forvar5617 = (forvar5617 + (1'h1)))
                    begin
                      reg5618 <= {reg599};
                      reg5619 <= $unsigned(forvar746);
                    end
                  for (forvar5620 = (1'h0); (forvar5620 < (2'h2)); forvar5620 = (forvar5620 + (1'h1)))
                    begin
                      reg5621 <= (reg5568 && reg647[(4'ha):(3'h5)]);
                      reg5622 <= reg694;
                      reg5623 <= $signed(({(reg5554 > forvar998)} ?
                          ((reg5605 ^~ reg915) ?
                              reg776[(1'h1):(1'h0)] : ((8'hb6) ?
                                  forvar828 : forvar631)) : reg788));
                      reg5624 <= (($unsigned({reg714}) ?
                              (~|(reg575 <= (8'h9f))) : {(~^(8'hb7))}) ?
                          reg900[(1'h1):(1'h0)] : $unsigned(($signed(reg611) & $unsigned(forvar5579))));
                    end
                end
              for (forvar5625 = (1'h0); (forvar5625 < (2'h3)); forvar5625 = (forvar5625 + (1'h1)))
                begin
                  if ((&$unsigned(reg890)))
                    begin
                      reg5626 <= (8'hb1);
                      reg5627 <= $signed(({(forvar960 ?
                                  forvar689 : forvar895)} ?
                          $signed(forvar671) : reg765[(4'h9):(3'h5)]));
                    end
                  else
                    begin
                      reg5626 <= forvar659[(4'ha):(3'h4)];
                      reg5627 <= $signed(reg964);
                      reg5628 <= $unsigned($signed($unsigned((~|wire558))));
                    end
                  if ({$unsigned($unsigned(reg639))})
                    begin
                      reg5629 <= ($unsigned($unsigned((~|reg1014))) + (((8'h9e) ?
                              forvar650 : $signed(reg597)) ?
                          $signed((~^(8'ha8))) : {reg795}));
                    end
                  else
                    begin
                      reg5629 <= ($unsigned(((reg5581 ? reg976 : (8'ha4)) ?
                              (reg676 || reg839) : (forvar704 >> reg5567))) ?
                          $signed($signed(forvar640[(4'hc):(1'h1)])) : forvar899[(1'h1):(1'h1)]);
                    end
                end
              if ($signed(reg678))
                begin
                  if (reg792[(1'h1):(1'h0)])
                    begin
                      reg5630 <= (8'hb1);
                      reg5631 <= (~&{((~reg5551) ?
                              (reg739 + forvar5583) : (^reg5593))});
                    end
                  else
                    begin
                      reg5630 <= (^~reg611);
                      reg5631 <= $signed(reg934[(3'h5):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar5630 = (1'h0); (forvar5630 < (2'h3)); forvar5630 = (forvar5630 + (1'h1)))
                    begin
                      reg5631 <= $signed($signed($signed(reg679[(3'h6):(1'h1)])));
                      reg5632 <= (^$unsigned($unsigned((reg639 << reg816))));
                      reg5633 <= reg759;
                      reg5634 <= (((|((8'hb1) + reg862)) ?
                          {forvar917} : $signed($signed(forvar924))) > ({$signed(reg774)} ?
                          reg566[(1'h0):(1'h0)] : {{forvar756}}));
                    end
                  if ($signed($signed(($signed(forvar688) <<< (reg5559 >>> forvar756)))))
                    begin
                      reg5635 <= (8'ha5);
                      reg5636 <= $unsigned({$signed({forvar775})});
                    end
                  else
                    begin
                      reg5635 <= (reg652[(2'h2):(1'h1)] <<< (((~|reg690) - (forvar5610 && forvar711)) >> forvar648));
                      reg5636 <= $unsigned(({forvar668} == reg581[(4'ha):(3'h6)]));
                      reg5637 <= reg684;
                    end
                  if (reg5584[(4'ha):(1'h0)])
                    begin
                      reg5638 <= $signed(forvar962[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg5638 <= $signed(({$unsigned(reg946)} ?
                          ((reg706 < reg736) ?
                              (^forvar887) : (forvar5572 && reg891)) : $signed($signed((8'hba)))));
                      reg5639 <= $unsigned(((reg570 ?
                              (~^reg929) : reg767[(3'h6):(3'h5)]) ?
                          reg5561 : reg5564[(3'h4):(2'h3)]));
                    end
                  if ((({(reg5588 ^~ forvar688)} ^ reg776[(2'h2):(1'h0)]) < (8'ha7)))
                    begin
                      reg5640 <= $unsigned(reg818);
                      reg5641 <= $unsigned((forvar633[(2'h3):(2'h2)] ?
                          (8'hab) : reg5599));
                      reg5642 <= ((8'hae) <= $signed($signed(wire5528[(3'h5):(1'h1)])));
                      reg5643 <= (reg5533[(3'h4):(1'h0)] + reg900);
                    end
                  else
                    begin
                      reg5640 <= $signed(reg884);
                    end
                end
            end
        end
      for (forvar5644 = (1'h0); (forvar5644 < (1'h0)); forvar5644 = (forvar5644 + (1'h1)))
        begin
          reg5645 <= (({(+forvar867)} ?
              forvar5572[(4'he):(2'h3)] : (+$unsigned(reg705))) >>> reg877[(3'h6):(1'h0)]);
          reg5646 <= reg889[(1'h1):(1'h1)];
        end
    end
  assign wire5647 = $unsigned($unsigned($unsigned((forvar644 << reg625))));
  always
    @(posedge clk) begin
      for (forvar5648 = (1'h0); (forvar5648 < (1'h1)); forvar5648 = (forvar5648 + (1'h1)))
        begin
          if ((|(&((reg749 < reg5618) <<< reg726))))
            begin
              if (reg5597)
                begin
                  if ((((!forvar5586[(3'h7):(3'h5)]) && $unsigned(((8'ha4) ?
                          reg900 : forvar626))) ?
                      forvar641[(4'hc):(3'h4)] : $unsigned(((forvar832 * reg757) >= (forvar595 ~^ reg5570)))))
                    begin
                      reg5649 <= (reg853[(2'h3):(1'h1)] <= (+reg865));
                      reg5650 <= ($unsigned(reg879[(1'h0):(1'h0)]) - $unsigned(forvar688));
                      reg5651 <= {$unsigned($unsigned(reg5574))};
                      reg5652 <= $unsigned($unsigned(reg591));
                    end
                  else
                    begin
                      reg5649 <= (^(&reg723[(2'h2):(1'h1)]));
                    end
                end
              else
                begin
                  reg5649 <= $unsigned((reg954[(1'h0):(1'h0)] ?
                      $unsigned(reg689) : ((reg739 >> reg5634) ?
                          (reg950 ? (8'haa) : (8'ha2)) : reg887)));
                  for (forvar5650 = (1'h0); (forvar5650 < (1'h1)); forvar5650 = (forvar5650 + (1'h1)))
                    begin
                      reg5651 <= reg676[(2'h3):(1'h1)];
                      reg5652 <= $unsigned((((reg5546 ~^ (8'h9e)) ?
                          $signed((8'hb1)) : reg889) ^ reg816[(4'h9):(1'h0)]));
                    end
                  reg5653 <= (($unsigned((!forvar819)) + reg5581[(1'h1):(1'h0)]) >= $unsigned((forvar669 < $signed(reg5561))));
                  for (forvar5654 = (1'h0); (forvar5654 < (1'h0)); forvar5654 = (forvar5654 + (1'h1)))
                    begin
                      reg5655 <= $signed(forvar620);
                      reg5656 <= reg977;
                      reg5657 <= reg678[(2'h3):(2'h3)];
                      reg5658 <= $unsigned((($signed(reg889) ?
                              $signed(forvar693) : {forvar668}) ?
                          $unsigned($signed(reg804)) : $unsigned(reg763[(1'h0):(1'h0)])));
                    end
                end
            end
          else
            begin
              for (forvar5649 = (1'h0); (forvar5649 < (1'h1)); forvar5649 = (forvar5649 + (1'h1)))
                begin
                  for (forvar5650 = (1'h0); (forvar5650 < (1'h1)); forvar5650 = (forvar5650 + (1'h1)))
                    begin
                      reg5651 <= (~reg850);
                      reg5652 <= (forvar954[(4'h9):(3'h4)] ^ $unsigned($unsigned($unsigned(reg5545))));
                      reg5653 <= reg1008[(4'hc):(2'h2)];
                      reg5654 <= (forvar926 >= reg725);
                    end
                end
            end
          reg5659 <= (~(~^(8'h9e)));
          if ({$signed($signed((reg886 != (8'hba))))})
            begin
              reg5660 <= reg859[(2'h3):(2'h3)];
              if (reg592)
                begin
                  if (($signed((forvar5555 - $signed(forvar648))) ?
                      forvar722 : $signed(reg5578)))
                    begin
                      reg5661 <= $signed(reg1006);
                    end
                  else
                    begin
                      reg5661 <= $unsigned($signed(reg872[(3'h7):(3'h5)]));
                      reg5662 <= (reg717[(4'ha):(3'h4)] ~^ ($unsigned(reg5537) ?
                          wire557[(2'h2):(1'h0)] : (|(reg654 || reg603))));
                    end
                  reg5663 <= (^$signed($unsigned((forvar790 || reg705))));
                  reg5664 <= $unsigned($signed((8'ha4)));
                  if (forvar689[(2'h3):(1'h1)])
                    begin
                      reg5665 <= (&$unsigned((|forvar894)));
                    end
                  else
                    begin
                      reg5665 <= ({(reg990 ?
                              {reg879} : (|reg853))} == forvar900);
                      reg5666 <= reg5557;
                    end
                end
              else
                begin
                  if ((|reg878[(3'h4):(1'h1)]))
                    begin
                      reg5661 <= $unsigned(reg898[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg5661 <= ($signed($unsigned($unsigned(reg597))) << (~^{$signed(reg878)}));
                      reg5662 <= (((|$unsigned(reg5628)) <= {$unsigned(reg810)}) ?
                          (^~$signed($signed(reg5665))) : reg5655[(2'h2):(2'h2)]);
                      reg5663 <= reg628;
                    end
                end
            end
          else
            begin
              for (forvar5660 = (1'h0); (forvar5660 < (2'h3)); forvar5660 = (forvar5660 + (1'h1)))
                begin
                  if ($unsigned((8'h9d)))
                    begin
                      reg5661 <= ((+reg656) | $signed($signed((reg949 ^~ reg5602))));
                      reg5662 <= (~$unsigned($unsigned($unsigned(reg5570))));
                    end
                  else
                    begin
                      reg5661 <= $unsigned((8'ha6));
                      reg5662 <= ((~^(reg757 && reg988[(2'h2):(2'h2)])) >>> reg591[(3'h4):(2'h3)]);
                      reg5663 <= reg941;
                      reg5664 <= (~|({reg990} <<< ({reg5658} ?
                          $unsigned(forvar702) : reg743[(4'hb):(1'h1)])));
                    end
                  reg5665 <= reg706;
                  if (reg628)
                    begin
                      reg5666 <= (~^$unsigned(((forvar711 - reg721) ?
                          (reg666 >>> reg919) : reg643)));
                    end
                  else
                    begin
                      reg5666 <= reg805;
                    end
                end
            end
          reg5667 <= reg678;
        end
      if ((|(8'hb0)))
        begin
          for (forvar5668 = (1'h0); (forvar5668 < (1'h1)); forvar5668 = (forvar5668 + (1'h1)))
            begin
              for (forvar5669 = (1'h0); (forvar5669 < (2'h3)); forvar5669 = (forvar5669 + (1'h1)))
                begin
                  if (reg907)
                    begin
                      reg5670 <= reg898[(4'h9):(1'h0)];
                    end
                  else
                    begin
                      reg5670 <= reg892;
                      reg5671 <= forvar5579[(4'hb):(3'h7)];
                      reg5672 <= $signed($signed(reg721));
                    end
                  if ({(forvar584 >= reg837[(1'h0):(1'h0)])})
                    begin
                      reg5673 <= (reg926 != $unsigned($unsigned(forvar975[(3'h4):(2'h3)])));
                      reg5674 <= (forvar689[(4'hb):(1'h0)] ?
                          $signed(((forvar5532 || reg572) ~^ reg789[(2'h2):(1'h0)])) : (!forvar641));
                      reg5675 <= (($unsigned($unsigned(reg801)) && {$signed(forvar693)}) < reg5642);
                      reg5676 <= (~^$signed((^$unsigned(reg828))));
                    end
                  else
                    begin
                      reg5673 <= (reg799[(3'h4):(1'h1)] >>> {$unsigned($signed(reg5670))});
                    end
                end
              for (forvar5677 = (1'h0); (forvar5677 < (2'h2)); forvar5677 = (forvar5677 + (1'h1)))
                begin
                  if ((-reg665[(1'h0):(1'h0)]))
                    begin
                      reg5678 <= forvar620[(1'h0):(1'h0)];
                      reg5679 <= $unsigned($signed($unsigned((reg808 != forvar893))));
                      reg5680 <= forvar824;
                      reg5681 <= ($signed((reg601[(3'h5):(3'h5)] ?
                          {reg637} : $unsigned(reg765))) >= ($signed((forvar746 ?
                          (8'h9f) : reg565)) > (&forvar893[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg5678 <= ((({reg567} ^ $signed(forvar5612)) ?
                          reg724 : $signed(reg5608)) && $unsigned(reg613));
                      reg5679 <= (($signed($unsigned(reg791)) >>> reg5535) >= {reg910[(3'h4):(2'h3)]});
                      reg5680 <= {($signed($unsigned(reg5645)) * wire5647[(3'h4):(3'h4)])};
                      reg5681 <= reg904[(3'h7):(3'h7)];
                    end
                  for (forvar5682 = (1'h0); (forvar5682 < (1'h1)); forvar5682 = (forvar5682 + (1'h1)))
                    begin
                      reg5683 <= (~forvar884);
                    end
                end
              for (forvar5684 = (1'h0); (forvar5684 < (2'h3)); forvar5684 = (forvar5684 + (1'h1)))
                begin
                  if ($signed({(((8'ha2) * reg5592) <<< {reg609})}))
                    begin
                      reg5685 <= $unsigned((!({reg995} ?
                          (|reg708) : $unsigned(reg5660))));
                      reg5686 <= {($unsigned({reg644}) ?
                              reg896 : (reg901 != (reg739 > reg915)))};
                      reg5687 <= forvar620[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg5685 <= reg708;
                      reg5686 <= $unsigned($signed($unsigned($unsigned(reg646))));
                      reg5687 <= forvar5564;
                      reg5688 <= ({{{reg740}}} >= forvar664);
                    end
                  if (reg905)
                    begin
                      reg5689 <= forvar768;
                    end
                  else
                    begin
                      reg5689 <= $signed($unsigned((reg887 ?
                          (~&forvar5648) : (reg752 ? (8'ha4) : reg603))));
                      reg5690 <= (((8'ha7) <<< $signed((!reg652))) * (((8'h9c) ?
                          $signed(reg623) : (reg684 + reg585)) ~^ {((8'hb6) ?
                              forvar5579 : reg5656)}));
                      reg5691 <= $signed(((|(reg5637 ^~ wire558)) ?
                          $signed(((8'ha9) ?
                              reg5683 : reg664)) : $unsigned({reg946})));
                      reg5692 <= ({(8'ha6)} < ((((8'hae) != reg961) + {reg592}) || reg971[(4'ha):(1'h1)]));
                    end
                  for (forvar5693 = (1'h0); (forvar5693 < (2'h2)); forvar5693 = (forvar5693 + (1'h1)))
                    begin
                      reg5694 <= $signed(($signed(forvar687) ?
                          {(^~forvar761)} : {reg952}));
                      reg5695 <= reg695;
                      reg5696 <= $unsigned((8'h9e));
                      reg5697 <= (!$signed(($signed(reg5611) ?
                          (reg602 ? forvar1005 : forvar895) : reg592)));
                    end
                  if (forvar953[(1'h0):(1'h0)])
                    begin
                      reg5698 <= reg5662;
                      reg5699 <= (~|reg5639[(1'h1):(1'h1)]);
                      reg5700 <= (|($unsigned((reg577 ?
                          reg806 : reg776)) * ($signed(reg635) ^~ (|reg791))));
                    end
                  else
                    begin
                      reg5698 <= {(~(~reg958))};
                      reg5699 <= $unsigned(((8'ha7) || ($unsigned(forvar900) ?
                          reg822[(3'h5):(1'h0)] : {forvar783})));
                      reg5700 <= (reg899[(1'h0):(1'h0)] ?
                          reg878 : $signed(((^~forvar851) ?
                              {reg617} : (reg670 >= reg734))));
                      reg5701 <= (reg5595 ? reg5556 : reg572[(2'h3):(2'h3)]);
                    end
                end
            end
          reg5702 <= (($signed($signed(reg849)) >= (!(reg832 ?
              reg658 : forvar608))) + forvar5615);
          for (forvar5703 = (1'h0); (forvar5703 < (2'h2)); forvar5703 = (forvar5703 + (1'h1)))
            begin
              reg5704 <= reg995;
            end
          for (forvar5705 = (1'h0); (forvar5705 < (1'h0)); forvar5705 = (forvar5705 + (1'h1)))
            begin
              reg5706 <= $unsigned($signed($unsigned(reg942)));
              for (forvar5707 = (1'h0); (forvar5707 < (2'h2)); forvar5707 = (forvar5707 + (1'h1)))
                begin
                  if ((~|((!{reg5580}) ? forvar886[(3'h4):(1'h0)] : {reg862})))
                    begin
                      reg5708 <= (reg988[(3'h7):(3'h4)] ?
                          {reg791[(1'h1):(1'h0)]} : (((reg628 ?
                                  reg831 : forvar824) ?
                              (reg968 ~^ reg752) : reg5534) ^ $unsigned(((8'hb9) ?
                              reg611 : (8'ha6)))));
                      reg5709 <= ($signed((reg5629 ~^ ((8'h9c) >= reg871))) >>> (&$unsigned(reg5552[(4'hc):(2'h2)])));
                      reg5710 <= $signed(reg801);
                      reg5711 <= reg732;
                    end
                  else
                    begin
                      reg5708 <= (($unsigned($unsigned((8'hb0))) ?
                          $signed((8'h9c)) : (~|(reg808 ?
                              forvar997 : (8'h9e)))) > forvar987);
                    end
                  for (forvar5712 = (1'h0); (forvar5712 < (1'h0)); forvar5712 = (forvar5712 + (1'h1)))
                    begin
                      reg5713 <= $unsigned(($unsigned((reg772 | forvar5712)) ?
                          {reg5582[(1'h1):(1'h0)]} : reg5638));
                    end
                end
              if ((forvar5581[(3'h5):(2'h3)] ?
                  reg786[(1'h0):(1'h0)] : ($signed((reg592 < reg625)) ^ (|reg916))))
                begin
                  reg5714 <= forvar562[(3'h6):(3'h5)];
                  for (forvar5715 = (1'h0); (forvar5715 < (1'h1)); forvar5715 = (forvar5715 + (1'h1)))
                    begin
                      reg5716 <= $unsigned($signed($signed($signed(reg942))));
                      reg5717 <= $unsigned(((!(8'haf)) ?
                          ($unsigned(wire555) ?
                              {forvar955} : {forvar927}) : ((forvar862 ^~ reg663) * {reg774})));
                    end
                end
              else
                begin
                  if (reg909)
                    begin
                      reg5714 <= $signed($signed({reg802}));
                      reg5715 <= ((^~(!reg832)) ?
                          reg915 : (&$signed((reg614 ? (8'hae) : reg675))));
                      reg5716 <= (^~((reg5643[(1'h1):(1'h0)] ?
                          reg874[(3'h4):(3'h4)] : $signed(reg680)) >= $unsigned(((8'ha0) ^ (8'ha4)))));
                    end
                  else
                    begin
                      reg5714 <= $unsigned(((~^reg678[(3'h6):(2'h2)]) || $signed((reg5571 ?
                          reg637 : (8'h9e)))));
                      reg5715 <= $signed((|reg813));
                      reg5716 <= $signed({forvar5615});
                      reg5717 <= reg803;
                    end
                  if ($signed((~&$unsigned({reg5692}))))
                    begin
                      reg5718 <= reg872[(1'h0):(1'h0)];
                      reg5719 <= $unsigned(reg984);
                      reg5720 <= (-$signed({(forvar893 && reg865)}));
                    end
                  else
                    begin
                      reg5718 <= forvar881[(4'ha):(3'h7)];
                      reg5719 <= (($signed(reg852[(3'h4):(2'h2)]) >>> $unsigned($signed(reg776))) & reg959[(1'h1):(1'h1)]);
                      reg5720 <= (reg605[(1'h0):(1'h0)] - ((^(forvar924 - reg602)) ?
                          $unsigned(reg5662[(2'h2):(1'h0)]) : $signed(forvar5541)));
                      reg5721 <= reg752;
                    end
                  for (forvar5722 = (1'h0); (forvar5722 < (2'h2)); forvar5722 = (forvar5722 + (1'h1)))
                    begin
                      reg5723 <= (|{((reg714 < reg578) ? (8'hb5) : reg914)});
                      reg5724 <= $unsigned(reg5674[(2'h2):(1'h1)]);
                      reg5725 <= ($unsigned((^~reg917[(1'h1):(1'h1)])) ~^ $unsigned(forvar567));
                    end
                  if ((($signed((~&forvar615)) ~^ (8'ha4)) ?
                      reg5597[(2'h2):(2'h2)] : {$signed((reg825 ?
                              forvar601 : reg938))}))
                    begin
                      reg5726 <= reg835[(4'h9):(1'h0)];
                      reg5727 <= $signed((~|((~|reg712) ~^ (-reg717))));
                      reg5728 <= forvar5591;
                      reg5729 <= $unsigned((&reg5718[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg5726 <= ((&(reg582[(3'h7):(2'h2)] + (reg825 < reg592))) | forvar5559[(4'hc):(3'h7)]);
                    end
                end
              reg5730 <= reg649;
            end
        end
      else
        begin
          for (forvar5668 = (1'h0); (forvar5668 < (1'h1)); forvar5668 = (forvar5668 + (1'h1)))
            begin
              reg5669 <= {(^((reg933 ? reg707 : (8'ha7)) ?
                      (8'had) : $signed(forvar991)))};
              if ($unsigned(($unsigned((reg872 ~^ forvar737)) || $signed($signed(reg895)))))
                begin
                  for (forvar5670 = (1'h0); (forvar5670 < (2'h2)); forvar5670 = (forvar5670 + (1'h1)))
                    begin
                      reg5671 <= reg715;
                      reg5672 <= forvar931;
                      reg5673 <= $signed($unsigned(($unsigned(reg5620) ?
                          $unsigned(forvar746) : $signed(reg869))));
                      reg5674 <= $signed((reg5545 <= ($unsigned(forvar899) ?
                          (+reg867) : (reg809 * reg690))));
                    end
                  if ($unsigned($unsigned((+$signed(reg690)))))
                    begin
                      reg5675 <= (($unsigned(reg900) ?
                          forvar5684[(1'h0):(1'h0)] : $signed(reg5544)) || {((reg5634 ?
                              forvar649 : (8'hb0)) <<< $unsigned(forvar942))});
                      reg5676 <= $signed(reg5695[(3'h4):(1'h0)]);
                      reg5677 <= (~((+reg689) * (reg906 ?
                          forvar952[(1'h0):(1'h0)] : (reg910 || forvar895))));
                    end
                  else
                    begin
                      reg5675 <= (^~reg731);
                      reg5676 <= ({forvar894[(2'h3):(1'h0)]} ^ (~reg5662));
                      reg5677 <= (~^((reg577 ?
                          (8'ha4) : $signed(forvar652)) < ((reg800 ?
                              (8'ha6) : reg821) ?
                          $unsigned(forvar647) : (reg769 ?
                              forvar713 : reg896))));
                    end
                end
              else
                begin
                  if ($unsigned($signed(reg979)))
                    begin
                      reg5670 <= (($signed(((8'hb2) & forvar5591)) ?
                          ({reg634} ?
                              $unsigned(reg901) : (~^reg838)) : reg5718[(2'h3):(2'h3)]) > (reg5613[(1'h1):(1'h1)] ^ (8'ha2)));
                      reg5671 <= (~|({reg5677} < $unsigned((forvar836 >>> reg749))));
                      reg5672 <= reg744[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg5670 <= reg5575[(4'h9):(3'h4)];
                      reg5671 <= forvar579[(4'hc):(2'h2)];
                    end
                  if ($signed({(|$unsigned(reg5597))}))
                    begin
                      reg5673 <= ($signed($unsigned(reg5539[(4'h8):(3'h5)])) ?
                          (+$unsigned(reg582[(2'h2):(1'h1)])) : (~$unsigned((~reg5618))));
                      reg5674 <= $unsigned(forvar595);
                      reg5675 <= $signed(($signed((-(8'ha8))) ?
                          reg5631 : ({forvar621} ?
                              (reg896 < forvar5610) : reg715)));
                    end
                  else
                    begin
                      reg5673 <= $unsigned((^(|reg5646)));
                      reg5674 <= $signed(forvar5722);
                      reg5675 <= reg750[(1'h1):(1'h1)];
                      reg5676 <= reg1018;
                    end
                  reg5677 <= reg575[(3'h6):(3'h6)];
                end
              for (forvar5678 = (1'h0); (forvar5678 < (2'h2)); forvar5678 = (forvar5678 + (1'h1)))
                begin
                  for (forvar5679 = (1'h0); (forvar5679 < (1'h0)); forvar5679 = (forvar5679 + (1'h1)))
                    begin
                      reg5680 <= $signed((~^{(reg5545 ? reg928 : reg907)}));
                      reg5681 <= $unsigned((reg910[(3'h4):(2'h2)] | reg5582[(2'h3):(2'h3)]));
                      reg5682 <= $unsigned({forvar620[(3'h5):(3'h5)]});
                      reg5683 <= $unsigned($signed($signed((forvar996 ^~ reg5726))));
                    end
                  for (forvar5684 = (1'h0); (forvar5684 < (1'h0)); forvar5684 = (forvar5684 + (1'h1)))
                    begin
                      reg5685 <= $unsigned(reg5623);
                    end
                  for (forvar5686 = (1'h0); (forvar5686 < (2'h2)); forvar5686 = (forvar5686 + (1'h1)))
                    begin
                      reg5687 <= $unsigned(wire5647);
                    end
                  for (forvar5688 = (1'h0); (forvar5688 < (2'h2)); forvar5688 = (forvar5688 + (1'h1)))
                    begin
                      reg5689 <= (reg1006[(3'h4):(1'h0)] ?
                          (8'hb6) : {(&$unsigned(forvar688))});
                      reg5690 <= reg5689;
                    end
                end
              reg5691 <= $signed((((!reg701) << $signed(reg616)) ?
                  $signed($unsigned(forvar911)) : $unsigned(((8'ha0) ^~ reg823))));
            end
          if (((reg973[(2'h3):(1'h1)] ^~ (((8'ha9) + forvar660) ?
              forvar5705[(2'h2):(2'h2)] : $unsigned((8'haf)))) <<< reg5724[(4'hb):(2'h2)]))
            begin
              for (forvar5692 = (1'h0); (forvar5692 < (2'h2)); forvar5692 = (forvar5692 + (1'h1)))
                begin
                  for (forvar5693 = (1'h0); (forvar5693 < (1'h1)); forvar5693 = (forvar5693 + (1'h1)))
                    begin
                      reg5694 <= {$unsigned(reg715[(3'h5):(1'h0)])};
                      reg5695 <= $signed(reg5723[(3'h4):(1'h1)]);
                      reg5696 <= reg972[(3'h4):(1'h1)];
                    end
                  for (forvar5697 = (1'h0); (forvar5697 < (2'h2)); forvar5697 = (forvar5697 + (1'h1)))
                    begin
                      reg5698 <= ((!$unsigned(reg5714)) ?
                          {(-$signed(reg5631))} : {reg635[(3'h5):(2'h2)]});
                      reg5699 <= reg5561[(4'h9):(1'h1)];
                      reg5700 <= {{(^~reg777)}};
                    end
                end
              if ((({reg680[(4'hc):(4'hb)]} ?
                      $unsigned((-reg5637)) : $signed($signed(reg5581))) ?
                  reg999 : ({(reg5632 ?
                          reg5539 : wire5524)} ~^ ($signed(reg610) + $unsigned(forvar831)))))
                begin
                  for (forvar5701 = (1'h0); (forvar5701 < (1'h0)); forvar5701 = (forvar5701 + (1'h1)))
                    begin
                      reg5702 <= $unsigned((forvar630 | $unsigned((~&reg826))));
                      reg5703 <= forvar770[(2'h3):(2'h3)];
                    end
                  if (reg5659)
                    begin
                      reg5704 <= (forvar895[(2'h2):(1'h1)] ?
                          (reg939 ?
                              reg566[(1'h1):(1'h0)] : {reg5660}) : reg915[(4'h8):(2'h2)]);
                      reg5705 <= ($unsigned({forvar638}) && (reg5653[(1'h1):(1'h0)] ?
                          (&$unsigned(reg701)) : (reg972 ?
                              (^~reg786) : reg1006)));
                      reg5706 <= forvar573;
                    end
                  else
                    begin
                      reg5704 <= (~&(((forvar886 != reg5676) & (^forvar629)) >> $signed((reg5556 >> reg900))));
                    end
                  for (forvar5707 = (1'h0); (forvar5707 < (1'h0)); forvar5707 = (forvar5707 + (1'h1)))
                    begin
                      reg5708 <= $signed((reg5724[(4'ha):(3'h6)] - (^~{forvar629})));
                      reg5709 <= $unsigned((+(forvar819[(1'h1):(1'h1)] ?
                          (8'hb7) : $signed((8'hac)))));
                      reg5710 <= $signed(reg5538);
                      reg5711 <= forvar5715;
                    end
                end
              else
                begin
                  for (forvar5701 = (1'h0); (forvar5701 < (1'h0)); forvar5701 = (forvar5701 + (1'h1)))
                    begin
                      reg5702 <= {($signed($unsigned(reg739)) ?
                              (!(~&wire557)) : (~&(reg5584 ?
                                  (8'hba) : (8'ha4))))};
                      reg5703 <= $signed((reg567[(3'h4):(2'h2)] ?
                          $signed(reg596) : (reg5730[(2'h2):(2'h2)] ?
                              (8'hac) : forvar659[(1'h0):(1'h0)])));
                    end
                  reg5704 <= forvar5707[(3'h4):(3'h4)];
                  for (forvar5705 = (1'h0); (forvar5705 < (1'h0)); forvar5705 = (forvar5705 + (1'h1)))
                    begin
                      reg5706 <= reg5559;
                      reg5707 <= (8'haa);
                      reg5708 <= (-$unsigned({{reg5636}}));
                    end
                end
            end
          else
            begin
              if ({forvar5555})
                begin
                  if (($signed($unsigned((reg5688 == (8'h9f)))) + {{(+forvar5583)}}))
                    begin
                      reg5692 <= {({$unsigned((8'hb7))} ?
                              $unsigned(reg801) : $signed((+(8'hae))))};
                      reg5693 <= wire560;
                      reg5694 <= $unsigned({(!$unsigned((8'haa)))});
                    end
                  else
                    begin
                      reg5692 <= $signed(($unsigned(forvar575) ?
                          reg886[(2'h3):(2'h2)] : $signed({(8'ha7)})));
                      reg5693 <= $unsigned((8'hae));
                    end
                  if (reg702)
                    begin
                      reg5695 <= {forvar607};
                      reg5696 <= (8'ha3);
                    end
                  else
                    begin
                      reg5695 <= ($unsigned(forvar722) >> reg614);
                    end
                end
              else
                begin
                  for (forvar5692 = (1'h0); (forvar5692 < (1'h1)); forvar5692 = (forvar5692 + (1'h1)))
                    begin
                      reg5693 <= ({(!$signed(forvar893))} != $unsigned(($signed(reg731) ?
                          $unsigned(reg670) : $unsigned(reg5676))));
                    end
                  for (forvar5694 = (1'h0); (forvar5694 < (2'h3)); forvar5694 = (forvar5694 + (1'h1)))
                    begin
                      reg5695 <= $unsigned(reg5723);
                      reg5696 <= forvar787;
                      reg5697 <= reg948[(1'h0):(1'h0)];
                    end
                  for (forvar5698 = (1'h0); (forvar5698 < (1'h0)); forvar5698 = (forvar5698 + (1'h1)))
                    begin
                      reg5699 <= forvar5550;
                      reg5700 <= $signed(((~|$signed(forvar567)) ?
                          $signed(reg662) : $unsigned($signed(reg5590))));
                      reg5701 <= reg5634;
                    end
                  for (forvar5702 = (1'h0); (forvar5702 < (2'h2)); forvar5702 = (forvar5702 + (1'h1)))
                    begin
                      reg5703 <= forvar931;
                      reg5704 <= forvar630[(3'h4):(3'h4)];
                      reg5705 <= (8'hae);
                    end
                end
              if ((8'hb0))
                begin
                  reg5706 <= (-reg5655);
                end
              else
                begin
                  if ($unsigned(forvar602[(1'h0):(1'h0)]))
                    begin
                      reg5706 <= (^{(8'hb7)});
                    end
                  else
                    begin
                      reg5706 <= ((~^$unsigned(reg5694)) ~^ $unsigned((~^(forvar588 ?
                          (8'hb4) : (8'ha3)))));
                      reg5707 <= reg5694[(3'h4):(2'h3)];
                      reg5708 <= $signed(reg597);
                    end
                  reg5709 <= reg5575[(3'h4):(2'h2)];
                  if ((reg673[(3'h6):(3'h4)] ~^ (~^reg601[(1'h0):(1'h0)])))
                    begin
                      reg5710 <= (~|reg5723);
                      reg5711 <= $unsigned($unsigned($unsigned((!wire5530))));
                      reg5712 <= $signed(($unsigned((reg573 ?
                          reg5723 : reg577)) >>> reg1000[(4'h8):(2'h2)]));
                    end
                  else
                    begin
                      reg5710 <= ({(^reg593[(3'h4):(2'h2)])} ?
                          (forvar5532 ?
                              {{(8'hb8)}} : $unsigned(reg703[(4'he):(3'h6)])) : ((reg655[(3'h6):(3'h5)] ?
                                  {reg694} : (|(8'ha9))) ?
                              {reg837} : {(reg936 ^~ reg851)}));
                    end
                  for (forvar5713 = (1'h0); (forvar5713 < (2'h3)); forvar5713 = (forvar5713 + (1'h1)))
                    begin
                      reg5714 <= {(-($unsigned(reg5562) ?
                              forvar5559 : $signed(reg955)))};
                      reg5715 <= reg5638[(2'h2):(1'h0)];
                      reg5716 <= (reg767 ?
                          $unsigned((&(forvar756 ?
                              reg797 : forvar688))) : ($signed((forvar5678 ?
                                  reg821 : reg906)) ?
                              forvar5705 : (~|(8'hb0))));
                    end
                end
              if ({(~forvar5588)})
                begin
                  reg5717 <= {reg663};
                  reg5718 <= (|(({forvar630} ?
                          (reg616 ?
                              reg5538 : forvar5703) : reg1010[(4'ha):(1'h0)]) ?
                      (~^(~&(8'hb3))) : $unsigned($signed((8'ha1)))));
                end
              else
                begin
                  for (forvar5717 = (1'h0); (forvar5717 < (2'h2)); forvar5717 = (forvar5717 + (1'h1)))
                    begin
                      reg5718 <= (~^(|(|(~|reg5677))));
                    end
                  if (forvar881[(4'h8):(2'h2)])
                    begin
                      reg5719 <= (8'hb3);
                    end
                  else
                    begin
                      reg5719 <= ($unsigned(((reg994 ? forvar922 : forvar643) ?
                              (forvar664 ?
                                  (8'hb9) : reg5717) : reg647[(4'h9):(4'h8)])) ?
                          (reg899 ?
                              {$signed((8'hb1))} : $unsigned((reg921 ?
                                  forvar702 : (8'haf)))) : $signed(($signed(reg869) < reg5643[(2'h3):(1'h1)])));
                      reg5720 <= (reg5589 ?
                          ({(reg5585 & forvar5678)} >>> forvar790) : reg838);
                    end
                  if ($unsigned((((reg870 - reg665) < $unsigned(forvar676)) & $signed(forvar704))))
                    begin
                      reg5721 <= reg912[(3'h6):(2'h3)];
                      reg5722 <= $signed({(~^reg916)});
                      reg5723 <= reg593;
                      reg5724 <= $unsigned($signed(((forvar987 | (8'hb4)) ?
                          reg739[(1'h1):(1'h0)] : $signed(forvar689))));
                    end
                  else
                    begin
                      reg5721 <= forvar602[(2'h2):(1'h1)];
                      reg5722 <= ($unsigned(($unsigned(reg704) ?
                          $unsigned(forvar5717) : forvar659)) - reg580[(3'h5):(3'h5)]);
                    end
                  for (forvar5725 = (1'h0); (forvar5725 < (2'h2)); forvar5725 = (forvar5725 + (1'h1)))
                    begin
                      reg5726 <= forvar996;
                      reg5727 <= ($signed({(reg830 ? reg1004 : reg660)}) ?
                          (forvar5588 ?
                              reg5551[(4'hd):(3'h6)] : ((reg862 ?
                                  (8'ha9) : reg791) - $signed(reg815))) : (&reg968));
                      reg5728 <= ({(reg686[(4'ha):(1'h0)] ?
                              $unsigned(forvar987) : (reg1012 * reg5560))} + (^~reg5638));
                    end
                end
              for (forvar5729 = (1'h0); (forvar5729 < (1'h1)); forvar5729 = (forvar5729 + (1'h1)))
                begin
                  for (forvar5730 = (1'h0); (forvar5730 < (2'h2)); forvar5730 = (forvar5730 + (1'h1)))
                    begin
                      reg5731 <= {(reg5711[(2'h2):(1'h1)] ?
                              reg943 : forvar806[(2'h2):(1'h0)])};
                      reg5732 <= ((^~$signed($unsigned(reg563))) ?
                          ((reg978 ?
                              $signed((8'ha0)) : {reg967}) >= (8'hb1)) : $unsigned({(+reg609)}));
                      reg5733 <= ($signed((reg704 ?
                              reg574 : (forvar5541 ? reg823 : (8'ha2)))) ?
                          (^(reg894 ?
                              $signed(reg992) : forvar906)) : ($unsigned((reg5669 ?
                              forvar5564 : (8'hb5))) <= (8'hb4)));
                      reg5734 <= ($unsigned($signed((reg5642 <<< forvar630))) ?
                          reg771 : $unsigned((reg655[(3'h4):(1'h1)] > $signed(forvar843))));
                    end
                end
            end
          reg5735 <= forvar620[(3'h4):(1'h1)];
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1021  (y, clk, wire1022, wire1023, wire1024, wire1025);
  output wire [(32'h170a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire1022;
  input wire [(5'h10):(1'h0)] wire1023;
  input wire [(3'h5):(1'h0)] wire1024;
  input wire signed [(3'h7):(1'h0)] wire1025;
  reg signed [(4'hb):(1'h0)] forvar5501 = (1'h0);
  reg [(3'h6):(1'h0)] reg5523 = (1'h0);
  reg [(4'hc):(1'h0)] reg5522 = (1'h0);
  reg [(2'h2):(1'h0)] reg5521 = (1'h0);
  reg [(4'h8):(1'h0)] reg5520 = (1'h0);
  reg [(4'hd):(1'h0)] reg5519 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5518 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5517 = (1'h0);
  reg [(5'h10):(1'h0)] reg5516 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5515 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5514 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5513 = (1'h0);
  reg [(3'h6):(1'h0)] reg5512 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5506 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5502 = (1'h0);
  reg [(2'h3):(1'h0)] reg5511 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5510 = (1'h0);
  reg [(4'he):(1'h0)] reg5509 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5508 = (1'h0);
  reg [(4'h9):(1'h0)] reg5507 = (1'h0);
  reg [(3'h4):(1'h0)] reg5506 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5505 = (1'h0);
  reg [(3'h4):(1'h0)] reg5504 = (1'h0);
  reg [(4'h9):(1'h0)] reg5503 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5502 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5501 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5500 = (1'h0);
  reg [(4'hd):(1'h0)] reg5499 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5491 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5495 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5493 = (1'h0);
  reg [(4'hf):(1'h0)] reg5489 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5480 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5488 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5478 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5469 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5468 = (1'h0);
  reg [(3'h6):(1'h0)] reg5498 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5497 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5496 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5495 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5494 = (1'h0);
  reg [(3'h6):(1'h0)] reg5493 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5492 = (1'h0);
  reg [(3'h5):(1'h0)] reg5491 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5490 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5489 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5488 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5487 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5484 = (1'h0);
  reg [(3'h7):(1'h0)] reg5486 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5485 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5484 = (1'h0);
  reg [(5'h10):(1'h0)] reg5483 = (1'h0);
  reg [(4'hf):(1'h0)] reg5482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5481 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5480 = (1'h0);
  reg [(4'hd):(1'h0)] reg5479 = (1'h0);
  reg [(2'h3):(1'h0)] reg5478 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5477 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5475 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5474 = (1'h0);
  reg [(5'h10):(1'h0)] reg5473 = (1'h0);
  reg [(4'h8):(1'h0)] reg5472 = (1'h0);
  reg [(3'h7):(1'h0)] reg5471 = (1'h0);
  reg [(3'h7):(1'h0)] reg5470 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5469 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5468 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5460 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5459 = (1'h0);
  reg [(4'h8):(1'h0)] reg5467 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5466 = (1'h0);
  reg [(4'hb):(1'h0)] reg5465 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5464 = (1'h0);
  reg [(4'hc):(1'h0)] reg5463 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5462 = (1'h0);
  reg [(2'h3):(1'h0)] reg5461 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5460 = (1'h0);
  reg [(4'hc):(1'h0)] reg5456 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5455 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5459 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5458 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5457 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5456 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5455 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5454 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5441 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5440 = (1'h0);
  reg [(3'h7):(1'h0)] reg5436 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5434 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5433 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5425 = (1'h0);
  reg [(4'hb):(1'h0)] reg5432 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5419 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5418 = (1'h0);
  reg [(4'ha):(1'h0)] reg5414 = (1'h0);
  reg [(4'hf):(1'h0)] reg5412 = (1'h0);
  reg [(4'he):(1'h0)] forvar5411 = (1'h0);
  reg [(4'h8):(1'h0)] reg5410 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5407 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5404 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5403 = (1'h0);
  reg [(3'h5):(1'h0)] reg5453 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5452 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5451 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5450 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5449 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5448 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5447 = (1'h0);
  reg [(2'h2):(1'h0)] reg5446 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5445 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5438 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5437 = (1'h0);
  reg [(3'h7):(1'h0)] reg5444 = (1'h0);
  reg [(4'hf):(1'h0)] reg5443 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5442 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5441 = (1'h0);
  reg [(4'he):(1'h0)] forvar5440 = (1'h0);
  reg [(4'hf):(1'h0)] reg5439 = (1'h0);
  reg [(4'he):(1'h0)] forvar5438 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5437 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5436 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5435 = (1'h0);
  reg [(3'h5):(1'h0)] reg5434 = (1'h0);
  reg [(4'hd):(1'h0)] reg5433 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5432 = (1'h0);
  reg [(4'h9):(1'h0)] reg5431 = (1'h0);
  reg [(4'hb):(1'h0)] reg5430 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5427 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5422 = (1'h0);
  reg [(4'h8):(1'h0)] reg5429 = (1'h0);
  reg [(3'h6):(1'h0)] reg5428 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5427 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5426 = (1'h0);
  reg [(3'h7):(1'h0)] reg5425 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5424 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5423 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5422 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5421 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5420 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5419 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5418 = (1'h0);
  reg [(4'hf):(1'h0)] reg5417 = (1'h0);
  reg [(5'h10):(1'h0)] reg5416 = (1'h0);
  reg [(3'h5):(1'h0)] reg5415 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5414 = (1'h0);
  reg [(4'hd):(1'h0)] reg5413 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5412 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5411 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5410 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5405 = (1'h0);
  reg [(2'h2):(1'h0)] reg5402 = (1'h0);
  reg [(3'h6):(1'h0)] reg5409 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5408 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5407 = (1'h0);
  reg [(5'h10):(1'h0)] reg5406 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5405 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5404 = (1'h0);
  reg [(3'h7):(1'h0)] reg5403 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5402 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5401 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5394 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5400 = (1'h0);
  reg [(2'h2):(1'h0)] reg5399 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5398 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5397 = (1'h0);
  reg [(3'h5):(1'h0)] reg5396 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5395 = (1'h0);
  reg [(5'h10):(1'h0)] reg5394 = (1'h0);
  reg [(3'h7):(1'h0)] reg5393 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5392 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5388 = (1'h0);
  reg [(4'hd):(1'h0)] reg5391 = (1'h0);
  reg [(3'h4):(1'h0)] reg5390 = (1'h0);
  reg [(3'h5):(1'h0)] reg5389 = (1'h0);
  reg [(4'he):(1'h0)] reg5388 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5387 = (1'h0);
  reg [(4'ha):(1'h0)] reg5386 = (1'h0);
  reg [(4'h8):(1'h0)] reg5385 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5383 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5382 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5381 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5380 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5379 = (1'h0);
  reg [(2'h3):(1'h0)] reg5379 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5378 = (1'h0);
  reg [(3'h7):(1'h0)] reg5377 = (1'h0);
  reg [(4'h8):(1'h0)] reg5376 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5375 = (1'h0);
  reg [(3'h7):(1'h0)] reg5374 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5373 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5372 = (1'h0);
  reg [(2'h3):(1'h0)] reg5371 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5369 = (1'h0);
  reg [(3'h4):(1'h0)] reg5368 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5367 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5366 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5365 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5364 = (1'h0);
  reg [(2'h2):(1'h0)] reg5363 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5362 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5361 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5360 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5359 = (1'h0);
  reg [(4'h9):(1'h0)] reg5358 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5357 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5356 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5355 = (1'h0);
  reg [(4'hd):(1'h0)] reg5354 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5353 = (1'h0);
  reg [(3'h7):(1'h0)] reg5352 = (1'h0);
  reg [(3'h4):(1'h0)] reg5351 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5349 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5346 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5341 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5347 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5343 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5339 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5338 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5350 = (1'h0);
  reg [(4'h9):(1'h0)] reg5349 = (1'h0);
  reg [(3'h5):(1'h0)] reg5348 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5347 = (1'h0);
  reg [(4'he):(1'h0)] reg5346 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5345 = (1'h0);
  reg [(4'ha):(1'h0)] reg5344 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5343 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5342 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5341 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5340 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5339 = (1'h0);
  reg [(5'h10):(1'h0)] reg5338 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5337 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire5336;
  reg [(3'h5):(1'h0)] reg5335 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5334 = (1'h0);
  reg [(4'ha):(1'h0)] reg5329 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5333 = (1'h0);
  reg [(3'h4):(1'h0)] reg5332 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5331 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5330 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5329 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5328 = (1'h0);
  reg [(4'hf):(1'h0)] reg5327 = (1'h0);
  reg [(5'h10):(1'h0)] reg5326 = (1'h0);
  reg [(4'h9):(1'h0)] reg5325 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5324 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5323 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5298 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5295 = (1'h0);
  reg [(3'h5):(1'h0)] reg5294 = (1'h0);
  reg [(4'hf):(1'h0)] reg5322 = (1'h0);
  reg [(2'h3):(1'h0)] reg5321 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5320 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5319 = (1'h0);
  reg [(4'hf):(1'h0)] reg5318 = (1'h0);
  reg [(3'h4):(1'h0)] reg5317 = (1'h0);
  reg [(4'h9):(1'h0)] reg5316 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5315 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5314 = (1'h0);
  reg [(2'h2):(1'h0)] reg5313 = (1'h0);
  reg [(3'h7):(1'h0)] reg5312 = (1'h0);
  reg [(4'he):(1'h0)] reg5311 = (1'h0);
  reg [(4'hf):(1'h0)] reg5310 = (1'h0);
  reg [(4'ha):(1'h0)] reg5309 = (1'h0);
  reg [(4'he):(1'h0)] reg5308 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5307 = (1'h0);
  reg [(4'hc):(1'h0)] reg5306 = (1'h0);
  reg [(4'he):(1'h0)] forvar5305 = (1'h0);
  reg [(4'hc):(1'h0)] reg5304 = (1'h0);
  reg [(3'h5):(1'h0)] reg5303 = (1'h0);
  reg [(4'h9):(1'h0)] reg5302 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5301 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5300 = (1'h0);
  reg [(4'hb):(1'h0)] reg5299 = (1'h0);
  reg [(3'h4):(1'h0)] reg5298 = (1'h0);
  reg [(4'hd):(1'h0)] reg5297 = (1'h0);
  reg [(2'h3):(1'h0)] reg5296 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5295 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5294 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5293 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5292 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire5291;
  wire [(3'h5):(1'h0)] wire5290;
  reg [(4'he):(1'h0)] reg5289 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5288 = (1'h0);
  reg [(4'he):(1'h0)] reg5287 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5286 = (1'h0);
  reg [(4'hf):(1'h0)] reg5285 = (1'h0);
  reg [(4'h9):(1'h0)] reg5284 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5282 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5278 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5271 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5270 = (1'h0);
  reg [(3'h5):(1'h0)] reg5281 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5276 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5272 = (1'h0);
  reg [(4'ha):(1'h0)] reg5283 = (1'h0);
  reg [(3'h6):(1'h0)] reg5282 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5281 = (1'h0);
  reg [(3'h6):(1'h0)] reg5280 = (1'h0);
  reg [(4'h8):(1'h0)] reg5279 = (1'h0);
  reg [(4'h9):(1'h0)] reg5278 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5277 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5276 = (1'h0);
  reg [(4'hd):(1'h0)] reg5275 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5274 = (1'h0);
  reg [(3'h6):(1'h0)] reg5273 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5272 = (1'h0);
  reg [(4'hf):(1'h0)] reg5271 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5270 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5269 = (1'h0);
  reg [(4'hc):(1'h0)] reg5268 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5267 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5260 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5255 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5266 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5265 = (1'h0);
  reg [(4'ha):(1'h0)] reg5264 = (1'h0);
  reg [(4'he):(1'h0)] reg5263 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5262 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5261 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5260 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5259 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5258 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5257 = (1'h0);
  reg [(4'he):(1'h0)] reg5256 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5255 = (1'h0);
  reg [(4'h9):(1'h0)] reg5254 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5253 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5252 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5251 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5250 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5249 = (1'h0);
  reg [(3'h6):(1'h0)] reg5248 = (1'h0);
  reg [(2'h2):(1'h0)] reg5247 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5246 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5245 = (1'h0);
  reg [(4'hf):(1'h0)] reg5244 = (1'h0);
  reg [(3'h5):(1'h0)] reg5243 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5242 = (1'h0);
  reg [(4'h9):(1'h0)] reg5241 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5240 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5239 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5238 = (1'h0);
  reg [(4'h9):(1'h0)] reg5237 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5236 = (1'h0);
  reg [(5'h10):(1'h0)] reg5235 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5234 = (1'h0);
  reg [(4'hc):(1'h0)] reg5233 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5232 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5231 = (1'h0);
  reg [(4'hd):(1'h0)] reg5230 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5229 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5228 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5227 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5226 = (1'h0);
  reg [(5'h10):(1'h0)] reg5225 = (1'h0);
  reg [(3'h7):(1'h0)] reg5224 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5223 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5222 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5221 = (1'h0);
  reg [(3'h7):(1'h0)] reg5220 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5219 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5218 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5217 = (1'h0);
  reg [(4'h9):(1'h0)] reg5216 = (1'h0);
  reg [(3'h4):(1'h0)] reg5215 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5214 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5213 = (1'h0);
  reg [(4'h9):(1'h0)] reg5212 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5211 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5210 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5209 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5208 = (1'h0);
  reg [(4'hd):(1'h0)] reg5192 = (1'h0);
  reg [(4'hf):(1'h0)] reg5187 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5185 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5182 = (1'h0);
  reg [(4'hd):(1'h0)] reg5207 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5206 = (1'h0);
  reg [(4'ha):(1'h0)] reg5205 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5204 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5203 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5202 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5201 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5200 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5199 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5198 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5197 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5196 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5195 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5194 = (1'h0);
  reg [(2'h2):(1'h0)] reg5193 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5192 = (1'h0);
  reg [(4'he):(1'h0)] reg5191 = (1'h0);
  reg [(3'h5):(1'h0)] reg5190 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5189 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5188 = (1'h0);
  reg [(4'he):(1'h0)] forvar5187 = (1'h0);
  reg [(4'hc):(1'h0)] reg5186 = (1'h0);
  reg [(3'h4):(1'h0)] reg5185 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5183 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5184 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5183 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5182 = (1'h0);
  reg [(4'h9):(1'h0)] reg5181 = (1'h0);
  reg [(2'h3):(1'h0)] reg5180 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5179 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5178 = (1'h0);
  reg [(2'h2):(1'h0)] reg5177 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5176 = (1'h0);
  reg [(4'he):(1'h0)] forvar5175 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5174 = (1'h0);
  reg [(3'h6):(1'h0)] reg5173 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5172 = (1'h0);
  reg [(4'h8):(1'h0)] reg5171 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5170 = (1'h0);
  reg [(5'h10):(1'h0)] reg5169 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5168 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5167 = (1'h0);
  reg [(4'he):(1'h0)] reg5166 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5165 = (1'h0);
  reg [(3'h7):(1'h0)] reg5164 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5163 = (1'h0);
  reg [(4'hf):(1'h0)] reg5162 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5161 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5160 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5159 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5158 = (1'h0);
  reg [(2'h2):(1'h0)] reg5157 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5156 = (1'h0);
  reg [(4'hb):(1'h0)] reg5155 = (1'h0);
  reg [(3'h7):(1'h0)] reg5154 = (1'h0);
  reg [(4'ha):(1'h0)] reg5153 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5152 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5151 = (1'h0);
  reg [(3'h6):(1'h0)] reg5150 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5149 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5148 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5147 = (1'h0);
  reg [(3'h5):(1'h0)] reg5146 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5141 = (1'h0);
  reg [(4'ha):(1'h0)] reg5139 = (1'h0);
  reg [(2'h2):(1'h0)] reg5145 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5144 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5143 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5142 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5141 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5140 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5139 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5138 = (1'h0);
  reg [(4'ha):(1'h0)] reg5137 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5136 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5117 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5116 = (1'h0);
  reg [(4'h8):(1'h0)] reg5135 = (1'h0);
  reg [(4'hb):(1'h0)] reg5134 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5133 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5132 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5131 = (1'h0);
  reg [(3'h6):(1'h0)] reg5130 = (1'h0);
  reg [(4'hb):(1'h0)] reg5129 = (1'h0);
  reg [(3'h4):(1'h0)] reg5128 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5127 = (1'h0);
  reg [(4'hb):(1'h0)] reg5126 = (1'h0);
  reg [(4'hc):(1'h0)] reg5125 = (1'h0);
  reg [(4'hb):(1'h0)] reg5124 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5123 = (1'h0);
  reg [(3'h5):(1'h0)] reg5122 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5121 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5120 = (1'h0);
  reg [(4'h9):(1'h0)] reg5119 = (1'h0);
  reg [(3'h4):(1'h0)] reg5118 = (1'h0);
  reg [(4'he):(1'h0)] forvar5117 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5116 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5115 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5109 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5106 = (1'h0);
  reg [(3'h4):(1'h0)] reg5114 = (1'h0);
  reg [(4'ha):(1'h0)] reg5113 = (1'h0);
  reg [(3'h5):(1'h0)] reg5112 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5111 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5110 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5109 = (1'h0);
  reg [(4'h8):(1'h0)] reg5108 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5107 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5106 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5105 = (1'h0);
  reg [(4'he):(1'h0)] reg5104 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5103 = (1'h0);
  reg [(4'hb):(1'h0)] reg5102 = (1'h0);
  reg [(4'hd):(1'h0)] reg5101 = (1'h0);
  reg [(3'h4):(1'h0)] reg5100 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5099 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5098 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5097 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5096 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5095 = (1'h0);
  reg [(4'hd):(1'h0)] reg5094 = (1'h0);
  reg [(4'hd):(1'h0)] reg5093 = (1'h0);
  reg [(2'h2):(1'h0)] reg5092 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5091 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5090 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5089 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5088 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5087 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5086 = (1'h0);
  reg [(5'h10):(1'h0)] reg5085 = (1'h0);
  reg [(3'h6):(1'h0)] reg5084 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5083 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5082 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5081 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5080 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5079 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5078 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5077 = (1'h0);
  reg [(4'hc):(1'h0)] reg5076 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5075 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5074 = (1'h0);
  reg [(4'he):(1'h0)] reg5073 = (1'h0);
  reg [(2'h3):(1'h0)] reg5072 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5071 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5070 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5069 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5068 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5067 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5066 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5065 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5064 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5063 = (1'h0);
  reg [(4'hd):(1'h0)] reg5062 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5061 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5060 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5059 = (1'h0);
  reg [(3'h5):(1'h0)] reg5058 = (1'h0);
  reg [(4'h9):(1'h0)] reg5057 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5056 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5055 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5054 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5053 = (1'h0);
  reg [(4'hc):(1'h0)] reg5052 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5051 = (1'h0);
  reg [(2'h2):(1'h0)] reg5050 = (1'h0);
  reg [(3'h5):(1'h0)] reg5049 = (1'h0);
  reg [(4'hd):(1'h0)] reg5048 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5047 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5046 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5045 = (1'h0);
  reg [(4'ha):(1'h0)] reg5044 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5043 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5042 = (1'h0);
  reg [(4'ha):(1'h0)] reg5041 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5040 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5033 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5030 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5039 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5038 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5037 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5036 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5035 = (1'h0);
  reg [(4'ha):(1'h0)] reg5034 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5033 = (1'h0);
  reg [(4'ha):(1'h0)] reg5032 = (1'h0);
  reg [(4'hd):(1'h0)] reg5031 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5030 = (1'h0);
  reg [(3'h4):(1'h0)] reg5029 = (1'h0);
  reg [(4'hd):(1'h0)] reg5028 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5027 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5026 = (1'h0);
  reg [(3'h4):(1'h0)] reg5025 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5024 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5023 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5022 = (1'h0);
  reg [(4'he):(1'h0)] reg5021 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5020 = (1'h0);
  reg [(4'he):(1'h0)] forvar5019 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5018 = (1'h0);
  reg [(4'hb):(1'h0)] reg5017 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5016 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5015 = (1'h0);
  reg [(4'hf):(1'h0)] reg5014 = (1'h0);
  reg [(3'h4):(1'h0)] reg5013 = (1'h0);
  reg [(4'h9):(1'h0)] reg5012 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5011 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5010 = (1'h0);
  reg [(4'h8):(1'h0)] reg5009 = (1'h0);
  reg [(4'ha):(1'h0)] reg5008 = (1'h0);
  reg [(3'h4):(1'h0)] reg5007 = (1'h0);
  reg [(3'h7):(1'h0)] reg5006 = (1'h0);
  reg [(3'h5):(1'h0)] reg5005 = (1'h0);
  reg [(5'h10):(1'h0)] reg5004 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5003 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5002 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5001 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5000 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4996 = (1'h0);
  reg [(4'h8):(1'h0)] reg4999 = (1'h0);
  reg [(4'ha):(1'h0)] reg4998 = (1'h0);
  reg [(4'ha):(1'h0)] reg4997 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4996 = (1'h0);
  reg [(3'h6):(1'h0)] reg4995 = (1'h0);
  reg [(4'hb):(1'h0)] reg4994 = (1'h0);
  reg [(2'h2):(1'h0)] reg4993 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4992 = (1'h0);
  reg [(3'h4):(1'h0)] reg4991 = (1'h0);
  reg [(5'h10):(1'h0)] reg4990 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4989 = (1'h0);
  reg [(2'h3):(1'h0)] reg4988 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4987 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4986 = (1'h0);
  reg [(4'ha):(1'h0)] reg4985 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4984 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4983 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4982 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4978 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4972 = (1'h0);
  reg [(4'hb):(1'h0)] reg4971 = (1'h0);
  reg [(4'hc):(1'h0)] reg4981 = (1'h0);
  reg [(4'h8):(1'h0)] reg4980 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4979 = (1'h0);
  reg [(3'h4):(1'h0)] reg4978 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4977 = (1'h0);
  reg [(2'h2):(1'h0)] reg4976 = (1'h0);
  reg [(4'hf):(1'h0)] reg4975 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4974 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4973 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4972 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4971 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4970 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire4969;
  wire [(3'h4):(1'h0)] wire4967;
  wire signed [(3'h5):(1'h0)] wire3538;
  reg [(5'h10):(1'h0)] reg1026 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire1027;
  wire signed [(4'hd):(1'h0)] wire1028;
  wire [(4'hb):(1'h0)] wire1029;
  wire [(5'h10):(1'h0)] wire1030;
  wire signed [(4'h9):(1'h0)] wire1031;
  wire [(5'h10):(1'h0)] wire3536;
  assign y = {forvar5501,
                 reg5523,
                 reg5522,
                 reg5521,
                 reg5520,
                 reg5519,
                 forvar5518,
                 reg5517,
                 reg5516,
                 reg5515,
                 reg5514,
                 reg5513,
                 reg5512,
                 forvar5506,
                 forvar5502,
                 reg5511,
                 reg5510,
                 reg5509,
                 forvar5508,
                 reg5507,
                 reg5506,
                 reg5505,
                 reg5504,
                 reg5503,
                 reg5502,
                 reg5501,
                 reg5500,
                 reg5499,
                 forvar5491,
                 reg5495,
                 forvar5493,
                 reg5489,
                 reg5480,
                 reg5488,
                 forvar5478,
                 forvar5469,
                 forvar5468,
                 reg5498,
                 reg5497,
                 reg5496,
                 forvar5495,
                 reg5494,
                 reg5493,
                 reg5492,
                 reg5491,
                 reg5490,
                 forvar5489,
                 forvar5488,
                 reg5487,
                 forvar5484,
                 reg5486,
                 reg5485,
                 reg5484,
                 reg5483,
                 reg5482,
                 reg5481,
                 forvar5480,
                 reg5479,
                 reg5478,
                 reg5477,
                 reg5476,
                 reg5475,
                 forvar5474,
                 reg5473,
                 reg5472,
                 reg5471,
                 reg5470,
                 reg5469,
                 reg5468,
                 reg5460,
                 forvar5459,
                 reg5467,
                 reg5466,
                 reg5465,
                 reg5464,
                 reg5463,
                 reg5462,
                 reg5461,
                 forvar5460,
                 reg5456,
                 forvar5455,
                 reg5459,
                 reg5458,
                 reg5457,
                 forvar5456,
                 reg5455,
                 forvar5454,
                 forvar5441,
                 reg5440,
                 reg5436,
                 forvar5434,
                 forvar5433,
                 forvar5425,
                 reg5432,
                 reg5419,
                 forvar5418,
                 reg5414,
                 reg5412,
                 forvar5411,
                 reg5410,
                 forvar5407,
                 forvar5404,
                 forvar5403,
                 reg5453,
                 reg5452,
                 forvar5451,
                 reg5450,
                 reg5449,
                 forvar5448,
                 forvar5447,
                 reg5446,
                 forvar5445,
                 reg5438,
                 forvar5437,
                 reg5444,
                 reg5443,
                 reg5442,
                 reg5441,
                 forvar5440,
                 reg5439,
                 forvar5438,
                 reg5437,
                 forvar5436,
                 reg5435,
                 reg5434,
                 reg5433,
                 forvar5432,
                 reg5431,
                 reg5430,
                 reg5427,
                 reg5422,
                 reg5429,
                 reg5428,
                 forvar5427,
                 reg5426,
                 reg5425,
                 reg5424,
                 reg5423,
                 forvar5422,
                 reg5421,
                 reg5420,
                 forvar5419,
                 reg5418,
                 reg5417,
                 reg5416,
                 reg5415,
                 forvar5414,
                 reg5413,
                 forvar5412,
                 reg5411,
                 forvar5410,
                 reg5405,
                 reg5402,
                 reg5409,
                 reg5408,
                 reg5407,
                 reg5406,
                 forvar5405,
                 reg5404,
                 reg5403,
                 forvar5402,
                 forvar5401,
                 forvar5394,
                 reg5400,
                 reg5399,
                 reg5398,
                 forvar5397,
                 reg5396,
                 reg5395,
                 reg5394,
                 reg5393,
                 reg5392,
                 forvar5388,
                 reg5391,
                 reg5390,
                 reg5389,
                 reg5388,
                 reg5387,
                 reg5386,
                 reg5385,
                 reg5384,
                 reg5383,
                 reg5382,
                 forvar5381,
                 reg5380,
                 forvar5379,
                 reg5379,
                 forvar5378,
                 reg5377,
                 reg5376,
                 forvar5375,
                 reg5374,
                 forvar5373,
                 reg5372,
                 reg5371,
                 reg5370,
                 reg5369,
                 reg5368,
                 reg5367,
                 reg5366,
                 reg5365,
                 forvar5364,
                 reg5363,
                 forvar5362,
                 reg5361,
                 forvar5360,
                 forvar5359,
                 reg5358,
                 forvar5357,
                 reg5356,
                 reg5355,
                 reg5354,
                 forvar5353,
                 reg5352,
                 reg5351,
                 forvar5349,
                 forvar5346,
                 forvar5341,
                 reg5347,
                 forvar5343,
                 reg5339,
                 forvar5338,
                 reg5350,
                 reg5349,
                 reg5348,
                 forvar5347,
                 reg5346,
                 reg5345,
                 reg5344,
                 reg5343,
                 reg5342,
                 reg5341,
                 reg5340,
                 forvar5339,
                 reg5338,
                 forvar5337,
                 wire5336,
                 reg5335,
                 reg5334,
                 reg5329,
                 reg5333,
                 reg5332,
                 reg5331,
                 reg5330,
                 forvar5329,
                 reg5328,
                 reg5327,
                 reg5326,
                 reg5325,
                 forvar5324,
                 forvar5323,
                 forvar5298,
                 reg5295,
                 reg5294,
                 reg5322,
                 reg5321,
                 reg5320,
                 forvar5319,
                 reg5318,
                 reg5317,
                 reg5316,
                 forvar5315,
                 forvar5314,
                 reg5313,
                 reg5312,
                 reg5311,
                 reg5310,
                 reg5309,
                 reg5308,
                 reg5307,
                 reg5306,
                 forvar5305,
                 reg5304,
                 reg5303,
                 reg5302,
                 forvar5301,
                 reg5300,
                 reg5299,
                 reg5298,
                 reg5297,
                 reg5296,
                 forvar5295,
                 forvar5294,
                 reg5293,
                 forvar5292,
                 wire5291,
                 wire5290,
                 reg5289,
                 forvar5288,
                 reg5287,
                 reg5286,
                 reg5285,
                 reg5284,
                 forvar5282,
                 forvar5278,
                 forvar5271,
                 forvar5270,
                 reg5281,
                 reg5276,
                 forvar5272,
                 reg5283,
                 reg5282,
                 forvar5281,
                 reg5280,
                 reg5279,
                 reg5278,
                 reg5277,
                 forvar5276,
                 reg5275,
                 reg5274,
                 reg5273,
                 reg5272,
                 reg5271,
                 reg5270,
                 reg5269,
                 reg5268,
                 forvar5267,
                 reg5260,
                 reg5255,
                 reg5266,
                 forvar5265,
                 reg5264,
                 reg5263,
                 reg5262,
                 reg5261,
                 forvar5260,
                 reg5259,
                 reg5258,
                 reg5257,
                 reg5256,
                 forvar5255,
                 reg5254,
                 reg5253,
                 forvar5252,
                 forvar5251,
                 reg5250,
                 forvar5249,
                 reg5248,
                 reg5247,
                 reg5246,
                 reg5245,
                 reg5244,
                 reg5243,
                 reg5242,
                 reg5241,
                 forvar5240,
                 forvar5239,
                 forvar5238,
                 reg5237,
                 forvar5236,
                 reg5235,
                 forvar5234,
                 reg5233,
                 reg5232,
                 reg5231,
                 reg5230,
                 reg5229,
                 reg5228,
                 forvar5227,
                 forvar5226,
                 reg5225,
                 reg5224,
                 forvar5223,
                 reg5222,
                 reg5221,
                 reg5220,
                 reg5219,
                 reg5218,
                 reg5217,
                 reg5216,
                 reg5215,
                 reg5214,
                 reg5213,
                 reg5212,
                 reg5211,
                 forvar5210,
                 forvar5209,
                 forvar5208,
                 reg5192,
                 reg5187,
                 forvar5185,
                 forvar5182,
                 reg5207,
                 forvar5206,
                 reg5205,
                 reg5204,
                 reg5203,
                 forvar5202,
                 forvar5201,
                 reg5200,
                 reg5199,
                 reg5198,
                 reg5197,
                 forvar5196,
                 reg5195,
                 reg5194,
                 reg5193,
                 forvar5192,
                 reg5191,
                 reg5190,
                 reg5189,
                 reg5188,
                 forvar5187,
                 reg5186,
                 reg5185,
                 reg5183,
                 reg5184,
                 forvar5183,
                 reg5182,
                 reg5181,
                 reg5180,
                 forvar5179,
                 reg5178,
                 reg5177,
                 reg5176,
                 forvar5175,
                 reg5174,
                 reg5173,
                 forvar5172,
                 reg5171,
                 reg5170,
                 reg5169,
                 reg5168,
                 forvar5167,
                 reg5166,
                 forvar5165,
                 reg5164,
                 reg5163,
                 reg5162,
                 forvar5161,
                 forvar5160,
                 forvar5159,
                 reg5158,
                 reg5157,
                 forvar5156,
                 reg5155,
                 reg5154,
                 reg5153,
                 reg5152,
                 reg5151,
                 reg5150,
                 reg5149,
                 reg5148,
                 forvar5147,
                 reg5146,
                 reg5141,
                 reg5139,
                 reg5145,
                 reg5144,
                 reg5143,
                 reg5142,
                 forvar5141,
                 reg5140,
                 forvar5139,
                 reg5138,
                 reg5137,
                 forvar5136,
                 reg5117,
                 reg5116,
                 reg5135,
                 reg5134,
                 reg5133,
                 reg5132,
                 forvar5131,
                 reg5130,
                 reg5129,
                 reg5128,
                 forvar5127,
                 reg5126,
                 reg5125,
                 reg5124,
                 reg5123,
                 reg5122,
                 reg5121,
                 reg5120,
                 reg5119,
                 reg5118,
                 forvar5117,
                 forvar5116,
                 reg5115,
                 reg5109,
                 reg5106,
                 reg5114,
                 reg5113,
                 reg5112,
                 reg5111,
                 reg5110,
                 forvar5109,
                 reg5108,
                 reg5107,
                 forvar5106,
                 reg5105,
                 reg5104,
                 forvar5103,
                 reg5102,
                 reg5101,
                 reg5100,
                 reg5099,
                 forvar5098,
                 forvar5097,
                 forvar5096,
                 forvar5095,
                 reg5094,
                 reg5093,
                 reg5092,
                 reg5091,
                 forvar5090,
                 forvar5089,
                 forvar5088,
                 forvar5087,
                 reg5086,
                 reg5085,
                 reg5084,
                 reg5083,
                 forvar5082,
                 forvar5081,
                 forvar5080,
                 forvar5079,
                 reg5078,
                 reg5077,
                 reg5076,
                 reg5075,
                 forvar5074,
                 reg5073,
                 reg5072,
                 reg5071,
                 forvar5070,
                 reg5069,
                 reg5068,
                 reg5067,
                 reg5066,
                 reg5065,
                 forvar5064,
                 reg5063,
                 reg5062,
                 forvar5061,
                 forvar5060,
                 reg5059,
                 reg5058,
                 reg5057,
                 reg5056,
                 forvar5055,
                 reg5054,
                 reg5053,
                 reg5052,
                 forvar5051,
                 reg5050,
                 reg5049,
                 reg5048,
                 forvar5047,
                 forvar5046,
                 forvar5045,
                 reg5044,
                 reg5043,
                 forvar5042,
                 reg5041,
                 forvar5040,
                 reg5033,
                 reg5030,
                 reg5039,
                 reg5038,
                 forvar5037,
                 reg5036,
                 reg5035,
                 reg5034,
                 forvar5033,
                 reg5032,
                 reg5031,
                 forvar5030,
                 reg5029,
                 reg5028,
                 reg5027,
                 reg5026,
                 reg5025,
                 forvar5024,
                 reg5023,
                 reg5022,
                 reg5021,
                 reg5020,
                 forvar5019,
                 forvar5018,
                 reg5017,
                 forvar5016,
                 reg5015,
                 reg5014,
                 reg5013,
                 reg5012,
                 forvar5011,
                 reg5010,
                 reg5009,
                 reg5008,
                 reg5007,
                 reg5006,
                 reg5005,
                 reg5004,
                 reg5003,
                 forvar5002,
                 forvar5001,
                 reg5000,
                 reg4996,
                 reg4999,
                 reg4998,
                 reg4997,
                 forvar4996,
                 reg4995,
                 reg4994,
                 reg4993,
                 reg4992,
                 reg4991,
                 reg4990,
                 forvar4989,
                 reg4988,
                 forvar4987,
                 forvar4986,
                 reg4985,
                 reg4984,
                 forvar4983,
                 forvar4982,
                 forvar4978,
                 forvar4972,
                 reg4971,
                 reg4981,
                 reg4980,
                 reg4979,
                 reg4978,
                 reg4977,
                 reg4976,
                 reg4975,
                 reg4974,
                 reg4973,
                 reg4972,
                 forvar4971,
                 forvar4970,
                 wire4969,
                 wire4967,
                 wire3538,
                 reg1026,
                 wire1027,
                 wire1028,
                 wire1029,
                 wire1030,
                 wire1031,
                 wire3536,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1026 <= ($unsigned(wire1025) ?
          (|wire1022[(4'h8):(1'h1)]) : {((+wire1024) >= $unsigned(wire1025))});
    end
  assign wire1027 = ($signed((wire1022[(3'h4):(1'h0)] ?
                        wire1023[(3'h7):(3'h4)] : (~^wire1024))) ^~ (!reg1026));
  assign wire1028 = $signed(reg1026);
  assign wire1029 = wire1025[(1'h1):(1'h0)];
  assign wire1030 = (wire1025[(3'h5):(1'h0)] << ((reg1026[(1'h1):(1'h0)] * ((8'h9f) ?
                        wire1029 : wire1029)) > (8'hb9)));
  assign wire1031 = wire1029;
  module1032 modinst3537 (wire3536, clk, wire1025, wire1027, wire1031, wire1028, wire1030);
  assign wire3538 = (wire1022 ?
                        (~&({(8'hac)} ?
                            wire1024 : (^~wire1024))) : ((~&(~wire1029)) ?
                            $unsigned((|wire1028)) : ((wire1024 > (8'hb2)) ?
                                (wire1027 ?
                                    wire1029 : wire1025) : (-wire1022))));
  module3539 modinst4968 (.y(wire4967), .wire3540(wire1023), .wire3543(wire3536), .wire3541(reg1026), .clk(clk), .wire3542(wire1029));
  assign wire4969 = wire3536;
  always
    @(posedge clk) begin
      for (forvar4970 = (1'h0); (forvar4970 < (1'h0)); forvar4970 = (forvar4970 + (1'h1)))
        begin
          if ($unsigned($signed($unsigned(wire4969))))
            begin
              if ($signed(wire1029[(1'h1):(1'h1)]))
                begin
                  for (forvar4971 = (1'h0); (forvar4971 < (1'h1)); forvar4971 = (forvar4971 + (1'h1)))
                    begin
                      reg4972 <= (wire1024[(2'h2):(2'h2)] ?
                          wire4969[(3'h7):(3'h7)] : (wire3536[(4'hc):(4'ha)] <= ((|wire1023) ?
                              $signed(forvar4971) : wire1024)));
                    end
                  if (((($unsigned(wire3536) ^~ (wire1030 - wire1031)) == wire1031) <= wire3538[(3'h5):(3'h4)]))
                    begin
                      reg4973 <= reg4972[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg4973 <= (((^$unsigned((8'hb2))) ~^ wire4969) ?
                          ((wire1022 ? $signed((8'hb9)) : $unsigned(wire3536)) ?
                              wire1025 : ({reg4972} >>> reg4972[(3'h5):(3'h4)])) : (reg1026[(4'hf):(3'h6)] >= (reg4972[(3'h6):(1'h0)] ?
                              (~wire1030) : ((8'hba) ? wire1028 : reg4973))));
                      reg4974 <= $unsigned(forvar4971[(3'h5):(2'h2)]);
                      reg4975 <= forvar4970;
                      reg4976 <= $unsigned((wire3538 ^~ reg4975[(1'h0):(1'h0)]));
                    end
                  if (wire1031)
                    begin
                      reg4977 <= $signed(((8'hb7) ?
                          ((~|wire1024) ?
                              (wire1024 ?
                                  reg4976 : wire1031) : $signed(wire3536)) : reg4972));
                      reg4978 <= wire3538;
                      reg4979 <= $signed(forvar4970);
                      reg4980 <= (-(~&{$signed(reg4974)}));
                    end
                  else
                    begin
                      reg4977 <= (~(wire1025[(3'h7):(3'h7)] <= $signed(wire1025)));
                      reg4978 <= (wire1030 ?
                          wire1022 : $signed({wire1025[(3'h6):(1'h1)]}));
                      reg4979 <= ($signed((wire1027[(4'ha):(4'ha)] ?
                          wire3538 : (~^wire1024))) != (8'hb5));
                      reg4980 <= wire1030;
                    end
                  reg4981 <= forvar4970[(3'h4):(1'h1)];
                end
              else
                begin
                  if (($unsigned(reg4972) ?
                      ($signed(reg4980) ?
                          reg4973 : ($unsigned(reg4981) ?
                              wire3536[(4'h9):(4'h8)] : $signed(wire1022))) : ((~(wire3538 ?
                          reg1026 : reg4981)) <= ((wire1028 ?
                          (8'ha1) : wire1027) << (wire1031 > wire1024)))))
                    begin
                      reg4971 <= wire3538;
                    end
                  else
                    begin
                      reg4971 <= wire1028;
                      reg4972 <= ((~&(~reg4974[(4'hf):(4'h8)])) ?
                          wire3538 : wire1025[(2'h3):(1'h1)]);
                    end
                end
            end
          else
            begin
              if ((|$unsigned((forvar4970[(2'h2):(1'h1)] << (wire1022 <= forvar4970)))))
                begin
                  reg4971 <= reg4974;
                  for (forvar4972 = (1'h0); (forvar4972 < (1'h0)); forvar4972 = (forvar4972 + (1'h1)))
                    begin
                      reg4973 <= $signed(reg4973);
                      reg4974 <= ($unsigned((+$unsigned(reg4980))) | ((^~(8'hb7)) || (reg4979[(1'h0):(1'h0)] >> $signed(wire1031))));
                      reg4975 <= reg4971;
                      reg4976 <= $signed((((~&wire1028) ?
                              wire1024[(3'h4):(1'h0)] : $unsigned(reg1026)) ?
                          ({reg1026} << (reg4977 >> reg4973)) : reg4972[(3'h4):(1'h1)]));
                    end
                  reg4977 <= wire1023;
                  for (forvar4978 = (1'h0); (forvar4978 < (1'h1)); forvar4978 = (forvar4978 + (1'h1)))
                    begin
                      reg4979 <= $unsigned(($signed(forvar4978[(1'h0):(1'h0)]) ^ ((^(8'ha9)) ?
                          (wire3538 ?
                              (8'hb0) : wire4969) : (wire1028 >>> reg1026))));
                      reg4980 <= ($unsigned(wire1030[(5'h10):(4'hb)]) >= reg4981[(2'h2):(1'h1)]);
                    end
                end
              else
                begin
                  if ($unsigned({$unsigned((~reg4978))}))
                    begin
                      reg4971 <= $signed((+$unsigned(((8'haf) > forvar4971))));
                      reg4972 <= {reg4977[(4'h9):(2'h3)]};
                    end
                  else
                    begin
                      reg4971 <= ($signed(forvar4971) - reg4980[(3'h6):(1'h1)]);
                      reg4972 <= $signed(wire3538[(1'h0):(1'h0)]);
                    end
                  if ($signed((|reg1026[(4'h8):(2'h3)])))
                    begin
                      reg4973 <= $signed((($signed(wire1029) | $unsigned(wire1022)) ?
                          (8'hb5) : wire3536));
                      reg4974 <= wire1028;
                      reg4975 <= (($unsigned((reg4973 ?
                              reg4973 : wire1029)) ~^ (-$signed(wire1022))) ?
                          $signed(wire1023[(3'h6):(2'h3)]) : $unsigned(((!reg4977) ?
                              (^~reg4981) : {reg4975})));
                    end
                  else
                    begin
                      reg4973 <= {{{wire3538}}};
                      reg4974 <= $signed($unsigned(wire3536[(3'h4):(1'h1)]));
                      reg4975 <= $signed(($signed($unsigned(reg1026)) ?
                          ((-(8'hb5)) & $unsigned(reg4975)) : ($signed((8'ha7)) ?
                              (reg1026 ?
                                  wire4967 : wire1024) : (reg4977 >>> wire1025))));
                      reg4976 <= {(8'ha0)};
                    end
                  reg4977 <= (($unsigned($unsigned(wire1028)) ?
                      {$unsigned(wire1030)} : (((8'hae) * reg4975) <= (~^wire3536))) <= (^$unsigned($unsigned(forvar4978))));
                end
            end
          for (forvar4982 = (1'h0); (forvar4982 < (1'h1)); forvar4982 = (forvar4982 + (1'h1)))
            begin
              for (forvar4983 = (1'h0); (forvar4983 < (2'h2)); forvar4983 = (forvar4983 + (1'h1)))
                begin
                  if (reg1026[(3'h5):(3'h5)])
                    begin
                      reg4984 <= $signed((wire1023 ?
                          {$signed(reg1026)} : {$unsigned(reg4981)}));
                      reg4985 <= $signed(forvar4971);
                    end
                  else
                    begin
                      reg4984 <= $unsigned((&(~reg4978)));
                      reg4985 <= (($signed((reg4974 >= forvar4983)) & reg4980) < $signed(forvar4978));
                    end
                end
              for (forvar4986 = (1'h0); (forvar4986 < (2'h2)); forvar4986 = (forvar4986 + (1'h1)))
                begin
                  for (forvar4987 = (1'h0); (forvar4987 < (1'h0)); forvar4987 = (forvar4987 + (1'h1)))
                    begin
                      reg4988 <= reg4972[(3'h6):(2'h2)];
                    end
                  for (forvar4989 = (1'h0); (forvar4989 < (1'h0)); forvar4989 = (forvar4989 + (1'h1)))
                    begin
                      reg4990 <= ($unsigned(forvar4978[(2'h3):(1'h0)]) ?
                          ($unsigned((+reg4980)) ?
                              ((^~reg4980) ?
                                  ((8'ha2) ?
                                      forvar4970 : reg4971) : {reg4981}) : $signed($signed(wire1025))) : (reg4984 * {((8'hac) ?
                                  wire3536 : reg4988)}));
                      reg4991 <= $unsigned({reg4979});
                    end
                  reg4992 <= $signed(reg4980);
                  reg4993 <= (forvar4978 ?
                      (^($signed(reg4985) ?
                          (|reg4971) : wire1025[(2'h2):(1'h1)])) : (|(8'h9e)));
                end
              if (({wire1025} & (~|(8'hac))))
                begin
                  if (wire1023[(4'hf):(4'h8)])
                    begin
                      reg4994 <= $signed(forvar4983[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg4994 <= reg4981;
                      reg4995 <= wire1031[(1'h1):(1'h1)];
                    end
                  for (forvar4996 = (1'h0); (forvar4996 < (1'h0)); forvar4996 = (forvar4996 + (1'h1)))
                    begin
                      reg4997 <= (($unsigned((+wire1031)) ?
                          $unsigned($signed(reg4992)) : {$signed(reg4995)}) >> forvar4971[(3'h7):(1'h1)]);
                      reg4998 <= (^{reg4990});
                      reg4999 <= forvar4987;
                    end
                end
              else
                begin
                  if ((wire1030[(1'h0):(1'h0)] ^~ $signed(reg4977)))
                    begin
                      reg4994 <= ($signed(reg4981[(4'hb):(2'h2)]) ?
                          $signed($unsigned({wire1022})) : (((8'hb1) << $unsigned(reg4977)) >>> ({wire1029} << (!(8'ha1)))));
                      reg4995 <= (8'hb3);
                      reg4996 <= $signed(wire1030);
                    end
                  else
                    begin
                      reg4994 <= (~reg4998);
                      reg4995 <= reg4981[(3'h4):(1'h0)];
                    end
                  if (forvar4970[(4'h9):(1'h1)])
                    begin
                      reg4997 <= reg4997;
                      reg4998 <= {(reg4998[(3'h5):(3'h4)] ?
                              reg4994 : $unsigned($unsigned(reg4979)))};
                      reg4999 <= $signed((forvar4972 ?
                          (-(forvar4972 ?
                              wire4969 : reg4978)) : $unsigned((reg4978 ?
                              reg4984 : wire1031))));
                    end
                  else
                    begin
                      reg4997 <= $unsigned(reg4976[(1'h0):(1'h0)]);
                      reg4998 <= {wire1025};
                      reg4999 <= $unsigned(reg4993);
                      reg5000 <= $unsigned($signed((+$signed(forvar4982))));
                    end
                end
              for (forvar5001 = (1'h0); (forvar5001 < (2'h2)); forvar5001 = (forvar5001 + (1'h1)))
                begin
                  for (forvar5002 = (1'h0); (forvar5002 < (1'h1)); forvar5002 = (forvar5002 + (1'h1)))
                    begin
                      reg5003 <= $signed((({forvar4983} ?
                              $signed((8'hb4)) : reg4977) ?
                          $unsigned((reg4975 * (8'ha3))) : reg4985[(3'h5):(3'h5)]));
                      reg5004 <= forvar4972[(3'h5):(2'h2)];
                      reg5005 <= $signed(($signed({reg4979}) << (+(forvar4987 ?
                          reg4990 : (8'haa)))));
                      reg5006 <= {reg5005};
                    end
                  if (((&$signed(wire1024[(2'h3):(2'h2)])) ?
                      {reg4993} : reg4999[(3'h6):(3'h6)]))
                    begin
                      reg5007 <= (!(($unsigned(reg4985) <= $signed(wire1031)) ?
                          $unsigned({wire4969}) : reg4981[(3'h6):(3'h5)]));
                      reg5008 <= (&($signed(wire1024) && ((reg4977 ?
                          reg1026 : wire1028) >> (8'ha3))));
                    end
                  else
                    begin
                      reg5007 <= reg4994;
                      reg5008 <= $unsigned($signed(reg4992[(1'h0):(1'h0)]));
                      reg5009 <= reg5004[(4'h9):(4'h8)];
                      reg5010 <= $signed(($signed(forvar4978[(1'h1):(1'h1)]) ?
                          ((forvar5001 ? reg4985 : reg4978) ?
                              reg4993 : reg4979) : reg4991[(2'h2):(2'h2)]));
                    end
                  for (forvar5011 = (1'h0); (forvar5011 < (2'h3)); forvar5011 = (forvar5011 + (1'h1)))
                    begin
                      reg5012 <= (~&((reg4984[(3'h4):(3'h4)] ?
                              (|reg4991) : (~reg4995)) ?
                          reg4976[(1'h1):(1'h0)] : {(~|forvar5001)}));
                      reg5013 <= $unsigned($unsigned((^~wire4967[(2'h3):(2'h2)])));
                      reg5014 <= reg4978[(2'h3):(2'h3)];
                      reg5015 <= $unsigned(($unsigned({forvar4996}) <<< wire1022[(4'h9):(1'h0)]));
                    end
                  for (forvar5016 = (1'h0); (forvar5016 < (2'h3)); forvar5016 = (forvar5016 + (1'h1)))
                    begin
                      reg5017 <= $unsigned((8'ha0));
                    end
                end
            end
          for (forvar5018 = (1'h0); (forvar5018 < (1'h0)); forvar5018 = (forvar5018 + (1'h1)))
            begin
              for (forvar5019 = (1'h0); (forvar5019 < (2'h2)); forvar5019 = (forvar5019 + (1'h1)))
                begin
                  if ({(+$signed(((8'ha2) ? forvar5016 : reg4976)))})
                    begin
                      reg5020 <= ($signed($unsigned(((8'hab) ?
                              wire1030 : wire1023))) ?
                          $signed($unsigned(reg4985[(2'h3):(2'h2)])) : (({reg5012} > $signed(reg4973)) ?
                              ($unsigned(forvar4971) ?
                                  (^reg4991) : reg4979) : ({wire4969} || (&reg4997))));
                      reg5021 <= reg4978[(3'h4):(1'h0)];
                      reg5022 <= (^($unsigned($signed(wire1030)) != $signed(forvar5002)));
                      reg5023 <= {wire1023};
                    end
                  else
                    begin
                      reg5020 <= ($signed((reg5007 <<< {reg4980})) ?
                          wire1024[(2'h3):(2'h2)] : forvar5018[(2'h2):(1'h0)]);
                      reg5021 <= (^$signed(forvar5016));
                    end
                  for (forvar5024 = (1'h0); (forvar5024 < (2'h2)); forvar5024 = (forvar5024 + (1'h1)))
                    begin
                      reg5025 <= ((reg1026[(1'h0):(1'h0)] ?
                          reg5017 : reg5012) * $unsigned(reg5013[(3'h4):(3'h4)]));
                    end
                  if ((((forvar5019[(4'he):(4'h8)] >>> $signed(reg4975)) ^ reg5010) - (~&$signed((!reg5013)))))
                    begin
                      reg5026 <= $unsigned($unsigned((&(reg5012 >> reg4995))));
                    end
                  else
                    begin
                      reg5026 <= (|((!forvar4978[(3'h4):(2'h3)]) <= (!(reg4991 == (8'hab)))));
                      reg5027 <= ((+(8'ha3)) ?
                          wire1031[(2'h3):(2'h2)] : {$signed($unsigned((8'hac)))});
                      reg5028 <= ($signed($unsigned($signed((8'had)))) ?
                          reg4999 : (reg4972 ?
                              reg5017[(2'h2):(1'h0)] : reg4981[(3'h4):(2'h2)]));
                      reg5029 <= {(&reg4984)};
                    end
                end
              if ($signed({(&{reg4975})}))
                begin
                  for (forvar5030 = (1'h0); (forvar5030 < (2'h3)); forvar5030 = (forvar5030 + (1'h1)))
                    begin
                      reg5031 <= $unsigned(forvar4970[(1'h0):(1'h0)]);
                      reg5032 <= ((!(8'hb8)) < $unsigned({wire4969}));
                    end
                  for (forvar5033 = (1'h0); (forvar5033 < (1'h1)); forvar5033 = (forvar5033 + (1'h1)))
                    begin
                      reg5034 <= $unsigned($signed((!reg5026)));
                      reg5035 <= forvar4986;
                      reg5036 <= (!((^(8'hb3)) ?
                          (-wire1029) : (reg5013 - ((8'ha6) ?
                              wire1030 : reg4991))));
                    end
                  for (forvar5037 = (1'h0); (forvar5037 < (2'h2)); forvar5037 = (forvar5037 + (1'h1)))
                    begin
                      reg5038 <= reg4977;
                    end
                  reg5039 <= (!wire4969[(4'hb):(1'h1)]);
                end
              else
                begin
                  if ((|($unsigned($unsigned(wire1023)) ~^ $signed((~(8'hb6))))))
                    begin
                      reg5030 <= ($unsigned($signed((forvar4986 || (8'h9e)))) ?
                          $signed((reg5025[(1'h1):(1'h0)] ?
                              $unsigned(reg4997) : $unsigned((8'h9d)))) : $signed(forvar4983[(1'h0):(1'h0)]));
                      reg5031 <= $signed((reg5035[(2'h2):(1'h0)] ?
                          ((^~(8'hb2)) >>> (forvar5001 == reg5013)) : {reg4977[(4'h8):(3'h6)]}));
                      reg5032 <= $signed(reg4995[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg5030 <= reg5008[(3'h6):(3'h6)];
                    end
                  reg5033 <= (^~{reg4978[(3'h4):(2'h3)]});
                end
              for (forvar5040 = (1'h0); (forvar5040 < (2'h3)); forvar5040 = (forvar5040 + (1'h1)))
                begin
                  reg5041 <= reg5028;
                  for (forvar5042 = (1'h0); (forvar5042 < (2'h3)); forvar5042 = (forvar5042 + (1'h1)))
                    begin
                      reg5043 <= (((reg5004[(4'hc):(4'hb)] ?
                              $unsigned(forvar5016) : ((8'hb8) && (8'hb6))) ?
                          forvar5002 : $unsigned(reg4979)) + reg4971[(4'hb):(3'h6)]);
                      reg5044 <= forvar5002[(4'ha):(4'h9)];
                    end
                end
            end
        end
      for (forvar5045 = (1'h0); (forvar5045 < (1'h1)); forvar5045 = (forvar5045 + (1'h1)))
        begin
          for (forvar5046 = (1'h0); (forvar5046 < (1'h1)); forvar5046 = (forvar5046 + (1'h1)))
            begin
              for (forvar5047 = (1'h0); (forvar5047 < (2'h2)); forvar5047 = (forvar5047 + (1'h1)))
                begin
                  if ((~{{$unsigned((8'hb5))}}))
                    begin
                      reg5048 <= (!({$signed(reg5044)} ^~ (|{reg5034})));
                      reg5049 <= forvar5045[(3'h5):(2'h3)];
                      reg5050 <= $signed(forvar4971[(3'h7):(3'h6)]);
                    end
                  else
                    begin
                      reg5048 <= (|$unsigned(reg5049));
                      reg5049 <= $unsigned($unsigned(reg4972));
                      reg5050 <= {(~&{$unsigned((8'hb5))})};
                    end
                end
              for (forvar5051 = (1'h0); (forvar5051 < (2'h3)); forvar5051 = (forvar5051 + (1'h1)))
                begin
                  if ((({wire1023[(4'h8):(2'h3)]} ?
                          (~(8'hac)) : $unsigned((reg5041 | (8'ha1)))) ?
                      forvar5045[(3'h4):(3'h4)] : (~$unsigned(wire1022[(1'h1):(1'h0)]))))
                    begin
                      reg5052 <= reg5027;
                      reg5053 <= reg5041[(4'ha):(1'h1)];
                    end
                  else
                    begin
                      reg5052 <= $unsigned((reg4978[(1'h0):(1'h0)] ?
                          (~(~^(8'h9e))) : ($unsigned(reg4996) >= $unsigned(reg5039))));
                      reg5053 <= $signed(($unsigned((reg4994 >= reg4997)) <<< reg5014[(1'h1):(1'h1)]));
                      reg5054 <= reg4972[(1'h1):(1'h1)];
                    end
                  for (forvar5055 = (1'h0); (forvar5055 < (1'h0)); forvar5055 = (forvar5055 + (1'h1)))
                    begin
                      reg5056 <= ((|forvar5019[(4'h8):(3'h4)]) ?
                          (|forvar5002[(4'ha):(3'h4)]) : reg4991);
                      reg5057 <= (~|{$unsigned((reg5027 < (8'ha5)))});
                      reg5058 <= forvar5016[(4'h8):(1'h1)];
                      reg5059 <= $signed((8'haf));
                    end
                end
              for (forvar5060 = (1'h0); (forvar5060 < (2'h3)); forvar5060 = (forvar5060 + (1'h1)))
                begin
                  for (forvar5061 = (1'h0); (forvar5061 < (1'h1)); forvar5061 = (forvar5061 + (1'h1)))
                    begin
                      reg5062 <= (reg4984 ?
                          $unsigned((+forvar4972)) : $signed((~^(&reg5054))));
                      reg5063 <= wire4969;
                    end
                  for (forvar5064 = (1'h0); (forvar5064 < (2'h3)); forvar5064 = (forvar5064 + (1'h1)))
                    begin
                      reg5065 <= (($unsigned((8'hb3)) ^ {{reg5014}}) ?
                          ({{reg5038}} ?
                              forvar4987 : forvar5047) : reg4994[(3'h6):(1'h1)]);
                      reg5066 <= $unsigned(reg5003[(3'h7):(3'h6)]);
                      reg5067 <= (~&$signed(reg5057[(3'h4):(3'h4)]));
                      reg5068 <= (reg5008 == (reg5033[(1'h1):(1'h1)] ?
                          forvar5033[(3'h4):(1'h0)] : ((forvar5040 ?
                              wire1027 : reg4999) * reg5028)));
                    end
                  reg5069 <= reg5012[(3'h7):(3'h7)];
                end
              for (forvar5070 = (1'h0); (forvar5070 < (1'h1)); forvar5070 = (forvar5070 + (1'h1)))
                begin
                  reg5071 <= (reg5044 > reg5063);
                  reg5072 <= (wire1031[(3'h5):(2'h2)] <<< $signed((^$signed(wire3538))));
                  reg5073 <= (reg4990[(4'hb):(3'h4)] >>> {{{(8'h9e)}}});
                  for (forvar5074 = (1'h0); (forvar5074 < (1'h1)); forvar5074 = (forvar5074 + (1'h1)))
                    begin
                      reg5075 <= reg5023;
                      reg5076 <= (forvar5019[(3'h5):(3'h5)] ^~ $unsigned(reg4971[(4'ha):(4'h8)]));
                    end
                end
            end
          reg5077 <= wire1022;
          reg5078 <= reg5014[(4'h8):(3'h4)];
        end
      for (forvar5079 = (1'h0); (forvar5079 < (2'h2)); forvar5079 = (forvar5079 + (1'h1)))
        begin
          for (forvar5080 = (1'h0); (forvar5080 < (1'h1)); forvar5080 = (forvar5080 + (1'h1)))
            begin
              for (forvar5081 = (1'h0); (forvar5081 < (1'h0)); forvar5081 = (forvar5081 + (1'h1)))
                begin
                  for (forvar5082 = (1'h0); (forvar5082 < (1'h1)); forvar5082 = (forvar5082 + (1'h1)))
                    begin
                      reg5083 <= ((+$unsigned(reg5039[(3'h6):(3'h4)])) ?
                          reg5039[(3'h6):(2'h2)] : (|(+(forvar4971 ?
                              reg5021 : (8'haf)))));
                    end
                  reg5084 <= ($signed((|$unsigned(forvar5081))) ~^ ($unsigned({reg5050}) ?
                      ({reg4972} | reg5012) : ((^reg5028) | {reg4988})));
                  reg5085 <= $unsigned((((8'hab) ?
                      (~^reg5033) : reg5063[(1'h1):(1'h0)]) ~^ $signed((8'h9e))));
                  reg5086 <= wire1031[(1'h0):(1'h0)];
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar5087 = (1'h0); (forvar5087 < (2'h2)); forvar5087 = (forvar5087 + (1'h1)))
        begin
          for (forvar5088 = (1'h0); (forvar5088 < (2'h2)); forvar5088 = (forvar5088 + (1'h1)))
            begin
              for (forvar5089 = (1'h0); (forvar5089 < (1'h1)); forvar5089 = (forvar5089 + (1'h1)))
                begin
                  for (forvar5090 = (1'h0); (forvar5090 < (1'h0)); forvar5090 = (forvar5090 + (1'h1)))
                    begin
                      reg5091 <= reg5005[(2'h3):(1'h0)];
                      reg5092 <= (reg5072 ? reg5009 : {reg5017[(3'h6):(3'h4)]});
                      reg5093 <= forvar4987[(1'h0):(1'h0)];
                      reg5094 <= reg5015[(3'h6):(1'h0)];
                    end
                end
            end
        end
      for (forvar5095 = (1'h0); (forvar5095 < (2'h2)); forvar5095 = (forvar5095 + (1'h1)))
        begin
          for (forvar5096 = (1'h0); (forvar5096 < (2'h3)); forvar5096 = (forvar5096 + (1'h1)))
            begin
              for (forvar5097 = (1'h0); (forvar5097 < (2'h3)); forvar5097 = (forvar5097 + (1'h1)))
                begin
                  for (forvar5098 = (1'h0); (forvar5098 < (2'h3)); forvar5098 = (forvar5098 + (1'h1)))
                    begin
                      reg5099 <= (~^(~|forvar4982[(1'h0):(1'h0)]));
                      reg5100 <= $signed(reg4999);
                      reg5101 <= (({{forvar4987}} - $unsigned({forvar5001})) ?
                          ((forvar5030 || (^reg5059)) > {forvar5095[(4'he):(3'h4)]}) : ({reg5043[(4'hb):(1'h0)]} ?
                              $unsigned($unsigned((8'hba))) : ($unsigned(reg5028) >= reg5027[(4'h8):(1'h0)])));
                      reg5102 <= {((((8'ha0) ?
                              (8'ha9) : reg5034) == {reg5058}) >= $unsigned((reg5050 ?
                              reg4985 : reg5000)))};
                    end
                end
              if ((|(8'hb5)))
                begin
                  for (forvar5103 = (1'h0); (forvar5103 < (2'h3)); forvar5103 = (forvar5103 + (1'h1)))
                    begin
                      reg5104 <= ({(~^$signed(reg5067))} <= (reg5068[(1'h1):(1'h1)] | (reg5071[(1'h0):(1'h0)] > $unsigned((8'hb6)))));
                      reg5105 <= reg5053;
                    end
                  for (forvar5106 = (1'h0); (forvar5106 < (2'h3)); forvar5106 = (forvar5106 + (1'h1)))
                    begin
                      reg5107 <= reg5022;
                      reg5108 <= $signed(reg4996);
                    end
                  for (forvar5109 = (1'h0); (forvar5109 < (1'h1)); forvar5109 = (forvar5109 + (1'h1)))
                    begin
                      reg5110 <= (~reg5100);
                    end
                  if (reg5059[(3'h7):(3'h5)])
                    begin
                      reg5111 <= {(reg5054[(3'h4):(2'h2)] ?
                              ($signed((8'hba)) <<< (reg5091 | forvar5109)) : (&$unsigned(forvar5089)))};
                      reg5112 <= $signed($unsigned((reg5036 >>> reg5021[(3'h5):(2'h3)])));
                      reg5113 <= $signed((($signed(reg4998) ?
                              (8'hb4) : (reg5085 ~^ reg5004)) ?
                          $signed(((8'hb3) >>> reg5054)) : $signed((8'hb7))));
                    end
                  else
                    begin
                      reg5111 <= {(~&reg5102)};
                      reg5112 <= $unsigned($signed(($signed(forvar4989) > {forvar4978})));
                      reg5113 <= $unsigned((^(forvar4989[(1'h1):(1'h1)] - reg5107)));
                      reg5114 <= (-$unsigned(($signed(reg5026) != (reg5032 & (8'ha3)))));
                    end
                end
              else
                begin
                  for (forvar5103 = (1'h0); (forvar5103 < (1'h0)); forvar5103 = (forvar5103 + (1'h1)))
                    begin
                      reg5104 <= ({$unsigned((reg5102 & (8'hae)))} != (~^($signed((8'ha1)) ?
                          reg5036 : wire1029)));
                      reg5105 <= $signed(wire1029);
                      reg5106 <= ((|(forvar5098[(1'h1):(1'h0)] ?
                              {reg5108} : (forvar5090 ?
                                  forvar5079 : (8'hb9)))) ?
                          $signed({$unsigned(reg4985)}) : $signed((forvar5033[(1'h1):(1'h0)] ?
                              $signed(reg4990) : $unsigned(wire4967))));
                    end
                  if ((~$signed({$signed((8'hba))})))
                    begin
                      reg5107 <= ({wire1023[(4'h8):(2'h2)]} ?
                          reg5054[(3'h6):(2'h3)] : reg5044[(3'h6):(2'h2)]);
                      reg5108 <= $signed(forvar5055[(3'h5):(3'h5)]);
                    end
                  else
                    begin
                      reg5107 <= $unsigned($unsigned($signed(reg5033[(1'h0):(1'h0)])));
                      reg5108 <= $unsigned($signed(($unsigned(reg4988) | $signed(forvar4970))));
                    end
                  if ((((|reg5029[(2'h2):(1'h0)]) <= ((+reg4978) ^ (reg5108 ?
                          forvar5011 : reg5058))) ?
                      ($signed((^~reg5000)) ?
                          ($unsigned(forvar5060) ?
                              (~^wire1022) : $signed((8'hb5))) : (reg5099[(2'h2):(1'h1)] != $signed(forvar5040))) : wire1025))
                    begin
                      reg5109 <= $unsigned($signed(forvar5037));
                      reg5110 <= (~{(~(reg5007 ? wire1027 : reg5014))});
                    end
                  else
                    begin
                      reg5109 <= ($unsigned(reg5099[(1'h1):(1'h0)]) ?
                          (~^wire1024) : {{reg5073}});
                      reg5110 <= reg5106[(1'h1):(1'h0)];
                      reg5111 <= reg4972;
                      reg5112 <= {$unsigned(wire3536[(1'h0):(1'h0)])};
                    end
                  if ((($unsigned($signed(forvar4982)) ^ {forvar5088}) << (&$signed(forvar5080))))
                    begin
                      reg5113 <= {forvar5042};
                      reg5114 <= (!$unsigned(((8'hb0) & ((8'h9e) ?
                          (8'hae) : reg5072))));
                      reg5115 <= (|(~{(forvar5024 ? reg5083 : reg5015)}));
                    end
                  else
                    begin
                      reg5113 <= $signed(reg5100[(3'h4):(1'h1)]);
                      reg5114 <= {(!((wire1025 ?
                              forvar4989 : forvar5018) >= reg4971[(3'h7):(1'h0)]))};
                    end
                end
            end
          if (reg5003[(1'h1):(1'h0)])
            begin
              for (forvar5116 = (1'h0); (forvar5116 < (1'h1)); forvar5116 = (forvar5116 + (1'h1)))
                begin
                  for (forvar5117 = (1'h0); (forvar5117 < (2'h2)); forvar5117 = (forvar5117 + (1'h1)))
                    begin
                      reg5118 <= (^$signed(((8'ha8) ^ $signed(reg4996))));
                      reg5119 <= (reg5027[(2'h3):(1'h1)] + {$signed(forvar4989)});
                      reg5120 <= ((forvar4971[(4'hd):(4'hc)] ?
                              (8'ha6) : (8'hb1)) ?
                          $unsigned((reg5030[(3'h5):(3'h5)] >> $signed(wire1022))) : ($signed({forvar5033}) || ((reg4996 ?
                              reg4977 : reg5091) ~^ $signed(forvar4987))));
                      reg5121 <= {(8'ha0)};
                    end
                  if (reg5043[(2'h3):(1'h1)])
                    begin
                      reg5122 <= reg4981[(3'h5):(2'h3)];
                      reg5123 <= $signed({$unsigned((&reg5071))});
                      reg5124 <= $unsigned(forvar5047[(4'hb):(4'ha)]);
                      reg5125 <= (reg5093[(4'hc):(4'hc)] ?
                          (({reg5052} & reg5052) != ({reg5119} ?
                              $unsigned(forvar5030) : reg5007)) : ((~^(forvar5109 & reg5049)) >>> $unsigned(reg5029)));
                    end
                  else
                    begin
                      reg5122 <= (+{$signed((reg5014 || wire3538))});
                      reg5123 <= reg5059[(2'h2):(1'h1)];
                      reg5124 <= {($signed($signed(forvar5060)) + forvar5033[(2'h2):(2'h2)])};
                      reg5125 <= ($signed(((8'ha2) <<< wire1027)) ?
                          (((^forvar5080) ?
                              (~^reg5012) : reg4993) <<< (-(reg5027 ^ reg5077))) : $unsigned((~^{reg4993})));
                    end
                  reg5126 <= {((8'ha3) < $unsigned($signed(reg5029)))};
                  for (forvar5127 = (1'h0); (forvar5127 < (2'h2)); forvar5127 = (forvar5127 + (1'h1)))
                    begin
                      reg5128 <= $unsigned($signed($signed(reg4990[(4'hf):(3'h7)])));
                      reg5129 <= (^(~|(forvar5040 ?
                          (~|forvar5079) : $unsigned(reg5020))));
                      reg5130 <= (forvar5016 * reg5105);
                    end
                end
              for (forvar5131 = (1'h0); (forvar5131 < (2'h3)); forvar5131 = (forvar5131 + (1'h1)))
                begin
                  if ((((-$signed(forvar5042)) ?
                          $signed((reg1026 ?
                              reg5028 : forvar5088)) : {reg5125[(2'h3):(1'h1)]}) ?
                      (^$signed((reg4980 ~^ reg5077))) : (-$unsigned({wire1023}))))
                    begin
                      reg5132 <= reg5105;
                      reg5133 <= (8'ha6);
                      reg5134 <= ((8'h9f) * (-(!(reg5004 >> forvar5097))));
                    end
                  else
                    begin
                      reg5132 <= $unsigned(({forvar4972[(2'h3):(2'h2)]} ?
                          ((reg5025 ? forvar5037 : forvar5001) ?
                              forvar5127[(1'h0):(1'h0)] : reg5027) : (wire1024[(2'h2):(1'h1)] ?
                              forvar4987 : {(8'ha3)})));
                    end
                end
              reg5135 <= $unsigned(($unsigned($signed(forvar5087)) >> reg5035[(2'h3):(1'h0)]));
            end
          else
            begin
              reg5116 <= {{$unsigned($signed((8'hb6)))}};
              reg5117 <= ((-{wire1030[(4'hd):(3'h7)]}) ?
                  (forvar5045[(1'h0):(1'h0)] > (+((8'hb9) ^~ (8'hac)))) : {((~(8'hb8)) ?
                          forvar5117[(3'h7):(2'h3)] : {reg4988})});
            end
          for (forvar5136 = (1'h0); (forvar5136 < (2'h2)); forvar5136 = (forvar5136 + (1'h1)))
            begin
              if (reg5085)
                begin
                  if ((~&reg5128[(2'h3):(2'h2)]))
                    begin
                      reg5137 <= $unsigned(reg5008[(4'h8):(4'h8)]);
                      reg5138 <= reg4974;
                    end
                  else
                    begin
                      reg5137 <= ($unsigned(reg5030[(2'h2):(1'h0)]) ?
                          (~$unsigned($signed(reg5036))) : $signed(((|reg5071) ?
                              (^forvar5136) : wire1023)));
                      reg5138 <= $signed(reg5056);
                    end
                  for (forvar5139 = (1'h0); (forvar5139 < (1'h0)); forvar5139 = (forvar5139 + (1'h1)))
                    begin
                      reg5140 <= reg4990[(2'h2):(1'h0)];
                    end
                  for (forvar5141 = (1'h0); (forvar5141 < (1'h1)); forvar5141 = (forvar5141 + (1'h1)))
                    begin
                      reg5142 <= (({(reg5112 ?
                                  reg4991 : reg5093)} | $signed((forvar5070 || (8'ha5)))) ?
                          {$unsigned(wire3538)} : ((|$unsigned(reg5137)) <= $unsigned($unsigned(reg4990))));
                    end
                  if ({$unsigned(((~|reg5073) ?
                          (8'had) : reg4977[(4'h9):(3'h6)]))})
                    begin
                      reg5143 <= $unsigned(reg4978);
                      reg5144 <= reg5025;
                      reg5145 <= $unsigned($signed(reg5050));
                    end
                  else
                    begin
                      reg5143 <= reg4975;
                    end
                end
              else
                begin
                  if ($unsigned((&$unsigned((forvar5095 | reg4981)))))
                    begin
                      reg5137 <= $signed($unsigned(((forvar4982 ?
                              (8'hb8) : forvar5040) ?
                          (reg5094 + forvar5139) : $signed(forvar5045))));
                      reg5138 <= {$unsigned($signed(reg5059[(3'h7):(2'h3)]))};
                      reg5139 <= ($signed(($signed(reg5100) ?
                          ((8'hba) ^ reg5023) : $signed(reg5092))) <<< $unsigned(reg5067[(1'h1):(1'h1)]));
                      reg5140 <= {$signed(reg5133[(3'h5):(2'h3)])};
                    end
                  else
                    begin
                      reg5137 <= ((reg5056 ?
                          $signed((reg5052 ^~ reg5076)) : (8'hb8)) | $unsigned((~{forvar5103})));
                      reg5138 <= (-($unsigned({reg5033}) ?
                          (&$signed((8'ha2))) : $signed({forvar5024})));
                      reg5139 <= reg5025[(1'h1):(1'h0)];
                      reg5140 <= (~&(reg4976[(1'h0):(1'h0)] ?
                          reg5027[(2'h3):(2'h2)] : $unsigned({reg5008})));
                    end
                  reg5141 <= wire1030[(5'h10):(3'h6)];
                end
              reg5146 <= (({$signed(reg5004)} >= ((~&forvar5074) - (forvar5033 ?
                      forvar5040 : (8'h9e)))) ?
                  $signed(reg4992[(1'h1):(1'h0)]) : (^$signed($unsigned((8'ha3)))));
              for (forvar5147 = (1'h0); (forvar5147 < (2'h3)); forvar5147 = (forvar5147 + (1'h1)))
                begin
                  if (((((reg4996 || forvar4970) ?
                          $signed(reg5007) : forvar5131[(2'h3):(1'h0)]) & $unsigned((~|(8'h9e)))) ?
                      (((reg5124 != (8'hae)) ?
                          reg5140[(1'h0):(1'h0)] : $unsigned(reg4994)) < (!$signed(reg5083))) : ((+wire3538) * forvar5061)))
                    begin
                      reg5148 <= $signed((8'had));
                      reg5149 <= forvar5131[(1'h0):(1'h0)];
                      reg5150 <= $unsigned((((reg5099 >>> forvar5018) | (reg4977 & wire1023)) ?
                          $signed({reg5123}) : forvar5098[(2'h3):(1'h1)]));
                      reg5151 <= (~(!((reg5122 ? forvar5040 : reg5150) ?
                          {reg5108} : forvar5079)));
                    end
                  else
                    begin
                      reg5148 <= $unsigned(((~&$unsigned(reg5009)) ?
                          $unsigned((reg5026 ?
                              (8'ha2) : reg4993)) : (~&reg5116[(2'h2):(2'h2)])));
                    end
                  if (((($signed(forvar4983) >>> ((8'ha6) ?
                      reg5039 : reg5151)) >> (^(reg5027 ^~ forvar5037))) >>> reg5000))
                    begin
                      reg5152 <= (wire3538[(3'h4):(1'h0)] ?
                          (((+forvar5024) ?
                                  reg4971[(1'h1):(1'h0)] : (reg4978 || reg5135)) ?
                              forvar5147[(1'h0):(1'h0)] : ((!reg5030) ?
                                  $unsigned(forvar5024) : (reg5107 & (8'hb1)))) : (((forvar5016 ?
                                  reg5124 : (8'hb7)) ?
                              reg4990 : $signed(reg5050)) | $signed($signed(reg5053))));
                    end
                  else
                    begin
                      reg5152 <= {$signed(({reg5108} ?
                              wire1031 : $signed(wire1022)))};
                      reg5153 <= $unsigned((reg5066 >>> ((reg5116 > reg5121) ?
                          $signed((8'haf)) : (reg5006 * reg4980))));
                      reg5154 <= (reg5065[(2'h3):(2'h2)] | ((!reg5030) ^~ $unsigned((^forvar4972))));
                    end
                end
            end
          reg5155 <= ($signed(reg5066) ? (reg5052 ~^ forvar5074) : forvar5074);
        end
      for (forvar5156 = (1'h0); (forvar5156 < (1'h1)); forvar5156 = (forvar5156 + (1'h1)))
        begin
          reg5157 <= $signed({($unsigned(reg5052) * reg4975[(4'hb):(1'h0)])});
          reg5158 <= wire1022;
          for (forvar5159 = (1'h0); (forvar5159 < (2'h3)); forvar5159 = (forvar5159 + (1'h1)))
            begin
              for (forvar5160 = (1'h0); (forvar5160 < (1'h0)); forvar5160 = (forvar5160 + (1'h1)))
                begin
                  for (forvar5161 = (1'h0); (forvar5161 < (1'h0)); forvar5161 = (forvar5161 + (1'h1)))
                    begin
                      reg5162 <= $signed(forvar5156);
                      reg5163 <= reg5125[(2'h2):(2'h2)];
                      reg5164 <= (!{reg4992});
                    end
                  for (forvar5165 = (1'h0); (forvar5165 < (1'h0)); forvar5165 = (forvar5165 + (1'h1)))
                    begin
                      reg5166 <= ($unsigned(reg5112[(3'h5):(1'h1)]) ?
                          reg5115[(4'hb):(3'h7)] : ((|$unsigned(reg4973)) | $unsigned($signed(forvar5082))));
                    end
                end
              for (forvar5167 = (1'h0); (forvar5167 < (1'h1)); forvar5167 = (forvar5167 + (1'h1)))
                begin
                  if (forvar5011)
                    begin
                      reg5168 <= $signed(reg5015[(1'h0):(1'h0)]);
                      reg5169 <= reg5058[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg5168 <= ((~&($unsigned(reg5053) != (reg5077 <<< reg4979))) || ((&(!(8'h9f))) == $unsigned(reg5084[(3'h5):(2'h3)])));
                      reg5169 <= ((reg4999[(4'h8):(2'h3)] ?
                          ((8'hac) >>> reg5000[(3'h4):(2'h3)]) : {(reg5144 ^~ reg5141)}) ^ $unsigned($unsigned((~&forvar5147))));
                      reg5170 <= ($signed({reg5100}) ?
                          {((reg5152 << reg4999) ?
                                  (forvar4970 ^ reg5163) : $unsigned(reg5069))} : $signed(reg5118[(1'h0):(1'h0)]));
                      reg5171 <= $unsigned($unsigned(($unsigned((8'h9c)) ?
                          reg5078 : (~^forvar5046))));
                    end
                end
              if ($unsigned((!(&(reg5030 ? reg5009 : reg5134)))))
                begin
                  for (forvar5172 = (1'h0); (forvar5172 < (2'h3)); forvar5172 = (forvar5172 + (1'h1)))
                    begin
                      reg5173 <= $signed(($unsigned((reg5004 ?
                          reg5071 : reg4975)) > $signed((~|reg5112))));
                      reg5174 <= $unsigned({$signed($unsigned((8'hb4)))});
                    end
                end
              else
                begin
                  for (forvar5172 = (1'h0); (forvar5172 < (2'h3)); forvar5172 = (forvar5172 + (1'h1)))
                    begin
                      reg5173 <= reg5122;
                    end
                end
              for (forvar5175 = (1'h0); (forvar5175 < (2'h3)); forvar5175 = (forvar5175 + (1'h1)))
                begin
                  if ((!$signed($unsigned(reg4979))))
                    begin
                      reg5176 <= $signed({(~&(reg4985 ? reg4985 : (8'hb3)))});
                      reg5177 <= forvar5156;
                      reg5178 <= reg5151;
                    end
                  else
                    begin
                      reg5176 <= (((forvar5161[(1'h1):(1'h0)] >= reg5116[(1'h0):(1'h0)]) ?
                          $signed((forvar5042 ?
                              forvar5018 : forvar5165)) : forvar5061) | (($signed(reg5059) <= forvar5047[(4'h8):(1'h1)]) == $signed($signed(forvar5167))));
                    end
                  for (forvar5179 = (1'h0); (forvar5179 < (1'h1)); forvar5179 = (forvar5179 + (1'h1)))
                    begin
                      reg5180 <= reg5066;
                      reg5181 <= ($unsigned(reg5122) >> {(reg5124[(3'h6):(1'h0)] ?
                              $unsigned(reg4988) : (reg5003 | (8'hb0)))});
                    end
                end
            end
          if (($unsigned(forvar4989[(2'h3):(1'h0)]) ?
              ((reg5072[(1'h1):(1'h0)] ?
                      $signed(reg5008) : forvar5159[(4'ha):(1'h1)]) ?
                  ($unsigned(forvar5141) ?
                      (reg5091 ^~ forvar5160) : (forvar5165 < reg4985)) : $unsigned((reg5093 && reg5120))) : $unsigned(reg5176)))
            begin
              if ((^(8'hb2)))
                begin
                  reg5182 <= reg5006;
                  for (forvar5183 = (1'h0); (forvar5183 < (2'h2)); forvar5183 = (forvar5183 + (1'h1)))
                    begin
                      reg5184 <= reg5101[(4'ha):(4'h9)];
                    end
                end
              else
                begin
                  if ((+($signed(((8'h9e) ? reg5138 : forvar5040)) ?
                      (8'hac) : wire1031[(1'h1):(1'h1)])))
                    begin
                      reg5182 <= reg5102[(3'h4):(1'h0)];
                      reg5183 <= reg5121;
                      reg5184 <= ((reg5049[(2'h2):(2'h2)] & ((8'ha2) ?
                          (!reg5145) : (~reg4981))) * ($signed({(8'ha9)}) ^~ ((!reg5102) & (forvar5088 ?
                          reg4971 : forvar5103))));
                    end
                  else
                    begin
                      reg5182 <= (forvar5061[(3'h6):(3'h6)] ?
                          (|((reg4997 >> reg5106) == reg4977)) : $signed($unsigned((!forvar5079))));
                      reg5183 <= ((+(8'ha2)) >= reg5014[(1'h1):(1'h1)]);
                      reg5184 <= (({reg5030} >> $unsigned((reg5092 <= reg5021))) ?
                          reg5066[(1'h1):(1'h0)] : reg5158);
                      reg5185 <= (reg5048 ?
                          ($unsigned((~&reg5057)) ^ (((8'hb1) < reg5033) ?
                              reg5054[(4'h8):(2'h2)] : reg4971[(1'h1):(1'h1)])) : $signed(forvar5001[(3'h7):(3'h4)]));
                    end
                  if (forvar5175)
                    begin
                      reg5186 <= {(~|(~(reg5108 ? reg5049 : reg5106)))};
                    end
                  else
                    begin
                      reg5186 <= forvar5030;
                    end
                  for (forvar5187 = (1'h0); (forvar5187 < (2'h2)); forvar5187 = (forvar5187 + (1'h1)))
                    begin
                      reg5188 <= $signed($signed(forvar5082));
                      reg5189 <= forvar4972[(2'h2):(1'h0)];
                      reg5190 <= (reg5114 - reg5144);
                      reg5191 <= $signed($signed($signed(forvar5060[(4'hb):(4'ha)])));
                    end
                end
              for (forvar5192 = (1'h0); (forvar5192 < (1'h0)); forvar5192 = (forvar5192 + (1'h1)))
                begin
                  reg5193 <= (^reg5010[(4'h8):(4'h8)]);
                  reg5194 <= reg5078[(3'h7):(3'h5)];
                  reg5195 <= ((((forvar4971 ? (8'hab) : reg5176) ?
                          $signed((8'h9f)) : reg5035[(2'h3):(2'h3)]) ~^ reg5069[(1'h0):(1'h0)]) ?
                      $signed(reg5077[(2'h3):(1'h0)]) : $signed((~&$unsigned((8'ha7)))));
                  for (forvar5196 = (1'h0); (forvar5196 < (2'h2)); forvar5196 = (forvar5196 + (1'h1)))
                    begin
                      reg5197 <= ($unsigned((reg5110[(3'h5):(2'h3)] ?
                          $signed(reg5109) : {forvar5109})) << $signed(((&forvar5131) ^ (reg5023 <<< (8'ha9)))));
                      reg5198 <= $unsigned((-($signed(reg5048) ^ reg5033)));
                      reg5199 <= (((8'hb0) ?
                              ({(8'hb9)} < $unsigned(forvar5024)) : reg5180) ?
                          ($unsigned($signed(reg4976)) ?
                              (&forvar5016) : $signed((reg5034 <= forvar5095))) : (+(~|$signed(reg5057))));
                      reg5200 <= forvar5159[(2'h2):(1'h1)];
                    end
                end
              for (forvar5201 = (1'h0); (forvar5201 < (2'h3)); forvar5201 = (forvar5201 + (1'h1)))
                begin
                  for (forvar5202 = (1'h0); (forvar5202 < (2'h2)); forvar5202 = (forvar5202 + (1'h1)))
                    begin
                      reg5203 <= forvar5160;
                      reg5204 <= $signed($signed(reg5041));
                      reg5205 <= $signed(($unsigned(forvar5082) * reg5041[(3'h6):(1'h0)]));
                    end
                  for (forvar5206 = (1'h0); (forvar5206 < (2'h3)); forvar5206 = (forvar5206 + (1'h1)))
                    begin
                      reg5207 <= (!(8'ha4));
                    end
                end
            end
          else
            begin
              if (forvar5064[(2'h2):(1'h1)])
                begin
                  for (forvar5182 = (1'h0); (forvar5182 < (1'h0)); forvar5182 = (forvar5182 + (1'h1)))
                    begin
                      reg5183 <= (+({$signed(reg5108)} - $signed(reg5054)));
                    end
                  reg5184 <= $unsigned(reg5063);
                  for (forvar5185 = (1'h0); (forvar5185 < (1'h0)); forvar5185 = (forvar5185 + (1'h1)))
                    begin
                      reg5186 <= (-(($unsigned((8'hb7)) || (reg5130 ?
                              reg4996 : forvar4972)) ?
                          reg5003 : {((8'hb8) ? forvar5047 : reg4990)}));
                      reg5187 <= $signed((!(|reg4981[(2'h3):(2'h3)])));
                      reg5188 <= (($unsigned((reg4972 ^ reg5093)) != forvar5095[(2'h2):(2'h2)]) > reg5072[(1'h1):(1'h1)]);
                    end
                  if (($signed({((8'hb6) ? reg5140 : reg5020)}) ?
                      $signed(($signed((8'hb8)) ?
                          forvar4989 : $signed(forvar5097))) : {(8'haf)}))
                    begin
                      reg5189 <= (~|(~&{(reg5013 || forvar5098)}));
                      reg5190 <= ($unsigned(forvar5060) && (reg5187[(4'hd):(2'h2)] <= (~|$signed((8'hab)))));
                      reg5191 <= (~&($signed($unsigned(wire1027)) ?
                          (forvar5030[(1'h1):(1'h1)] ?
                              $unsigned(reg5071) : reg5144) : reg5108[(3'h5):(1'h0)]));
                      reg5192 <= forvar5160;
                    end
                  else
                    begin
                      reg5189 <= ((&reg5033[(1'h1):(1'h1)]) <<< forvar5074[(3'h4):(2'h3)]);
                      reg5190 <= (reg5169 >> wire3538);
                      reg5191 <= $signed($signed(reg4994[(3'h7):(3'h4)]));
                      reg5192 <= reg5110;
                    end
                end
              else
                begin
                  if ((^~reg5177))
                    begin
                      reg5182 <= $signed($signed((8'hb3)));
                    end
                  else
                    begin
                      reg5182 <= reg5203[(3'h7):(2'h3)];
                    end
                end
              reg5193 <= {$unsigned(forvar5087)};
            end
        end
      for (forvar5208 = (1'h0); (forvar5208 < (2'h2)); forvar5208 = (forvar5208 + (1'h1)))
        begin
          for (forvar5209 = (1'h0); (forvar5209 < (2'h2)); forvar5209 = (forvar5209 + (1'h1)))
            begin
              if ($unsigned((reg5110[(2'h3):(2'h3)] ^~ ({forvar5081} ?
                  $signed(forvar5141) : (^reg5014)))))
                begin
                  for (forvar5210 = (1'h0); (forvar5210 < (2'h2)); forvar5210 = (forvar5210 + (1'h1)))
                    begin
                      reg5211 <= forvar5037;
                      reg5212 <= $signed(reg5030);
                    end
                  reg5213 <= ((reg5207 ?
                          {forvar5096[(2'h3):(1'h1)]} : $signed((reg5188 || (8'hb2)))) ?
                      $signed(forvar5167[(2'h2):(1'h0)]) : ({(forvar5210 != (8'hb2))} & (((8'ha2) ?
                          (8'h9e) : reg5211) && (reg5166 ?
                          forvar5087 : reg5048))));
                end
              else
                begin
                  for (forvar5210 = (1'h0); (forvar5210 < (1'h0)); forvar5210 = (forvar5210 + (1'h1)))
                    begin
                      reg5211 <= (~&forvar5088[(3'h4):(3'h4)]);
                      reg5212 <= reg5023[(2'h2):(2'h2)];
                      reg5213 <= $unsigned($signed({{reg5170}}));
                      reg5214 <= (($signed(forvar5201) ?
                              (~{reg4977}) : (|{reg5092})) ?
                          $signed((&$unsigned(reg4978))) : reg5033[(1'h1):(1'h1)]);
                    end
                  if ((!({$signed(reg5191)} ?
                      $unsigned(reg5025[(3'h4):(2'h3)]) : $signed($unsigned(reg5168)))))
                    begin
                      reg5215 <= {(+((reg5140 ? reg5057 : reg5137) ?
                              (forvar4982 ?
                                  reg5140 : forvar5024) : $unsigned((8'haf))))};
                      reg5216 <= {(^reg5065[(4'hd):(4'hc)])};
                      reg5217 <= ((|{(reg4991 || reg5207)}) ?
                          $unsigned(wire1030[(4'h8):(3'h5)]) : ((forvar5089 ?
                                  {(8'ha5)} : reg5174[(3'h7):(1'h1)]) ?
                              reg4995 : $signed(forvar4986)));
                      reg5218 <= $unsigned(((((8'hb0) < reg5176) ?
                          (+forvar5045) : {forvar5060}) << reg5003));
                    end
                  else
                    begin
                      reg5215 <= reg5146;
                      reg5216 <= ((~&($signed(wire1024) - forvar5064[(1'h1):(1'h0)])) ?
                          (((8'ha3) != (!reg5112)) >> $unsigned((forvar5061 * reg5114))) : $signed({$unsigned(reg5164)}));
                    end
                  if (reg5067[(2'h3):(2'h3)])
                    begin
                      reg5219 <= $signed(reg5180[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg5219 <= {(reg5170[(1'h1):(1'h0)] ?
                              {reg5138[(1'h1):(1'h1)]} : reg5091[(3'h5):(3'h5)])};
                      reg5220 <= (~^reg5031);
                      reg5221 <= {reg5204[(1'h1):(1'h0)]};
                      reg5222 <= (!$unsigned((reg5190[(1'h0):(1'h0)] ?
                          ((8'h9d) >> (8'hac)) : (wire1022 <<< reg5151))));
                    end
                  for (forvar5223 = (1'h0); (forvar5223 < (1'h0)); forvar5223 = (forvar5223 + (1'h1)))
                    begin
                      reg5224 <= (((-$unsigned(reg5066)) - ((forvar5051 != reg5066) ?
                              (reg5067 & reg5166) : reg5059[(3'h6):(1'h1)])) ?
                          ($unsigned($signed(reg5118)) <= ({forvar4983} - (reg5062 ?
                              reg5057 : reg5143))) : (+reg4973[(3'h5):(2'h3)]));
                      reg5225 <= ({$signed({reg5104})} ?
                          ($unsigned(((8'hb8) ? forvar5179 : forvar4989)) ?
                              (~reg5029[(1'h1):(1'h1)]) : reg5203[(4'h8):(3'h7)]) : $signed(($signed((8'hb0)) ?
                              reg5158 : $signed(reg5166))));
                    end
                end
              for (forvar5226 = (1'h0); (forvar5226 < (2'h2)); forvar5226 = (forvar5226 + (1'h1)))
                begin
                  for (forvar5227 = (1'h0); (forvar5227 < (1'h0)); forvar5227 = (forvar5227 + (1'h1)))
                    begin
                      reg5228 <= forvar5082;
                      reg5229 <= reg5212;
                    end
                  if (reg5004)
                    begin
                      reg5230 <= {reg5086};
                      reg5231 <= reg5166;
                      reg5232 <= (|{reg5204[(1'h0):(1'h0)]});
                      reg5233 <= ((~&reg5191[(4'hc):(2'h2)]) ?
                          wire1029[(3'h4):(2'h3)] : (~^$unsigned(forvar5037[(3'h5):(3'h4)])));
                    end
                  else
                    begin
                      reg5230 <= $unsigned($unsigned((8'hb7)));
                      reg5231 <= reg5126[(4'ha):(4'h8)];
                      reg5232 <= (~|((-(forvar5127 ~^ reg5232)) ?
                          (reg5086[(3'h5):(3'h4)] ?
                              ((8'h9f) - reg4980) : (reg5078 ?
                                  reg5195 : reg5008)) : (~(reg5221 ?
                              reg5199 : forvar5060))));
                    end
                  for (forvar5234 = (1'h0); (forvar5234 < (2'h2)); forvar5234 = (forvar5234 + (1'h1)))
                    begin
                      reg5235 <= $signed(forvar5055);
                    end
                  for (forvar5236 = (1'h0); (forvar5236 < (2'h3)); forvar5236 = (forvar5236 + (1'h1)))
                    begin
                      reg5237 <= $unsigned((-reg5008[(4'ha):(2'h2)]));
                    end
                end
            end
          for (forvar5238 = (1'h0); (forvar5238 < (2'h2)); forvar5238 = (forvar5238 + (1'h1)))
            begin
              for (forvar5239 = (1'h0); (forvar5239 < (2'h2)); forvar5239 = (forvar5239 + (1'h1)))
                begin
                  for (forvar5240 = (1'h0); (forvar5240 < (2'h2)); forvar5240 = (forvar5240 + (1'h1)))
                    begin
                      reg5241 <= ($unsigned($unsigned($unsigned(forvar5236))) ?
                          reg5153 : {((-reg5154) + $unsigned(reg5030))});
                      reg5242 <= $unsigned(((!$unsigned(reg4977)) ?
                          $signed((!(8'ha6))) : reg5178[(1'h0):(1'h0)]));
                      reg5243 <= $signed(reg5121[(4'hb):(1'h1)]);
                      reg5244 <= (~&(reg5229 >>> (8'h9e)));
                    end
                  reg5245 <= $signed($unsigned(($unsigned((8'hb6)) ?
                      $unsigned((8'ha6)) : $signed(reg5157))));
                  if ((-(reg5104 ? reg4975 : {{reg5180}})))
                    begin
                      reg5246 <= (~forvar5208[(4'ha):(3'h7)]);
                      reg5247 <= $signed(forvar5106[(1'h0):(1'h0)]);
                      reg5248 <= $signed(reg5063[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg5246 <= ((({wire1023} < $unsigned(reg5191)) >= (!$signed(reg5086))) ?
                          ((&reg5000[(1'h1):(1'h0)]) * (~$signed(forvar5079))) : $unsigned(($unsigned(reg5107) ?
                              (reg5117 ?
                                  reg5235 : reg5038) : $signed((8'haf)))));
                    end
                  for (forvar5249 = (1'h0); (forvar5249 < (2'h3)); forvar5249 = (forvar5249 + (1'h1)))
                    begin
                      reg5250 <= reg5163;
                    end
                end
              for (forvar5251 = (1'h0); (forvar5251 < (2'h2)); forvar5251 = (forvar5251 + (1'h1)))
                begin
                  for (forvar5252 = (1'h0); (forvar5252 < (2'h3)); forvar5252 = (forvar5252 + (1'h1)))
                    begin
                      reg5253 <= ($unsigned((~$signed(reg5029))) - forvar5109[(2'h3):(2'h2)]);
                      reg5254 <= ({((reg5035 == reg5049) ?
                                  reg5185[(2'h3):(1'h1)] : reg5169)} ?
                          $unsigned((+$signed(forvar4978))) : (-($signed(forvar5208) & $signed(reg5222))));
                    end
                end
              if ((reg5073 ?
                  $unsigned(((reg5109 > wire1022) ?
                      {reg5244} : $unsigned(reg5199))) : (~&($unsigned(reg5141) << ((8'ha5) ?
                      reg5178 : reg5242)))))
                begin
                  for (forvar5255 = (1'h0); (forvar5255 < (1'h1)); forvar5255 = (forvar5255 + (1'h1)))
                    begin
                      reg5256 <= ($unsigned(((8'ha9) ?
                              {reg4977} : $unsigned(reg5123))) ?
                          {$signed({reg5245})} : {reg5182[(2'h2):(2'h2)]});
                      reg5257 <= reg5053;
                      reg5258 <= ((~|$unsigned((reg5114 ?
                          reg5138 : reg5164))) >>> reg5068[(3'h6):(3'h5)]);
                    end
                  reg5259 <= (({{forvar5095}} ?
                      reg5192 : (reg5187 == reg5141[(4'ha):(2'h2)])) && ((8'ha3) + (^~$signed(forvar5037))));
                  for (forvar5260 = (1'h0); (forvar5260 < (1'h1)); forvar5260 = (forvar5260 + (1'h1)))
                    begin
                      reg5261 <= reg4996;
                      reg5262 <= ($signed((-(reg5135 < (8'hb0)))) ?
                          (&reg5144) : ($signed(reg5057) ?
                              $signed(reg5067[(4'ha):(2'h2)]) : forvar5161));
                      reg5263 <= (^~$signed(reg5145[(2'h2):(2'h2)]));
                      reg5264 <= reg4994;
                    end
                  for (forvar5265 = (1'h0); (forvar5265 < (1'h1)); forvar5265 = (forvar5265 + (1'h1)))
                    begin
                      reg5266 <= ((($signed(forvar5037) >>> $signed(reg5215)) ?
                              reg4976[(1'h0):(1'h0)] : ($unsigned(forvar5117) * (wire1028 ?
                                  reg5261 : reg5132))) ?
                          $unsigned($unsigned((!(8'ha7)))) : ((~|{reg5204}) >= (reg5186[(4'hb):(1'h0)] >>> reg5109[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  if (((($unsigned(forvar5060) ?
                          (8'hba) : reg5084[(3'h4):(1'h1)]) == ((~^forvar5080) ?
                          (~|reg5139) : (~|reg5266))) ?
                      ($signed(reg5110) ?
                          $signed(forvar5082) : (-(|forvar5051))) : reg5142[(2'h2):(2'h2)]))
                    begin
                      reg5255 <= reg1026[(4'h8):(2'h2)];
                      reg5256 <= {(-$unsigned((forvar5201 ^~ reg5032)))};
                    end
                  else
                    begin
                      reg5255 <= reg4990[(3'h7):(3'h6)];
                      reg5256 <= ($signed((|(forvar5179 ?
                          reg4971 : wire4967))) * $unsigned(({forvar5024} ?
                          (reg5185 ? reg5017 : reg5003) : (-reg5025))));
                      reg5257 <= (&$signed(forvar4972[(2'h3):(2'h3)]));
                      reg5258 <= {{reg5043[(4'h8):(4'h8)]}};
                    end
                  if (reg5220[(2'h3):(2'h3)])
                    begin
                      reg5259 <= (wire1023[(4'he):(2'h2)] != reg5077);
                      reg5260 <= reg5116[(1'h1):(1'h1)];
                      reg5261 <= (^~reg5169);
                      reg5262 <= {(+reg5182[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg5259 <= forvar5209[(2'h2):(1'h1)];
                      reg5260 <= reg5059;
                      reg5261 <= (~|(forvar4971[(1'h1):(1'h0)] ?
                          $signed(forvar5095) : (~^$unsigned(reg5190))));
                    end
                  if ($unsigned(reg5194))
                    begin
                      reg5263 <= {(^reg5182[(3'h6):(1'h0)])};
                    end
                  else
                    begin
                      reg5263 <= ((~&({reg5177} ?
                              $signed(reg5176) : $signed((8'haa)))) ?
                          (reg5105 ?
                              $unsigned((reg5184 | (8'hb2))) : (^~$unsigned(reg5083))) : (forvar5079[(2'h2):(1'h1)] ?
                              ((forvar5251 >>> reg5068) && $unsigned(reg5243)) : forvar5160));
                      reg5264 <= wire1029[(4'h9):(3'h7)];
                    end
                end
            end
          if (({{$signed(reg5192)}} ?
              forvar5074[(3'h4):(2'h3)] : $unsigned($signed((forvar5033 <<< reg5221)))))
            begin
              for (forvar5267 = (1'h0); (forvar5267 < (2'h2)); forvar5267 = (forvar5267 + (1'h1)))
                begin
                  reg5268 <= reg5170[(1'h1):(1'h1)];
                  reg5269 <= $unsigned(((&{(8'h9f)}) == ($signed(reg5029) || {forvar5223})));
                  if (reg1026)
                    begin
                      reg5270 <= forvar5179[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg5270 <= (((|reg5200[(2'h2):(2'h2)]) ?
                              (&(reg5120 ?
                                  (8'hb5) : reg5102)) : ($unsigned(forvar5210) > ((8'hac) ?
                                  reg5233 : reg5049))) ?
                          $unsigned(reg5194[(4'ha):(4'h9)]) : (!{(8'ha1)}));
                    end
                end
              reg5271 <= ($signed(reg5149) ^~ $unsigned($signed((reg4974 * reg5124))));
              if ({wire1025[(2'h3):(2'h3)]})
                begin
                  if ({{(~|(-reg5154))}})
                    begin
                      reg5272 <= reg5044;
                      reg5273 <= ($signed((|forvar5047)) ^ (^~{reg5000}));
                      reg5274 <= $signed($unsigned($unsigned($signed(forvar5131))));
                      reg5275 <= (~&(!(reg5030 ?
                          (forvar5098 < forvar5080) : reg5119)));
                    end
                  else
                    begin
                      reg5272 <= (~reg4977[(2'h3):(2'h2)]);
                      reg5273 <= (~|reg5028);
                    end
                  for (forvar5276 = (1'h0); (forvar5276 < (2'h3)); forvar5276 = (forvar5276 + (1'h1)))
                    begin
                      reg5277 <= ($unsigned(forvar5096[(3'h4):(3'h4)]) == $signed((reg5137 <= (reg5182 ~^ forvar5276))));
                      reg5278 <= reg5273;
                      reg5279 <= $signed(reg5262[(1'h0):(1'h0)]);
                    end
                  reg5280 <= (forvar4970 + (~^reg5242[(1'h0):(1'h0)]));
                  for (forvar5281 = (1'h0); (forvar5281 < (2'h2)); forvar5281 = (forvar5281 + (1'h1)))
                    begin
                      reg5282 <= ($unsigned(((~|reg5132) ?
                          {reg5263} : $signed(reg5043))) & $signed($signed($signed((8'ha8)))));
                      reg5283 <= ($unsigned($unsigned((~reg5033))) * ((!reg5138[(1'h0):(1'h0)]) & (!reg5187)));
                    end
                end
              else
                begin
                  for (forvar5272 = (1'h0); (forvar5272 < (2'h3)); forvar5272 = (forvar5272 + (1'h1)))
                    begin
                      reg5273 <= ((({reg5137} << $unsigned(reg5104)) <= forvar5206) && $unsigned(((reg4985 ?
                          reg5092 : forvar5251) + (&reg5034))));
                      reg5274 <= $signed(forvar5002[(4'hc):(3'h4)]);
                    end
                  if ($unsigned((reg5279[(3'h5):(1'h1)] ?
                      reg5091[(3'h5):(2'h2)] : (forvar5209 ^ {reg5118}))))
                    begin
                      reg5275 <= forvar5234[(4'h9):(3'h7)];
                      reg5276 <= (reg1026[(4'hc):(4'ha)] <<< (~reg5230));
                      reg5277 <= {($unsigned($unsigned(reg5230)) ?
                              (8'ha4) : $signed((~&reg4999)))};
                    end
                  else
                    begin
                      reg5275 <= forvar5060;
                    end
                  if (reg4979)
                    begin
                      reg5278 <= ($unsigned(((reg5000 ?
                          (8'hba) : forvar5018) ~^ (8'hb8))) ^~ $signed(reg5025));
                      reg5279 <= $signed($unsigned(($signed(forvar5179) ?
                          {reg5150} : (reg5152 ? forvar5160 : (8'hba)))));
                      reg5280 <= $unsigned($signed(wire1022[(4'hb):(1'h1)]));
                      reg5281 <= (({$signed(reg5243)} == ({forvar5210} ?
                              (reg5132 ? reg5191 : reg5242) : {reg5149})) ?
                          $unsigned($unsigned($unsigned(reg5205))) : (&forvar5095));
                    end
                  else
                    begin
                      reg5278 <= {reg5021[(4'he):(2'h3)]};
                    end
                end
            end
          else
            begin
              for (forvar5267 = (1'h0); (forvar5267 < (1'h1)); forvar5267 = (forvar5267 + (1'h1)))
                begin
                  reg5268 <= (^~(~|forvar5234[(1'h1):(1'h0)]));
                  reg5269 <= $unsigned($unsigned($unsigned(reg5276[(1'h0):(1'h0)])));
                end
              for (forvar5270 = (1'h0); (forvar5270 < (1'h0)); forvar5270 = (forvar5270 + (1'h1)))
                begin
                  for (forvar5271 = (1'h0); (forvar5271 < (2'h3)); forvar5271 = (forvar5271 + (1'h1)))
                    begin
                      reg5272 <= $signed(forvar5024[(3'h7):(2'h3)]);
                      reg5273 <= reg5246;
                    end
                  reg5274 <= $signed(reg5216[(3'h5):(1'h1)]);
                  if ((&(-(reg5203[(3'h4):(1'h1)] >>> $signed(wire4969)))))
                    begin
                      reg5275 <= $signed({$signed(reg5162)});
                      reg5276 <= reg5145[(1'h0):(1'h0)];
                      reg5277 <= ((&reg4974) ~^ ($unsigned($unsigned(forvar5182)) ?
                          $unsigned((reg4981 ?
                              reg5187 : reg5258)) : (-{reg5013})));
                    end
                  else
                    begin
                      reg5275 <= $signed((((reg5140 + (8'ha5)) ?
                          reg5015[(3'h4):(3'h4)] : reg5116) && ((~reg5244) ?
                          ((8'haf) - wire1031) : (reg5269 <= reg5164))));
                      reg5276 <= $signed($signed((^(forvar5208 >> reg5144))));
                    end
                  for (forvar5278 = (1'h0); (forvar5278 < (2'h3)); forvar5278 = (forvar5278 + (1'h1)))
                    begin
                      reg5279 <= $signed((&($unsigned(forvar5070) ?
                          $signed(reg5104) : $unsigned(forvar5001))));
                      reg5280 <= (!$unsigned((^$unsigned(reg5235))));
                    end
                end
              for (forvar5281 = (1'h0); (forvar5281 < (2'h2)); forvar5281 = (forvar5281 + (1'h1)))
                begin
                  for (forvar5282 = (1'h0); (forvar5282 < (1'h0)); forvar5282 = (forvar5282 + (1'h1)))
                    begin
                      reg5283 <= ((~^(^~(~^reg5104))) == ({reg5195} ?
                          ($unsigned(forvar5037) ^~ (8'ha6)) : forvar5255));
                      reg5284 <= (^(({reg5003} == (reg5004 - (8'hb4))) || ($signed(reg5124) ?
                          (reg5091 & wire1031) : {reg5166})));
                      reg5285 <= ((!(&reg5100)) > reg5093[(3'h6):(3'h4)]);
                      reg5286 <= forvar5051;
                    end
                  reg5287 <= $unsigned({((reg5085 ~^ (8'hab)) ?
                          $unsigned(reg5142) : reg5007[(2'h2):(1'h1)])});
                  for (forvar5288 = (1'h0); (forvar5288 < (2'h2)); forvar5288 = (forvar5288 + (1'h1)))
                    begin
                      reg5289 <= $unsigned(((forvar5239 ?
                          (forvar5175 ?
                              reg5181 : wire1024) : $unsigned(wire1024)) ~^ ($signed(reg5247) + (8'ha3))));
                    end
                end
            end
        end
    end
  assign wire5290 = $signed($unsigned((^~forvar5239)));
  assign wire5291 = reg5152;
  always
    @(posedge clk) begin
      for (forvar5292 = (1'h0); (forvar5292 < (1'h1)); forvar5292 = (forvar5292 + (1'h1)))
        begin
          reg5293 <= $unsigned((~&$signed(wire1025)));
          if ((forvar5070 ?
              (-($unsigned(wire1027) ?
                  (^forvar5082) : reg5129[(4'hb):(3'h4)])) : (((+reg5261) ?
                      (reg4976 <= reg5121) : $signed(reg5263)) ?
                  ($signed((8'ha8)) || reg5115[(3'h4):(1'h1)]) : {$signed(forvar5208)})))
            begin
              for (forvar5294 = (1'h0); (forvar5294 < (1'h0)); forvar5294 = (forvar5294 + (1'h1)))
                begin
                  for (forvar5295 = (1'h0); (forvar5295 < (2'h3)); forvar5295 = (forvar5295 + (1'h1)))
                    begin
                      reg5296 <= $signed((^((reg5186 ?
                              forvar5206 : forvar4970) ?
                          $unsigned(forvar5051) : $unsigned(reg5228))));
                      reg5297 <= (forvar5249 ?
                          forvar4971 : ((reg5157 ?
                                  reg5148[(4'h8):(3'h7)] : ((8'h9f) ?
                                      (8'ha4) : reg5286)) ?
                              reg5164[(1'h1):(1'h0)] : ({(8'hae)} ~^ (forvar5033 ?
                                  (8'hb0) : reg5133))));
                      reg5298 <= $signed((((reg5005 ? forvar5226 : forvar5106) ?
                          $signed(reg5261) : $unsigned((8'haf))) == {$unsigned(reg5211)}));
                      reg5299 <= $signed((~|$signed(reg5274[(4'ha):(3'h6)])));
                    end
                  reg5300 <= (~|{$signed((reg5050 ? reg5266 : (8'hab)))});
                  for (forvar5301 = (1'h0); (forvar5301 < (1'h1)); forvar5301 = (forvar5301 + (1'h1)))
                    begin
                      reg5302 <= $signed(forvar5255[(4'h8):(3'h5)]);
                      reg5303 <= $signed($unsigned(reg5027));
                      reg5304 <= {(^$unsigned(reg5035))};
                    end
                  for (forvar5305 = (1'h0); (forvar5305 < (2'h2)); forvar5305 = (forvar5305 + (1'h1)))
                    begin
                      reg5306 <= $unsigned(forvar5016[(4'h8):(1'h1)]);
                    end
                end
              reg5307 <= wire4969;
              if (reg1026)
                begin
                  if ((+(reg5012 ?
                      (&(wire1029 ?
                          reg5039 : reg5189)) : $unsigned((~&reg5274)))))
                    begin
                      reg5308 <= (8'hb4);
                      reg5309 <= reg5183;
                      reg5310 <= reg5049;
                      reg5311 <= forvar5109[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg5308 <= $signed(forvar5047[(3'h4):(2'h2)]);
                      reg5309 <= $unsigned($signed((~|(8'h9e))));
                    end
                end
              else
                begin
                  if ($unsigned((-({reg5262} ?
                      forvar5095[(4'he):(2'h3)] : $signed(reg5222)))))
                    begin
                      reg5308 <= $unsigned((forvar5260 ^ reg5230[(4'hd):(4'hc)]));
                      reg5309 <= (~|({reg5178[(2'h3):(2'h3)]} <= reg5143));
                      reg5310 <= reg5176[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg5308 <= $signed(($unsigned(reg5077) ?
                          forvar5208[(3'h5):(1'h0)] : reg5126));
                    end
                  reg5311 <= $unsigned((forvar5103 == (reg5211 == {forvar5196})));
                  if (reg5177[(1'h1):(1'h1)])
                    begin
                      reg5312 <= (8'hb9);
                      reg5313 <= ($signed((~^wire4969)) ? reg5271 : reg5015);
                    end
                  else
                    begin
                      reg5312 <= forvar5001[(2'h3):(1'h1)];
                      reg5313 <= (~&reg5306[(2'h2):(1'h0)]);
                    end
                end
              for (forvar5314 = (1'h0); (forvar5314 < (2'h2)); forvar5314 = (forvar5314 + (1'h1)))
                begin
                  for (forvar5315 = (1'h0); (forvar5315 < (1'h0)); forvar5315 = (forvar5315 + (1'h1)))
                    begin
                      reg5316 <= reg5078[(3'h7):(2'h2)];
                      reg5317 <= reg5191[(2'h2):(2'h2)];
                      reg5318 <= (forvar5046 + (($unsigned(forvar5282) ?
                              (8'hb8) : forvar5051) ?
                          $unsigned($unsigned(reg5015)) : $signed(reg5048[(2'h2):(1'h0)])));
                    end
                  for (forvar5319 = (1'h0); (forvar5319 < (1'h0)); forvar5319 = (forvar5319 + (1'h1)))
                    begin
                      reg5320 <= (8'hb0);
                      reg5321 <= ({(reg5307 ^ $signed(forvar5209))} ?
                          (reg5225[(2'h2):(1'h0)] >> ($signed(reg5110) ?
                              reg5268 : (&(8'hb5)))) : $unsigned($signed(reg5132[(2'h3):(2'h2)])));
                      reg5322 <= reg5107;
                    end
                end
            end
          else
            begin
              if (forvar5185[(2'h2):(2'h2)])
                begin
                  reg5294 <= $unsigned($signed({(&forvar5096)}));
                  for (forvar5295 = (1'h0); (forvar5295 < (2'h2)); forvar5295 = (forvar5295 + (1'h1)))
                    begin
                      reg5296 <= reg5313;
                    end
                  reg5297 <= (^($signed((^reg5248)) - ({(8'hb6)} ?
                      (reg5116 ?
                          forvar5156 : reg5059) : reg5145[(1'h0):(1'h0)])));
                end
              else
                begin
                  for (forvar5294 = (1'h0); (forvar5294 < (2'h2)); forvar5294 = (forvar5294 + (1'h1)))
                    begin
                      reg5295 <= (~^(~&((!reg5277) ~^ reg5038)));
                      reg5296 <= reg5215;
                    end
                  reg5297 <= (~|(^~forvar5040[(3'h7):(3'h4)]));
                  for (forvar5298 = (1'h0); (forvar5298 < (2'h2)); forvar5298 = (forvar5298 + (1'h1)))
                    begin
                      reg5299 <= ({$unsigned((reg5286 <= reg5021))} ^~ (($unsigned((8'ha7)) ?
                              reg5217 : reg4994) ?
                          ((reg5266 <= reg5304) ?
                              (reg5154 ^ (8'ha8)) : {reg1026}) : ((reg5084 > wire1023) ?
                              reg5205 : (reg5076 == reg5311))));
                    end
                end
            end
          if (forvar5011[(3'h4):(2'h3)])
            begin
              for (forvar5323 = (1'h0); (forvar5323 < (2'h2)); forvar5323 = (forvar5323 + (1'h1)))
                begin
                  for (forvar5324 = (1'h0); (forvar5324 < (2'h3)); forvar5324 = (forvar5324 + (1'h1)))
                    begin
                      reg5325 <= (((-forvar5210) ?
                              forvar4986 : {((8'hac) ? reg5214 : reg5192)}) ?
                          $signed({(reg5207 >>> reg5093)}) : ($unsigned($unsigned((8'hb0))) ?
                              forvar5011[(1'h1):(1'h0)] : $signed(reg5072[(2'h2):(1'h1)])));
                    end
                  reg5326 <= ($signed($unsigned(reg5054)) ?
                      reg5289[(4'hb):(1'h1)] : ($signed($unsigned(reg5187)) | $signed((forvar5314 | (8'ha7)))));
                  if ((({$signed(reg5049)} ^~ $signed($signed(reg5150))) ?
                      reg5067 : $unsigned((^{forvar5047}))))
                    begin
                      reg5327 <= (^~(($unsigned(forvar5270) && $signed(reg5153)) ?
                          $signed($unsigned(forvar5267)) : (!forvar5175)));
                      reg5328 <= reg5326[(4'ha):(1'h0)];
                    end
                  else
                    begin
                      reg5327 <= (reg5280 ?
                          (!$signed($signed((8'ha1)))) : (((8'hb0) <= forvar5206) ?
                              reg5211[(3'h6):(3'h5)] : {reg5168[(1'h1):(1'h1)]}));
                      reg5328 <= ((8'h9e) < forvar5265[(4'hb):(3'h7)]);
                    end
                end
              for (forvar5329 = (1'h0); (forvar5329 < (2'h3)); forvar5329 = (forvar5329 + (1'h1)))
                begin
                  if ($unsigned(($unsigned($unsigned(forvar5276)) != {$signed(reg5318)})))
                    begin
                      reg5330 <= ($unsigned(($unsigned(reg5155) * $unsigned(reg5084))) ?
                          ((|(reg5162 ?
                              (8'ha3) : (8'ha6))) <<< ((reg5200 ~^ reg5326) < $unsigned(forvar5040))) : ($signed((forvar5202 ?
                              reg4976 : reg5119)) >= {(~(8'hab))}));
                      reg5331 <= $unsigned($unsigned(reg5282[(3'h5):(3'h4)]));
                      reg5332 <= $unsigned({{reg5008[(4'ha):(4'h8)]}});
                      reg5333 <= reg5123[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg5330 <= forvar5117[(2'h3):(2'h2)];
                      reg5331 <= $unsigned($signed((+$signed(reg5322))));
                      reg5332 <= ((&$unsigned(forvar5227[(3'h7):(3'h7)])) >= $unsigned($signed((^~forvar5175))));
                    end
                end
            end
          else
            begin
              for (forvar5323 = (1'h0); (forvar5323 < (2'h3)); forvar5323 = (forvar5323 + (1'h1)))
                begin
                  for (forvar5324 = (1'h0); (forvar5324 < (2'h2)); forvar5324 = (forvar5324 + (1'h1)))
                    begin
                      reg5325 <= forvar5046;
                      reg5326 <= ($signed(reg5114) != ($unsigned($unsigned(forvar5074)) ?
                          reg5312[(2'h2):(1'h1)] : ((reg5085 ?
                              forvar5238 : reg5271) < (reg5145 ?
                              forvar5098 : forvar5070))));
                      reg5327 <= (8'hb6);
                    end
                  reg5328 <= (($signed(forvar5208[(4'h8):(1'h1)]) <= $unsigned((+reg5231))) - (reg5092 != $unsigned($signed(wire1028))));
                  if ($unsigned(reg5145[(1'h0):(1'h0)]))
                    begin
                      reg5329 <= reg5100[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg5329 <= ((~^forvar5030[(4'h8):(3'h4)]) > $unsigned(reg5188));
                      reg5330 <= {$unsigned((forvar5192[(3'h6):(2'h3)] ?
                              reg5293 : (forvar5116 != forvar5106)))};
                      reg5331 <= $signed((^$signed(reg5258[(4'h9):(3'h7)])));
                    end
                end
            end
          reg5334 <= (~{$unsigned((reg5327 ? reg5182 : reg5148))});
        end
      reg5335 <= {$signed($signed(forvar5251))};
    end
  assign wire5336 = (^~$unsigned(((&reg5071) ^~ reg5306[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      for (forvar5337 = (1'h0); (forvar5337 < (2'h2)); forvar5337 = (forvar5337 + (1'h1)))
        begin
          if (forvar5249)
            begin
              reg5338 <= reg5225[(4'h9):(3'h5)];
              for (forvar5339 = (1'h0); (forvar5339 < (2'h2)); forvar5339 = (forvar5339 + (1'h1)))
                begin
                  if (reg5141)
                    begin
                      reg5340 <= ((((forvar5079 ^~ reg5144) - (8'ha4)) ?
                          $signed((^(8'ha6))) : ($signed((8'h9f)) ?
                              {reg5295} : (|reg5274))) < forvar5087[(4'h9):(3'h7)]);
                    end
                  else
                    begin
                      reg5340 <= reg5000[(1'h1):(1'h0)];
                      reg5341 <= {$unsigned(((~^forvar5055) ?
                              (reg5243 + reg4975) : (forvar5096 > reg5035)))};
                      reg5342 <= reg5116;
                    end
                  reg5343 <= reg5108;
                  if ($unsigned({((+forvar5301) * $unsigned(reg5318))}))
                    begin
                      reg5344 <= (8'hb9);
                    end
                  else
                    begin
                      reg5344 <= $unsigned($unsigned(reg5192[(3'h5):(1'h1)]));
                    end
                  if (reg5057[(3'h5):(1'h1)])
                    begin
                      reg5345 <= (reg5142[(4'hd):(4'hb)] ?
                          ((reg4988[(1'h0):(1'h0)] ?
                              (&reg4997) : $unsigned(reg5007)) << {(~&forvar5156)}) : reg5269[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg5345 <= ($signed(($unsigned((8'ha9)) ?
                              $signed(reg5338) : (reg5137 ?
                                  reg5312 : reg5139))) ?
                          reg5282[(1'h1):(1'h0)] : ((((8'haa) ?
                                  reg5264 : reg5225) > (reg5255 ?
                                  reg5278 : reg5246)) ?
                              reg5067[(3'h4):(1'h0)] : {reg5012}));
                      reg5346 <= $unsigned(($unsigned(((8'h9f) ~^ (8'ha3))) ^ $unsigned(forvar5183)));
                    end
                end
              for (forvar5347 = (1'h0); (forvar5347 < (1'h1)); forvar5347 = (forvar5347 + (1'h1)))
                begin
                  if (((&((forvar5042 ?
                      reg5330 : (8'hb5)) | $unsigned(reg5077))) > (+$signed(reg5099[(1'h1):(1'h1)]))))
                    begin
                      reg5348 <= {(&((!wire1023) ?
                              reg5035[(3'h4):(2'h2)] : forvar5088[(2'h2):(1'h0)]))};
                      reg5349 <= ({{(^forvar5239)}} ?
                          {(((8'ha4) ?
                                  forvar5103 : reg5129) < (8'hb6))} : (^~((8'had) ?
                              $signed(forvar5175) : {reg5012})));
                    end
                  else
                    begin
                      reg5348 <= (forvar5251[(4'h9):(3'h4)] ?
                          $signed({reg5183[(3'h6):(3'h5)]}) : $signed((~(reg5077 ?
                              reg5237 : reg5153))));
                      reg5349 <= $unsigned($signed((&reg5067)));
                      reg5350 <= wire1023[(4'he):(4'hb)];
                    end
                end
            end
          else
            begin
              if (reg5232)
                begin
                  for (forvar5338 = (1'h0); (forvar5338 < (1'h1)); forvar5338 = (forvar5338 + (1'h1)))
                    begin
                      reg5339 <= (($unsigned(forvar5156) * ((~reg5150) ^ $signed(reg5049))) >>> (^(8'h9f)));
                      reg5340 <= (+$signed(reg5000[(3'h4):(3'h4)]));
                    end
                  if ($unsigned({(+{forvar5249})}))
                    begin
                      reg5341 <= (((forvar5095[(2'h2):(2'h2)] >= (~forvar5172)) ?
                              ((+reg5322) >= {reg5005}) : {$signed(reg4973)}) ?
                          ($signed((!reg5274)) ?
                              (|{reg5215}) : {$signed(reg5217)}) : ($unsigned($signed(reg5152)) || {{forvar5282}}));
                      reg5342 <= reg5218[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg5341 <= reg5078[(2'h2):(1'h0)];
                    end
                  for (forvar5343 = (1'h0); (forvar5343 < (1'h1)); forvar5343 = (forvar5343 + (1'h1)))
                    begin
                      reg5344 <= ({$signed((|(8'h9d)))} || reg4972);
                      reg5345 <= forvar5226;
                      reg5346 <= $signed($signed($unsigned((reg5177 || reg5110))));
                    end
                  if (reg5026[(3'h4):(2'h2)])
                    begin
                      reg5347 <= reg5198;
                    end
                  else
                    begin
                      reg5347 <= ((|((forvar5234 ?
                              reg5154 : reg5054) >= $signed(forvar5251))) ?
                          {{$signed(reg5144)}} : $unsigned((|(reg5113 ?
                              reg5152 : reg5318))));
                      reg5348 <= {$signed((+(reg5221 ? reg5004 : (8'ha8))))};
                    end
                end
              else
                begin
                  reg5338 <= forvar5002[(4'ha):(1'h1)];
                  if (reg5132)
                    begin
                      reg5339 <= $unsigned(forvar5185);
                      reg5340 <= ((reg5326 ?
                          (~|(-reg4980)) : {forvar5209[(5'h10):(4'ha)]}) == $unsigned({(reg5278 ^~ forvar5090)}));
                    end
                  else
                    begin
                      reg5339 <= $signed($signed(($unsigned(reg4999) ?
                          ((8'ha8) ? reg5347 : reg4985) : (reg5339 ?
                              (8'hb0) : forvar5315))));
                    end
                  for (forvar5341 = (1'h0); (forvar5341 < (2'h2)); forvar5341 = (forvar5341 + (1'h1)))
                    begin
                      reg5342 <= ($unsigned(reg4992) ?
                          (-forvar5288) : (reg5344[(3'h7):(3'h5)] ?
                              (~(^~forvar5329)) : wire4967[(2'h2):(1'h1)]));
                      reg5343 <= $unsigned({{forvar5047[(2'h2):(2'h2)]}});
                      reg5344 <= reg5207;
                      reg5345 <= (reg5284 ? reg5263 : $unsigned(reg4984));
                    end
                  for (forvar5346 = (1'h0); (forvar5346 < (1'h1)); forvar5346 = (forvar5346 + (1'h1)))
                    begin
                      reg5347 <= reg5327;
                    end
                end
              for (forvar5349 = (1'h0); (forvar5349 < (1'h0)); forvar5349 = (forvar5349 + (1'h1)))
                begin
                  if ($signed(forvar5019))
                    begin
                      reg5350 <= (forvar5337[(1'h0):(1'h0)] ?
                          (8'ha9) : (|($signed(reg5062) == (+(8'h9d)))));
                    end
                  else
                    begin
                      reg5350 <= (($signed((^forvar5074)) >> $signed($unsigned(reg5068))) ?
                          $signed(((8'hab) ?
                              $unsigned(forvar5265) : (8'hb3))) : (!{(reg5318 == forvar5060)}));
                      reg5351 <= $signed((8'ha5));
                      reg5352 <= (8'hb3);
                    end
                  for (forvar5353 = (1'h0); (forvar5353 < (1'h1)); forvar5353 = (forvar5353 + (1'h1)))
                    begin
                      reg5354 <= (&(~|(forvar5226 < $signed(reg5248))));
                    end
                  if (({(reg5067[(3'h7):(1'h1)] ?
                          (forvar5329 ?
                              reg5044 : forvar5272) : $unsigned(reg5237))} >= $unsigned((~&$signed((8'h9e))))))
                    begin
                      reg5355 <= $signed(((&(reg5003 + reg5218)) ?
                          forvar5019 : (!(~&(8'ha8)))));
                      reg5356 <= (((forvar5227 ?
                          (reg5355 ?
                              (8'ha7) : forvar5206) : (forvar5141 ^~ reg5295)) << forvar5202) ^~ reg5176);
                    end
                  else
                    begin
                      reg5355 <= reg5309;
                      reg5356 <= (^~reg5163[(1'h1):(1'h1)]);
                    end
                end
            end
          for (forvar5357 = (1'h0); (forvar5357 < (1'h1)); forvar5357 = (forvar5357 + (1'h1)))
            begin
              reg5358 <= reg5149[(3'h7):(2'h3)];
              for (forvar5359 = (1'h0); (forvar5359 < (2'h3)); forvar5359 = (forvar5359 + (1'h1)))
                begin
                  for (forvar5360 = (1'h0); (forvar5360 < (1'h1)); forvar5360 = (forvar5360 + (1'h1)))
                    begin
                      reg5361 <= $unsigned((|reg1026));
                    end
                  for (forvar5362 = (1'h0); (forvar5362 < (1'h0)); forvar5362 = (forvar5362 + (1'h1)))
                    begin
                      reg5363 <= (($unsigned((~&wire5291)) ?
                              $signed((~reg5221)) : reg5113[(1'h0):(1'h0)]) ?
                          ($unsigned($unsigned(reg5264)) ?
                              $unsigned(reg5013[(2'h3):(2'h3)]) : reg5163[(2'h2):(2'h2)]) : reg5004);
                    end
                end
              for (forvar5364 = (1'h0); (forvar5364 < (1'h1)); forvar5364 = (forvar5364 + (1'h1)))
                begin
                  if (reg5351[(1'h0):(1'h0)])
                    begin
                      reg5365 <= $unsigned(reg5184);
                      reg5366 <= $unsigned(({{(8'ha8)}} ?
                          (8'had) : (forvar5349 <= (reg5245 ?
                              forvar4989 : reg4995))));
                      reg5367 <= reg5078[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg5365 <= (-reg4995[(3'h5):(2'h3)]);
                      reg5366 <= (8'hb2);
                    end
                  reg5368 <= $unsigned(forvar5070);
                  reg5369 <= {((8'hae) == (forvar5040[(4'h8):(1'h0)] ?
                          $signed((8'hb0)) : (reg5296 ^~ forvar5080)))};
                  if ($unsigned($signed(reg5329[(2'h3):(2'h3)])))
                    begin
                      reg5370 <= $signed($unsigned(((-(8'hb2)) ?
                          (reg5358 + reg5065) : ((8'hb0) ?
                              reg5245 : forvar5357))));
                      reg5371 <= ((8'ha8) | $unsigned($signed({reg5345})));
                    end
                  else
                    begin
                      reg5370 <= reg5012;
                      reg5371 <= reg5350[(2'h3):(1'h0)];
                      reg5372 <= (($unsigned((wire1025 | (8'hb1))) - $unsigned(forvar5347)) ?
                          $unsigned(({reg4999} >> $unsigned(reg5133))) : {$unsigned((reg5153 ?
                                  forvar5074 : reg5010))});
                    end
                end
              for (forvar5373 = (1'h0); (forvar5373 < (2'h2)); forvar5373 = (forvar5373 + (1'h1)))
                begin
                  reg5374 <= $unsigned(reg5058);
                  for (forvar5375 = (1'h0); (forvar5375 < (2'h2)); forvar5375 = (forvar5375 + (1'h1)))
                    begin
                      reg5376 <= reg4975[(3'h4):(2'h2)];
                      reg5377 <= (~|{(reg5145 >= (|forvar5281))});
                    end
                end
            end
          for (forvar5378 = (1'h0); (forvar5378 < (1'h1)); forvar5378 = (forvar5378 + (1'h1)))
            begin
              if ((~&{($signed(forvar5055) * $signed(reg5303))}))
                begin
                  reg5379 <= $signed(reg5085);
                end
              else
                begin
                  for (forvar5379 = (1'h0); (forvar5379 < (1'h1)); forvar5379 = (forvar5379 + (1'h1)))
                    begin
                      reg5380 <= (($signed((reg5325 >> forvar5337)) ?
                              (|$unsigned(reg5298)) : (!(|reg5205))) ?
                          $unsigned(((-reg5293) ~^ wire4969)) : (^(^~reg5057)));
                    end
                  for (forvar5381 = (1'h0); (forvar5381 < (1'h0)); forvar5381 = (forvar5381 + (1'h1)))
                    begin
                      reg5382 <= reg5275[(4'hd):(4'hc)];
                    end
                  if ($signed(($unsigned($unsigned(forvar5165)) ?
                      $signed(reg5118) : ($signed(reg5343) ~^ $unsigned((8'h9e))))))
                    begin
                      reg5383 <= (-(!((reg5008 ?
                          reg5173 : forvar5033) + reg5300)));
                      reg5384 <= $unsigned({(reg5259[(3'h6):(3'h6)] ^~ $signed((8'hab)))});
                      reg5385 <= (^(^{(8'h9f)}));
                    end
                  else
                    begin
                      reg5383 <= (reg5123[(2'h2):(1'h1)] ~^ forvar5278);
                      reg5384 <= reg5058[(2'h2):(1'h0)];
                    end
                end
              if ($signed($signed(forvar5341[(1'h1):(1'h0)])))
                begin
                  if ($signed(((|$unsigned(reg5297)) != $signed(reg5282))))
                    begin
                      reg5386 <= $signed((reg5286 > $unsigned((^~(8'ha0)))));
                    end
                  else
                    begin
                      reg5386 <= (~|reg5010[(4'he):(3'h7)]);
                      reg5387 <= ($signed((~forvar5329)) ? (8'h9d) : reg5281);
                      reg5388 <= (((-(reg5283 ?
                              reg5221 : reg5306)) <= (+$unsigned(forvar5252))) ?
                          reg5072 : ($signed((forvar5051 ? reg5350 : reg5280)) ?
                              (^(+(8'ha0))) : (+$unsigned(reg5032))));
                    end
                  if ($unsigned((|{(reg5099 ? forvar5375 : reg5108)})))
                    begin
                      reg5389 <= {$signed(reg5385)};
                      reg5390 <= (|(reg5078 * $unsigned($signed(reg5298))));
                      reg5391 <= (+(8'ha4));
                    end
                  else
                    begin
                      reg5389 <= $signed(reg4976);
                      reg5390 <= reg5355;
                    end
                end
              else
                begin
                  if (reg4976[(1'h0):(1'h0)])
                    begin
                      reg5386 <= ($unsigned(($signed((8'hac)) ?
                              $unsigned(forvar5202) : (reg5091 >= (8'hab)))) ?
                          reg5093 : reg4996);
                      reg5387 <= (!$unsigned($unsigned(reg5173[(3'h4):(1'h0)])));
                    end
                  else
                    begin
                      reg5386 <= {($signed((forvar5040 ?
                              (8'h9f) : reg5352)) ~^ forvar5343)};
                      reg5387 <= (^wire1024[(3'h4):(1'h0)]);
                    end
                  for (forvar5388 = (1'h0); (forvar5388 < (1'h0)); forvar5388 = (forvar5388 + (1'h1)))
                    begin
                      reg5389 <= $unsigned((~$unsigned($signed(forvar5379))));
                      reg5390 <= {(-((wire4967 ? reg5325 : forvar5236) ?
                              reg4976[(1'h0):(1'h0)] : reg5215[(3'h4):(2'h2)]))};
                      reg5391 <= (8'hb8);
                      reg5392 <= $signed(((|$signed(reg5214)) == $unsigned((&reg5162))));
                    end
                  reg5393 <= $unsigned(($unsigned(((8'ha8) != reg5332)) << ((reg5067 != reg5026) ?
                      (reg5271 != reg5168) : reg5219)));
                end
              if (reg5390[(2'h3):(2'h2)])
                begin
                  if (reg5297[(3'h7):(3'h7)])
                    begin
                      reg5394 <= (-$signed(forvar5201));
                      reg5395 <= (8'h9f);
                    end
                  else
                    begin
                      reg5394 <= ((((reg5133 ? forvar5033 : reg5299) ?
                              $signed(reg5356) : $unsigned(forvar5295)) ?
                          $unsigned({forvar5378}) : $signed((~&forvar5234))) - (((reg5383 ?
                              forvar5033 : reg5146) ?
                          $signed(reg5349) : (8'hb7)) + (((8'hb5) ?
                              reg5352 : reg5298) ?
                          reg5244 : wire1029)));
                    end
                  reg5396 <= $signed(reg5387[(1'h1):(1'h1)]);
                  for (forvar5397 = (1'h0); (forvar5397 < (2'h2)); forvar5397 = (forvar5397 + (1'h1)))
                    begin
                      reg5398 <= (-((+reg5093[(2'h3):(1'h0)]) ?
                          reg5183 : (reg5241 ? reg5316 : (reg5296 * reg4976))));
                      reg5399 <= ({({(8'hb3)} & ((8'ha2) ?
                                  reg5241 : reg5212))} ?
                          $signed($unsigned({(8'ha5)})) : ($unsigned(reg5281[(2'h2):(2'h2)]) ?
                              $signed(reg5105[(1'h0):(1'h0)]) : ((reg5213 | reg5248) ?
                                  forvar5098[(1'h1):(1'h0)] : ((8'ha0) ?
                                      reg5150 : reg5062))));
                    end
                  reg5400 <= (reg5112[(1'h0):(1'h0)] ?
                      reg5356 : reg5317[(2'h3):(1'h0)]);
                end
              else
                begin
                  for (forvar5394 = (1'h0); (forvar5394 < (1'h0)); forvar5394 = (forvar5394 + (1'h1)))
                    begin
                      reg5395 <= $unsigned(forvar5249);
                      reg5396 <= $unsigned((reg5255 << (-(~|forvar5210))));
                    end
                end
            end
        end
      if (reg5274[(4'h8):(2'h3)])
        begin
          for (forvar5401 = (1'h0); (forvar5401 < (1'h0)); forvar5401 = (forvar5401 + (1'h1)))
            begin
              if ((~&reg5334[(2'h2):(2'h2)]))
                begin
                  for (forvar5402 = (1'h0); (forvar5402 < (2'h3)); forvar5402 = (forvar5402 + (1'h1)))
                    begin
                      reg5403 <= ((^~(((8'hb5) ?
                              reg5393 : (8'hb0)) >>> (forvar5095 ?
                              (8'hb4) : forvar5227))) ?
                          $signed({(reg5245 ?
                                  forvar5061 : reg5389)}) : forvar5397[(1'h0):(1'h0)]);
                      reg5404 <= reg5107;
                    end
                  for (forvar5405 = (1'h0); (forvar5405 < (2'h3)); forvar5405 = (forvar5405 + (1'h1)))
                    begin
                      reg5406 <= ((((forvar5227 != reg5389) + reg5289[(4'hc):(1'h1)]) != (((8'h9c) >>> reg5102) >> $signed(reg5250))) ?
                          {(((8'ha2) ?
                                  (8'hb6) : reg5192) <= reg5151)} : $signed(reg5008[(3'h6):(2'h2)]));
                      reg5407 <= (8'hac);
                      reg5408 <= $unsigned((+(forvar5187 ?
                          $unsigned((8'hb1)) : (~|reg5148))));
                      reg5409 <= (forvar5298 * (($signed(forvar5081) ^~ $signed((8'ha7))) <<< (((8'ha6) + (8'ha7)) - (&forvar5187))));
                    end
                end
              else
                begin
                  if (forvar5272[(2'h3):(2'h2)])
                    begin
                      reg5402 <= forvar5037[(1'h0):(1'h0)];
                      reg5403 <= reg5402;
                      reg5404 <= $unsigned($unsigned((~&$unsigned(reg5250))));
                    end
                  else
                    begin
                      reg5402 <= (({(^reg4978)} + reg5008[(3'h6):(2'h3)]) - reg5130[(1'h1):(1'h1)]);
                      reg5403 <= $signed(forvar4970);
                      reg5404 <= reg5125;
                      reg5405 <= reg5100;
                    end
                  if ($signed(reg5142[(4'h9):(3'h6)]))
                    begin
                      reg5406 <= (({(reg5262 ? forvar5238 : reg5371)} ?
                              reg5025[(2'h3):(1'h0)] : $signed((reg5188 ?
                                  forvar4972 : (8'hb6)))) ?
                          $unsigned($unsigned(reg5140[(1'h1):(1'h0)])) : $signed($unsigned(reg5329)));
                      reg5407 <= reg5030[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg5406 <= reg5352;
                      reg5407 <= reg5118[(2'h3):(2'h3)];
                      reg5408 <= $signed(reg5113[(2'h3):(2'h2)]);
                    end
                end
              for (forvar5410 = (1'h0); (forvar5410 < (1'h1)); forvar5410 = (forvar5410 + (1'h1)))
                begin
                  reg5411 <= $signed(reg5075);
                  for (forvar5412 = (1'h0); (forvar5412 < (1'h1)); forvar5412 = (forvar5412 + (1'h1)))
                    begin
                      reg5413 <= reg5232[(3'h6):(2'h2)];
                    end
                end
              for (forvar5414 = (1'h0); (forvar5414 < (1'h0)); forvar5414 = (forvar5414 + (1'h1)))
                begin
                  if ((reg5244[(4'hb):(4'h8)] <= $signed((-forvar4996[(1'h1):(1'h0)]))))
                    begin
                      reg5415 <= (-{{$unsigned(reg5311)}});
                      reg5416 <= ($signed(reg5271) ?
                          $signed((^(|(8'h9e)))) : forvar5227[(3'h7):(3'h6)]);
                      reg5417 <= ((~|reg5148[(3'h4):(1'h1)]) != ($unsigned(((8'ha2) ?
                              forvar5234 : reg5382)) ?
                          forvar5260[(3'h6):(2'h3)] : $signed((~|reg5187))));
                      reg5418 <= (~(~$unsigned($signed((8'ha3)))));
                    end
                  else
                    begin
                      reg5415 <= (($signed($signed(reg5218)) * ((reg5129 + reg5263) > $signed((8'ha0)))) | $signed($signed((reg5233 ?
                          reg5168 : reg5107))));
                      reg5416 <= reg5086;
                      reg5417 <= reg5303;
                      reg5418 <= $unsigned($signed($unsigned((&reg5304))));
                    end
                end
              if ({((8'ha1) >>> {(+forvar4986)})})
                begin
                  for (forvar5419 = (1'h0); (forvar5419 < (1'h1)); forvar5419 = (forvar5419 + (1'h1)))
                    begin
                      reg5420 <= $signed(forvar5183[(1'h1):(1'h0)]);
                      reg5421 <= $signed(reg5049[(2'h3):(1'h1)]);
                    end
                  for (forvar5422 = (1'h0); (forvar5422 < (2'h3)); forvar5422 = (forvar5422 + (1'h1)))
                    begin
                      reg5423 <= {wire1025};
                      reg5424 <= (8'ha8);
                      reg5425 <= (reg5224 ? reg5169[(3'h7):(1'h0)] : reg5246);
                      reg5426 <= {{reg4975}};
                    end
                  for (forvar5427 = (1'h0); (forvar5427 < (1'h0)); forvar5427 = (forvar5427 + (1'h1)))
                    begin
                      reg5428 <= $unsigned(reg5004);
                      reg5429 <= ((+$unsigned((^reg5108))) ?
                          reg5369[(1'h0):(1'h0)] : $signed($signed({reg5115})));
                    end
                end
              else
                begin
                  for (forvar5419 = (1'h0); (forvar5419 < (2'h3)); forvar5419 = (forvar5419 + (1'h1)))
                    begin
                      reg5420 <= ($unsigned((~(reg5059 <<< reg5015))) ?
                          reg5035 : (8'hb6));
                      reg5421 <= (reg5335[(3'h4):(2'h3)] ?
                          (reg5117 ?
                              ((reg5407 || wire5336) ?
                                  wire3538[(3'h5):(1'h1)] : (&reg5329)) : reg5130[(3'h4):(1'h1)]) : ((~&$unsigned(reg5133)) <<< ((~^forvar5236) * $unsigned(reg5361))));
                      reg5422 <= $signed((|(8'hba)));
                      reg5423 <= reg5310[(4'hf):(3'h7)];
                    end
                  if (reg5244)
                    begin
                      reg5424 <= (forvar5082 ?
                          (forvar5323 < reg5085[(4'hd):(1'h0)]) : {((reg5294 ?
                                      reg4972 : (8'hac)) ?
                                  (reg5122 ?
                                      reg5243 : reg5296) : (~&reg5137))});
                    end
                  else
                    begin
                      reg5424 <= $unsigned($signed(reg5379[(2'h2):(1'h1)]));
                      reg5425 <= $unsigned(reg5341);
                      reg5426 <= $signed((-(reg5104 >> (~reg5246))));
                      reg5427 <= $signed($unsigned((((8'hb9) ?
                              reg5058 : reg5332) ?
                          $unsigned(reg5140) : ((8'hba) ^ reg5303))));
                    end
                  if ($unsigned($signed($unsigned($unsigned(forvar5240)))))
                    begin
                      reg5428 <= ($signed($unsigned($signed(reg5166))) & $signed(reg5054));
                      reg5429 <= $unsigned((-forvar5055));
                      reg5430 <= forvar5141[(3'h4):(1'h1)];
                      reg5431 <= (reg5077 ?
                          reg5108 : ({(reg4984 ?
                                  forvar5288 : reg5086)} ^ $signed($unsigned(reg5093))));
                    end
                  else
                    begin
                      reg5428 <= reg5351[(3'h4):(1'h1)];
                      reg5429 <= reg5153[(3'h5):(2'h2)];
                      reg5430 <= reg5072[(2'h3):(2'h2)];
                    end
                  for (forvar5432 = (1'h0); (forvar5432 < (2'h2)); forvar5432 = (forvar5432 + (1'h1)))
                    begin
                      reg5433 <= ($unsigned($unsigned($unsigned(reg5318))) ^~ $unsigned(((reg5264 >= reg5221) ^ (reg5126 ?
                          reg5427 : (8'ha1)))));
                      reg5434 <= $unsigned((8'ha9));
                      reg5435 <= (reg5216[(3'h5):(1'h1)] <= $unsigned($signed(reg5109)));
                    end
                end
            end
          for (forvar5436 = (1'h0); (forvar5436 < (1'h1)); forvar5436 = (forvar5436 + (1'h1)))
            begin
              if ({($unsigned(forvar5160) ?
                      {forvar5362} : $unsigned((forvar5074 ?
                          reg5271 : forvar5109)))})
                begin
                  reg5437 <= (&(reg5396[(2'h2):(2'h2)] <<< $signed({forvar5397})));
                  for (forvar5438 = (1'h0); (forvar5438 < (2'h3)); forvar5438 = (forvar5438 + (1'h1)))
                    begin
                      reg5439 <= (^$signed($unsigned((reg5203 ?
                          forvar5183 : reg5308))));
                    end
                  for (forvar5440 = (1'h0); (forvar5440 < (2'h2)); forvar5440 = (forvar5440 + (1'h1)))
                    begin
                      reg5441 <= reg5346;
                      reg5442 <= (reg5188 + $signed($unsigned($unsigned(reg5395))));
                      reg5443 <= ((-{(8'had)}) ?
                          (~|$unsigned((reg5316 >> reg5344))) : $signed((reg5312[(3'h7):(1'h1)] ?
                              (reg5367 << reg5271) : $signed((8'h9c)))));
                      reg5444 <= $unsigned(reg5117[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar5437 = (1'h0); (forvar5437 < (2'h3)); forvar5437 = (forvar5437 + (1'h1)))
                    begin
                      reg5438 <= {$unsigned(reg5356[(1'h1):(1'h1)])};
                      reg5439 <= (reg5003[(3'h4):(3'h4)] ^~ (8'ha4));
                    end
                  for (forvar5440 = (1'h0); (forvar5440 < (2'h2)); forvar5440 = (forvar5440 + (1'h1)))
                    begin
                      reg5441 <= reg5029[(2'h3):(2'h3)];
                      reg5442 <= forvar4972[(1'h1):(1'h0)];
                      reg5443 <= $signed($signed({$unsigned(reg5348)}));
                    end
                end
            end
          for (forvar5445 = (1'h0); (forvar5445 < (1'h1)); forvar5445 = (forvar5445 + (1'h1)))
            begin
              reg5446 <= {$unsigned($signed(reg5399[(2'h2):(1'h0)]))};
            end
          for (forvar5447 = (1'h0); (forvar5447 < (1'h1)); forvar5447 = (forvar5447 + (1'h1)))
            begin
              for (forvar5448 = (1'h0); (forvar5448 < (2'h3)); forvar5448 = (forvar5448 + (1'h1)))
                begin
                  reg5449 <= (~(~^reg5056[(1'h0):(1'h0)]));
                  reg5450 <= reg5328;
                  for (forvar5451 = (1'h0); (forvar5451 < (2'h2)); forvar5451 = (forvar5451 + (1'h1)))
                    begin
                      reg5452 <= (|{(~^reg5184)});
                      reg5453 <= (reg4971 ?
                          ($signed($signed(reg5350)) * (&$signed(forvar5030))) : (forvar5410 || $signed(reg5186[(3'h4):(2'h3)])));
                    end
                end
            end
        end
      else
        begin
          for (forvar5401 = (1'h0); (forvar5401 < (1'h1)); forvar5401 = (forvar5401 + (1'h1)))
            begin
              reg5402 <= (8'hb8);
              for (forvar5403 = (1'h0); (forvar5403 < (1'h1)); forvar5403 = (forvar5403 + (1'h1)))
                begin
                  for (forvar5404 = (1'h0); (forvar5404 < (2'h3)); forvar5404 = (forvar5404 + (1'h1)))
                    begin
                      reg5405 <= (($unsigned((forvar5090 <<< (8'hb2))) ~^ $signed((&reg5105))) << $signed(forvar5088[(3'h4):(1'h1)]));
                      reg5406 <= {(reg5333 ?
                              reg5335 : (~|$unsigned(forvar5227)))};
                    end
                  for (forvar5407 = (1'h0); (forvar5407 < (1'h0)); forvar5407 = (forvar5407 + (1'h1)))
                    begin
                      reg5408 <= reg5062;
                      reg5409 <= ((^~{(forvar4982 ?
                              forvar5347 : forvar5089)}) & {forvar5227});
                      reg5410 <= ($unsigned($unsigned((reg5109 >= reg5205))) || forvar5324);
                    end
                end
              if (reg4984[(4'hb):(2'h3)])
                begin
                  for (forvar5411 = (1'h0); (forvar5411 < (2'h3)); forvar5411 = (forvar5411 + (1'h1)))
                    begin
                      reg5412 <= reg5215;
                      reg5413 <= (~&reg5356[(2'h3):(2'h2)]);
                    end
                  if (($unsigned(((reg4981 ?
                      reg5366 : reg5059) == forvar5047)) | ((8'ha2) ^~ (8'ha4))))
                    begin
                      reg5414 <= ($unsigned(({reg5274} < $signed(reg5335))) ?
                          ({(~^reg5311)} || $unsigned($signed((8'h9e)))) : (8'h9d));
                      reg5415 <= ({((reg5027 ? forvar5236 : reg5274) ?
                              reg5235[(3'h6):(2'h2)] : reg5367)} ^~ (reg5032 ?
                          $signed($unsigned(reg5355)) : $signed((^~reg5187))));
                      reg5416 <= ((~|((reg5371 + forvar5404) - $unsigned(reg4993))) ?
                          (((8'hb3) ? wire1025 : reg5057[(4'h9):(3'h5)]) ?
                              $signed($signed(forvar5051)) : reg5415[(3'h5):(3'h4)]) : $unsigned($unsigned(reg5310[(4'h9):(3'h7)])));
                      reg5417 <= {forvar5403[(2'h3):(2'h2)]};
                    end
                  else
                    begin
                      reg5414 <= $signed({(8'h9e)});
                      reg5415 <= ({reg5370[(2'h3):(1'h1)]} == (^({reg5308} ?
                          reg5342[(1'h0):(1'h0)] : $signed(reg5363))));
                      reg5416 <= (&$unsigned(forvar5271[(1'h0):(1'h0)]));
                    end
                  for (forvar5418 = (1'h0); (forvar5418 < (2'h2)); forvar5418 = (forvar5418 + (1'h1)))
                    begin
                      reg5419 <= reg5149;
                      reg5420 <= reg5296;
                      reg5421 <= reg5263[(2'h2):(1'h1)];
                      reg5422 <= reg4998;
                    end
                  reg5423 <= (!(~|((forvar4971 ^~ forvar5172) & reg5408)));
                end
              else
                begin
                  if (forvar5001)
                    begin
                      reg5411 <= ({((~reg5232) ?
                              forvar5165 : ((8'ha5) ?
                                  forvar5179 : forvar5360))} << (!(!$unsigned(reg5426))));
                      reg5412 <= $unsigned(reg5034[(2'h2):(2'h2)]);
                      reg5413 <= ($unsigned($unsigned(((8'ha2) << reg5355))) ?
                          {($signed((8'h9f)) << reg5093)} : {$unsigned(forvar5260[(1'h1):(1'h0)])});
                    end
                  else
                    begin
                      reg5411 <= reg5077[(2'h2):(1'h0)];
                    end
                end
            end
          if ({(reg5006 <<< reg5392)})
            begin
              if ({(~{$signed((8'hab))})})
                begin
                  reg5424 <= $signed(forvar5364);
                  if (forvar5305[(4'h9):(4'h9)])
                    begin
                      reg5425 <= ($signed($signed((reg5028 | reg5428))) | (~^{(~&forvar5182)}));
                      reg5426 <= $signed((reg5369 ^~ (|(reg5303 ?
                          reg5242 : forvar5095))));
                    end
                  else
                    begin
                      reg5425 <= reg5250;
                    end
                  if ({((~^$signed(reg5421)) >> reg5004)})
                    begin
                      reg5427 <= ($unsigned($unsigned(reg5413)) ?
                          ({(^~forvar5159)} && {$unsigned(reg5427)}) : forvar5001);
                      reg5428 <= reg5442;
                      reg5429 <= reg5320;
                    end
                  else
                    begin
                      reg5427 <= {reg5269[(1'h0):(1'h0)]};
                      reg5428 <= reg5032[(4'h8):(4'h8)];
                    end
                  if (forvar5379[(1'h0):(1'h0)])
                    begin
                      reg5430 <= (8'hb8);
                    end
                  else
                    begin
                      reg5430 <= (+(((~|forvar5360) <<< (reg5180 ^ reg5344)) >> forvar5339[(2'h3):(1'h1)]));
                      reg5431 <= reg5093[(1'h0):(1'h0)];
                      reg5432 <= ((reg5258 <= (reg5274[(4'ha):(3'h4)] ?
                              (^~reg5154) : reg5446)) ?
                          {forvar5192} : ((((8'h9c) ^~ forvar5281) ?
                              forvar5404 : $signed(forvar5394)) + (-(reg5446 <= (8'haf)))));
                    end
                end
              else
                begin
                  if ((+((((8'ha6) << reg5430) && $unsigned(reg5155)) ?
                      (reg5344 ?
                          wire3536 : (~^reg5101)) : $signed($unsigned((8'ha3))))))
                    begin
                      reg5424 <= reg5390[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg5424 <= ((reg5328[(2'h3):(2'h2)] ?
                              {(forvar5131 ?
                                      reg5035 : (8'hb2))} : $signed((^~(8'hb9)))) ?
                          forvar4987 : $unsigned(($unsigned(reg5195) ?
                              reg5358[(4'h9):(1'h0)] : $signed(reg5231))));
                    end
                  for (forvar5425 = (1'h0); (forvar5425 < (1'h1)); forvar5425 = (forvar5425 + (1'h1)))
                    begin
                      reg5426 <= (((reg5119[(2'h3):(1'h0)] <= reg5076) ?
                              ({(8'had)} ~^ (reg5168 & reg5371)) : ($unsigned((8'ha9)) * (reg5022 == reg5141))) ?
                          $unsigned(reg5250[(4'h8):(3'h7)]) : forvar5087[(4'h8):(1'h0)]);
                      reg5427 <= (^~(forvar5223 | (|((8'hba) ?
                          reg5109 : reg5389))));
                      reg5428 <= (~|$signed($signed(reg5217)));
                    end
                end
              for (forvar5433 = (1'h0); (forvar5433 < (1'h1)); forvar5433 = (forvar5433 + (1'h1)))
                begin
                  for (forvar5434 = (1'h0); (forvar5434 < (2'h2)); forvar5434 = (forvar5434 + (1'h1)))
                    begin
                      reg5435 <= ($unsigned($unsigned((forvar4972 ?
                              reg5152 : reg5370))) ?
                          reg5442 : (({reg5285} * (reg5122 >= reg5446)) ?
                              ($signed(forvar5432) == $signed(forvar5315)) : $signed($unsigned(reg5433))));
                    end
                  if (forvar5337)
                    begin
                      reg5436 <= $signed((-(^~reg5350[(1'h0):(1'h0)])));
                      reg5437 <= reg5316;
                      reg5438 <= reg5409;
                    end
                  else
                    begin
                      reg5436 <= ((8'h9c) != ($signed(reg5218) ?
                          ((reg5126 ?
                              reg5149 : wire3536) & reg5219[(1'h0):(1'h0)]) : ((reg5392 ?
                                  reg5214 : forvar5281) ?
                              forvar5103 : (8'hb4))));
                      reg5437 <= (($signed((forvar4983 ?
                              (8'hba) : reg5260)) || $unsigned((~&reg4992))) ?
                          (&$unsigned({forvar5347})) : (+(^~forvar5172)));
                      reg5438 <= {(forvar5405[(1'h0):(1'h0)] ?
                              ((^forvar5047) ?
                                  $unsigned(reg5108) : (forvar5016 <<< (8'ha7))) : (|((8'hb7) ?
                                  reg5281 : forvar5033)))};
                      reg5439 <= (reg5348 ?
                          (reg5148[(3'h5):(1'h0)] >= $signed(reg1026)) : $signed($signed((reg5444 ^ reg4975))));
                    end
                end
              reg5440 <= reg5379;
              for (forvar5441 = (1'h0); (forvar5441 < (1'h1)); forvar5441 = (forvar5441 + (1'h1)))
                begin
                  if (reg5063)
                    begin
                      reg5442 <= reg5148;
                      reg5443 <= reg5193[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg5442 <= (&$unsigned({((8'ha7) ~^ (8'h9d))}));
                    end
                end
            end
          else
            begin
              reg5424 <= reg5380;
            end
        end
      for (forvar5454 = (1'h0); (forvar5454 < (2'h3)); forvar5454 = (forvar5454 + (1'h1)))
        begin
          if ((reg5185 ?
              (~($signed(reg5365) ?
                  (reg4975 && (8'haa)) : (|reg5211))) : (+reg5176)))
            begin
              if ((&{reg5366[(2'h3):(2'h3)]}))
                begin
                  reg5455 <= $signed((~|((8'ha2) <<< {reg5120})));
                  for (forvar5456 = (1'h0); (forvar5456 < (2'h2)); forvar5456 = (forvar5456 + (1'h1)))
                    begin
                      reg5457 <= (($unsigned($signed((8'ha1))) ?
                              forvar4989[(4'hb):(4'hb)] : (~&{reg5279})) ?
                          (((|forvar5037) << reg5420) << forvar4972[(4'h9):(1'h0)]) : (8'hb4));
                    end
                  if (forvar4983[(1'h0):(1'h0)])
                    begin
                      reg5458 <= $signed(reg5100);
                    end
                  else
                    begin
                      reg5458 <= reg5003[(4'h8):(1'h0)];
                    end
                  reg5459 <= $unsigned(((8'ha5) <= ((reg5303 ?
                          (8'ha9) : forvar5182) ?
                      $unsigned(reg5150) : (~reg5302))));
                end
              else
                begin
                  for (forvar5455 = (1'h0); (forvar5455 < (2'h2)); forvar5455 = (forvar5455 + (1'h1)))
                    begin
                      reg5456 <= $unsigned((reg5253[(1'h0):(1'h0)] ?
                          $unsigned(reg5351[(2'h2):(1'h0)]) : $unsigned($unsigned(forvar5082))));
                      reg5457 <= $signed(reg5285);
                      reg5458 <= $unsigned($unsigned((~^(~^reg5152))));
                      reg5459 <= $unsigned((((^reg5299) ?
                              ((8'hb0) ?
                                  wire1025 : (8'haf)) : reg4973[(3'h5):(2'h2)]) ?
                          $unsigned((~|reg4997)) : forvar5226[(1'h0):(1'h0)]));
                    end
                  for (forvar5460 = (1'h0); (forvar5460 < (2'h3)); forvar5460 = (forvar5460 + (1'h1)))
                    begin
                      reg5461 <= forvar5270[(2'h3):(1'h1)];
                      reg5462 <= {reg5152[(3'h4):(2'h3)]};
                      reg5463 <= $signed({$signed((reg5333 ?
                              reg5145 : reg5415))});
                      reg5464 <= (!forvar5210[(1'h1):(1'h0)]);
                    end
                end
              reg5465 <= reg5348[(3'h4):(1'h1)];
              reg5466 <= (+$unsigned(((reg5382 ?
                  (8'h9e) : reg5218) && (-(8'hba)))));
              reg5467 <= ($unsigned((^(8'h9c))) ?
                  ($unsigned(reg5356) ?
                      ($signed(forvar5323) >>> (forvar5460 ?
                          (8'hb7) : reg5118)) : $unsigned({reg5450})) : reg5026[(1'h0):(1'h0)]);
            end
          else
            begin
              if ((~forvar5270[(1'h1):(1'h0)]))
                begin
                  for (forvar5455 = (1'h0); (forvar5455 < (1'h1)); forvar5455 = (forvar5455 + (1'h1)))
                    begin
                      reg5456 <= (!forvar5117);
                      reg5457 <= ((((reg5214 - reg5449) && forvar5175) ?
                              reg5431 : reg5044[(3'h7):(3'h5)]) ?
                          ((|{reg5466}) ?
                              (&(^reg5170)) : reg5467[(2'h2):(1'h1)]) : forvar5018);
                      reg5458 <= reg5067;
                    end
                  reg5459 <= (((reg5120[(4'h8):(2'h2)] << $signed((8'ha1))) != $unsigned((!reg5069))) >= (((forvar5270 > reg5344) * (!reg4997)) ^ (~|reg5182)));
                end
              else
                begin
                  for (forvar5455 = (1'h0); (forvar5455 < (2'h2)); forvar5455 = (forvar5455 + (1'h1)))
                    begin
                      reg5456 <= $unsigned((^~wire1029));
                      reg5457 <= reg5298;
                      reg5458 <= (((^~((8'hb2) >= reg5341)) + reg5125) ?
                          (~($unsigned(reg5345) & $unsigned(forvar5139))) : (~|forvar5375[(2'h3):(2'h3)]));
                    end
                  for (forvar5459 = (1'h0); (forvar5459 < (1'h0)); forvar5459 = (forvar5459 + (1'h1)))
                    begin
                      reg5460 <= $signed((!(^(forvar5252 ?
                          reg5217 : (8'hac)))));
                      reg5461 <= forvar5196[(3'h5):(3'h4)];
                    end
                end
            end
          if ($signed((8'ha3)))
            begin
              if ((({reg5204[(2'h3):(1'h1)]} + reg5383) ?
                  {$signed((reg5409 && (8'hb8)))} : {reg5347}))
                begin
                  if ($signed(forvar4978))
                    begin
                      reg5468 <= ($signed({$unsigned(forvar5046)}) ?
                          (({(8'ha7)} >= reg5440) << ($unsigned(reg5346) + $unsigned(reg5166))) : reg5225);
                      reg5469 <= $signed(($unsigned({reg5100}) ?
                          $signed((^reg5200)) : (&(8'hae))));
                      reg5470 <= $unsigned($signed(($unsigned(reg5276) + $unsigned(reg5331))));
                    end
                  else
                    begin
                      reg5468 <= (~&(^~$signed((8'h9f))));
                      reg5469 <= (forvar5046[(4'ha):(4'ha)] ?
                          reg5043 : {($unsigned(reg5269) ?
                                  reg5028 : (reg5271 >= forvar5117))});
                    end
                end
              else
                begin
                  if ((~&$unsigned($unsigned((reg5216 ?
                      reg5416 : forvar5338)))))
                    begin
                      reg5468 <= (+($unsigned($signed(forvar5210)) ?
                          $unsigned((~(8'h9f))) : forvar5223[(3'h7):(2'h3)]));
                      reg5469 <= (&((&(reg5036 != forvar5088)) ?
                          (forvar5364[(4'hc):(3'h6)] >>> (forvar5278 ?
                              reg5073 : reg5013)) : (((8'ha4) >= reg5091) ?
                              (forvar5082 == reg5428) : (forvar5079 > (8'hb4)))));
                      reg5470 <= $signed($signed((~|(reg5031 >> forvar5447))));
                      reg5471 <= (8'hb4);
                    end
                  else
                    begin
                      reg5468 <= (reg5026[(4'h9):(3'h4)] & $unsigned(($unsigned((8'hb4)) ?
                          (forvar5045 != (8'ha3)) : $unsigned(reg4980))));
                      reg5469 <= $signed(reg4980[(1'h1):(1'h1)]);
                      reg5470 <= (reg5094 ?
                          reg5063[(2'h2):(1'h0)] : $signed(((!forvar5208) ?
                              (8'hb2) : reg5168[(3'h6):(3'h6)])));
                    end
                  if ($signed((reg5446 != {(~&reg5049)})))
                    begin
                      reg5472 <= ((^(-reg4991)) ?
                          ((~&reg5331) ?
                              $signed((~&reg5417)) : ((reg5367 ?
                                  forvar5455 : wire1030) > $signed(forvar5412))) : reg5221);
                      reg5473 <= (reg5329 ?
                          ($signed(forvar5255[(4'hf):(4'h9)]) <<< forvar5201) : $unsigned($unsigned(reg5114)));
                    end
                  else
                    begin
                      reg5472 <= $signed(reg5200);
                    end
                  for (forvar5474 = (1'h0); (forvar5474 < (2'h2)); forvar5474 = (forvar5474 + (1'h1)))
                    begin
                      reg5475 <= {$unsigned(((forvar5051 >> reg5217) ^~ (reg5386 ^ forvar5156)))};
                      reg5476 <= wire4969[(4'ha):(4'ha)];
                      reg5477 <= (-$signed(reg4975[(3'h7):(1'h1)]));
                      reg5478 <= $unsigned($unsigned(((reg5100 | reg5340) | (reg5100 ?
                          reg5246 : forvar5419))));
                    end
                  reg5479 <= $signed(((forvar4971[(3'h5):(2'h2)] & wire5336) * $unsigned(((8'hb0) ?
                      reg5124 : (8'hb5)))));
                end
              if ($unsigned(forvar5474[(3'h5):(1'h0)]))
                begin
                  for (forvar5480 = (1'h0); (forvar5480 < (2'h3)); forvar5480 = (forvar5480 + (1'h1)))
                    begin
                      reg5481 <= $unsigned((!$unsigned(forvar5016[(3'h6):(1'h1)])));
                      reg5482 <= (8'ha7);
                    end
                  if ($signed(($signed((forvar5460 ?
                      forvar4972 : reg4971)) >> ({reg5171} || (reg5261 && reg5411)))))
                    begin
                      reg5483 <= (~|($unsigned((reg5215 == (8'haa))) > (reg5038[(2'h3):(2'h2)] || ((8'ha2) ?
                          forvar5447 : forvar5359))));
                      reg5484 <= reg5479[(4'hb):(4'h8)];
                      reg5485 <= reg5259;
                      reg5486 <= (+(((8'hb3) == (reg5313 >>> reg5012)) && (^~(8'hb0))));
                    end
                  else
                    begin
                      reg5483 <= $unsigned($signed($unsigned((reg5077 ?
                          reg5129 : reg5483))));
                      reg5484 <= (reg5228[(3'h4):(1'h0)] * ($signed((reg5189 ?
                          forvar5117 : forvar5238)) * forvar5042));
                      reg5485 <= {$signed((8'ha7))};
                    end
                end
              else
                begin
                  for (forvar5480 = (1'h0); (forvar5480 < (1'h0)); forvar5480 = (forvar5480 + (1'h1)))
                    begin
                      reg5481 <= ((($signed(reg5403) ?
                                  $signed(forvar5407) : reg5382) ?
                              $signed(reg5032) : $unsigned(reg5346[(4'ha):(3'h5)])) ?
                          {reg5344} : $unsigned({(|(8'haa))}));
                      reg5482 <= $unsigned($unsigned($signed(reg5456)));
                      reg5483 <= ((~|((^forvar5480) << (reg5363 <<< reg5467))) ?
                          $signed(forvar5373[(1'h1):(1'h1)]) : ((!$signed(forvar4996)) ?
                              $unsigned((forvar5440 ?
                                  reg5113 : (8'hba))) : reg5371[(1'h1):(1'h1)]));
                    end
                  for (forvar5484 = (1'h0); (forvar5484 < (1'h0)); forvar5484 = (forvar5484 + (1'h1)))
                    begin
                      reg5485 <= reg5406[(1'h1):(1'h1)];
                      reg5486 <= $signed((|$unsigned($unsigned(reg5176))));
                      reg5487 <= (8'hb3);
                    end
                end
              for (forvar5488 = (1'h0); (forvar5488 < (1'h0)); forvar5488 = (forvar5488 + (1'h1)))
                begin
                  for (forvar5489 = (1'h0); (forvar5489 < (2'h3)); forvar5489 = (forvar5489 + (1'h1)))
                    begin
                      reg5490 <= wire1022[(4'h8):(2'h3)];
                      reg5491 <= (reg5424 && $signed(((~&reg5129) ^ reg5012[(1'h0):(1'h0)])));
                      reg5492 <= forvar5292;
                      reg5493 <= ($signed($unsigned((forvar5319 >= (8'hac)))) ?
                          $unsigned($signed($signed(reg5180))) : $unsigned(((&wire5291) == (forvar5298 != reg5463))));
                    end
                  reg5494 <= forvar5161[(1'h1):(1'h0)];
                  for (forvar5495 = (1'h0); (forvar5495 < (2'h3)); forvar5495 = (forvar5495 + (1'h1)))
                    begin
                      reg5496 <= {$signed(reg5321)};
                      reg5497 <= reg5413[(3'h7):(3'h6)];
                      reg5498 <= (reg5071[(1'h1):(1'h0)] ?
                          {forvar4987[(2'h2):(1'h0)]} : forvar5271);
                    end
                end
            end
          else
            begin
              for (forvar5468 = (1'h0); (forvar5468 < (1'h0)); forvar5468 = (forvar5468 + (1'h1)))
                begin
                  for (forvar5469 = (1'h0); (forvar5469 < (2'h3)); forvar5469 = (forvar5469 + (1'h1)))
                    begin
                      reg5470 <= {$signed(reg5142)};
                      reg5471 <= {{reg5485}};
                      reg5472 <= (~&$signed(($signed(forvar5338) ?
                          reg5152[(3'h7):(3'h4)] : (8'ha9))));
                      reg5473 <= $unsigned($signed((8'hb7)));
                    end
                  for (forvar5474 = (1'h0); (forvar5474 < (2'h2)); forvar5474 = (forvar5474 + (1'h1)))
                    begin
                      reg5475 <= {(((wire1025 ?
                              (8'haa) : forvar5480) & (8'ha5)) * $unsigned(reg5494))};
                      reg5476 <= forvar5402;
                      reg5477 <= ((8'hb4) + forvar5407);
                    end
                end
              for (forvar5478 = (1'h0); (forvar5478 < (1'h0)); forvar5478 = (forvar5478 + (1'h1)))
                begin
                  reg5479 <= $unsigned((forvar5427 ^~ forvar5037[(3'h4):(3'h4)]));
                end
              if ((forvar5159 != (8'h9f)))
                begin
                  for (forvar5480 = (1'h0); (forvar5480 < (2'h3)); forvar5480 = (forvar5480 + (1'h1)))
                    begin
                      reg5481 <= ((~^(^((8'hb8) ?
                          (8'ha0) : (8'haf)))) > reg5427);
                      reg5482 <= $signed((forvar5410[(4'h9):(3'h7)] ?
                          reg5189[(3'h7):(1'h0)] : {reg5004[(2'h3):(2'h2)]}));
                      reg5483 <= reg5112[(1'h0):(1'h0)];
                      reg5484 <= $unsigned((~|$unsigned((^~(8'hba)))));
                    end
                  if (reg5004)
                    begin
                      reg5485 <= ($signed(reg5049[(3'h4):(1'h1)]) <= $unsigned(({forvar5484} ?
                          reg5439[(2'h2):(1'h0)] : ((8'ha2) ?
                              reg5369 : forvar5468))));
                      reg5486 <= $unsigned(($signed({reg5119}) ?
                          ((reg5310 ^~ reg5197) ?
                              (^forvar5165) : (reg5135 != reg5459)) : forvar5160[(4'hb):(3'h6)]));
                      reg5487 <= ($unsigned($unsigned($signed((8'h9e)))) <= {$signed((reg5486 == reg5347))});
                      reg5488 <= reg5278;
                    end
                  else
                    begin
                      reg5485 <= forvar5172;
                      reg5486 <= {$signed(reg5438[(3'h4):(1'h1)])};
                      reg5487 <= forvar5167[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  if ((wire3538 ~^ forvar5422))
                    begin
                      reg5480 <= ((~&$signed(reg5133[(2'h2):(2'h2)])) <<< (8'haa));
                      reg5481 <= (^~(+forvar5488[(3'h6):(2'h3)]));
                      reg5482 <= {{reg5282}};
                      reg5483 <= (reg1026 ?
                          $signed($unsigned(((8'hab) << reg5197))) : (~^(!$unsigned((8'ha5)))));
                    end
                  else
                    begin
                      reg5480 <= ($unsigned(reg5193) ?
                          (~((forvar5276 ? reg5333 : forvar5255) ?
                              (^~reg5403) : (^~reg5162))) : reg5387);
                      reg5481 <= ($unsigned(reg5469[(1'h1):(1'h1)]) << forvar4971[(4'ha):(3'h6)]);
                      reg5482 <= (&($signed((reg5195 <<< reg5052)) != (-reg4974)));
                      reg5483 <= ($signed((forvar4996 ?
                              forvar4970 : forvar5037[(3'h4):(1'h0)])) ?
                          reg5263[(1'h1):(1'h0)] : (8'hab));
                    end
                  reg5484 <= (~|(~^(-(~^reg5083))));
                  if (reg5141)
                    begin
                      reg5485 <= {(~^reg5271[(4'hc):(4'ha)])};
                      reg5486 <= ((8'hb9) >>> ((^~forvar5454) == forvar5448));
                      reg5487 <= (+($unsigned($signed(forvar5489)) ?
                          $signed((reg5358 ^~ reg5124)) : $unsigned((reg5286 == reg5465))));
                      reg5488 <= $unsigned(reg5425);
                    end
                  else
                    begin
                      reg5485 <= (($signed((reg5056 ? forvar5109 : (8'ha9))) ?
                          (reg5455 + forvar5001) : {(reg5237 == reg5366)}) | (reg5169[(2'h3):(2'h2)] ?
                          $unsigned((reg5273 && reg5473)) : ((8'haf) ?
                              (reg4997 ?
                                  reg5456 : (8'hb9)) : reg5204[(2'h3):(1'h1)])));
                      reg5486 <= $signed($unsigned((8'h9c)));
                    end
                  if ($unsigned($unsigned(($unsigned((8'ha7)) ?
                      (reg5486 >>> reg5405) : ((8'ha0) ^ (8'ha5))))))
                    begin
                      reg5489 <= (^~forvar5375[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg5489 <= {$signed($signed(reg5285[(4'h8):(1'h0)]))};
                    end
                end
              if ({($unsigned($signed(forvar5251)) ?
                      (+reg4998) : (((8'hb1) ? reg5232 : reg5189) ?
                          reg5488[(4'h9):(4'h8)] : reg5477))})
                begin
                  if ({(^~{forvar5271[(2'h3):(1'h1)]})})
                    begin
                      reg5490 <= (($unsigned(reg5416[(4'hd):(2'h2)]) ?
                              reg5012[(2'h3):(1'h0)] : ((forvar5011 ~^ forvar5468) >= (forvar5401 & reg5052))) ?
                          $signed({(!(8'hb2))}) : $unsigned($signed((reg5158 ?
                              reg5259 : reg5307))));
                      reg5491 <= (+(+((reg5459 ?
                          (8'ha5) : (8'h9c)) >>> reg5158)));
                      reg5492 <= $unsigned(reg5490[(3'h5):(2'h3)]);
                    end
                  else
                    begin
                      reg5490 <= reg5104;
                    end
                  for (forvar5493 = (1'h0); (forvar5493 < (1'h1)); forvar5493 = (forvar5493 + (1'h1)))
                    begin
                      reg5494 <= reg5464[(3'h5):(1'h0)];
                      reg5495 <= {$signed($signed(reg5310))};
                      reg5496 <= (~|$signed((+reg5038)));
                      reg5497 <= {(&$signed($signed(wire1024)))};
                    end
                end
              else
                begin
                  reg5490 <= reg5482[(4'hd):(3'h6)];
                  for (forvar5491 = (1'h0); (forvar5491 < (2'h2)); forvar5491 = (forvar5491 + (1'h1)))
                    begin
                      reg5492 <= $unsigned($signed(reg5183));
                      reg5493 <= (-forvar5474[(4'h8):(3'h4)]);
                      reg5494 <= $unsigned(($signed(reg5121[(4'hb):(1'h0)]) ?
                          $signed(reg5340[(4'hb):(1'h1)]) : reg5164));
                      reg5495 <= {($signed((forvar5394 <<< reg5463)) >= reg5134[(3'h5):(2'h2)])};
                    end
                  if ({reg5094})
                    begin
                      reg5496 <= reg5462;
                      reg5497 <= {($signed((reg4984 ? (8'ha3) : reg5402)) ?
                              reg5349 : {reg5388})};
                      reg5498 <= $unsigned($signed(($signed(reg5304) ?
                          reg5304[(4'ha):(2'h2)] : $signed(reg5053))));
                      reg5499 <= reg5225;
                    end
                  else
                    begin
                      reg5496 <= (reg5044 - reg5459[(1'h0):(1'h0)]);
                      reg5497 <= (~|forvar5468[(3'h6):(2'h3)]);
                    end
                end
            end
          reg5500 <= $signed((forvar5404[(1'h0):(1'h0)] & forvar5427));
          if (reg5303)
            begin
              if (reg5143[(4'hb):(1'h1)])
                begin
                  if ($signed(((((8'ha6) < reg5275) ?
                      reg5121[(3'h4):(1'h1)] : $signed(reg5125)) << {{reg5010}})))
                    begin
                      reg5501 <= ($signed({(reg5421 ?
                              forvar5175 : reg5182)}) & reg5328[(3'h4):(1'h0)]);
                      reg5502 <= (((~&(^reg5277)) > ($signed((8'hb3)) ?
                          {(8'ha2)} : $signed(reg5491))) ^ $unsigned((|reg4995[(3'h5):(1'h0)])));
                      reg5503 <= (($unsigned((wire1022 > reg5325)) ?
                              ({reg5420} ?
                                  (-reg5408) : (forvar5061 || forvar5227)) : (~&{reg5033})) ?
                          (!reg5211) : reg5017);
                      reg5504 <= ((|(|{reg5044})) ^~ wire3536[(4'h9):(3'h4)]);
                    end
                  else
                    begin
                      reg5501 <= $signed((8'ha0));
                      reg5502 <= (+$unsigned((&(-forvar5484))));
                      reg5503 <= $signed((~$signed((reg5053 - (8'hae)))));
                    end
                  if ($unsigned($unsigned($signed($unsigned(wire3538)))))
                    begin
                      reg5505 <= forvar5089[(1'h1):(1'h1)];
                      reg5506 <= {(&(~|(reg5295 ^~ forvar5088)))};
                      reg5507 <= $signed({forvar5117});
                    end
                  else
                    begin
                      reg5505 <= reg5027;
                      reg5506 <= reg5394[(4'h9):(1'h0)];
                    end
                  for (forvar5508 = (1'h0); (forvar5508 < (1'h0)); forvar5508 = (forvar5508 + (1'h1)))
                    begin
                      reg5509 <= ($unsigned({$unsigned(reg5085)}) && (reg5442 && (&$unsigned(reg5191))));
                      reg5510 <= (reg5494 ?
                          ((((8'hb9) ? reg5091 : (8'had)) ?
                                  reg5459[(1'h1):(1'h0)] : $signed(forvar5419)) ?
                              (8'hb4) : reg5105[(1'h0):(1'h0)]) : (($unsigned(reg5138) ?
                              $signed(reg5109) : {reg5385}) - $unsigned((forvar4986 ^~ reg5482))));
                    end
                  reg5511 <= {$unsigned(($signed(forvar5223) ?
                          (reg5033 || reg5044) : reg4992))};
                end
              else
                begin
                  reg5501 <= $unsigned({reg5294[(1'h1):(1'h0)]});
                  for (forvar5502 = (1'h0); (forvar5502 < (2'h3)); forvar5502 = (forvar5502 + (1'h1)))
                    begin
                      reg5503 <= $unsigned($signed(reg5278));
                      reg5504 <= $signed($unsigned($unsigned({forvar5441})));
                      reg5505 <= reg4975;
                    end
                  for (forvar5506 = (1'h0); (forvar5506 < (1'h0)); forvar5506 = (forvar5506 + (1'h1)))
                    begin
                      reg5507 <= (reg5279 ?
                          $signed((|(reg5498 || (8'hb3)))) : (|$signed({reg5216})));
                    end
                end
              if (reg5470[(2'h2):(1'h1)])
                begin
                  reg5512 <= $unsigned(($signed(((8'hb3) >>> (8'ha1))) && ($signed(forvar5001) ?
                      reg5285 : (8'ha3))));
                end
              else
                begin
                  if ((+(-forvar4983)))
                    begin
                      reg5512 <= $unsigned(forvar5337[(1'h0):(1'h0)]);
                      reg5513 <= $signed(reg5199[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg5512 <= (~|$signed(reg5313));
                      reg5513 <= $signed({forvar5448[(3'h5):(2'h3)]});
                    end
                  if ((+forvar5156))
                    begin
                      reg5514 <= (|reg5112);
                      reg5515 <= forvar5478;
                    end
                  else
                    begin
                      reg5514 <= ($unsigned($unsigned({(8'hac)})) <= reg5247);
                      reg5515 <= ((((reg5482 ^ reg5472) >> wire1030) - reg5471) ?
                          $unsigned(reg5383) : $signed($signed((reg5233 ?
                              forvar5480 : forvar5011))));
                      reg5516 <= (forvar5116 && forvar5418[(2'h2):(1'h0)]);
                      reg5517 <= $signed({reg5272});
                    end
                  for (forvar5518 = (1'h0); (forvar5518 < (2'h2)); forvar5518 = (forvar5518 + (1'h1)))
                    begin
                      reg5519 <= reg5355[(3'h4):(3'h4)];
                      reg5520 <= $unsigned(forvar5070[(1'h1):(1'h1)]);
                    end
                  if (reg5199)
                    begin
                      reg5521 <= (reg5213[(1'h0):(1'h0)] + $unsigned({forvar5410}));
                      reg5522 <= ((reg5406[(2'h3):(1'h1)] ?
                              {(-reg4975)} : $signed($signed(reg5106))) ?
                          $unsigned(forvar5488) : {((forvar5046 ?
                                  reg5264 : (8'ha2)) || $signed(reg5340))});
                      reg5523 <= ((|reg5421) ? reg5432 : $signed(reg5094));
                    end
                  else
                    begin
                      reg5521 <= forvar5109;
                    end
                end
            end
          else
            begin
              for (forvar5501 = (1'h0); (forvar5501 < (2'h3)); forvar5501 = (forvar5501 + (1'h1)))
                begin
                  if ((reg5346[(4'ha):(3'h7)] || (forvar5070 ~^ $signed((&reg5187)))))
                    begin
                      reg5502 <= $signed((((^~(8'h9d)) >> $unsigned(reg5068)) == $signed(forvar5046)));
                      reg5503 <= $unsigned((8'ha0));
                      reg5504 <= $signed(reg5178);
                      reg5505 <= reg5107;
                    end
                  else
                    begin
                      reg5502 <= (~&(&$signed(((8'ha4) ? reg5395 : (8'ha6)))));
                    end
                end
              reg5506 <= $signed(forvar5414);
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3539
#( parameter param4966 = (+((((8'hac) ? (8'ha3) : (8'h9e)) ? ((8'ha4) ~^ (8'h9e)) : (&(8'hb2))) + (~|((8'ha3) ? (8'ha5) : (8'ha8))))) )
(y, clk, wire3543, wire3542, wire3541, wire3540);
  output wire [(32'h1295):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire3543;
  input wire [(2'h3):(1'h0)] wire3542;
  input wire signed [(4'he):(1'h0)] wire3541;
  input wire [(4'h8):(1'h0)] wire3540;
  wire [(4'h9):(1'h0)] wire4965;
  wire signed [(3'h6):(1'h0)] wire4964;
  reg signed [(4'hc):(1'h0)] forvar4891 = (1'h0);
  reg [(3'h6):(1'h0)] reg4879 = (1'h0);
  reg [(3'h6):(1'h0)] reg4878 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4906 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4901 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4902 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4892 = (1'h0);
  reg [(3'h4):(1'h0)] reg4899 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4897 = (1'h0);
  reg [(4'h8):(1'h0)] reg4896 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4895 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4894 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4890 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4963 = (1'h0);
  reg [(2'h3):(1'h0)] reg4962 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4961 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4960 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4959 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4958 = (1'h0);
  reg [(2'h3):(1'h0)] reg4957 = (1'h0);
  reg [(4'hd):(1'h0)] reg4956 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4955 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4954 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4953 = (1'h0);
  reg [(4'h8):(1'h0)] reg4952 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4951 = (1'h0);
  reg [(4'h8):(1'h0)] reg4950 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4949 = (1'h0);
  reg [(4'h8):(1'h0)] reg4948 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4947 = (1'h0);
  reg [(4'ha):(1'h0)] reg4946 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4945 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4944 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4943 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4942 = (1'h0);
  reg [(4'h8):(1'h0)] reg4941 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4940 = (1'h0);
  reg [(4'ha):(1'h0)] reg4939 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4938 = (1'h0);
  reg [(3'h7):(1'h0)] reg4937 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4936 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4935 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4934 = (1'h0);
  reg [(4'hf):(1'h0)] reg4928 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4927 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4926 = (1'h0);
  reg [(2'h2):(1'h0)] reg4925 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4933 = (1'h0);
  reg [(4'hf):(1'h0)] reg4932 = (1'h0);
  reg [(4'hc):(1'h0)] reg4931 = (1'h0);
  reg [(4'hf):(1'h0)] reg4930 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4929 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4928 = (1'h0);
  reg [(3'h5):(1'h0)] reg4927 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4926 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4925 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4924 = (1'h0);
  reg [(2'h2):(1'h0)] reg4923 = (1'h0);
  reg [(3'h5):(1'h0)] reg4922 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4921 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4920 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4919 = (1'h0);
  reg [(4'hd):(1'h0)] reg4918 = (1'h0);
  reg [(3'h7):(1'h0)] reg4917 = (1'h0);
  reg [(4'ha):(1'h0)] reg4916 = (1'h0);
  reg [(4'hb):(1'h0)] reg4915 = (1'h0);
  reg [(2'h3):(1'h0)] reg4914 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4911 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4907 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4904 = (1'h0);
  reg [(4'h9):(1'h0)] reg4900 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4898 = (1'h0);
  reg [(5'h10):(1'h0)] reg4913 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4912 = (1'h0);
  reg [(4'he):(1'h0)] reg4911 = (1'h0);
  reg [(4'hd):(1'h0)] reg4910 = (1'h0);
  reg [(4'h8):(1'h0)] reg4909 = (1'h0);
  reg [(3'h5):(1'h0)] reg4908 = (1'h0);
  reg [(4'h9):(1'h0)] reg4907 = (1'h0);
  reg [(3'h4):(1'h0)] reg4906 = (1'h0);
  reg [(3'h4):(1'h0)] reg4905 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4904 = (1'h0);
  reg [(3'h5):(1'h0)] reg4903 = (1'h0);
  reg [(4'ha):(1'h0)] reg4902 = (1'h0);
  reg [(3'h6):(1'h0)] reg4901 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4900 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4899 = (1'h0);
  reg [(4'h9):(1'h0)] reg4898 = (1'h0);
  reg [(3'h7):(1'h0)] reg4897 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4896 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4895 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4894 = (1'h0);
  reg [(4'hd):(1'h0)] reg4893 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4892 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4891 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4889 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4888 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4886 = (1'h0);
  reg [(4'h9):(1'h0)] reg4890 = (1'h0);
  reg [(4'hf):(1'h0)] reg4889 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4888 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4887 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4886 = (1'h0);
  reg [(3'h5):(1'h0)] reg4885 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4884 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4883 = (1'h0);
  reg [(2'h3):(1'h0)] reg4882 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4881 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4880 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4879 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4878 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4877 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4876 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4875 = (1'h0);
  reg [(4'hf):(1'h0)] reg4874 = (1'h0);
  reg [(2'h2):(1'h0)] reg4873 = (1'h0);
  reg [(2'h2):(1'h0)] reg4872 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4868 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4867 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4871 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4870 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4869 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4868 = (1'h0);
  reg [(3'h6):(1'h0)] reg4867 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4866 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4865 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire4864;
  reg [(4'ha):(1'h0)] reg4863 = (1'h0);
  reg [(4'hf):(1'h0)] reg4862 = (1'h0);
  reg [(4'hb):(1'h0)] reg4861 = (1'h0);
  reg [(4'ha):(1'h0)] reg4860 = (1'h0);
  reg [(4'ha):(1'h0)] reg4859 = (1'h0);
  reg [(4'hc):(1'h0)] reg4858 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4857 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4856 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4855 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4854 = (1'h0);
  reg [(3'h5):(1'h0)] reg4853 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4852 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4851 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4850 = (1'h0);
  reg [(5'h10):(1'h0)] reg4850 = (1'h0);
  reg [(3'h6):(1'h0)] reg4849 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4848 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4839 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4830 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4824 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4823 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4819 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4814 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4813 = (1'h0);
  reg [(2'h3):(1'h0)] reg4810 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4808 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4802 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4798 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4803 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4801 = (1'h0);
  reg [(3'h7):(1'h0)] reg4797 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4796 = (1'h0);
  reg [(4'h8):(1'h0)] reg4834 = (1'h0);
  reg [(5'h10):(1'h0)] reg4829 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4826 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4825 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4822 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4843 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4842 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4847 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4846 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4845 = (1'h0);
  reg [(4'hc):(1'h0)] reg4844 = (1'h0);
  reg [(4'h9):(1'h0)] reg4843 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4842 = (1'h0);
  reg [(4'ha):(1'h0)] reg4841 = (1'h0);
  reg [(5'h10):(1'h0)] reg4840 = (1'h0);
  reg [(4'hf):(1'h0)] reg4839 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4838 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4837 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4836 = (1'h0);
  reg [(3'h7):(1'h0)] reg4835 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4834 = (1'h0);
  reg [(4'h8):(1'h0)] reg4833 = (1'h0);
  reg [(4'hb):(1'h0)] reg4832 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4831 = (1'h0);
  reg [(3'h7):(1'h0)] reg4830 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4829 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4828 = (1'h0);
  reg [(2'h3):(1'h0)] reg4827 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4826 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4825 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4824 = (1'h0);
  reg [(4'h8):(1'h0)] reg4823 = (1'h0);
  reg [(4'hb):(1'h0)] reg4822 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4821 = (1'h0);
  reg [(4'hd):(1'h0)] reg4820 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4819 = (1'h0);
  reg [(4'hb):(1'h0)] reg4818 = (1'h0);
  reg [(4'h9):(1'h0)] reg4817 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4816 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4815 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4814 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4813 = (1'h0);
  reg [(4'h8):(1'h0)] reg4812 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4811 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4810 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4809 = (1'h0);
  reg [(3'h7):(1'h0)] reg4808 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4807 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4806 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4805 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4804 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4803 = (1'h0);
  reg [(4'ha):(1'h0)] reg4802 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4801 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4800 = (1'h0);
  reg [(4'hb):(1'h0)] reg4799 = (1'h0);
  reg [(4'ha):(1'h0)] reg4798 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4797 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4796 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4795 = (1'h0);
  wire [(3'h4):(1'h0)] wire4794;
  wire signed [(4'hb):(1'h0)] wire4793;
  reg [(3'h4):(1'h0)] reg4792 = (1'h0);
  reg [(4'ha):(1'h0)] reg4791 = (1'h0);
  reg [(3'h5):(1'h0)] reg4790 = (1'h0);
  reg [(4'ha):(1'h0)] reg4789 = (1'h0);
  reg [(4'hd):(1'h0)] reg4788 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4787 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4786 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4785 = (1'h0);
  reg [(3'h6):(1'h0)] reg4784 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4783 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4782 = (1'h0);
  reg [(2'h2):(1'h0)] reg4781 = (1'h0);
  reg [(5'h10):(1'h0)] reg4780 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4779 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4777 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4773 = (1'h0);
  reg [(3'h6):(1'h0)] reg4764 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4763 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4761 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4760 = (1'h0);
  reg [(4'ha):(1'h0)] reg4758 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4752 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4750 = (1'h0);
  reg [(4'ha):(1'h0)] reg4746 = (1'h0);
  reg [(3'h4):(1'h0)] reg4745 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4743 = (1'h0);
  reg [(4'hb):(1'h0)] reg4738 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4736 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4778 = (1'h0);
  reg [(4'hc):(1'h0)] reg4777 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4776 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4775 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4774 = (1'h0);
  reg [(4'he):(1'h0)] reg4773 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4772 = (1'h0);
  reg [(2'h3):(1'h0)] reg4771 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4770 = (1'h0);
  reg [(4'hd):(1'h0)] reg4769 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4768 = (1'h0);
  reg [(3'h6):(1'h0)] reg4767 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4766 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4765 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4764 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4763 = (1'h0);
  reg [(2'h2):(1'h0)] reg4762 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4761 = (1'h0);
  reg [(4'h8):(1'h0)] reg4760 = (1'h0);
  reg [(4'hf):(1'h0)] reg4759 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4758 = (1'h0);
  reg [(3'h7):(1'h0)] reg4757 = (1'h0);
  reg [(3'h4):(1'h0)] reg4756 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4755 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4754 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4753 = (1'h0);
  reg [(4'h9):(1'h0)] reg4749 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4752 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4751 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4750 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4749 = (1'h0);
  reg [(4'hb):(1'h0)] reg4748 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4747 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4746 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4745 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4744 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4743 = (1'h0);
  reg [(3'h5):(1'h0)] reg4742 = (1'h0);
  reg [(4'hb):(1'h0)] reg4741 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4740 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4739 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4738 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4737 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4736 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4735 = (1'h0);
  reg [(3'h5):(1'h0)] reg4734 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire4733;
  wire signed [(3'h7):(1'h0)] wire4732;
  wire signed [(4'hc):(1'h0)] wire4730;
  wire signed [(4'hc):(1'h0)] wire3768;
  wire signed [(4'hd):(1'h0)] wire3767;
  wire [(4'hb):(1'h0)] wire3766;
  reg signed [(4'h9):(1'h0)] reg3765 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3764 = (1'h0);
  reg [(3'h4):(1'h0)] reg3763 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3762 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3761 = (1'h0);
  reg [(2'h3):(1'h0)] reg3760 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3759 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3758 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3757 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3756 = (1'h0);
  reg [(2'h3):(1'h0)] reg3755 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3754 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3753 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3752 = (1'h0);
  reg [(5'h10):(1'h0)] reg3751 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3750 = (1'h0);
  reg [(3'h6):(1'h0)] reg3749 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3748 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3747 = (1'h0);
  reg [(2'h3):(1'h0)] reg3746 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3745 = (1'h0);
  reg [(4'hf):(1'h0)] reg3744 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3742 = (1'h0);
  reg [(4'he):(1'h0)] reg3740 = (1'h0);
  reg [(5'h10):(1'h0)] reg3743 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3742 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3741 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3740 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3739 = (1'h0);
  reg [(3'h5):(1'h0)] reg3734 = (1'h0);
  reg [(3'h5):(1'h0)] reg3738 = (1'h0);
  reg [(4'hb):(1'h0)] reg3737 = (1'h0);
  reg [(2'h3):(1'h0)] reg3736 = (1'h0);
  reg [(2'h3):(1'h0)] reg3735 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3734 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3733 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3732 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3731 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3730 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3729 = (1'h0);
  reg [(3'h5):(1'h0)] reg3728 = (1'h0);
  reg [(4'he):(1'h0)] reg3727 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3726 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3725 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3724 = (1'h0);
  reg [(3'h4):(1'h0)] reg3723 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3722 = (1'h0);
  reg [(4'hf):(1'h0)] reg3721 = (1'h0);
  reg [(2'h3):(1'h0)] reg3720 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3719 = (1'h0);
  reg [(2'h2):(1'h0)] reg3718 = (1'h0);
  reg [(4'he):(1'h0)] forvar3717 = (1'h0);
  reg [(4'hf):(1'h0)] reg3716 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3715 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3714 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3713 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3712 = (1'h0);
  reg [(4'he):(1'h0)] forvar3711 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3710 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3709 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3708 = (1'h0);
  reg [(2'h3):(1'h0)] reg3707 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3706 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3705 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3704 = (1'h0);
  reg [(3'h5):(1'h0)] reg3703 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3702 = (1'h0);
  reg [(4'ha):(1'h0)] reg3701 = (1'h0);
  reg [(3'h4):(1'h0)] reg3700 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3699 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3698 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3697 = (1'h0);
  reg [(3'h7):(1'h0)] reg3696 = (1'h0);
  reg [(3'h7):(1'h0)] reg3695 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3694 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3693 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3692 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3691 = (1'h0);
  reg [(4'hb):(1'h0)] reg3690 = (1'h0);
  reg [(4'h9):(1'h0)] reg3689 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3688 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3687 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3686 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3685 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3684 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3683 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3682 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3681 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3676 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3672 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3671 = (1'h0);
  reg [(4'h8):(1'h0)] reg3669 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3660 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3657 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3656 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3655 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3654 = (1'h0);
  reg [(2'h2):(1'h0)] reg3652 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3646 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3645 = (1'h0);
  reg [(4'hc):(1'h0)] reg3680 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3679 = (1'h0);
  reg [(3'h4):(1'h0)] reg3678 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3677 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3676 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3675 = (1'h0);
  reg [(2'h3):(1'h0)] reg3674 = (1'h0);
  reg [(3'h5):(1'h0)] reg3673 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3672 = (1'h0);
  reg [(5'h10):(1'h0)] reg3671 = (1'h0);
  reg [(3'h5):(1'h0)] reg3670 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3669 = (1'h0);
  reg [(4'h8):(1'h0)] reg3668 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3667 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3666 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3665 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3664 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3663 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3662 = (1'h0);
  reg [(4'h9):(1'h0)] reg3661 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3660 = (1'h0);
  reg [(4'h8):(1'h0)] reg3659 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3658 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3657 = (1'h0);
  reg [(4'h9):(1'h0)] reg3656 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3655 = (1'h0);
  reg [(4'hb):(1'h0)] reg3654 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3653 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3652 = (1'h0);
  reg [(2'h3):(1'h0)] reg3651 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3650 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3649 = (1'h0);
  reg [(3'h5):(1'h0)] reg3648 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3647 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3646 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3645 = (1'h0);
  reg [(3'h5):(1'h0)] reg3644 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3643 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3642 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3641 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3640 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3639 = (1'h0);
  reg [(4'hc):(1'h0)] reg3638 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3637 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3636 = (1'h0);
  reg [(4'hc):(1'h0)] reg3635 = (1'h0);
  reg [(4'hc):(1'h0)] reg3634 = (1'h0);
  reg [(3'h6):(1'h0)] reg3633 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3632 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3631 = (1'h0);
  reg [(3'h5):(1'h0)] reg3630 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3628 = (1'h0);
  reg [(3'h5):(1'h0)] reg3627 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3626 = (1'h0);
  reg [(5'h10):(1'h0)] reg3625 = (1'h0);
  reg [(3'h4):(1'h0)] reg3624 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3623 = (1'h0);
  reg [(4'ha):(1'h0)] reg3622 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3619 = (1'h0);
  reg [(4'he):(1'h0)] reg3621 = (1'h0);
  reg [(5'h10):(1'h0)] reg3620 = (1'h0);
  reg [(3'h4):(1'h0)] reg3619 = (1'h0);
  reg [(3'h6):(1'h0)] reg3615 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3618 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3617 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3616 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3615 = (1'h0);
  reg [(4'ha):(1'h0)] reg3614 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3613 = (1'h0);
  reg [(5'h10):(1'h0)] reg3612 = (1'h0);
  reg [(4'ha):(1'h0)] reg3611 = (1'h0);
  reg [(2'h3):(1'h0)] reg3610 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3609 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3608 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3607 = (1'h0);
  reg [(4'hb):(1'h0)] reg3606 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3605 = (1'h0);
  reg [(4'ha):(1'h0)] reg3604 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3603 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3602 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3601 = (1'h0);
  reg [(4'ha):(1'h0)] reg3593 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3600 = (1'h0);
  reg [(3'h7):(1'h0)] reg3599 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3598 = (1'h0);
  reg [(4'hd):(1'h0)] reg3597 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3596 = (1'h0);
  reg [(4'h9):(1'h0)] reg3595 = (1'h0);
  reg [(4'he):(1'h0)] reg3594 = (1'h0);
  reg [(4'he):(1'h0)] forvar3593 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3592 = (1'h0);
  reg [(4'h9):(1'h0)] reg3591 = (1'h0);
  reg [(4'hb):(1'h0)] reg3590 = (1'h0);
  reg [(4'he):(1'h0)] forvar3589 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3588 = (1'h0);
  reg [(4'hf):(1'h0)] reg3587 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3586 = (1'h0);
  reg [(4'he):(1'h0)] reg3585 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3584 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3583 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3582 = (1'h0);
  reg [(3'h6):(1'h0)] reg3581 = (1'h0);
  reg [(4'hb):(1'h0)] reg3580 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3579 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3578 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3577 = (1'h0);
  reg [(5'h10):(1'h0)] reg3576 = (1'h0);
  reg [(4'h9):(1'h0)] reg3575 = (1'h0);
  reg [(4'ha):(1'h0)] reg3574 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3573 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3572 = (1'h0);
  reg [(3'h4):(1'h0)] reg3571 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3570 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3569 = (1'h0);
  reg [(4'hc):(1'h0)] reg3568 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3567 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3566 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3565 = (1'h0);
  reg [(3'h4):(1'h0)] reg3564 = (1'h0);
  reg [(5'h10):(1'h0)] reg3563 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3562 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3561 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3560 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3559 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3558 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3552 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3545 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3553 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3549 = (1'h0);
  reg [(5'h10):(1'h0)] reg3548 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3547 = (1'h0);
  reg [(4'h8):(1'h0)] reg3559 = (1'h0);
  reg [(3'h5):(1'h0)] reg3544 = (1'h0);
  reg [(4'hf):(1'h0)] reg3558 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3557 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3556 = (1'h0);
  reg [(4'hb):(1'h0)] reg3555 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3554 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3553 = (1'h0);
  reg [(3'h6):(1'h0)] reg3552 = (1'h0);
  reg [(5'h10):(1'h0)] reg3551 = (1'h0);
  reg [(4'hc):(1'h0)] reg3550 = (1'h0);
  reg [(3'h7):(1'h0)] reg3549 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3548 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3547 = (1'h0);
  reg [(4'hd):(1'h0)] reg3546 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3545 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3544 = (1'h0);
  assign y = {wire4965,
                 wire4964,
                 forvar4891,
                 reg4879,
                 reg4878,
                 forvar4906,
                 forvar4901,
                 forvar4902,
                 forvar4892,
                 reg4899,
                 forvar4897,
                 reg4896,
                 reg4895,
                 forvar4894,
                 forvar4890,
                 reg4963,
                 reg4962,
                 reg4961,
                 reg4960,
                 forvar4959,
                 reg4958,
                 reg4957,
                 reg4956,
                 reg4955,
                 forvar4954,
                 reg4953,
                 reg4952,
                 reg4951,
                 reg4950,
                 forvar4949,
                 reg4948,
                 reg4947,
                 reg4946,
                 reg4945,
                 forvar4944,
                 reg4943,
                 reg4942,
                 reg4941,
                 forvar4940,
                 reg4939,
                 reg4938,
                 reg4937,
                 reg4936,
                 forvar4935,
                 forvar4934,
                 reg4928,
                 forvar4927,
                 forvar4926,
                 reg4925,
                 reg4933,
                 reg4932,
                 reg4931,
                 reg4930,
                 reg4929,
                 forvar4928,
                 reg4927,
                 reg4926,
                 forvar4925,
                 reg4924,
                 reg4923,
                 reg4922,
                 forvar4921,
                 forvar4920,
                 reg4919,
                 reg4918,
                 reg4917,
                 reg4916,
                 reg4915,
                 reg4914,
                 forvar4911,
                 forvar4907,
                 reg4904,
                 reg4900,
                 forvar4898,
                 reg4913,
                 reg4912,
                 reg4911,
                 reg4910,
                 reg4909,
                 reg4908,
                 reg4907,
                 reg4906,
                 reg4905,
                 forvar4904,
                 reg4903,
                 reg4902,
                 reg4901,
                 forvar4900,
                 forvar4899,
                 reg4898,
                 reg4897,
                 forvar4896,
                 forvar4895,
                 reg4894,
                 reg4893,
                 reg4892,
                 reg4891,
                 forvar4889,
                 forvar4888,
                 reg4886,
                 reg4890,
                 reg4889,
                 reg4888,
                 reg4887,
                 forvar4886,
                 reg4885,
                 reg4884,
                 reg4883,
                 reg4882,
                 reg4881,
                 reg4880,
                 forvar4879,
                 forvar4878,
                 reg4877,
                 reg4876,
                 reg4875,
                 reg4874,
                 reg4873,
                 reg4872,
                 reg4868,
                 forvar4867,
                 reg4871,
                 reg4870,
                 reg4869,
                 forvar4868,
                 reg4867,
                 forvar4866,
                 forvar4865,
                 wire4864,
                 reg4863,
                 reg4862,
                 reg4861,
                 reg4860,
                 reg4859,
                 reg4858,
                 reg4857,
                 reg4856,
                 forvar4855,
                 reg4854,
                 reg4853,
                 forvar4852,
                 reg4851,
                 forvar4850,
                 reg4850,
                 reg4849,
                 forvar4848,
                 forvar4839,
                 forvar4830,
                 forvar4824,
                 forvar4823,
                 forvar4819,
                 reg4814,
                 forvar4813,
                 reg4810,
                 forvar4808,
                 forvar4802,
                 forvar4798,
                 reg4803,
                 forvar4801,
                 reg4797,
                 forvar4796,
                 reg4834,
                 reg4829,
                 forvar4826,
                 forvar4825,
                 forvar4822,
                 forvar4843,
                 reg4842,
                 reg4847,
                 reg4846,
                 reg4845,
                 reg4844,
                 reg4843,
                 forvar4842,
                 reg4841,
                 reg4840,
                 reg4839,
                 reg4838,
                 reg4837,
                 reg4836,
                 reg4835,
                 forvar4834,
                 reg4833,
                 reg4832,
                 reg4831,
                 reg4830,
                 forvar4829,
                 reg4828,
                 reg4827,
                 reg4826,
                 reg4825,
                 reg4824,
                 reg4823,
                 reg4822,
                 reg4821,
                 reg4820,
                 reg4819,
                 reg4818,
                 reg4817,
                 reg4816,
                 forvar4815,
                 forvar4814,
                 reg4813,
                 reg4812,
                 reg4811,
                 forvar4810,
                 forvar4809,
                 reg4808,
                 reg4807,
                 reg4806,
                 reg4805,
                 reg4804,
                 forvar4803,
                 reg4802,
                 reg4801,
                 reg4800,
                 reg4799,
                 reg4798,
                 forvar4797,
                 reg4796,
                 forvar4795,
                 wire4794,
                 wire4793,
                 reg4792,
                 reg4791,
                 reg4790,
                 reg4789,
                 reg4788,
                 reg4787,
                 reg4786,
                 reg4785,
                 reg4784,
                 forvar4783,
                 forvar4782,
                 reg4781,
                 reg4780,
                 reg4779,
                 forvar4777,
                 forvar4773,
                 reg4764,
                 reg4763,
                 reg4761,
                 forvar4760,
                 reg4758,
                 forvar4752,
                 forvar4750,
                 reg4746,
                 reg4745,
                 reg4743,
                 reg4738,
                 reg4736,
                 reg4778,
                 reg4777,
                 reg4776,
                 reg4775,
                 reg4774,
                 reg4773,
                 reg4772,
                 reg4771,
                 forvar4770,
                 reg4769,
                 reg4768,
                 reg4767,
                 reg4766,
                 forvar4765,
                 forvar4764,
                 forvar4763,
                 reg4762,
                 forvar4761,
                 reg4760,
                 reg4759,
                 forvar4758,
                 reg4757,
                 reg4756,
                 reg4755,
                 reg4754,
                 forvar4753,
                 reg4749,
                 reg4752,
                 reg4751,
                 reg4750,
                 forvar4749,
                 reg4748,
                 reg4747,
                 forvar4746,
                 forvar4745,
                 reg4744,
                 forvar4743,
                 reg4742,
                 reg4741,
                 reg4740,
                 reg4739,
                 forvar4738,
                 reg4737,
                 forvar4736,
                 forvar4735,
                 reg4734,
                 wire4733,
                 wire4732,
                 wire4730,
                 wire3768,
                 wire3767,
                 wire3766,
                 reg3765,
                 reg3764,
                 reg3763,
                 reg3762,
                 reg3761,
                 reg3760,
                 reg3759,
                 reg3758,
                 reg3757,
                 reg3756,
                 reg3755,
                 forvar3754,
                 forvar3753,
                 reg3752,
                 reg3751,
                 reg3750,
                 reg3749,
                 forvar3748,
                 reg3747,
                 reg3746,
                 forvar3745,
                 reg3744,
                 forvar3742,
                 reg3740,
                 reg3743,
                 reg3742,
                 reg3741,
                 forvar3740,
                 forvar3739,
                 reg3734,
                 reg3738,
                 reg3737,
                 reg3736,
                 reg3735,
                 forvar3734,
                 reg3733,
                 reg3732,
                 reg3731,
                 reg3730,
                 reg3729,
                 reg3728,
                 reg3727,
                 reg3726,
                 forvar3725,
                 reg3724,
                 reg3723,
                 forvar3722,
                 reg3721,
                 reg3720,
                 forvar3719,
                 reg3718,
                 forvar3717,
                 reg3716,
                 forvar3715,
                 reg3714,
                 reg3713,
                 reg3712,
                 forvar3711,
                 forvar3710,
                 reg3709,
                 reg3708,
                 reg3707,
                 forvar3706,
                 reg3705,
                 reg3704,
                 reg3703,
                 forvar3702,
                 reg3701,
                 reg3700,
                 forvar3699,
                 forvar3698,
                 forvar3697,
                 reg3696,
                 reg3695,
                 reg3694,
                 reg3693,
                 reg3692,
                 reg3691,
                 reg3690,
                 reg3689,
                 reg3688,
                 reg3687,
                 forvar3686,
                 reg3685,
                 reg3684,
                 reg3683,
                 forvar3682,
                 forvar3681,
                 reg3676,
                 forvar3672,
                 forvar3671,
                 reg3669,
                 reg3660,
                 reg3657,
                 forvar3656,
                 reg3655,
                 forvar3654,
                 reg3652,
                 reg3646,
                 forvar3645,
                 reg3680,
                 reg3679,
                 reg3678,
                 reg3677,
                 forvar3676,
                 reg3675,
                 reg3674,
                 reg3673,
                 reg3672,
                 reg3671,
                 reg3670,
                 forvar3669,
                 reg3668,
                 reg3667,
                 reg3666,
                 reg3665,
                 forvar3664,
                 reg3663,
                 reg3662,
                 reg3661,
                 forvar3660,
                 reg3659,
                 reg3658,
                 forvar3657,
                 reg3656,
                 forvar3655,
                 reg3654,
                 reg3653,
                 forvar3652,
                 reg3651,
                 reg3650,
                 reg3649,
                 reg3648,
                 forvar3647,
                 forvar3646,
                 reg3645,
                 reg3644,
                 reg3643,
                 reg3642,
                 forvar3641,
                 reg3640,
                 reg3639,
                 reg3638,
                 reg3637,
                 forvar3636,
                 reg3635,
                 reg3634,
                 reg3633,
                 reg3632,
                 forvar3631,
                 reg3630,
                 reg3629,
                 reg3628,
                 reg3627,
                 forvar3626,
                 reg3625,
                 reg3624,
                 forvar3623,
                 reg3622,
                 forvar3619,
                 reg3621,
                 reg3620,
                 reg3619,
                 reg3615,
                 reg3618,
                 reg3617,
                 reg3616,
                 forvar3615,
                 reg3614,
                 forvar3613,
                 reg3612,
                 reg3611,
                 reg3610,
                 forvar3609,
                 reg3608,
                 forvar3607,
                 reg3606,
                 reg3605,
                 reg3604,
                 reg3603,
                 forvar3602,
                 forvar3601,
                 reg3593,
                 reg3600,
                 reg3599,
                 forvar3598,
                 reg3597,
                 reg3596,
                 reg3595,
                 reg3594,
                 forvar3593,
                 reg3592,
                 reg3591,
                 reg3590,
                 forvar3589,
                 reg3588,
                 reg3587,
                 reg3586,
                 reg3585,
                 reg3584,
                 reg3583,
                 reg3582,
                 reg3581,
                 reg3580,
                 forvar3579,
                 forvar3578,
                 forvar3577,
                 reg3576,
                 reg3575,
                 reg3574,
                 forvar3573,
                 reg3572,
                 reg3571,
                 reg3570,
                 reg3569,
                 reg3568,
                 forvar3567,
                 forvar3566,
                 reg3565,
                 reg3564,
                 reg3563,
                 reg3562,
                 reg3561,
                 forvar3560,
                 forvar3559,
                 forvar3558,
                 forvar3552,
                 forvar3545,
                 reg3553,
                 forvar3549,
                 reg3548,
                 forvar3547,
                 reg3559,
                 reg3544,
                 reg3558,
                 reg3557,
                 reg3556,
                 reg3555,
                 reg3554,
                 forvar3553,
                 reg3552,
                 reg3551,
                 reg3550,
                 reg3549,
                 forvar3548,
                 reg3547,
                 reg3546,
                 reg3545,
                 forvar3544,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned((~|$signed($signed(wire3541)))))
        begin
          if ((8'ha5))
            begin
              if ($unsigned((wire3540 == wire3542[(1'h1):(1'h1)])))
                begin
                  for (forvar3544 = (1'h0); (forvar3544 < (2'h2)); forvar3544 = (forvar3544 + (1'h1)))
                    begin
                      reg3545 <= $signed(wire3542[(1'h0):(1'h0)]);
                      reg3546 <= ({forvar3544} ?
                          (($unsigned(wire3541) ?
                              wire3543[(2'h2):(2'h2)] : $unsigned(wire3541)) * wire3542) : $signed($unsigned({reg3545})));
                      reg3547 <= ($signed((reg3545[(2'h3):(2'h3)] >= (wire3540 ~^ reg3546))) - ($unsigned({reg3546}) ?
                          $signed($unsigned(reg3545)) : wire3543[(4'h8):(3'h5)]));
                    end
                  for (forvar3548 = (1'h0); (forvar3548 < (2'h2)); forvar3548 = (forvar3548 + (1'h1)))
                    begin
                      reg3549 <= reg3547;
                      reg3550 <= wire3541;
                      reg3551 <= $signed($signed(((reg3549 ?
                              reg3550 : reg3546) ?
                          (reg3545 | reg3550) : $unsigned(reg3546))));
                      reg3552 <= $unsigned(forvar3544[(2'h2):(1'h1)]);
                    end
                  for (forvar3553 = (1'h0); (forvar3553 < (2'h2)); forvar3553 = (forvar3553 + (1'h1)))
                    begin
                      reg3554 <= (-reg3546);
                      reg3555 <= reg3552;
                      reg3556 <= forvar3544;
                      reg3557 <= (reg3551 & (~&reg3545[(4'ha):(3'h6)]));
                    end
                  reg3558 <= {(8'ha4)};
                end
              else
                begin
                  if ($signed(wire3540))
                    begin
                      reg3544 <= ($unsigned((~&((8'h9f) != reg3552))) ?
                          ({reg3555[(4'hb):(3'h7)]} ?
                              $signed((~&reg3557)) : ((reg3549 ?
                                      reg3550 : forvar3548) ?
                                  reg3556[(4'ha):(4'h9)] : (forvar3553 <= reg3557))) : reg3556);
                      reg3545 <= (|(|$unsigned((reg3551 << forvar3544))));
                    end
                  else
                    begin
                      reg3544 <= (~^wire3541);
                      reg3545 <= reg3551;
                    end
                end
              reg3559 <= (&reg3555);
            end
          else
            begin
              for (forvar3544 = (1'h0); (forvar3544 < (1'h1)); forvar3544 = (forvar3544 + (1'h1)))
                begin
                  if ($signed(forvar3548))
                    begin
                      reg3545 <= (~{((8'ha6) ?
                              forvar3553 : (forvar3548 ? reg3546 : reg3549))});
                      reg3546 <= ((+(~&{(8'hb8)})) ?
                          reg3558[(3'h6):(1'h1)] : $unsigned(($signed(reg3550) ?
                              {reg3557} : reg3545[(4'hf):(2'h2)])));
                    end
                  else
                    begin
                      reg3545 <= ({(~(|reg3552))} <= $signed(wire3542));
                    end
                end
              for (forvar3547 = (1'h0); (forvar3547 < (2'h3)); forvar3547 = (forvar3547 + (1'h1)))
                begin
                  reg3548 <= reg3557;
                  for (forvar3549 = (1'h0); (forvar3549 < (1'h0)); forvar3549 = (forvar3549 + (1'h1)))
                    begin
                      reg3550 <= ((~reg3558[(3'h6):(1'h1)]) ?
                          $unsigned($signed((wire3542 & reg3557))) : (&reg3547));
                      reg3551 <= {reg3550[(3'h6):(3'h5)]};
                      reg3552 <= $signed((~$signed(wire3542)));
                      reg3553 <= reg3548;
                    end
                end
            end
        end
      else
        begin
          for (forvar3544 = (1'h0); (forvar3544 < (1'h1)); forvar3544 = (forvar3544 + (1'h1)))
            begin
              if ((reg3545 ?
                  $signed({(reg3546 ?
                          (8'hb7) : reg3552)}) : (+reg3559[(2'h3):(1'h0)])))
                begin
                  for (forvar3545 = (1'h0); (forvar3545 < (1'h0)); forvar3545 = (forvar3545 + (1'h1)))
                    begin
                      reg3546 <= (($unsigned(((8'hac) - forvar3553)) >>> $unsigned($unsigned(forvar3545))) ?
                          wire3543 : (^reg3554[(4'h9):(3'h7)]));
                      reg3547 <= ($unsigned((~|{wire3541})) ?
                          reg3554[(2'h3):(1'h0)] : forvar3544);
                    end
                  if ($signed(reg3548[(4'hb):(2'h3)]))
                    begin
                      reg3548 <= $signed(((reg3547[(4'hc):(4'h8)] * $unsigned(reg3554)) ?
                          (+reg3551) : reg3544[(1'h0):(1'h0)]));
                      reg3549 <= wire3543[(4'he):(3'h5)];
                      reg3550 <= (wire3543 ?
                          $signed((reg3554[(4'hb):(2'h2)] ?
                              {wire3540} : (wire3540 & forvar3547))) : forvar3548);
                    end
                  else
                    begin
                      reg3548 <= reg3555;
                      reg3549 <= (|{forvar3553});
                      reg3550 <= $unsigned($signed(({reg3559} > $unsigned(reg3552))));
                      reg3551 <= reg3549;
                    end
                  for (forvar3552 = (1'h0); (forvar3552 < (2'h2)); forvar3552 = (forvar3552 + (1'h1)))
                    begin
                      reg3553 <= $unsigned({{(wire3543 ?
                                  reg3550 : forvar3544)}});
                    end
                end
              else
                begin
                  for (forvar3545 = (1'h0); (forvar3545 < (2'h3)); forvar3545 = (forvar3545 + (1'h1)))
                    begin
                      reg3546 <= $signed((+$signed({reg3559})));
                      reg3547 <= ((8'had) <<< {reg3545});
                      reg3548 <= forvar3552[(1'h0):(1'h0)];
                      reg3549 <= {$signed(forvar3553[(1'h1):(1'h0)])};
                    end
                  if ((+(forvar3552 == (~(reg3552 ? reg3549 : wire3541)))))
                    begin
                      reg3550 <= reg3550[(3'h6):(1'h1)];
                      reg3551 <= ($unsigned($signed($unsigned(forvar3549))) ?
                          reg3548[(4'he):(2'h3)] : ($signed(forvar3552[(3'h6):(3'h6)]) ?
                              {forvar3547[(4'hd):(4'ha)]} : ((|reg3555) ?
                                  $signed(reg3546) : $unsigned((8'hb1)))));
                    end
                  else
                    begin
                      reg3550 <= wire3541[(3'h6):(3'h4)];
                      reg3551 <= ($unsigned($signed($unsigned(reg3552))) ?
                          (~^{forvar3552[(1'h1):(1'h1)]}) : ($signed(forvar3552) & $unsigned({forvar3548})));
                      reg3552 <= reg3544[(1'h0):(1'h0)];
                    end
                  for (forvar3553 = (1'h0); (forvar3553 < (2'h2)); forvar3553 = (forvar3553 + (1'h1)))
                    begin
                      reg3554 <= reg3553;
                      reg3555 <= ($unsigned((wire3541 && (8'hb5))) >> (((+forvar3548) >= $unsigned(reg3558)) ?
                          {(forvar3545 ?
                                  forvar3553 : forvar3545)} : $unsigned(reg3547[(3'h4):(2'h2)])));
                      reg3556 <= $unsigned(forvar3547);
                    end
                end
              reg3557 <= (reg3545 ?
                  (((reg3552 == reg3555) ?
                          ((8'hae) ?
                              reg3556 : forvar3544) : (reg3549 == reg3549)) ?
                      $signed(reg3550) : (forvar3549[(4'h8):(3'h5)] > forvar3545)) : (reg3551[(1'h0):(1'h0)] + $unsigned((reg3550 * reg3556))));
            end
          for (forvar3558 = (1'h0); (forvar3558 < (1'h1)); forvar3558 = (forvar3558 + (1'h1)))
            begin
              for (forvar3559 = (1'h0); (forvar3559 < (1'h0)); forvar3559 = (forvar3559 + (1'h1)))
                begin
                  for (forvar3560 = (1'h0); (forvar3560 < (1'h1)); forvar3560 = (forvar3560 + (1'h1)))
                    begin
                      reg3561 <= {(($unsigned(forvar3544) ?
                                  (~|(8'hb3)) : $signed((8'h9c))) ?
                              (8'hb0) : reg3546[(1'h0):(1'h0)])};
                      reg3562 <= reg3558;
                      reg3563 <= (~|(~reg3548));
                    end
                  if ($unsigned($unsigned(({wire3540} <<< $signed(reg3563)))))
                    begin
                      reg3564 <= $unsigned(forvar3552[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg3564 <= $unsigned(reg3546[(4'h9):(1'h0)]);
                    end
                end
              reg3565 <= (~|(8'ha9));
              for (forvar3566 = (1'h0); (forvar3566 < (2'h3)); forvar3566 = (forvar3566 + (1'h1)))
                begin
                  for (forvar3567 = (1'h0); (forvar3567 < (1'h0)); forvar3567 = (forvar3567 + (1'h1)))
                    begin
                      reg3568 <= (~^forvar3552[(3'h7):(2'h2)]);
                      reg3569 <= $signed((~&(^$signed(wire3543))));
                      reg3570 <= forvar3548[(2'h3):(1'h0)];
                      reg3571 <= ($signed(((~^forvar3559) > $signed(reg3556))) ?
                          (~&(~&(8'h9d))) : $signed($signed($signed((8'hac)))));
                    end
                  reg3572 <= reg3553[(1'h0):(1'h0)];
                  for (forvar3573 = (1'h0); (forvar3573 < (1'h1)); forvar3573 = (forvar3573 + (1'h1)))
                    begin
                      reg3574 <= forvar3560;
                      reg3575 <= reg3546[(3'h5):(2'h3)];
                      reg3576 <= ($unsigned(reg3557[(4'h9):(3'h4)]) && (forvar3573 * $unsigned(reg3549[(1'h1):(1'h1)])));
                    end
                end
            end
          for (forvar3577 = (1'h0); (forvar3577 < (2'h2)); forvar3577 = (forvar3577 + (1'h1)))
            begin
              for (forvar3578 = (1'h0); (forvar3578 < (1'h0)); forvar3578 = (forvar3578 + (1'h1)))
                begin
                  for (forvar3579 = (1'h0); (forvar3579 < (1'h0)); forvar3579 = (forvar3579 + (1'h1)))
                    begin
                      reg3580 <= ((8'haa) | {forvar3560});
                      reg3581 <= {(((reg3572 ? forvar3545 : reg3569) ?
                              $unsigned(reg3565) : (forvar3547 ~^ forvar3559)) == reg3562)};
                      reg3582 <= (((reg3570[(3'h5):(1'h1)] ?
                              forvar3558[(3'h6):(3'h4)] : forvar3545) <= reg3576) ?
                          forvar3553[(2'h2):(1'h0)] : forvar3545[(3'h4):(1'h0)]);
                      reg3583 <= {forvar3577};
                    end
                  reg3584 <= reg3554[(4'hb):(2'h2)];
                  if ({(&((reg3549 < reg3548) - (8'haf)))})
                    begin
                      reg3585 <= reg3584[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3585 <= {(8'h9e)};
                      reg3586 <= (~($unsigned($unsigned(reg3581)) + (forvar3552[(4'h9):(3'h7)] ?
                          ((8'ha0) ?
                              reg3564 : reg3568) : (forvar3560 <= reg3571))));
                      reg3587 <= reg3548[(1'h0):(1'h0)];
                      reg3588 <= {((~|(reg3550 - reg3553)) ?
                              reg3550 : $unsigned(((8'haa) ?
                                  reg3585 : forvar3552)))};
                    end
                end
              if ((reg3586 ?
                  reg3570[(4'h9):(3'h4)] : (($unsigned((8'hb2)) ?
                          (forvar3573 | reg3583) : (!forvar3567)) ?
                      (|$signed(reg3576)) : ((-(8'hb2)) != (&forvar3547)))))
                begin
                  for (forvar3589 = (1'h0); (forvar3589 < (2'h3)); forvar3589 = (forvar3589 + (1'h1)))
                    begin
                      reg3590 <= wire3542;
                      reg3591 <= ($signed(reg3569) != $signed(wire3543[(4'hc):(4'h9)]));
                      reg3592 <= reg3576[(4'hb):(3'h4)];
                    end
                  for (forvar3593 = (1'h0); (forvar3593 < (2'h3)); forvar3593 = (forvar3593 + (1'h1)))
                    begin
                      reg3594 <= $signed(reg3551[(1'h0):(1'h0)]);
                      reg3595 <= $signed($signed($signed(reg3591[(1'h1):(1'h0)])));
                      reg3596 <= ({(forvar3558[(3'h4):(1'h0)] > reg3562)} ?
                          $unsigned($signed({reg3555})) : reg3591[(4'h9):(1'h0)]);
                      reg3597 <= {reg3562[(4'hc):(1'h0)]};
                    end
                  for (forvar3598 = (1'h0); (forvar3598 < (1'h0)); forvar3598 = (forvar3598 + (1'h1)))
                    begin
                      reg3599 <= (!reg3563[(4'hd):(4'h9)]);
                      reg3600 <= (({(reg3568 || reg3556)} - (reg3575 ^~ (forvar3545 << reg3551))) ?
                          (^~$unsigned(reg3562[(3'h4):(3'h4)])) : wire3543[(4'hc):(4'hb)]);
                    end
                end
              else
                begin
                  for (forvar3589 = (1'h0); (forvar3589 < (2'h3)); forvar3589 = (forvar3589 + (1'h1)))
                    begin
                      reg3590 <= $signed((((forvar3544 > reg3549) || (reg3584 << (8'hb7))) ?
                          ((forvar3559 ? forvar3598 : reg3558) ?
                              $unsigned((8'haa)) : reg3599) : ((reg3549 <<< reg3575) + $signed(reg3586))));
                      reg3591 <= $signed(reg3564);
                      reg3592 <= (($signed((8'h9c)) ?
                              forvar3545 : $signed(reg3587[(3'h4):(2'h2)])) ?
                          reg3594[(4'ha):(3'h5)] : {((~forvar3560) ?
                                  reg3556 : reg3581[(2'h2):(2'h2)])});
                    end
                  if ((~|reg3585))
                    begin
                      reg3593 <= $unsigned(($unsigned(reg3556[(3'h7):(1'h0)]) ?
                          (reg3551 ?
                              reg3584 : $unsigned(reg3574)) : {{reg3554}}));
                      reg3594 <= $signed((-$unsigned(reg3555)));
                    end
                  else
                    begin
                      reg3593 <= $signed((reg3585[(4'hd):(4'ha)] << {$signed(reg3595)}));
                      reg3594 <= $signed(forvar3598);
                      reg3595 <= reg3565[(1'h1):(1'h0)];
                      reg3596 <= (~^forvar3547);
                    end
                  reg3597 <= (&(^~wire3540));
                end
              for (forvar3601 = (1'h0); (forvar3601 < (2'h3)); forvar3601 = (forvar3601 + (1'h1)))
                begin
                  for (forvar3602 = (1'h0); (forvar3602 < (2'h2)); forvar3602 = (forvar3602 + (1'h1)))
                    begin
                      reg3603 <= (^wire3543[(3'h7):(3'h5)]);
                      reg3604 <= forvar3544;
                      reg3605 <= $unsigned(($signed((reg3570 ?
                              reg3599 : forvar3558)) ?
                          $unsigned((~&forvar3602)) : (!$signed(reg3548))));
                      reg3606 <= (((reg3580[(4'h9):(3'h6)] ?
                              $unsigned(forvar3559) : $unsigned(reg3553)) ^ $signed((reg3586 >= reg3565))) ?
                          forvar3601 : (+reg3596));
                    end
                  for (forvar3607 = (1'h0); (forvar3607 < (1'h1)); forvar3607 = (forvar3607 + (1'h1)))
                    begin
                      reg3608 <= $unsigned((~reg3551));
                    end
                  for (forvar3609 = (1'h0); (forvar3609 < (1'h0)); forvar3609 = (forvar3609 + (1'h1)))
                    begin
                      reg3610 <= ((((forvar3553 ^ reg3550) << (reg3575 || forvar3601)) ?
                              $unsigned((reg3581 <= reg3569)) : forvar3601[(1'h1):(1'h0)]) ?
                          $unsigned((forvar3547 ?
                              $unsigned((8'ha8)) : (+(8'ha6)))) : (reg3576 ?
                              (|forvar3609) : {$signed(wire3542)}));
                      reg3611 <= (^~(&$signed((forvar3559 ?
                          reg3595 : forvar3548))));
                      reg3612 <= (~&{$signed((!(8'haf)))});
                    end
                end
            end
        end
      if ($signed($unsigned(($unsigned(reg3595) ?
          forvar3548[(4'ha):(4'h9)] : (!reg3557)))))
        begin
          for (forvar3613 = (1'h0); (forvar3613 < (1'h1)); forvar3613 = (forvar3613 + (1'h1)))
            begin
              if ($signed(reg3610[(1'h0):(1'h0)]))
                begin
                  if ($unsigned(({$unsigned(reg3544)} ?
                      $signed((+wire3542)) : $signed($unsigned((8'hb2))))))
                    begin
                      reg3614 <= {forvar3601};
                    end
                  else
                    begin
                      reg3614 <= (reg3603[(4'h9):(4'h8)] ?
                          ($signed((forvar3558 < wire3541)) ?
                              ({reg3568} ?
                                  (reg3592 ?
                                      (8'hb2) : reg3563) : forvar3613[(2'h2):(2'h2)]) : reg3587) : ((^~$unsigned(forvar3552)) ?
                              ($unsigned(reg3590) == $signed(reg3550)) : ((^forvar3598) ?
                                  $unsigned(reg3563) : (+reg3562))));
                    end
                  for (forvar3615 = (1'h0); (forvar3615 < (2'h2)); forvar3615 = (forvar3615 + (1'h1)))
                    begin
                      reg3616 <= reg3557;
                      reg3617 <= $signed((forvar3566[(1'h0):(1'h0)] ?
                          forvar3548[(2'h2):(1'h1)] : $signed($unsigned(reg3608))));
                      reg3618 <= ({($unsigned(forvar3566) == (^~forvar3578))} ?
                          $signed($unsigned((reg3562 ?
                              reg3570 : reg3582))) : $signed({(forvar3615 && forvar3615)}));
                    end
                end
              else
                begin
                  reg3614 <= (8'h9c);
                  if ((&forvar3573[(4'h9):(4'h8)]))
                    begin
                      reg3615 <= $signed(($signed((reg3561 + reg3616)) || $unsigned((reg3610 ^ (8'haa)))));
                      reg3616 <= $signed(reg3599[(3'h5):(1'h1)]);
                      reg3617 <= {(((forvar3547 ?
                                  reg3547 : (8'h9e)) ~^ {reg3544}) ?
                              wire3543 : (|$unsigned(forvar3577)))};
                      reg3618 <= (|(((8'haa) ?
                              reg3563[(2'h3):(1'h1)] : (reg3575 >>> reg3610)) ?
                          $signed(forvar3593[(3'h4):(3'h4)]) : (forvar3559 - (~&forvar3615))));
                    end
                  else
                    begin
                      reg3615 <= reg3593;
                    end
                end
              reg3619 <= ((forvar3566 - reg3552[(2'h2):(1'h1)]) ?
                  ($signed((^~reg3616)) ?
                      (^~reg3585[(4'hd):(3'h6)]) : reg3572) : $unsigned($signed((reg3562 ~^ reg3608))));
              reg3620 <= $signed((forvar3615[(3'h5):(3'h4)] && (^~wire3540)));
            end
          reg3621 <= ((((forvar3593 == reg3608) | {(8'hae)}) ^~ (-$unsigned(reg3585))) == reg3588);
        end
      else
        begin
          for (forvar3613 = (1'h0); (forvar3613 < (1'h1)); forvar3613 = (forvar3613 + (1'h1)))
            begin
              if ($signed((~((-reg3550) ? (forvar3607 ^ reg3545) : {(8'hb3)}))))
                begin
                  if (({reg3549[(3'h7):(3'h6)]} ?
                      ((reg3620[(3'h5):(1'h0)] + reg3568) ?
                          (^(reg3586 ?
                              reg3558 : (8'hac))) : reg3575[(2'h3):(1'h1)]) : ((reg3590 - reg3553) + $unsigned(reg3548[(3'h6):(3'h4)]))))
                    begin
                      reg3614 <= (8'hb0);
                      reg3615 <= reg3593;
                      reg3616 <= (($signed(((8'ha2) < (8'ha3))) == {(reg3585 < forvar3566)}) ?
                          ((8'hb8) ^~ {forvar3558}) : (($unsigned(reg3592) + (!forvar3559)) <<< (~&{forvar3552})));
                      reg3617 <= {$unsigned($unsigned((~(8'hae))))};
                    end
                  else
                    begin
                      reg3614 <= $unsigned(({reg3588[(1'h0):(1'h0)]} ?
                          $unsigned((reg3591 ?
                              (8'hac) : reg3550)) : forvar3578[(1'h0):(1'h0)]));
                      reg3615 <= ((forvar3553[(1'h1):(1'h1)] >>> forvar3544) ?
                          reg3596[(3'h5):(1'h1)] : $unsigned(($unsigned(reg3561) | forvar3567[(3'h4):(3'h4)])));
                      reg3616 <= (forvar3552[(3'h7):(3'h4)] & $signed((reg3548[(1'h0):(1'h0)] ?
                          reg3599 : $unsigned(reg3593))));
                    end
                  reg3618 <= $unsigned(((forvar3601[(3'h4):(1'h1)] ?
                      ((8'ha3) != reg3603) : $unsigned(reg3581)) & reg3586));
                  for (forvar3619 = (1'h0); (forvar3619 < (2'h2)); forvar3619 = (forvar3619 + (1'h1)))
                    begin
                      reg3620 <= reg3597[(1'h1):(1'h1)];
                      reg3621 <= reg3615;
                      reg3622 <= (8'haf);
                    end
                  for (forvar3623 = (1'h0); (forvar3623 < (1'h1)); forvar3623 = (forvar3623 + (1'h1)))
                    begin
                      reg3624 <= forvar3566[(3'h6):(3'h6)];
                      reg3625 <= ($signed((+$signed(forvar3552))) ?
                          reg3576[(3'h6):(3'h5)] : ((&reg3594[(3'h4):(2'h2)]) ?
                              ((8'ha3) ?
                                  (~^forvar3579) : $unsigned(reg3612)) : ($unsigned((8'ha3)) ?
                                  (forvar3609 ?
                                      reg3599 : reg3548) : reg3619[(2'h3):(1'h1)])));
                    end
                end
              else
                begin
                  if (forvar3553[(1'h0):(1'h0)])
                    begin
                      reg3614 <= {(8'hb3)};
                    end
                  else
                    begin
                      reg3614 <= ($unsigned($signed(forvar3598[(1'h1):(1'h1)])) ?
                          (({(8'ha3)} > (forvar3589 || reg3604)) ?
                              ((~reg3611) || $unsigned(wire3541)) : (~(~|reg3561))) : $signed(reg3619));
                      reg3615 <= (8'hb9);
                      reg3616 <= {reg3611};
                      reg3617 <= ($signed(reg3550[(3'h5):(1'h1)]) <<< {wire3542});
                    end
                  reg3618 <= (forvar3593 ^ reg3587[(2'h3):(2'h3)]);
                  if (forvar3547)
                    begin
                      reg3619 <= {$unsigned(reg3564[(2'h2):(2'h2)])};
                      reg3620 <= forvar3558;
                      reg3621 <= reg3545;
                      reg3622 <= reg3608;
                    end
                  else
                    begin
                      reg3619 <= (-reg3570[(3'h5):(3'h4)]);
                      reg3620 <= $unsigned((&forvar3593[(3'h4):(1'h1)]));
                      reg3621 <= forvar3545[(4'h9):(3'h7)];
                      reg3622 <= (8'hba);
                    end
                end
              for (forvar3626 = (1'h0); (forvar3626 < (2'h3)); forvar3626 = (forvar3626 + (1'h1)))
                begin
                  if ($unsigned($signed({forvar3553[(1'h0):(1'h0)]})))
                    begin
                      reg3627 <= reg3565;
                      reg3628 <= (&reg3548[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg3627 <= {reg3595[(4'h9):(3'h4)]};
                      reg3628 <= reg3593[(4'h9):(3'h4)];
                      reg3629 <= $unsigned($signed(forvar3573[(2'h2):(1'h1)]));
                      reg3630 <= ({reg3611} >> ((!$signed((8'haa))) ?
                          wire3541[(4'hb):(1'h1)] : ((reg3544 > reg3565) ?
                              (forvar3593 ?
                                  reg3603 : reg3610) : $unsigned(reg3595))));
                    end
                  for (forvar3631 = (1'h0); (forvar3631 < (2'h3)); forvar3631 = (forvar3631 + (1'h1)))
                    begin
                      reg3632 <= $signed($signed(($signed(reg3620) ?
                          reg3612[(3'h4):(2'h2)] : (forvar3601 ?
                              reg3548 : reg3617))));
                      reg3633 <= {(forvar3623 ^~ (!reg3592))};
                      reg3634 <= (forvar3573 ?
                          $signed((+((8'ha9) ^ reg3569))) : $signed((~reg3568[(2'h2):(2'h2)])));
                      reg3635 <= reg3615[(3'h4):(3'h4)];
                    end
                  for (forvar3636 = (1'h0); (forvar3636 < (2'h3)); forvar3636 = (forvar3636 + (1'h1)))
                    begin
                      reg3637 <= $unsigned((~^reg3590[(4'h9):(3'h6)]));
                      reg3638 <= (reg3622[(3'h6):(3'h6)] <= forvar3573);
                      reg3639 <= $unsigned($signed((reg3584 || (forvar3567 ?
                          reg3585 : (8'hb3)))));
                      reg3640 <= reg3603;
                    end
                  for (forvar3641 = (1'h0); (forvar3641 < (2'h2)); forvar3641 = (forvar3641 + (1'h1)))
                    begin
                      reg3642 <= reg3591;
                      reg3643 <= $signed($unsigned(({forvar3609} + (8'ha6))));
                      reg3644 <= ($unsigned({(!reg3576)}) ?
                          reg3570[(3'h5):(3'h4)] : {(-$signed(reg3627))});
                    end
                end
            end
          if ($unsigned($signed(reg3639[(1'h1):(1'h0)])))
            begin
              reg3645 <= $signed($signed(reg3557[(3'h5):(1'h0)]));
              for (forvar3646 = (1'h0); (forvar3646 < (1'h0)); forvar3646 = (forvar3646 + (1'h1)))
                begin
                  for (forvar3647 = (1'h0); (forvar3647 < (2'h3)); forvar3647 = (forvar3647 + (1'h1)))
                    begin
                      reg3648 <= reg3594[(1'h0):(1'h0)];
                      reg3649 <= $unsigned(reg3621[(4'h8):(3'h5)]);
                      reg3650 <= $unsigned(forvar3545[(1'h1):(1'h1)]);
                      reg3651 <= (+(($unsigned(reg3550) ?
                          {reg3568} : reg3611) > ({forvar3636} != {forvar3559})));
                    end
                  for (forvar3652 = (1'h0); (forvar3652 < (1'h0)); forvar3652 = (forvar3652 + (1'h1)))
                    begin
                      reg3653 <= ($unsigned($unsigned((^reg3563))) ?
                          forvar3559[(1'h1):(1'h0)] : (~reg3570[(2'h3):(2'h2)]));
                      reg3654 <= $signed((~|$signed($signed((8'hae)))));
                    end
                  for (forvar3655 = (1'h0); (forvar3655 < (1'h0)); forvar3655 = (forvar3655 + (1'h1)))
                    begin
                      reg3656 <= (~^$signed({(reg3583 || reg3650)}));
                    end
                  for (forvar3657 = (1'h0); (forvar3657 < (1'h1)); forvar3657 = (forvar3657 + (1'h1)))
                    begin
                      reg3658 <= (&reg3620[(1'h0):(1'h0)]);
                      reg3659 <= (+((!forvar3549[(1'h1):(1'h0)]) ?
                          ($unsigned(reg3593) ?
                              ((8'h9d) <<< forvar3613) : $signed(reg3622)) : ($signed(reg3594) ?
                              reg3643[(1'h0):(1'h0)] : $signed(forvar3647))));
                    end
                end
              for (forvar3660 = (1'h0); (forvar3660 < (1'h0)); forvar3660 = (forvar3660 + (1'h1)))
                begin
                  if (reg3640)
                    begin
                      reg3661 <= ($unsigned(((reg3635 && forvar3646) != $unsigned(reg3597))) ^~ (reg3644 ^~ $signed((reg3559 ^~ forvar3619))));
                      reg3662 <= ((reg3651[(2'h3):(2'h2)] != $unsigned($unsigned(reg3656))) ?
                          $signed(reg3603[(4'hc):(4'h8)]) : {$unsigned($unsigned(reg3605))});
                      reg3663 <= $unsigned($unsigned(forvar3660));
                    end
                  else
                    begin
                      reg3661 <= $signed(((~|reg3544[(2'h2):(1'h0)]) && {(reg3554 && (8'ha2))}));
                    end
                end
              for (forvar3664 = (1'h0); (forvar3664 < (2'h2)); forvar3664 = (forvar3664 + (1'h1)))
                begin
                  if ((~(-($signed(reg3632) & (forvar3601 ?
                      reg3653 : reg3562)))))
                    begin
                      reg3665 <= reg3662[(1'h0):(1'h0)];
                      reg3666 <= $unsigned(($unsigned($signed(reg3665)) ?
                          $unsigned((~^reg3555)) : $signed((reg3584 << reg3653))));
                      reg3667 <= ({(^~reg3656)} ?
                          $unsigned(((8'ha7) ^~ reg3571[(1'h1):(1'h0)])) : $signed($unsigned((reg3605 ?
                              forvar3544 : reg3637))));
                      reg3668 <= ($signed($signed(reg3612)) ?
                          (($unsigned(forvar3573) <<< (reg3651 && (8'ha0))) ?
                              reg3555[(1'h1):(1'h1)] : ((forvar3589 ?
                                  forvar3652 : reg3558) < (^~reg3610))) : (!$unsigned((~^forvar3578))));
                    end
                  else
                    begin
                      reg3665 <= $signed((-($unsigned(reg3668) ?
                          $signed(forvar3566) : $unsigned(forvar3607))));
                    end
                  for (forvar3669 = (1'h0); (forvar3669 < (1'h0)); forvar3669 = (forvar3669 + (1'h1)))
                    begin
                      reg3670 <= {reg3628[(1'h0):(1'h0)]};
                      reg3671 <= reg3597[(4'h8):(3'h6)];
                      reg3672 <= {{{(~reg3651)}}};
                      reg3673 <= $signed(($signed(forvar3547) ?
                          $unsigned((reg3606 >> reg3556)) : reg3588[(1'h0):(1'h0)]));
                    end
                  if (($unsigned($signed((&(8'hb4)))) < $signed($unsigned(reg3580[(1'h1):(1'h1)]))))
                    begin
                      reg3674 <= ($signed(({reg3555} >>> (forvar3566 ?
                              reg3562 : reg3658))) ?
                          $signed($signed(reg3575[(3'h6):(3'h5)])) : {(!$unsigned((8'ha8)))});
                    end
                  else
                    begin
                      reg3674 <= reg3605[(3'h6):(2'h3)];
                      reg3675 <= $unsigned(forvar3602[(4'hb):(3'h4)]);
                    end
                  for (forvar3676 = (1'h0); (forvar3676 < (2'h2)); forvar3676 = (forvar3676 + (1'h1)))
                    begin
                      reg3677 <= forvar3602[(4'hc):(1'h1)];
                      reg3678 <= reg3614[(1'h1):(1'h1)];
                      reg3679 <= $unsigned(reg3643[(1'h1):(1'h1)]);
                      reg3680 <= reg3624;
                    end
                end
            end
          else
            begin
              for (forvar3645 = (1'h0); (forvar3645 < (2'h3)); forvar3645 = (forvar3645 + (1'h1)))
                begin
                  reg3646 <= reg3575[(4'h9):(2'h2)];
                  for (forvar3647 = (1'h0); (forvar3647 < (1'h1)); forvar3647 = (forvar3647 + (1'h1)))
                    begin
                      reg3648 <= reg3635;
                      reg3649 <= forvar3560[(4'hc):(3'h7)];
                      reg3650 <= (8'ha5);
                      reg3651 <= (reg3550 ?
                          (~|$signed($signed(reg3659))) : $signed($unsigned((reg3585 <<< (8'had)))));
                    end
                  reg3652 <= {({reg3656[(1'h1):(1'h1)]} ?
                          $unsigned(reg3673) : ({reg3545} ?
                              reg3646[(3'h4):(1'h0)] : $unsigned(reg3640)))};
                  reg3653 <= ({{$signed(reg3630)}} <<< forvar3664);
                end
              for (forvar3654 = (1'h0); (forvar3654 < (2'h3)); forvar3654 = (forvar3654 + (1'h1)))
                begin
                  if ($unsigned({{(reg3568 >= reg3675)}}))
                    begin
                      reg3655 <= forvar3641[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg3655 <= $unsigned($unsigned(forvar3559[(2'h2):(2'h2)]));
                    end
                  for (forvar3656 = (1'h0); (forvar3656 < (2'h2)); forvar3656 = (forvar3656 + (1'h1)))
                    begin
                      reg3657 <= {forvar3548[(2'h2):(1'h0)]};
                      reg3658 <= ((reg3555 >= $signed((reg3615 >>> reg3580))) ?
                          $signed((((8'ha9) >> (8'hae)) ?
                              reg3564 : (~&reg3597))) : (((8'hae) << reg3627[(2'h3):(1'h1)]) >= ($unsigned(reg3657) ?
                              forvar3553 : reg3590)));
                      reg3659 <= $unsigned(reg3571);
                    end
                  if (($signed((reg3661 ^ reg3611)) ?
                      $signed((-(8'hb5))) : ($unsigned($unsigned(reg3595)) ?
                          $signed($unsigned(reg3624)) : ((forvar3645 ?
                                  (8'hb5) : reg3582) ?
                              ((8'haa) << reg3576) : {(8'hb8)}))))
                    begin
                      reg3660 <= ((~reg3670) ?
                          $signed(({reg3562} ?
                              reg3590 : {(8'had)})) : $unsigned(reg3580));
                      reg3661 <= forvar3558[(4'h9):(4'h9)];
                    end
                  else
                    begin
                      reg3660 <= $unsigned($signed((!{(8'hb6)})));
                      reg3661 <= $unsigned($signed($unsigned((|forvar3656))));
                      reg3662 <= ((8'ha3) ?
                          ($signed(((8'hb8) ?
                              reg3667 : reg3580)) + forvar3553) : (|forvar3598));
                      reg3663 <= reg3550[(3'h5):(1'h0)];
                    end
                end
              for (forvar3664 = (1'h0); (forvar3664 < (2'h2)); forvar3664 = (forvar3664 + (1'h1)))
                begin
                  if ((~&$signed($unsigned($signed(reg3611)))))
                    begin
                      reg3665 <= {$signed($unsigned((forvar3579 != reg3570)))};
                      reg3666 <= reg3611;
                      reg3667 <= $signed((((reg3656 >>> reg3629) ?
                          forvar3560 : (~&forvar3598)) || $unsigned($signed(forvar3645))));
                    end
                  else
                    begin
                      reg3665 <= {(~|$unsigned({reg3574}))};
                    end
                  if (forvar3602[(2'h3):(1'h1)])
                    begin
                      reg3668 <= forvar3656[(2'h3):(2'h2)];
                      reg3669 <= reg3603;
                      reg3670 <= reg3605[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg3668 <= reg3595[(3'h5):(2'h3)];
                      reg3669 <= reg3679;
                      reg3670 <= reg3627[(1'h1):(1'h1)];
                    end
                end
              for (forvar3671 = (1'h0); (forvar3671 < (2'h3)); forvar3671 = (forvar3671 + (1'h1)))
                begin
                  for (forvar3672 = (1'h0); (forvar3672 < (1'h1)); forvar3672 = (forvar3672 + (1'h1)))
                    begin
                      reg3673 <= (reg3658[(3'h7):(3'h7)] + ($signed($signed(forvar3593)) ?
                          ($unsigned(reg3549) ?
                              (reg3606 ?
                                  reg3610 : reg3606) : reg3648) : (-reg3663)));
                      reg3674 <= ($unsigned((|reg3642[(5'h10):(3'h7)])) == (&((&reg3572) ?
                          (forvar3577 ?
                              reg3673 : (8'ha6)) : $signed((8'ha3)))));
                      reg3675 <= {reg3660[(3'h5):(3'h4)]};
                      reg3676 <= (|((8'ha2) > forvar3613[(4'h9):(3'h6)]));
                    end
                  reg3677 <= $signed(reg3666);
                end
            end
          for (forvar3681 = (1'h0); (forvar3681 < (1'h0)); forvar3681 = (forvar3681 + (1'h1)))
            begin
              for (forvar3682 = (1'h0); (forvar3682 < (2'h2)); forvar3682 = (forvar3682 + (1'h1)))
                begin
                  if ($unsigned((~&reg3584[(2'h3):(1'h1)])))
                    begin
                      reg3683 <= $signed((forvar3615[(1'h1):(1'h1)] ?
                          $unsigned((~&forvar3623)) : $unsigned($signed((8'h9c)))));
                      reg3684 <= $signed($unsigned({forvar3598}));
                      reg3685 <= (^forvar3646);
                    end
                  else
                    begin
                      reg3683 <= $unsigned($signed(forvar3567[(3'h5):(3'h4)]));
                      reg3684 <= forvar3601[(3'h6):(2'h3)];
                      reg3685 <= forvar3544;
                    end
                  for (forvar3686 = (1'h0); (forvar3686 < (1'h0)); forvar3686 = (forvar3686 + (1'h1)))
                    begin
                      reg3687 <= $signed(reg3572[(4'h8):(2'h3)]);
                    end
                  reg3688 <= ((~&$signed(reg3570)) ?
                      (~|(!(~|reg3637))) : $unsigned((reg3618 ?
                          reg3552 : (~reg3658))));
                end
              if (reg3588[(2'h2):(1'h1)])
                begin
                  if (($signed(reg3648[(1'h0):(1'h0)]) ^ ($signed({reg3620}) ?
                      $unsigned((reg3608 >= reg3620)) : $signed($signed(reg3633)))))
                    begin
                      reg3689 <= $unsigned({$signed($signed(reg3611))});
                      reg3690 <= ($unsigned(({forvar3613} ?
                          reg3662 : {forvar3664})) + wire3543);
                    end
                  else
                    begin
                      reg3689 <= reg3593[(3'h6):(2'h2)];
                      reg3690 <= (^~{reg3621});
                      reg3691 <= $signed(forvar3623);
                    end
                end
              else
                begin
                  if ($unsigned({$unsigned($signed((8'hb3)))}))
                    begin
                      reg3689 <= ($signed(reg3616[(1'h0):(1'h0)]) ~^ (reg3619[(1'h1):(1'h0)] ?
                          $signed((reg3576 ?
                              reg3583 : reg3656)) : ((wire3542 - reg3597) ?
                              $signed(reg3547) : (reg3627 ?
                                  reg3684 : (8'hb6)))));
                      reg3690 <= reg3620;
                    end
                  else
                    begin
                      reg3689 <= ((reg3611 ?
                          (|reg3612) : reg3679[(2'h2):(1'h1)]) | (!reg3620));
                      reg3690 <= forvar3573;
                      reg3691 <= {{$signed($signed(reg3670))}};
                    end
                  if ($signed($unsigned((-{forvar3560}))))
                    begin
                      reg3692 <= ((((^reg3587) <= {reg3580}) == $signed((~|reg3605))) ?
                          reg3687[(1'h0):(1'h0)] : (+$signed($signed(reg3653))));
                      reg3693 <= $unsigned(((~|{(8'hb6)}) != (reg3615[(3'h4):(2'h2)] ?
                          (!forvar3660) : {reg3671})));
                      reg3694 <= forvar3579;
                      reg3695 <= (reg3614[(3'h5):(1'h0)] == wire3542[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg3692 <= $unsigned($unsigned(({reg3629} ?
                          forvar3559[(3'h4):(1'h1)] : (reg3544 ?
                              reg3611 : (8'hab)))));
                    end
                end
              reg3696 <= (8'hac);
            end
          for (forvar3697 = (1'h0); (forvar3697 < (1'h1)); forvar3697 = (forvar3697 + (1'h1)))
            begin
              for (forvar3698 = (1'h0); (forvar3698 < (2'h3)); forvar3698 = (forvar3698 + (1'h1)))
                begin
                  for (forvar3699 = (1'h0); (forvar3699 < (1'h1)); forvar3699 = (forvar3699 + (1'h1)))
                    begin
                      reg3700 <= reg3671[(3'h5):(3'h5)];
                    end
                  reg3701 <= (8'ha7);
                end
              for (forvar3702 = (1'h0); (forvar3702 < (1'h0)); forvar3702 = (forvar3702 + (1'h1)))
                begin
                  if (($unsigned((^$signed(reg3676))) ?
                      forvar3601[(2'h3):(2'h3)] : {reg3552[(2'h3):(2'h2)]}))
                    begin
                      reg3703 <= forvar3660;
                    end
                  else
                    begin
                      reg3703 <= $signed($signed((((8'hae) ?
                              reg3570 : reg3600) ?
                          (~|reg3591) : (forvar3560 ? reg3592 : forvar3645))));
                      reg3704 <= ((reg3608[(3'h7):(2'h2)] ?
                              forvar3631[(2'h2):(1'h0)] : ((~^forvar3623) + (reg3651 ^~ forvar3645))) ?
                          ((forvar3602[(1'h0):(1'h0)] ?
                                  $signed(reg3656) : reg3559) ?
                              {(8'hae)} : reg3608[(4'h8):(3'h5)]) : $unsigned($signed((~|reg3680))));
                      reg3705 <= forvar3641[(1'h0):(1'h0)];
                    end
                  for (forvar3706 = (1'h0); (forvar3706 < (2'h2)); forvar3706 = (forvar3706 + (1'h1)))
                    begin
                      reg3707 <= reg3570;
                    end
                  if ($signed(forvar3626[(2'h2):(1'h1)]))
                    begin
                      reg3708 <= (^reg3637);
                    end
                  else
                    begin
                      reg3708 <= (forvar3657 ?
                          $unsigned($signed((reg3550 != reg3606))) : {($signed(reg3692) < $unsigned(reg3575))});
                      reg3709 <= reg3585[(4'hb):(2'h2)];
                    end
                end
              for (forvar3710 = (1'h0); (forvar3710 < (2'h3)); forvar3710 = (forvar3710 + (1'h1)))
                begin
                  for (forvar3711 = (1'h0); (forvar3711 < (1'h1)); forvar3711 = (forvar3711 + (1'h1)))
                    begin
                      reg3712 <= ((|reg3669) ?
                          $signed($signed($signed(reg3587))) : ($signed((!reg3658)) ?
                              reg3629 : $unsigned((forvar3647 ?
                                  reg3549 : reg3692))));
                      reg3713 <= (~&$signed((~|$signed(reg3667))));
                      reg3714 <= $unsigned((forvar3549 ?
                          $unsigned((~|forvar3697)) : {(reg3625 >> reg3586)}));
                    end
                end
            end
        end
      for (forvar3715 = (1'h0); (forvar3715 < (1'h0)); forvar3715 = (forvar3715 + (1'h1)))
        begin
          reg3716 <= reg3550;
          for (forvar3717 = (1'h0); (forvar3717 < (2'h2)); forvar3717 = (forvar3717 + (1'h1)))
            begin
              reg3718 <= reg3630[(3'h5):(2'h3)];
              for (forvar3719 = (1'h0); (forvar3719 < (1'h1)); forvar3719 = (forvar3719 + (1'h1)))
                begin
                  if (reg3659[(1'h1):(1'h1)])
                    begin
                      reg3720 <= $signed((~&((~&forvar3647) ?
                          $unsigned((8'hac)) : (reg3675 ?
                              (8'ha4) : forvar3579))));
                      reg3721 <= (reg3625 ? (+$unsigned(reg3615)) : reg3653);
                    end
                  else
                    begin
                      reg3720 <= reg3580[(4'h8):(2'h3)];
                      reg3721 <= ($unsigned($unsigned({(8'haa)})) ?
                          reg3703 : ((((8'had) > reg3557) ?
                              $unsigned(reg3575) : (&reg3624)) - ($unsigned(reg3640) ?
                              (reg3622 ?
                                  reg3637 : forvar3664) : reg3583[(1'h0):(1'h0)])));
                    end
                  for (forvar3722 = (1'h0); (forvar3722 < (2'h3)); forvar3722 = (forvar3722 + (1'h1)))
                    begin
                      reg3723 <= $unsigned(forvar3589[(2'h3):(1'h0)]);
                      reg3724 <= forvar3676;
                    end
                  for (forvar3725 = (1'h0); (forvar3725 < (2'h2)); forvar3725 = (forvar3725 + (1'h1)))
                    begin
                      reg3726 <= $unsigned($signed((+(reg3610 ?
                          (8'ha1) : reg3552))));
                      reg3727 <= $signed({({reg3630} ?
                              $signed(reg3612) : ((8'haf) ?
                                  (8'ha6) : reg3615))});
                    end
                end
              if ($unsigned((+$signed(reg3658))))
                begin
                  if ((forvar3560[(3'h7):(2'h3)] && reg3606[(4'h8):(2'h2)]))
                    begin
                      reg3728 <= (($signed($signed(reg3668)) ?
                          reg3723[(1'h1):(1'h0)] : $signed((reg3617 >> reg3708))) == forvar3598);
                      reg3729 <= (~$signed(forvar3699[(3'h5):(3'h4)]));
                      reg3730 <= ($unsigned(reg3703[(3'h4):(1'h0)]) ?
                          (^(^$signed(reg3572))) : ($unsigned(((8'had) ?
                                  (8'h9c) : reg3610)) ?
                              $unsigned((reg3673 ?
                                  forvar3623 : forvar3609)) : ($signed(reg3677) > $signed(reg3721))));
                      reg3731 <= (forvar3626[(1'h0):(1'h0)] ?
                          (~^((reg3696 ~^ forvar3646) ?
                              $unsigned(forvar3645) : forvar3619)) : reg3724[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg3728 <= $unsigned((reg3709[(4'h9):(1'h0)] ~^ $signed($unsigned(reg3650))));
                      reg3729 <= {reg3593[(3'h6):(1'h0)]};
                    end
                  if ($unsigned(forvar3699[(2'h3):(1'h0)]))
                    begin
                      reg3732 <= $signed(forvar3558[(4'ha):(3'h5)]);
                    end
                  else
                    begin
                      reg3732 <= $signed((~^{reg3663}));
                      reg3733 <= (&(((reg3668 ? reg3654 : reg3712) ?
                              (forvar3607 ?
                                  reg3596 : (8'ha1)) : $signed(reg3569)) ?
                          $signed((~&forvar3656)) : (!(reg3693 | (8'ha4)))));
                    end
                  for (forvar3734 = (1'h0); (forvar3734 < (1'h0)); forvar3734 = (forvar3734 + (1'h1)))
                    begin
                      reg3735 <= ((((reg3701 >> (8'haf)) == {reg3660}) >>> {$unsigned(reg3568)}) > reg3658[(3'h5):(3'h5)]);
                      reg3736 <= (&forvar3734[(2'h2):(1'h1)]);
                      reg3737 <= {$signed({(^~reg3656)})};
                      reg3738 <= $signed({((wire3542 >> reg3646) + reg3620[(3'h4):(2'h2)])});
                    end
                end
              else
                begin
                  if ($unsigned($unsigned(({forvar3573} ?
                      {(8'ha6)} : $signed(forvar3734)))))
                    begin
                      reg3728 <= $signed(((~&{wire3543}) - (8'h9e)));
                      reg3729 <= reg3718[(1'h0):(1'h0)];
                      reg3730 <= $signed(((8'h9f) ?
                          $unsigned($unsigned(forvar3722)) : ((8'haf) ^~ (~^reg3672))));
                    end
                  else
                    begin
                      reg3728 <= reg3638;
                      reg3729 <= $signed(($unsigned(reg3545[(4'h8):(3'h4)]) && forvar3719[(2'h2):(1'h0)]));
                      reg3730 <= reg3663[(2'h3):(2'h2)];
                      reg3731 <= {$unsigned($signed($signed(reg3663)))};
                    end
                  reg3732 <= reg3574;
                  if (((reg3718 ?
                      reg3614[(1'h0):(1'h0)] : (~^(~&reg3732))) ~^ $signed(reg3569)))
                    begin
                      reg3733 <= ($signed($signed($unsigned(forvar3641))) ?
                          ((&{(8'hae)}) || ($signed(forvar3558) ?
                              $signed(reg3668) : $unsigned(reg3676))) : (((8'ha5) ^~ reg3582[(4'ha):(3'h4)]) ?
                              reg3732[(1'h0):(1'h0)] : $unsigned($unsigned(reg3569))));
                      reg3734 <= (((reg3592 >> forvar3593) ?
                          reg3622[(3'h7):(1'h0)] : $signed((reg3633 > forvar3552))) - (^reg3691[(3'h4):(1'h0)]));
                      reg3735 <= ($signed(((reg3649 ? forvar3682 : reg3673) ?
                              (forvar3601 & reg3630) : reg3708[(3'h6):(2'h2)])) ?
                          {$unsigned($signed(reg3707))} : (forvar3636 ?
                              reg3595[(1'h1):(1'h0)] : (reg3603[(5'h10):(3'h4)] ?
                                  ((8'ha6) ?
                                      forvar3710 : (8'h9c)) : (reg3629 < forvar3567))));
                      reg3736 <= ($signed(reg3637[(1'h0):(1'h0)]) ?
                          (^~$unsigned($signed(reg3624))) : forvar3560[(4'hd):(3'h6)]);
                    end
                  else
                    begin
                      reg3733 <= ($unsigned(forvar3615) ^ (($signed(forvar3544) ~^ $unsigned(reg3632)) ?
                          forvar3645 : (~&(forvar3626 ?
                              reg3564 : forvar3654))));
                    end
                end
            end
          for (forvar3739 = (1'h0); (forvar3739 < (2'h2)); forvar3739 = (forvar3739 + (1'h1)))
            begin
              if ($unsigned((&$unsigned($signed(reg3620)))))
                begin
                  for (forvar3740 = (1'h0); (forvar3740 < (2'h3)); forvar3740 = (forvar3740 + (1'h1)))
                    begin
                      reg3741 <= reg3653[(3'h5):(1'h0)];
                    end
                  if ((forvar3669[(1'h1):(1'h0)] ^~ ((^~(|forvar3669)) | ({(8'hb4)} ?
                      (reg3718 ? reg3546 : reg3611) : (reg3610 + (8'hb0))))))
                    begin
                      reg3742 <= $unsigned((((reg3687 | (8'h9e)) | forvar3672[(1'h0):(1'h0)]) ?
                          $unsigned($unsigned((8'hb0))) : (^~(8'ha5))));
                      reg3743 <= {$unsigned($signed((reg3714 << reg3728)))};
                    end
                  else
                    begin
                      reg3742 <= reg3614;
                    end
                end
              else
                begin
                  reg3740 <= (-(((reg3652 + forvar3544) ?
                          forvar3710 : forvar3636) ?
                      $unsigned($unsigned(reg3554)) : $signed((~&forvar3647))));
                  reg3741 <= forvar3654;
                  for (forvar3742 = (1'h0); (forvar3742 < (1'h1)); forvar3742 = (forvar3742 + (1'h1)))
                    begin
                      reg3743 <= (reg3592 ?
                          reg3723 : $signed(forvar3598[(2'h3):(1'h0)]));
                      reg3744 <= (8'hb4);
                    end
                end
              for (forvar3745 = (1'h0); (forvar3745 < (1'h0)); forvar3745 = (forvar3745 + (1'h1)))
                begin
                  if ($signed(({$unsigned(reg3617)} ?
                      (~|$unsigned(forvar3686)) : ((-reg3740) ?
                          $unsigned(forvar3706) : (forvar3647 ?
                              forvar3553 : forvar3547)))))
                    begin
                      reg3746 <= forvar3671[(4'ha):(2'h2)];
                      reg3747 <= forvar3676[(3'h7):(3'h5)];
                    end
                  else
                    begin
                      reg3746 <= ($unsigned($signed((reg3718 <<< (8'h9e)))) ?
                          (8'h9e) : reg3616[(2'h2):(2'h2)]);
                      reg3747 <= {{forvar3631}};
                    end
                  for (forvar3748 = (1'h0); (forvar3748 < (1'h1)); forvar3748 = (forvar3748 + (1'h1)))
                    begin
                      reg3749 <= ($signed(reg3671) && ((!((8'hb2) ?
                              forvar3660 : reg3660)) ?
                          ($signed(reg3663) ?
                              ((8'ha9) ~^ reg3658) : $unsigned(forvar3654)) : $signed(reg3670[(2'h2):(2'h2)])));
                      reg3750 <= (reg3651 >>> $unsigned($unsigned((+forvar3710))));
                      reg3751 <= reg3597;
                      reg3752 <= reg3747;
                    end
                end
              for (forvar3753 = (1'h0); (forvar3753 < (2'h2)); forvar3753 = (forvar3753 + (1'h1)))
                begin
                  for (forvar3754 = (1'h0); (forvar3754 < (2'h2)); forvar3754 = (forvar3754 + (1'h1)))
                    begin
                      reg3755 <= (!(~&{(reg3624 ~^ reg3590)}));
                      reg3756 <= reg3572[(4'hb):(3'h5)];
                      reg3757 <= $unsigned($signed((+forvar3615[(1'h0):(1'h0)])));
                    end
                  if (reg3640[(2'h2):(1'h0)])
                    begin
                      reg3758 <= {(reg3576 ?
                              reg3689 : ($signed(reg3568) ?
                                  (~^reg3695) : (forvar3740 && reg3749)))};
                      reg3759 <= (((~&{reg3665}) >>> $unsigned((8'h9c))) <= forvar3609);
                      reg3760 <= $unsigned((8'ha9));
                      reg3761 <= reg3670[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3758 <= {reg3746};
                    end
                  if (forvar3631)
                    begin
                      reg3762 <= $signed(reg3581[(1'h1):(1'h0)]);
                      reg3763 <= reg3568;
                      reg3764 <= (-reg3550);
                      reg3765 <= reg3639[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg3762 <= $unsigned(reg3659[(3'h5):(3'h4)]);
                    end
                end
            end
        end
    end
  assign wire3766 = {reg3594[(4'h8):(3'h5)]};
  assign wire3767 = (&reg3673);
  assign wire3768 = ((+$signed(reg3752)) << reg3583);
  module3769 modinst4731 (.wire3772(reg3689), .y(wire4730), .clk(clk), .wire3770(forvar3753), .wire3773(reg3600), .wire3771(reg3660));
  assign wire4732 = (((reg3684[(2'h2):(1'h1)] ?
                                $unsigned(reg3733) : (&reg3662)) ?
                            ($unsigned((8'ha6)) && $signed((8'hb5))) : $unsigned($signed(reg3557))) ?
                        reg3546[(3'h6):(3'h6)] : (forvar3607[(2'h2):(1'h1)] | reg3671));
  assign wire4733 = (~^{reg3688[(2'h2):(1'h1)]});
  always
    @(posedge clk) begin
      reg4734 <= ((8'hb6) && ($unsigned((reg3721 <= (8'hb2))) + ((~reg3559) ?
          reg3582 : (reg3724 ? forvar3734 : forvar3717))));
      if ({($signed((^reg3740)) * forvar3647)})
        begin
          for (forvar4735 = (1'h0); (forvar4735 < (2'h2)); forvar4735 = (forvar4735 + (1'h1)))
            begin
              for (forvar4736 = (1'h0); (forvar4736 < (1'h1)); forvar4736 = (forvar4736 + (1'h1)))
                begin
                  reg4737 <= $signed($unsigned({(forvar3636 ?
                          forvar3548 : reg3644)}));
                  for (forvar4738 = (1'h0); (forvar4738 < (2'h2)); forvar4738 = (forvar4738 + (1'h1)))
                    begin
                      reg4739 <= $signed(($signed(reg3683) + {forvar3656}));
                      reg4740 <= reg3562;
                      reg4741 <= $unsigned($unsigned({(reg3605 ?
                              reg3568 : forvar3719)}));
                      reg4742 <= forvar3578;
                    end
                  for (forvar4743 = (1'h0); (forvar4743 < (2'h2)); forvar4743 = (forvar4743 + (1'h1)))
                    begin
                      reg4744 <= $unsigned(($unsigned((reg3558 ?
                          reg4740 : forvar3697)) != (|$signed(reg3759))));
                    end
                end
              for (forvar4745 = (1'h0); (forvar4745 < (1'h0)); forvar4745 = (forvar4745 + (1'h1)))
                begin
                  for (forvar4746 = (1'h0); (forvar4746 < (2'h3)); forvar4746 = (forvar4746 + (1'h1)))
                    begin
                      reg4747 <= $unsigned((~&$signed(reg4742)));
                      reg4748 <= $signed((({forvar3553} ?
                          (~&reg3618) : ((8'haa) | wire3767)) && $signed((reg3645 ?
                          reg3660 : reg3605))));
                    end
                end
              if ((!reg3596))
                begin
                  for (forvar4749 = (1'h0); (forvar4749 < (2'h2)); forvar4749 = (forvar4749 + (1'h1)))
                    begin
                      reg4750 <= $signed($unsigned(forvar3660[(1'h0):(1'h0)]));
                      reg4751 <= (reg3557 ?
                          reg3749 : ({(reg3619 && forvar3656)} > reg3644));
                    end
                  reg4752 <= {((-(-reg4740)) ?
                          (reg3553[(3'h7):(1'h0)] >= (&forvar3671)) : ($signed(forvar3725) ?
                              $unsigned((8'hb3)) : (&reg3693)))};
                end
              else
                begin
                  if (reg4740)
                    begin
                      reg4749 <= {((~wire4733) ^~ forvar3609[(1'h0):(1'h0)])};
                      reg4750 <= (({reg3652[(1'h1):(1'h1)]} ?
                              $unsigned(reg3595) : reg3761) ?
                          forvar3549[(3'h4):(1'h1)] : forvar3734);
                      reg4751 <= ((8'hb1) == forvar3577);
                    end
                  else
                    begin
                      reg4749 <= ($signed(forvar3711[(4'h8):(4'h8)]) ^ ($unsigned({reg4749}) ?
                          ((~wire3768) < (!reg3662)) : (forvar3636 ?
                              (^reg3689) : (forvar3579 == reg3723))));
                      reg4750 <= $unsigned(reg3685);
                    end
                  reg4752 <= (reg3738[(2'h3):(2'h3)] == ((reg3556 << reg3572) | forvar3544));
                  for (forvar4753 = (1'h0); (forvar4753 < (2'h3)); forvar4753 = (forvar4753 + (1'h1)))
                    begin
                      reg4754 <= $unsigned($signed($signed($signed(forvar3706))));
                      reg4755 <= $signed(forvar3602[(4'hb):(4'h9)]);
                      reg4756 <= $signed($signed(reg4755[(2'h2):(1'h1)]));
                      reg4757 <= ((~(reg3570 ? $signed(forvar3657) : reg3627)) ?
                          (|{$unsigned((8'ha9))}) : reg3642);
                    end
                  for (forvar4758 = (1'h0); (forvar4758 < (1'h0)); forvar4758 = (forvar4758 + (1'h1)))
                    begin
                      reg4759 <= reg3562[(4'hd):(3'h6)];
                      reg4760 <= (reg3758[(1'h0):(1'h0)] + (~&reg3563));
                    end
                end
            end
          for (forvar4761 = (1'h0); (forvar4761 < (2'h3)); forvar4761 = (forvar4761 + (1'h1)))
            begin
              reg4762 <= (reg3741[(3'h5):(2'h2)] && ((reg3708 ?
                      reg3763 : (&forvar3722)) ?
                  (wire4733[(3'h6):(1'h0)] == (8'ha9)) : $signed($unsigned((8'hb2)))));
            end
          for (forvar4763 = (1'h0); (forvar4763 < (1'h1)); forvar4763 = (forvar4763 + (1'h1)))
            begin
              for (forvar4764 = (1'h0); (forvar4764 < (2'h3)); forvar4764 = (forvar4764 + (1'h1)))
                begin
                  for (forvar4765 = (1'h0); (forvar4765 < (2'h2)); forvar4765 = (forvar4765 + (1'h1)))
                    begin
                      reg4766 <= $signed($unsigned((^(reg3628 ?
                          reg3627 : (8'hab)))));
                      reg4767 <= (wire3540 ?
                          (reg3741 ?
                              (!$unsigned(forvar3682)) : $signed($signed(forvar4765))) : $unsigned((reg3741[(3'h4):(1'h1)] ?
                              (!(8'h9d)) : $unsigned(forvar3589))));
                      reg4768 <= ((((reg3646 | reg4762) ?
                              (reg3691 ?
                                  (8'hba) : forvar3547) : forvar3676[(3'h4):(1'h0)]) ?
                          (~^$unsigned(forvar3686)) : $unsigned({reg3597})) - $unsigned($unsigned($unsigned(reg3576))));
                      reg4769 <= {(~&((|reg3621) ^~ (reg3750 ?
                              reg3701 : reg3639)))};
                    end
                  for (forvar4770 = (1'h0); (forvar4770 < (1'h1)); forvar4770 = (forvar4770 + (1'h1)))
                    begin
                      reg4771 <= (~|reg3548[(4'h8):(2'h2)]);
                      reg4772 <= $unsigned(reg3593);
                      reg4773 <= $signed(reg3724[(2'h2):(2'h2)]);
                      reg4774 <= $signed($signed(forvar3593[(4'hd):(4'h8)]));
                    end
                  reg4775 <= $signed($unsigned(((forvar3547 ~^ forvar3706) <<< (reg3597 ?
                      reg3653 : forvar3681))));
                  if ($unsigned($signed(forvar4758[(3'h6):(1'h0)])))
                    begin
                      reg4776 <= $unsigned({reg3561});
                      reg4777 <= $signed((8'hba));
                    end
                  else
                    begin
                      reg4776 <= reg3555[(1'h0):(1'h0)];
                      reg4777 <= $signed((-((reg3659 ?
                          forvar3710 : reg3639) > $unsigned((8'ha6)))));
                      reg4778 <= $unsigned($unsigned(reg4744[(2'h2):(1'h0)]));
                    end
                end
            end
        end
      else
        begin
          for (forvar4735 = (1'h0); (forvar4735 < (2'h3)); forvar4735 = (forvar4735 + (1'h1)))
            begin
              if ((^(!$unsigned((reg3741 >= forvar3553)))))
                begin
                  reg4736 <= reg3594[(3'h6):(3'h5)];
                end
              else
                begin
                  if (reg3642)
                    begin
                      reg4736 <= $unsigned($unsigned(($signed(reg3735) * $signed(reg3743))));
                      reg4737 <= {$unsigned((forvar4745[(2'h2):(1'h1)] ?
                              (reg3737 ?
                                  forvar4770 : reg3585) : (-forvar3544)))};
                    end
                  else
                    begin
                      reg4736 <= reg3544;
                      reg4737 <= $signed(reg3638[(2'h2):(2'h2)]);
                      reg4738 <= ((((!reg3662) ?
                              {reg3744} : $unsigned(forvar3577)) ?
                          $signed((!forvar3631)) : forvar4749[(2'h2):(1'h1)]) >> (!$unsigned((reg4774 ?
                          forvar3710 : forvar3672))));
                      reg4739 <= reg3645[(2'h2):(1'h0)];
                    end
                  if (reg3617[(3'h6):(3'h5)])
                    begin
                      reg4740 <= reg3632[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg4740 <= $unsigned((+((reg3705 ?
                          forvar3655 : (8'ha5)) <<< $unsigned(reg3738))));
                      reg4741 <= $unsigned($unsigned(reg4773[(4'hc):(4'hb)]));
                      reg4742 <= $unsigned((!forvar3697));
                      reg4743 <= ((reg3689[(2'h3):(1'h0)] * (~|$signed(reg3556))) * forvar3598);
                    end
                end
              if (((^(~|reg4742[(3'h5):(1'h0)])) ?
                  $signed((^forvar3706[(2'h2):(1'h0)])) : reg3634[(4'h8):(1'h1)]))
                begin
                  if ($unsigned((^~{forvar3641[(3'h6):(3'h4)]})))
                    begin
                      reg4744 <= reg3742;
                      reg4745 <= $signed(forvar3682);
                      reg4746 <= reg3676[(4'h8):(3'h7)];
                      reg4747 <= (reg3645[(1'h1):(1'h1)] || forvar4745);
                    end
                  else
                    begin
                      reg4744 <= $signed((~$unsigned((+reg3595))));
                    end
                  if (reg3595)
                    begin
                      reg4748 <= (8'haa);
                      reg4749 <= ((reg3610 && $signed((forvar3672 || reg3737))) ?
                          (reg3627[(2'h3):(1'h0)] ?
                              (((8'ha1) ? forvar3711 : forvar3698) ?
                                  $unsigned(reg4750) : $unsigned((8'h9c))) : reg3550) : $unsigned(reg3740));
                    end
                  else
                    begin
                      reg4748 <= ((((reg4736 - reg3727) ^~ $unsigned(forvar4758)) >>> (reg3693[(1'h1):(1'h0)] ?
                          $signed(reg3564) : (|reg3594))) > (((~|forvar3742) < (^~(8'hab))) ?
                          $signed($unsigned(forvar3623)) : {reg3625[(4'hc):(3'h6)]}));
                    end
                  for (forvar4750 = (1'h0); (forvar4750 < (2'h2)); forvar4750 = (forvar4750 + (1'h1)))
                    begin
                      reg4751 <= (reg4774 ^ $signed(forvar3646[(3'h6):(2'h2)]));
                    end
                end
              else
                begin
                  reg4744 <= reg3691;
                  reg4745 <= ($signed(((forvar3544 <= wire3766) ?
                      ((8'ha0) ?
                          reg3549 : (8'ha3)) : $signed((8'haa)))) & $signed($unsigned($unsigned(reg4745))));
                  reg4746 <= $signed((reg3666 ?
                      $unsigned((8'hb1)) : forvar3754));
                end
              for (forvar4752 = (1'h0); (forvar4752 < (1'h0)); forvar4752 = (forvar4752 + (1'h1)))
                begin
                  for (forvar4753 = (1'h0); (forvar4753 < (1'h1)); forvar4753 = (forvar4753 + (1'h1)))
                    begin
                      reg4754 <= reg3736[(1'h1):(1'h0)];
                      reg4755 <= $signed($unsigned(wire3542));
                    end
                  if ({({$signed(reg3723)} ?
                          $unsigned($unsigned(forvar4765)) : (+(!reg4734)))})
                    begin
                      reg4756 <= reg3741;
                    end
                  else
                    begin
                      reg4756 <= (~|(!(reg3760 ?
                          reg3595[(2'h2):(1'h0)] : ((8'ha8) >> (8'hb1)))));
                    end
                  if (forvar3552[(1'h0):(1'h0)])
                    begin
                      reg4757 <= ((reg4747 ?
                          $signed(reg4769) : forvar4736) ^~ ((wire3543[(4'hd):(4'ha)] < reg4767) ?
                          reg3617[(4'h8):(2'h2)] : (8'hb4)));
                      reg4758 <= (($unsigned((reg3684 ?
                              reg3723 : reg3731)) * (!(reg3720 ?
                              wire4732 : reg3659))) ?
                          (^~($signed(reg3691) - (reg3662 && reg3732))) : forvar4749[(4'h9):(3'h6)]);
                      reg4759 <= $unsigned(wire3540);
                    end
                  else
                    begin
                      reg4757 <= reg3727;
                    end
                  for (forvar4760 = (1'h0); (forvar4760 < (1'h0)); forvar4760 = (forvar4760 + (1'h1)))
                    begin
                      reg4761 <= $unsigned($unsigned({$signed((8'hab))}));
                      reg4762 <= (-{(forvar4735 >> (reg3675 ?
                              (8'h9d) : (8'hb1)))});
                    end
                end
            end
          if ($unsigned(reg4758[(4'h9):(2'h2)]))
            begin
              reg4763 <= (|(8'hb8));
            end
          else
            begin
              for (forvar4763 = (1'h0); (forvar4763 < (2'h2)); forvar4763 = (forvar4763 + (1'h1)))
                begin
                  if ($unsigned((!($unsigned(forvar3601) > $signed(reg3675)))))
                    begin
                      reg4764 <= forvar3636;
                    end
                  else
                    begin
                      reg4764 <= (|(|$unsigned($signed(reg3615))));
                    end
                  for (forvar4765 = (1'h0); (forvar4765 < (1'h0)); forvar4765 = (forvar4765 + (1'h1)))
                    begin
                      reg4766 <= ((8'ha4) ?
                          (forvar3626[(2'h2):(1'h1)] ?
                              reg3594 : $unsigned(forvar4752[(1'h0):(1'h0)])) : (-$signed($signed(reg3627))));
                      reg4767 <= (reg3649[(3'h7):(1'h0)] ?
                          {$unsigned($signed(reg4777))} : $unsigned((forvar3734[(5'h10):(3'h6)] ?
                              reg3572[(4'h8):(3'h5)] : {reg3735})));
                      reg4768 <= forvar3698;
                      reg4769 <= ($unsigned($unsigned(reg3587)) << {(^~$unsigned(reg3628))});
                    end
                  for (forvar4770 = (1'h0); (forvar4770 < (2'h3)); forvar4770 = (forvar4770 + (1'h1)))
                    begin
                      reg4771 <= ($unsigned($unsigned(reg4752)) || $signed((|(~&forvar3669))));
                    end
                  if ($unsigned(forvar3734[(4'h9):(1'h0)]))
                    begin
                      reg4772 <= ((+(reg3632[(1'h0):(1'h0)] ^ (reg3730 <<< reg3756))) + $signed(reg3667[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg4772 <= $signed($signed(reg3734[(1'h0):(1'h0)]));
                    end
                end
              for (forvar4773 = (1'h0); (forvar4773 < (2'h3)); forvar4773 = (forvar4773 + (1'h1)))
                begin
                  if ({(!(!$unsigned((8'hb8))))})
                    begin
                      reg4774 <= $signed(($unsigned($unsigned(reg4771)) ^ (((8'ha0) >> reg4747) ?
                          forvar3547[(4'h8):(4'h8)] : $unsigned(reg3600))));
                      reg4775 <= reg3587[(4'h8):(2'h3)];
                      reg4776 <= ((((!forvar3613) > (-(8'ha0))) > $unsigned(forvar4752[(2'h3):(1'h1)])) >= (reg3763 ?
                          $unsigned($unsigned(wire3540)) : $unsigned({reg3563})));
                    end
                  else
                    begin
                      reg4774 <= reg3736[(2'h3):(1'h0)];
                      reg4775 <= (forvar3739[(3'h4):(1'h1)] ?
                          (^~forvar3601[(1'h1):(1'h1)]) : $unsigned(($signed(forvar3559) + forvar3566[(3'h6):(3'h5)])));
                      reg4776 <= {{$unsigned((forvar3739 >= forvar4745))}};
                    end
                  for (forvar4777 = (1'h0); (forvar4777 < (1'h1)); forvar4777 = (forvar4777 + (1'h1)))
                    begin
                      reg4778 <= (reg3672[(1'h1):(1'h0)] >> (~&($signed(reg3736) + reg4747[(3'h7):(3'h5)])));
                      reg4779 <= $unsigned({(~|{reg3586})});
                      reg4780 <= forvar3548;
                      reg4781 <= reg3688;
                    end
                end
              for (forvar4782 = (1'h0); (forvar4782 < (1'h1)); forvar4782 = (forvar4782 + (1'h1)))
                begin
                  for (forvar4783 = (1'h0); (forvar4783 < (2'h3)); forvar4783 = (forvar4783 + (1'h1)))
                    begin
                      reg4784 <= (^forvar3706);
                    end
                  if (forvar3626[(1'h1):(1'h0)])
                    begin
                      reg4785 <= {(-forvar3748)};
                      reg4786 <= $unsigned(reg3761[(1'h1):(1'h1)]);
                      reg4787 <= ((8'hb1) << $signed((reg3668 - $signed(reg3662))));
                      reg4788 <= {$unsigned($signed((forvar3660 <<< reg3752)))};
                    end
                  else
                    begin
                      reg4785 <= reg3653;
                      reg4786 <= reg3621;
                      reg4787 <= reg3605[(4'ha):(1'h0)];
                    end
                  if ((+$signed(((-reg4771) ? (^reg3694) : $signed((8'hb7))))))
                    begin
                      reg4789 <= {$signed(reg3595[(3'h7):(3'h5)])};
                      reg4790 <= ((&reg3763) ~^ (-(|forvar3578)));
                      reg4791 <= {reg4740};
                      reg4792 <= (({{forvar3698}} && (8'h9e)) ?
                          (~(8'ha0)) : (~|$signed((reg4740 >> forvar3681))));
                    end
                  else
                    begin
                      reg4789 <= {((~|(forvar3669 >> reg4750)) && {$unsigned(forvar4770)})};
                      reg4790 <= (reg4768[(3'h7):(1'h0)] ?
                          forvar3699 : (|$unsigned(((8'ha4) ?
                              reg4771 : forvar3567))));
                    end
                end
            end
        end
    end
  assign wire4793 = $signed(reg4738[(1'h1):(1'h0)]);
  assign wire4794 = $signed(reg4763[(3'h6):(1'h1)]);
  always
    @(posedge clk) begin
      if ((reg4759 ?
          {($unsigned(forvar4750) ?
                  reg3644 : reg3736[(1'h1):(1'h1)])} : ($signed(reg3658) ?
              $signed(reg3549) : $signed($signed(forvar4736)))))
        begin
          for (forvar4795 = (1'h0); (forvar4795 < (2'h3)); forvar4795 = (forvar4795 + (1'h1)))
            begin
              reg4796 <= reg3637;
              for (forvar4797 = (1'h0); (forvar4797 < (2'h2)); forvar4797 = (forvar4797 + (1'h1)))
                begin
                  if (reg3591)
                    begin
                      reg4798 <= $signed($signed((((8'hae) && forvar4797) ?
                          reg3629 : (reg4740 >> reg3690))));
                      reg4799 <= $signed((reg3646[(2'h2):(1'h1)] >= (+$signed(reg3720))));
                      reg4800 <= wire3540[(3'h7):(1'h1)];
                      reg4801 <= $signed($signed((reg3572[(4'hf):(3'h6)] ?
                          forvar4753 : ((8'ha8) ? reg3655 : wire4733))));
                    end
                  else
                    begin
                      reg4798 <= $unsigned((|(reg3611[(1'h0):(1'h0)] ?
                          ((8'haf) ^~ reg4779) : (-reg3604))));
                      reg4799 <= (((((8'hb6) ? reg3703 : (8'hb5)) ?
                              (reg3558 < forvar3655) : $unsigned(reg3701)) - (!$signed(forvar3742))) ?
                          reg3742[(3'h4):(1'h0)] : ($signed({(8'hb6)}) && {reg3546}));
                      reg4800 <= ((!(8'hb9)) ?
                          (^(reg3553[(2'h2):(1'h0)] << (forvar3672 ?
                              (8'ha1) : reg3721))) : ((reg3743 && reg3642[(4'ha):(3'h5)]) - $signed($signed(reg3701))));
                      reg4801 <= (!(reg4790[(1'h0):(1'h0)] || forvar3740[(2'h3):(2'h3)]));
                    end
                  if ((~{(~$unsigned(reg3622))}))
                    begin
                      reg4802 <= $unsigned(reg4785[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg4802 <= reg3707[(2'h2):(1'h1)];
                    end
                  for (forvar4803 = (1'h0); (forvar4803 < (1'h1)); forvar4803 = (forvar4803 + (1'h1)))
                    begin
                      reg4804 <= {(forvar3623 ?
                              reg4758 : $unsigned((reg4790 ?
                                  reg3627 : reg4772)))};
                    end
                  if ($unsigned({reg4785}))
                    begin
                      reg4805 <= (reg3700 ?
                          {(+$unsigned(forvar3681))} : (^~(~&$signed(forvar3682))));
                      reg4806 <= ((8'haa) ?
                          (8'ha8) : $unsigned((reg3646 >> (~&reg3744))));
                      reg4807 <= forvar4736[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg4805 <= (({$signed((8'hb0))} << $signed($unsigned(reg3583))) ?
                          reg4756 : (~&((~|reg3696) >>> forvar3589[(4'hc):(4'ha)])));
                      reg4806 <= ({$unsigned($signed(reg4762))} ?
                          $signed(reg4756) : (((reg3557 < reg4743) ~^ forvar3669) <<< $signed((reg3683 == (8'h9d)))));
                      reg4807 <= $unsigned(reg3716[(3'h4):(1'h1)]);
                      reg4808 <= (~^(+reg4764));
                    end
                end
              for (forvar4809 = (1'h0); (forvar4809 < (1'h1)); forvar4809 = (forvar4809 + (1'h1)))
                begin
                  for (forvar4810 = (1'h0); (forvar4810 < (2'h3)); forvar4810 = (forvar4810 + (1'h1)))
                    begin
                      reg4811 <= {reg3572[(2'h3):(2'h2)]};
                      reg4812 <= $signed(($signed(reg4754) ?
                          $unsigned($signed(forvar4770)) : {(~&reg4805)}));
                      reg4813 <= $signed(reg3572[(4'hf):(1'h0)]);
                    end
                end
              for (forvar4814 = (1'h0); (forvar4814 < (2'h2)); forvar4814 = (forvar4814 + (1'h1)))
                begin
                  for (forvar4815 = (1'h0); (forvar4815 < (1'h1)); forvar4815 = (forvar4815 + (1'h1)))
                    begin
                      reg4816 <= reg4792;
                      reg4817 <= $unsigned(((~&(~^reg3709)) <<< reg3571));
                      reg4818 <= {reg3660[(1'h1):(1'h1)]};
                    end
                  reg4819 <= {$unsigned($signed((reg4744 > reg4751)))};
                  if ((+{$unsigned(reg3735[(2'h3):(1'h0)])}))
                    begin
                      reg4820 <= (8'hb3);
                    end
                  else
                    begin
                      reg4820 <= $signed(forvar3686);
                      reg4821 <= (($signed({(8'ha8)}) && ((~^reg4756) ?
                              $signed(reg4756) : (reg3635 | reg3568))) ?
                          forvar3660[(2'h2):(1'h1)] : reg3726[(1'h1):(1'h1)]);
                    end
                end
            end
          if (forvar4803)
            begin
              if ((reg3688 <<< reg4773[(3'h6):(1'h0)]))
                begin
                  reg4822 <= $unsigned($signed({(reg3548 || reg3750)}));
                end
              else
                begin
                  if ((reg3742 ?
                      (reg3557 == reg3720[(1'h1):(1'h1)]) : reg4796[(1'h0):(1'h0)]))
                    begin
                      reg4822 <= (wire3768[(2'h2):(1'h1)] ?
                          $signed(wire3766) : (reg3599[(3'h7):(3'h7)] ?
                              $unsigned($signed(reg4749)) : (reg3680[(3'h4):(3'h4)] <<< reg3571)));
                      reg4823 <= forvar3602[(3'h4):(2'h3)];
                      reg4824 <= $signed((~&(reg3650[(2'h3):(2'h3)] | $unsigned(reg3545))));
                      reg4825 <= ($signed($signed($signed((8'h9e)))) ?
                          ((8'hae) ?
                              reg3634[(4'hc):(1'h1)] : $unsigned(reg3658[(3'h6):(3'h5)])) : ((reg3734 << reg3563[(2'h2):(1'h1)]) ?
                              forvar3715[(1'h1):(1'h0)] : $signed({reg3685})));
                    end
                  else
                    begin
                      reg4822 <= {reg3611};
                    end
                end
              if ((8'hb6))
                begin
                  reg4826 <= reg3709[(4'h8):(3'h4)];
                end
              else
                begin
                  if ({{$unsigned($signed(reg4777))}})
                    begin
                      reg4826 <= {($unsigned((8'hba)) <= ((reg3587 ?
                              forvar3697 : reg4796) - (reg4819 && reg3691)))};
                      reg4827 <= reg4737;
                    end
                  else
                    begin
                      reg4826 <= (reg3634 ? reg3713[(1'h1):(1'h0)] : reg3734);
                    end
                  reg4828 <= (($signed($signed(reg4741)) ?
                      ((forvar4782 ? reg3553 : forvar4770) ?
                          (forvar4753 & reg3723) : reg4787[(3'h4):(2'h2)]) : reg3670) <= ((^((8'hb3) ?
                          wire3766 : reg4800)) ?
                      ({reg4775} ? {reg4788} : wire3540) : ((^~forvar3646) ?
                          $unsigned(reg3683) : (8'hae))));
                end
              for (forvar4829 = (1'h0); (forvar4829 < (1'h0)); forvar4829 = (forvar4829 + (1'h1)))
                begin
                  if ($signed((&(reg3615 > ((8'hb5) ^~ forvar4809)))))
                    begin
                      reg4830 <= {(~^$signed($signed(reg3759)))};
                      reg4831 <= forvar3660;
                    end
                  else
                    begin
                      reg4830 <= (^reg3689[(4'h8):(3'h4)]);
                      reg4831 <= $signed({$signed(reg3687[(2'h2):(1'h0)])});
                      reg4832 <= $signed(reg4768);
                      reg4833 <= $unsigned((8'hb4));
                    end
                  for (forvar4834 = (1'h0); (forvar4834 < (1'h1)); forvar4834 = (forvar4834 + (1'h1)))
                    begin
                      reg4835 <= $unsigned($unsigned(reg3763[(2'h3):(1'h0)]));
                      reg4836 <= reg3687;
                      reg4837 <= $unsigned(((reg3696[(3'h4):(1'h1)] || reg4763) ?
                          $unsigned((reg4737 ?
                              reg3709 : forvar4738)) : reg4781));
                    end
                  reg4838 <= (({{forvar3589}} ?
                          $unsigned(forvar3613) : (reg3679[(3'h7):(3'h5)] <<< (~^reg4816))) ?
                      $unsigned(reg3618) : ((|$unsigned(reg4734)) & $unsigned(reg3648[(2'h2):(1'h1)])));
                end
              if ($unsigned($signed($unsigned($signed((8'hb7))))))
                begin
                  if (((~(reg3705 ? reg3635 : reg3720[(1'h1):(1'h1)])) ?
                      $signed($signed(reg3674)) : $unsigned($unsigned($signed((8'ha5))))))
                    begin
                      reg4839 <= forvar3655[(4'h9):(3'h6)];
                    end
                  else
                    begin
                      reg4839 <= {(8'hb3)};
                      reg4840 <= (~reg3736[(2'h3):(1'h0)]);
                      reg4841 <= $signed(((reg3569 ?
                          {reg4804} : ((8'hb5) == reg4737)) * {{reg4840}}));
                    end
                  for (forvar4842 = (1'h0); (forvar4842 < (1'h0)); forvar4842 = (forvar4842 + (1'h1)))
                    begin
                      reg4843 <= $signed((reg4804[(2'h2):(1'h0)] << (+(reg3656 ?
                          reg4800 : reg3690))));
                      reg4844 <= (8'h9d);
                      reg4845 <= $signed({reg3552[(2'h3):(2'h2)]});
                      reg4846 <= {(-reg4768)};
                    end
                  reg4847 <= {$unsigned(($unsigned(reg3590) ?
                          (reg3629 ?
                              forvar4761 : forvar3545) : $signed(forvar3698)))};
                end
              else
                begin
                  if ((&$signed($unsigned(forvar3552[(1'h0):(1'h0)]))))
                    begin
                      reg4839 <= (~^forvar3623);
                    end
                  else
                    begin
                      reg4839 <= (reg3651 < reg3610);
                      reg4840 <= forvar3615[(3'h5):(2'h3)];
                      reg4841 <= reg4763[(1'h0):(1'h0)];
                      reg4842 <= (!reg4819);
                    end
                  for (forvar4843 = (1'h0); (forvar4843 < (1'h1)); forvar4843 = (forvar4843 + (1'h1)))
                    begin
                      reg4844 <= (((&reg3746[(1'h1):(1'h1)]) && (reg3617 ~^ reg3683)) ?
                          $unsigned((reg3581[(1'h0):(1'h0)] <<< {reg3763})) : $unsigned(reg3657));
                      reg4845 <= reg3738[(2'h2):(1'h0)];
                    end
                end
            end
          else
            begin
              if ($signed(reg4796))
                begin
                  for (forvar4822 = (1'h0); (forvar4822 < (1'h1)); forvar4822 = (forvar4822 + (1'h1)))
                    begin
                      reg4823 <= ($unsigned((reg3581 >>> $unsigned(reg4767))) ?
                          {(+reg4781[(1'h1):(1'h0)])} : reg4774[(4'hd):(2'h2)]);
                      reg4824 <= $unsigned(reg4825[(1'h1):(1'h0)]);
                    end
                  for (forvar4825 = (1'h0); (forvar4825 < (2'h3)); forvar4825 = (forvar4825 + (1'h1)))
                    begin
                      reg4826 <= ((8'hae) ?
                          (-reg4843) : {reg3634[(4'hc):(4'hc)]});
                      reg4827 <= reg3737;
                      reg4828 <= reg3564[(2'h2):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar4822 = (1'h0); (forvar4822 < (1'h1)); forvar4822 = (forvar4822 + (1'h1)))
                    begin
                      reg4823 <= $unsigned($signed(forvar3593));
                      reg4824 <= $signed(reg3765[(3'h5):(2'h3)]);
                      reg4825 <= (^~reg3760);
                    end
                  for (forvar4826 = (1'h0); (forvar4826 < (1'h0)); forvar4826 = (forvar4826 + (1'h1)))
                    begin
                      reg4827 <= (reg4749[(4'h8):(4'h8)] ?
                          reg4773[(4'h9):(1'h1)] : (forvar3647[(4'h8):(3'h4)] && $signed(reg3742[(1'h0):(1'h0)])));
                      reg4828 <= ((8'haf) ?
                          $signed(reg4752) : forvar4765[(3'h6):(3'h4)]);
                      reg4829 <= reg3608[(3'h7):(2'h2)];
                      reg4830 <= reg4801[(2'h3):(1'h1)];
                    end
                  reg4831 <= $signed((|$unsigned(forvar4842[(2'h3):(1'h1)])));
                  if ((8'h9e))
                    begin
                      reg4832 <= (8'h9c);
                      reg4833 <= {reg3685};
                      reg4834 <= (~^$unsigned({((8'hb8) ?
                              (8'ha0) : forvar3549)}));
                    end
                  else
                    begin
                      reg4832 <= ($unsigned((|(reg3679 ~^ reg3594))) >>> (forvar3636[(3'h4):(3'h4)] ?
                          ((~^reg3586) <<< {wire4733}) : {forvar4825[(3'h5):(2'h3)]}));
                      reg4833 <= $unsigned($unsigned(($signed((8'ha6)) ?
                          ((8'h9f) <<< reg3721) : $signed(reg3615))));
                      reg4834 <= reg3550[(2'h2):(2'h2)];
                    end
                end
            end
        end
      else
        begin
          for (forvar4795 = (1'h0); (forvar4795 < (1'h1)); forvar4795 = (forvar4795 + (1'h1)))
            begin
              if (($signed((reg4754 ? reg3618[(1'h1):(1'h0)] : {reg3628})) ?
                  $unsigned((reg3730 ?
                      (forvar4735 * wire3540) : reg3667[(4'hb):(3'h7)])) : (|($signed(reg3639) ?
                      forvar4834[(1'h0):(1'h0)] : (reg3759 >>> (8'haa))))))
                begin
                  for (forvar4796 = (1'h0); (forvar4796 < (1'h0)); forvar4796 = (forvar4796 + (1'h1)))
                    begin
                      reg4797 <= ((((reg3705 <= reg4792) != $unsigned(reg3683)) ?
                          reg3677[(2'h3):(2'h2)] : (forvar3573[(2'h3):(2'h2)] << $signed((8'ha1)))) == (reg3624[(3'h4):(2'h2)] ?
                          $signed($signed(reg3759)) : $signed((reg3594 < (8'h9d)))));
                      reg4798 <= forvar3656[(2'h3):(2'h3)];
                      reg4799 <= ($signed((~^(reg3716 ?
                          (8'hab) : reg4843))) && (forvar4761[(2'h2):(2'h2)] < (reg4813[(3'h4):(1'h1)] ?
                          reg3684[(3'h4):(2'h3)] : ((8'hb7) >>> reg3553))));
                      reg4800 <= reg3572[(4'hd):(4'h8)];
                    end
                  for (forvar4801 = (1'h0); (forvar4801 < (1'h1)); forvar4801 = (forvar4801 + (1'h1)))
                    begin
                      reg4802 <= reg4791[(2'h2):(2'h2)];
                      reg4803 <= $signed(($signed(forvar3676[(3'h7):(2'h2)]) ?
                          reg3568[(4'ha):(3'h4)] : (!$unsigned((8'ha8)))));
                    end
                  if ((~^$unsigned($unsigned({forvar3607}))))
                    begin
                      reg4804 <= ({forvar3725} != reg4740[(1'h1):(1'h0)]);
                      reg4805 <= $unsigned($signed(((-reg3727) ?
                          reg3705[(2'h3):(2'h3)] : reg3554[(4'hb):(2'h2)])));
                      reg4806 <= $signed(reg3628);
                    end
                  else
                    begin
                      reg4804 <= (~|(^(reg3724[(3'h4):(2'h3)] ?
                          reg3628[(1'h0):(1'h0)] : ((8'hb3) ?
                              forvar3681 : (8'ha4)))));
                      reg4805 <= ((reg4791 ~^ $unsigned((~&reg3637))) ^~ reg3703[(3'h5):(3'h5)]);
                      reg4806 <= (~^((&reg4805[(1'h0):(1'h0)]) ?
                          ((-forvar3682) ^ (reg3629 * (8'hb1))) : {(forvar3706 ?
                                  reg3622 : forvar4796)}));
                      reg4807 <= $signed((~&(-(!forvar3598))));
                    end
                end
              else
                begin
                  for (forvar4796 = (1'h0); (forvar4796 < (1'h1)); forvar4796 = (forvar4796 + (1'h1)))
                    begin
                      reg4797 <= (-((&(forvar3559 ?
                          reg3553 : reg3558)) << $unsigned((wire3543 ?
                          forvar3623 : (8'had)))));
                    end
                  for (forvar4798 = (1'h0); (forvar4798 < (2'h2)); forvar4798 = (forvar4798 + (1'h1)))
                    begin
                      reg4799 <= {reg3764[(3'h7):(3'h4)]};
                      reg4800 <= (reg3652[(1'h1):(1'h1)] * (!{$unsigned(reg4791)}));
                      reg4801 <= (reg4787[(4'h9):(1'h0)] ?
                          (^~reg4830) : $unsigned((8'hae)));
                    end
                  for (forvar4802 = (1'h0); (forvar4802 < (2'h3)); forvar4802 = (forvar4802 + (1'h1)))
                    begin
                      reg4803 <= $signed((8'ha2));
                    end
                end
              for (forvar4808 = (1'h0); (forvar4808 < (2'h2)); forvar4808 = (forvar4808 + (1'h1)))
                begin
                  for (forvar4809 = (1'h0); (forvar4809 < (2'h2)); forvar4809 = (forvar4809 + (1'h1)))
                    begin
                      reg4810 <= {reg4834};
                      reg4811 <= reg3645[(3'h4):(1'h0)];
                      reg4812 <= forvar3656;
                    end
                end
              for (forvar4813 = (1'h0); (forvar4813 < (2'h2)); forvar4813 = (forvar4813 + (1'h1)))
                begin
                  reg4814 <= $unsigned(((~{reg3737}) ?
                      ($signed(reg4767) ^~ (reg4768 ?
                          forvar3567 : reg4748)) : forvar3573[(3'h5):(2'h3)]));
                  for (forvar4815 = (1'h0); (forvar4815 < (2'h3)); forvar4815 = (forvar4815 + (1'h1)))
                    begin
                      reg4816 <= $unsigned($unsigned($unsigned(((8'ha1) ~^ reg4737))));
                      reg4817 <= reg3740;
                      reg4818 <= (reg4766[(4'ha):(2'h3)] ?
                          forvar4809[(1'h0):(1'h0)] : reg3716[(3'h6):(1'h0)]);
                    end
                  for (forvar4819 = (1'h0); (forvar4819 < (1'h0)); forvar4819 = (forvar4819 + (1'h1)))
                    begin
                      reg4820 <= reg4842[(3'h6):(3'h4)];
                      reg4821 <= reg4758;
                      reg4822 <= $signed(({(forvar4834 <= forvar4843)} + reg4842[(4'hc):(2'h2)]));
                    end
                end
            end
          for (forvar4823 = (1'h0); (forvar4823 < (2'h2)); forvar4823 = (forvar4823 + (1'h1)))
            begin
              for (forvar4824 = (1'h0); (forvar4824 < (1'h0)); forvar4824 = (forvar4824 + (1'h1)))
                begin
                  for (forvar4825 = (1'h0); (forvar4825 < (2'h3)); forvar4825 = (forvar4825 + (1'h1)))
                    begin
                      reg4826 <= (forvar3619[(1'h0):(1'h0)] ?
                          (^~({reg3645} ?
                              $unsigned(reg3747) : {reg3548})) : (^~reg3546));
                      reg4827 <= $signed(({{reg3679}} >= (((8'hab) ^~ reg3652) ~^ (wire3766 ^~ forvar4842))));
                      reg4828 <= reg4798;
                      reg4829 <= (8'haa);
                    end
                  for (forvar4830 = (1'h0); (forvar4830 < (1'h0)); forvar4830 = (forvar4830 + (1'h1)))
                    begin
                      reg4831 <= (reg3746 ^ ($signed(reg4844[(4'hc):(3'h7)]) ?
                          ((^reg4841) <= reg3724) : $unsigned((|reg4747))));
                      reg4832 <= (($unsigned($unsigned(reg4768)) > reg3743[(4'h8):(3'h5)]) ?
                          ((&(reg3651 < reg3763)) == $unsigned(reg3657[(2'h3):(2'h2)])) : (reg3600[(2'h2):(1'h1)] >> reg3591));
                      reg4833 <= reg3733[(1'h0):(1'h0)];
                    end
                  for (forvar4834 = (1'h0); (forvar4834 < (1'h1)); forvar4834 = (forvar4834 + (1'h1)))
                    begin
                      reg4835 <= reg4817[(3'h4):(2'h2)];
                      reg4836 <= $signed({$signed(forvar4819[(4'h8):(1'h0)])});
                      reg4837 <= {reg3677[(3'h6):(2'h3)]};
                      reg4838 <= (~&($signed((reg3559 * reg3583)) | (~^reg3750)));
                    end
                end
              if ((forvar4736 == $signed(forvar3593)))
                begin
                  for (forvar4839 = (1'h0); (forvar4839 < (1'h1)); forvar4839 = (forvar4839 + (1'h1)))
                    begin
                      reg4840 <= ((^((~|reg4746) ?
                          (reg4756 << reg3677) : $signed(forvar3544))) * reg3576[(3'h6):(2'h2)]);
                      reg4841 <= {$signed({(reg3692 * forvar3686)})};
                    end
                  for (forvar4842 = (1'h0); (forvar4842 < (1'h1)); forvar4842 = (forvar4842 + (1'h1)))
                    begin
                      reg4843 <= forvar4842;
                    end
                  reg4844 <= ((^~(reg3606 < forvar3654)) ?
                      {$unsigned($unsigned(reg4827))} : $unsigned((((8'hb5) ?
                          reg4822 : reg4814) > reg3685[(4'h9):(3'h7)])));
                end
              else
                begin
                  reg4839 <= $unsigned(($unsigned($unsigned(reg3701)) ?
                      $unsigned(reg3705[(2'h2):(2'h2)]) : $signed((forvar3742 <<< forvar4753))));
                end
              reg4845 <= (forvar3753[(2'h3):(1'h1)] ^~ $signed($signed((&(8'h9e)))));
            end
        end
      for (forvar4848 = (1'h0); (forvar4848 < (1'h1)); forvar4848 = (forvar4848 + (1'h1)))
        begin
          reg4849 <= $unsigned(forvar3686[(2'h3):(1'h1)]);
          if (($signed({(~&reg3619)}) >>> {reg3761}))
            begin
              reg4850 <= $unsigned({$signed($signed(reg3675))});
            end
          else
            begin
              for (forvar4850 = (1'h0); (forvar4850 < (2'h2)); forvar4850 = (forvar4850 + (1'h1)))
                begin
                  reg4851 <= reg4819;
                  for (forvar4852 = (1'h0); (forvar4852 < (2'h3)); forvar4852 = (forvar4852 + (1'h1)))
                    begin
                      reg4853 <= reg4843[(3'h5):(2'h2)];
                      reg4854 <= ({$signed($unsigned((8'hb0)))} ?
                          $unsigned(reg4774) : (8'ha7));
                    end
                  for (forvar4855 = (1'h0); (forvar4855 < (1'h1)); forvar4855 = (forvar4855 + (1'h1)))
                    begin
                      reg4856 <= $signed($signed(reg3597));
                      reg4857 <= reg3645;
                      reg4858 <= ((&$signed(reg3624[(3'h4):(2'h3)])) >= reg3701);
                    end
                  if (reg3661[(4'h8):(2'h2)])
                    begin
                      reg4859 <= (~^reg4850);
                      reg4860 <= (({$unsigned(reg3676)} ~^ (forvar4802[(1'h1):(1'h0)] < (forvar3664 && reg4738))) == {forvar3566});
                      reg4861 <= $unsigned(($signed(reg4798) ?
                          (((8'ha2) ?
                              reg4844 : forvar3615) ^~ $signed(reg4763)) : reg3761));
                    end
                  else
                    begin
                      reg4859 <= (reg4837 || reg3727);
                      reg4860 <= reg3705;
                    end
                end
            end
          reg4862 <= (8'had);
          reg4863 <= reg3635;
        end
    end
  assign wire4864 = (~|reg4748[(4'ha):(2'h2)]);
  always
    @(posedge clk) begin
      for (forvar4865 = (1'h0); (forvar4865 < (1'h0)); forvar4865 = (forvar4865 + (1'h1)))
        begin
          for (forvar4866 = (1'h0); (forvar4866 < (1'h0)); forvar4866 = (forvar4866 + (1'h1)))
            begin
              if (reg3742[(3'h4):(1'h1)])
                begin
                  reg4867 <= (&$unsigned(reg3616));
                  for (forvar4868 = (1'h0); (forvar4868 < (2'h2)); forvar4868 = (forvar4868 + (1'h1)))
                    begin
                      reg4869 <= (reg3620 ? (~&(!$signed((8'ha2)))) : reg3707);
                    end
                  if (reg3738)
                    begin
                      reg4870 <= $unsigned($unsigned((~^$unsigned(reg4772))));
                    end
                  else
                    begin
                      reg4870 <= $unsigned((+((forvar3601 <<< wire4730) ?
                          ((8'had) ~^ forvar4868) : {(8'hb8)})));
                      reg4871 <= reg4811;
                    end
                end
              else
                begin
                  for (forvar4867 = (1'h0); (forvar4867 < (1'h0)); forvar4867 = (forvar4867 + (1'h1)))
                    begin
                      reg4868 <= reg4777[(4'h9):(1'h1)];
                    end
                  if ((-(^$unsigned($unsigned(forvar4823)))))
                    begin
                      reg4869 <= ($signed(reg3559) ?
                          (-reg3582[(1'h1):(1'h1)]) : (|$signed(reg4736[(3'h7):(3'h5)])));
                    end
                  else
                    begin
                      reg4869 <= (-(~(&(reg4822 ? reg4843 : (8'h9d)))));
                      reg4870 <= (forvar3579[(4'hd):(4'hc)] & reg3666);
                      reg4871 <= reg3755;
                      reg4872 <= ((^$signed((+(8'ha1)))) ?
                          reg3604 : reg3599[(2'h3):(2'h2)]);
                    end
                  if ($unsigned(forvar3753[(4'he):(4'h8)]))
                    begin
                      reg4873 <= (~(~$signed((~forvar3669))));
                      reg4874 <= (&$signed($unsigned((^~reg4828))));
                    end
                  else
                    begin
                      reg4873 <= reg3659[(3'h5):(1'h1)];
                      reg4874 <= $unsigned((~^reg3624[(2'h3):(1'h0)]));
                      reg4875 <= (~((^~reg3741) ? wire4793 : (8'ha1)));
                    end
                end
              reg4876 <= forvar4752[(2'h2):(1'h0)];
            end
        end
      reg4877 <= forvar3748;
      if (((~(-(reg3557 ? reg4876 : (8'hac)))) ?
          ((^reg4748) | ($unsigned(reg4796) >>> (&(8'hac)))) : (8'ha0)))
        begin
          if (($signed(((forvar3722 >> reg3603) && (reg4871 ~^ reg3591))) ?
              $signed((reg3707[(1'h0):(1'h0)] ?
                  (reg4835 ^~ wire3542) : ((8'hb5) ^ reg3612))) : forvar4801[(3'h7):(3'h7)]))
            begin
              for (forvar4878 = (1'h0); (forvar4878 < (1'h0)); forvar4878 = (forvar4878 + (1'h1)))
                begin
                  for (forvar4879 = (1'h0); (forvar4879 < (1'h0)); forvar4879 = (forvar4879 + (1'h1)))
                    begin
                      reg4880 <= reg3692[(2'h2):(2'h2)];
                      reg4881 <= ((($unsigned(reg3615) ?
                              (reg3726 << forvar3636) : reg4740[(1'h0):(1'h0)]) ?
                          (&(forvar3589 << (8'ha4))) : reg3667[(1'h0):(1'h0)]) * ($signed($signed(forvar4743)) ?
                          ((8'ha8) == (+reg3724)) : $unsigned($signed(reg4740))));
                      reg4882 <= (~|$signed((+(forvar3544 ?
                          forvar4797 : reg3600))));
                      reg4883 <= (reg3757 ~^ (8'hb2));
                    end
                  if ((forvar4765[(1'h1):(1'h0)] <= (^reg3610[(1'h0):(1'h0)])))
                    begin
                      reg4884 <= (reg3633[(2'h2):(2'h2)] > reg3606);
                      reg4885 <= (reg3695[(2'h2):(1'h0)] ?
                          forvar3647[(3'h5):(3'h4)] : forvar3657[(4'h9):(1'h1)]);
                    end
                  else
                    begin
                      reg4884 <= {(($signed((8'had)) ?
                              forvar3748[(1'h1):(1'h0)] : forvar4782[(3'h7):(2'h3)]) << reg3750)};
                    end
                  for (forvar4886 = (1'h0); (forvar4886 < (1'h0)); forvar4886 = (forvar4886 + (1'h1)))
                    begin
                      reg4887 <= {$signed($signed(forvar3697))};
                      reg4888 <= (($unsigned(reg3564) ?
                              ($unsigned(reg3692) <<< forvar4842) : $signed({reg4780})) ?
                          {forvar4735[(4'h8):(1'h1)]} : $signed((^(reg4801 ?
                              reg3619 : forvar4752))));
                    end
                end
              reg4889 <= $unsigned(reg3761[(1'h0):(1'h0)]);
              reg4890 <= ($signed((forvar3740[(1'h1):(1'h0)] ^ (reg4826 & forvar4866))) ?
                  (!$unsigned((|reg4828))) : reg4862[(4'hf):(4'hf)]);
            end
          else
            begin
              for (forvar4878 = (1'h0); (forvar4878 < (2'h3)); forvar4878 = (forvar4878 + (1'h1)))
                begin
                  for (forvar4879 = (1'h0); (forvar4879 < (1'h1)); forvar4879 = (forvar4879 + (1'h1)))
                    begin
                      reg4880 <= reg3659[(4'h8):(2'h2)];
                      reg4881 <= $signed($signed(((reg3734 ?
                          (8'ha7) : (8'ha6)) ^ (forvar3645 ?
                          forvar3742 : reg3728))));
                    end
                  reg4882 <= forvar4823;
                  reg4883 <= (|$signed((~|reg4779[(1'h0):(1'h0)])));
                  if ($unsigned((&$signed((8'hb4)))))
                    begin
                      reg4884 <= (forvar3553[(1'h1):(1'h1)] + (forvar3656 ?
                          $unsigned(forvar3706) : {reg3608}));
                      reg4885 <= $unsigned($signed((reg3746[(2'h2):(1'h0)] ?
                          ((8'ha3) && reg4880) : $unsigned(forvar3636))));
                      reg4886 <= reg3552;
                      reg4887 <= $unsigned($unsigned({reg3730}));
                    end
                  else
                    begin
                      reg4884 <= (^~($signed($signed(forvar4842)) ?
                          reg4764[(1'h1):(1'h0)] : (+(~forvar4852))));
                    end
                end
              for (forvar4888 = (1'h0); (forvar4888 < (1'h1)); forvar4888 = (forvar4888 + (1'h1)))
                begin
                  for (forvar4889 = (1'h0); (forvar4889 < (1'h0)); forvar4889 = (forvar4889 + (1'h1)))
                    begin
                      reg4890 <= (^~(&{(reg3696 ? reg3600 : forvar3740)}));
                      reg4891 <= reg3716[(4'he):(4'hc)];
                    end
                  if (reg3673[(3'h4):(3'h4)])
                    begin
                      reg4892 <= (-$signed(reg4842[(1'h0):(1'h0)]));
                      reg4893 <= $unsigned(($unsigned(reg3639[(1'h1):(1'h1)]) ?
                          reg4819 : reg3605));
                      reg4894 <= $signed((($signed((8'hb7)) ?
                              ((8'had) ?
                                  forvar4796 : reg3675) : reg3615[(2'h3):(1'h1)]) ?
                          forvar3645[(1'h1):(1'h1)] : reg4846[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg4892 <= (~|((reg3556 ?
                          reg4819[(4'h8):(1'h1)] : $unsigned((8'ha1))) ^ (reg4860[(3'h4):(3'h4)] ~^ reg4742)));
                      reg4893 <= $unsigned((reg3582 ?
                          (8'hab) : reg4741[(1'h0):(1'h0)]));
                      reg4894 <= (8'ha1);
                    end
                end
            end
          if (reg3569[(4'hc):(1'h0)])
            begin
              for (forvar4895 = (1'h0); (forvar4895 < (2'h2)); forvar4895 = (forvar4895 + (1'h1)))
                begin
                  for (forvar4896 = (1'h0); (forvar4896 < (1'h0)); forvar4896 = (forvar4896 + (1'h1)))
                    begin
                      reg4897 <= reg3668[(3'h7):(3'h5)];
                      reg4898 <= (reg3729[(1'h0):(1'h0)] ?
                          (((|reg4779) && (|reg3558)) << $signed({reg3605})) : {$unsigned($unsigned(forvar3722))});
                    end
                end
              for (forvar4899 = (1'h0); (forvar4899 < (2'h2)); forvar4899 = (forvar4899 + (1'h1)))
                begin
                  for (forvar4900 = (1'h0); (forvar4900 < (2'h3)); forvar4900 = (forvar4900 + (1'h1)))
                    begin
                      reg4901 <= (($signed((|reg3758)) ?
                              $signed($signed(forvar4796)) : ($signed(reg3734) ?
                                  (&forvar4814) : {reg3669})) ?
                          reg4844 : reg4789[(2'h2):(1'h0)]);
                      reg4902 <= ((((8'hb7) ?
                              $signed(reg3558) : (reg4788 ?
                                  forvar3645 : forvar4801)) ?
                          $unsigned(reg4792) : $unsigned(reg3660)) ~^ (reg3572 ?
                          forvar3547 : $signed((reg3564 ? reg3742 : reg4840))));
                      reg4903 <= (({((8'ha4) == reg3738)} ?
                              $signed($signed(reg4869)) : {reg4766[(4'hb):(4'h9)]}) ?
                          (|$unsigned((reg3721 <<< reg4842))) : $unsigned({reg4893[(4'h8):(2'h3)]}));
                    end
                  for (forvar4904 = (1'h0); (forvar4904 < (1'h0)); forvar4904 = (forvar4904 + (1'h1)))
                    begin
                      reg4905 <= forvar4879[(3'h6):(1'h1)];
                      reg4906 <= $unsigned(reg4898);
                      reg4907 <= {(((reg4876 ?
                                  forvar3710 : forvar4850) ^ reg3724) ?
                              $signed(reg4845) : $unsigned((reg3673 ?
                                  forvar4758 : (8'ha2))))};
                    end
                  if ((reg4755[(2'h2):(1'h1)] >= $unsigned($signed($unsigned(wire3767)))))
                    begin
                      reg4908 <= (+$unsigned($unsigned((reg3569 - forvar4797))));
                    end
                  else
                    begin
                      reg4908 <= {reg3729};
                      reg4909 <= ((-(((8'h9e) ? reg4759 : (8'ha1)) ?
                              $unsigned(reg3700) : forvar4825[(2'h3):(1'h1)])) ?
                          (&$signed((&reg4870))) : (~|reg3571));
                    end
                  if (reg3733[(1'h0):(1'h0)])
                    begin
                      reg4910 <= forvar4750;
                    end
                  else
                    begin
                      reg4910 <= (reg3635[(4'h9):(3'h4)] ?
                          (&(reg3652 <= {reg3743})) : reg4862[(3'h7):(1'h1)]);
                      reg4911 <= (^~reg4810);
                      reg4912 <= forvar4824[(3'h4):(1'h0)];
                      reg4913 <= ($signed(reg4871[(3'h5):(2'h2)]) ?
                          reg3659[(4'h8):(1'h0)] : ({(forvar3654 ?
                                  wire4730 : forvar4895)} << (^~((8'hba) ?
                              forvar3545 : forvar4865))));
                    end
                end
            end
          else
            begin
              for (forvar4895 = (1'h0); (forvar4895 < (1'h1)); forvar4895 = (forvar4895 + (1'h1)))
                begin
                  for (forvar4896 = (1'h0); (forvar4896 < (1'h0)); forvar4896 = (forvar4896 + (1'h1)))
                    begin
                      reg4897 <= reg3731[(4'ha):(3'h6)];
                    end
                end
              for (forvar4898 = (1'h0); (forvar4898 < (2'h3)); forvar4898 = (forvar4898 + (1'h1)))
                begin
                  for (forvar4899 = (1'h0); (forvar4899 < (1'h1)); forvar4899 = (forvar4899 + (1'h1)))
                    begin
                      reg4900 <= reg4746[(2'h2):(1'h1)];
                      reg4901 <= (({reg4789} ?
                              $signed(reg3550[(4'hc):(3'h7)]) : reg3569) ?
                          (((8'hae) ?
                              (~reg3655) : reg3723[(1'h1):(1'h1)]) * (~reg4789[(4'h8):(3'h7)])) : (reg3620[(2'h3):(1'h1)] ?
                              $unsigned($signed(reg4746)) : $unsigned((8'hb3))));
                    end
                  if ($unsigned($unsigned($unsigned({forvar3601}))))
                    begin
                      reg4902 <= reg4796;
                      reg4903 <= reg4828;
                      reg4904 <= $unsigned((((^~(8'h9e)) >>> $signed(reg3550)) - reg4740));
                      reg4905 <= $unsigned(forvar4900[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg4902 <= reg3554[(4'ha):(1'h1)];
                    end
                end
              reg4906 <= ($signed(($signed(reg3652) ? (~|(8'hb9)) : reg4874)) ?
                  forvar4829[(1'h0):(1'h0)] : ($unsigned($unsigned((8'ha2))) ?
                      $signed((reg4734 ?
                          reg4818 : (8'hba))) : (+$unsigned(forvar3745))));
              for (forvar4907 = (1'h0); (forvar4907 < (2'h3)); forvar4907 = (forvar4907 + (1'h1)))
                begin
                  if ({reg3616[(1'h0):(1'h0)]})
                    begin
                      reg4908 <= reg3555[(3'h7):(3'h7)];
                      reg4909 <= ({{$signed(reg3670)}} ^~ ((~&{reg4891}) ?
                          reg3550 : $unsigned((~reg3645))));
                      reg4910 <= reg4743[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg4908 <= reg3574;
                      reg4909 <= reg3709;
                      reg4910 <= reg3648[(2'h2):(2'h2)];
                    end
                  for (forvar4911 = (1'h0); (forvar4911 < (1'h1)); forvar4911 = (forvar4911 + (1'h1)))
                    begin
                      reg4912 <= forvar4848;
                    end
                  if (($signed(reg4856[(1'h1):(1'h1)]) * $signed(reg3671)))
                    begin
                      reg4913 <= (8'hb7);
                      reg4914 <= (~&(&($unsigned(reg3600) ?
                          (reg3746 ^~ reg3557) : forvar4808[(1'h1):(1'h0)])));
                      reg4915 <= {{(~{reg4904})}};
                    end
                  else
                    begin
                      reg4913 <= ({(+$signed((8'hb2)))} == reg3660);
                      reg4914 <= $unsigned(($unsigned($unsigned(reg4811)) ?
                          reg4870[(4'hc):(3'h6)] : $signed(forvar4895[(2'h3):(2'h2)])));
                    end
                  if ({forvar3702})
                    begin
                      reg4916 <= (((~|(reg3712 ?
                              reg3630 : reg4870)) >>> reg4889) ?
                          reg3568[(2'h3):(2'h3)] : reg3750[(1'h1):(1'h1)]);
                      reg4917 <= forvar4760;
                      reg4918 <= ($signed($signed((wire4793 >= reg3687))) ?
                          (((~forvar4907) ?
                              $unsigned(reg4902) : (reg3582 * wire4794)) ^~ forvar4911) : (forvar4736[(1'h0):(1'h0)] ?
                              (forvar3613 ?
                                  $signed(reg4884) : {reg3568}) : wire4733));
                      reg4919 <= ($signed(({reg4792} ?
                              $signed(reg4831) : forvar3601)) ?
                          $unsigned($unsigned((~&reg3597))) : reg4749);
                    end
                  else
                    begin
                      reg4916 <= wire4794[(1'h1):(1'h0)];
                    end
                end
            end
          if ($signed(reg4870))
            begin
              for (forvar4920 = (1'h0); (forvar4920 < (2'h2)); forvar4920 = (forvar4920 + (1'h1)))
                begin
                  for (forvar4921 = (1'h0); (forvar4921 < (2'h3)); forvar4921 = (forvar4921 + (1'h1)))
                    begin
                      reg4922 <= ($unsigned($unsigned(forvar4886)) & ($signed(forvar4810) * {(^~reg3561)}));
                      reg4923 <= (-(8'hb7));
                      reg4924 <= $unsigned(((~$signed(forvar3558)) ?
                          {$signed(reg4806)} : (~&$signed(reg4902))));
                    end
                  for (forvar4925 = (1'h0); (forvar4925 < (2'h3)); forvar4925 = (forvar4925 + (1'h1)))
                    begin
                      reg4926 <= $unsigned(reg4842[(4'hc):(3'h7)]);
                      reg4927 <= reg3629;
                    end
                  for (forvar4928 = (1'h0); (forvar4928 < (2'h3)); forvar4928 = (forvar4928 + (1'h1)))
                    begin
                      reg4929 <= (&({{reg4917}} * $signed((~&reg4791))));
                      reg4930 <= {reg4919};
                      reg4931 <= $signed(reg4868);
                      reg4932 <= $unsigned($signed(reg4850[(4'h8):(2'h3)]));
                    end
                  reg4933 <= (~&(^reg3661));
                end
            end
          else
            begin
              for (forvar4920 = (1'h0); (forvar4920 < (2'h3)); forvar4920 = (forvar4920 + (1'h1)))
                begin
                  for (forvar4921 = (1'h0); (forvar4921 < (2'h3)); forvar4921 = (forvar4921 + (1'h1)))
                    begin
                      reg4922 <= reg3676[(3'h4):(1'h0)];
                      reg4923 <= ((($signed(forvar4760) ?
                              reg3581[(1'h0):(1'h0)] : $unsigned((8'ha0))) >>> (reg3684 < (reg4819 == forvar3593))) ?
                          ($unsigned($unsigned(reg3665)) ?
                              (reg3703[(1'h1):(1'h1)] == (reg4797 ?
                                  reg3576 : forvar3753)) : reg3646[(1'h0):(1'h0)]) : forvar3676);
                      reg4924 <= (($unsigned($signed(forvar3641)) ^ (((8'ha3) ?
                              reg4906 : reg4813) ?
                          (forvar3549 ?
                              (8'ha8) : reg4906) : forvar4842)) - ($unsigned(reg3564) ?
                          reg3558[(3'h7):(2'h2)] : $unsigned((reg3714 * reg4755))));
                      reg4925 <= {$unsigned({$unsigned(reg4894)})};
                    end
                end
              for (forvar4926 = (1'h0); (forvar4926 < (1'h0)); forvar4926 = (forvar4926 + (1'h1)))
                begin
                  for (forvar4927 = (1'h0); (forvar4927 < (2'h3)); forvar4927 = (forvar4927 + (1'h1)))
                    begin
                      reg4928 <= ($unsigned(reg3673[(1'h0):(1'h0)]) ?
                          reg4800[(1'h0):(1'h0)] : reg3677[(4'ha):(2'h2)]);
                      reg4929 <= reg3676;
                    end
                  if (forvar3710)
                    begin
                      reg4930 <= (($unsigned($unsigned(reg3630)) ?
                          ((forvar4822 ? reg3705 : reg4761) ?
                              (&(8'hb4)) : reg4751[(1'h1):(1'h1)]) : (^~{reg3730})) <<< $unsigned(($unsigned(reg4844) + reg3689[(2'h2):(1'h1)])));
                      reg4931 <= $unsigned((+{$unsigned((8'h9c))}));
                    end
                  else
                    begin
                      reg4930 <= ((forvar3558 != reg3764[(3'h7):(3'h5)]) ?
                          $signed(((8'ha8) ?
                              $signed((8'ha4)) : $signed(reg4801))) : $unsigned(reg4750));
                      reg4931 <= (forvar4826[(1'h0):(1'h0)] ?
                          reg3552 : {(&(reg3701 && reg4749))});
                      reg4932 <= reg4854;
                      reg4933 <= (forvar3619[(2'h3):(1'h1)] ?
                          $signed(((reg3617 ? reg3618 : reg3583) > (reg3570 ?
                              reg3600 : (8'h9f)))) : reg3549);
                    end
                end
            end
          for (forvar4934 = (1'h0); (forvar4934 < (2'h3)); forvar4934 = (forvar4934 + (1'h1)))
            begin
              if ((reg4824 << {($unsigned(forvar3645) ?
                      (~|reg3741) : (~|reg3557))}))
                begin
                  for (forvar4935 = (1'h0); (forvar4935 < (1'h1)); forvar4935 = (forvar4935 + (1'h1)))
                    begin
                      reg4936 <= $unsigned(((wire3767[(3'h4):(1'h1)] ?
                              (reg3620 ?
                                  reg3584 : reg3638) : $unsigned(reg3640)) ?
                          forvar4839[(1'h0):(1'h0)] : ((+reg4828) ?
                              (reg3621 ?
                                  (8'hb3) : wire4864) : (~&forvar3607))));
                      reg4937 <= forvar4773[(2'h3):(2'h3)];
                      reg4938 <= $unsigned($unsigned(reg4910[(2'h3):(1'h0)]));
                      reg4939 <= {$unsigned($signed((-reg3709)))};
                    end
                  for (forvar4940 = (1'h0); (forvar4940 < (2'h2)); forvar4940 = (forvar4940 + (1'h1)))
                    begin
                      reg4941 <= ((({forvar4736} < reg3639) ~^ forvar4796) * (($unsigned(reg4851) - forvar4839) == forvar4777));
                      reg4942 <= $signed((forvar3706[(1'h0):(1'h0)] ?
                          (reg4759 ^~ $signed(reg3751)) : reg3546[(4'h9):(3'h6)]));
                    end
                end
              else
                begin
                  for (forvar4935 = (1'h0); (forvar4935 < (1'h0)); forvar4935 = (forvar4935 + (1'h1)))
                    begin
                      reg4936 <= (reg3580[(3'h5):(2'h2)] > reg3559[(3'h7):(1'h1)]);
                      reg4937 <= ((+reg3635) ?
                          (~^$unsigned(reg4826[(2'h3):(2'h3)])) : (8'hb8));
                      reg4938 <= forvar4802;
                      reg4939 <= $unsigned($signed($signed(reg3612)));
                    end
                end
              reg4943 <= $signed(reg4811[(3'h4):(2'h2)]);
              for (forvar4944 = (1'h0); (forvar4944 < (2'h3)); forvar4944 = (forvar4944 + (1'h1)))
                begin
                  if (forvar3672)
                    begin
                      reg4945 <= {((&{reg4807}) | (forvar3547 ?
                              $signed((8'hab)) : reg4850[(4'hd):(3'h7)]))};
                      reg4946 <= forvar4746;
                      reg4947 <= $unsigned(forvar3711);
                      reg4948 <= ($signed({forvar3681[(3'h4):(1'h0)]}) ?
                          (^((-reg4873) >= (reg3752 ^ reg3614))) : reg4810);
                    end
                  else
                    begin
                      reg4945 <= ((^(reg3618[(3'h4):(3'h4)] + ((8'hb5) ?
                              reg4757 : reg4863))) ?
                          forvar3626 : $unsigned(((forvar4803 ?
                              reg3596 : reg3732) < (reg3712 << reg4915))));
                      reg4946 <= {(8'hb4)};
                    end
                  for (forvar4949 = (1'h0); (forvar4949 < (2'h3)); forvar4949 = (forvar4949 + (1'h1)))
                    begin
                      reg4950 <= (((~|(8'ha7)) ~^ $unsigned((reg4768 ?
                          forvar4758 : reg3691))) ^~ (reg4767[(1'h0):(1'h0)] ?
                          (~|reg4779[(1'h1):(1'h1)]) : forvar3549));
                      reg4951 <= reg4751;
                      reg4952 <= reg4882[(2'h3):(2'h3)];
                      reg4953 <= $signed(($unsigned(reg4762[(2'h2):(1'h1)]) > (reg3750[(2'h2):(1'h0)] < forvar4829)));
                    end
                  for (forvar4954 = (1'h0); (forvar4954 < (2'h2)); forvar4954 = (forvar4954 + (1'h1)))
                    begin
                      reg4955 <= reg3596[(3'h6):(2'h3)];
                      reg4956 <= {reg3625};
                      reg4957 <= ((+(8'hb4)) ?
                          ((8'ha8) ?
                              (8'h9f) : reg3683) : forvar4810[(1'h1):(1'h1)]);
                      reg4958 <= $unsigned(reg4845[(4'h9):(2'h2)]);
                    end
                  for (forvar4959 = (1'h0); (forvar4959 < (1'h0)); forvar4959 = (forvar4959 + (1'h1)))
                    begin
                      reg4960 <= reg3599[(2'h2):(1'h1)];
                      reg4961 <= ((|reg4862[(2'h3):(1'h1)]) <<< $unsigned((reg4957[(1'h1):(1'h0)] >> (forvar3579 ?
                          reg4792 : reg3727))));
                      reg4962 <= ({reg3723[(1'h1):(1'h0)]} ?
                          (~^$signed(reg4948[(4'h8):(1'h0)])) : $unsigned($unsigned(reg4805[(3'h4):(2'h2)])));
                      reg4963 <= ($unsigned($unsigned((~&reg3620))) ?
                          $unsigned(((&reg4773) && wire3540[(1'h0):(1'h0)])) : {((^~(8'h9d)) | (forvar4855 ?
                                  reg4871 : reg3620))});
                    end
                end
            end
        end
      else
        begin
          if ($unsigned(forvar3739[(2'h2):(1'h0)]))
            begin
              for (forvar4878 = (1'h0); (forvar4878 < (2'h3)); forvar4878 = (forvar4878 + (1'h1)))
                begin
                  for (forvar4879 = (1'h0); (forvar4879 < (1'h1)); forvar4879 = (forvar4879 + (1'h1)))
                    begin
                      reg4880 <= $unsigned($unsigned($signed($unsigned(reg4762))));
                      reg4881 <= ({$unsigned({reg3568})} ?
                          (!reg4799) : forvar4773[(2'h2):(2'h2)]);
                    end
                  if ($signed($unsigned(forvar4834)))
                    begin
                      reg4882 <= (~^$signed(reg4937[(3'h7):(1'h1)]));
                      reg4883 <= $signed((!(8'had)));
                      reg4884 <= {forvar4824[(1'h1):(1'h1)]};
                      reg4885 <= (~{reg4880});
                    end
                  else
                    begin
                      reg4882 <= (~^reg3568[(4'hc):(3'h4)]);
                      reg4883 <= {$signed(forvar3636[(4'h9):(3'h6)])};
                      reg4884 <= $unsigned($unsigned($signed(reg4749)));
                    end
                  for (forvar4886 = (1'h0); (forvar4886 < (2'h3)); forvar4886 = (forvar4886 + (1'h1)))
                    begin
                      reg4887 <= $signed(forvar3607[(3'h5):(3'h4)]);
                      reg4888 <= reg4876;
                    end
                  reg4889 <= (((|((8'ha6) >> wire3766)) < $unsigned($unsigned(forvar4735))) != (^reg4907));
                end
              if (($signed(($signed(reg3665) >= $unsigned((8'ha4)))) ^~ (reg4882 ?
                  reg3605[(2'h3):(2'h3)] : {(!forvar4911)})))
                begin
                  for (forvar4890 = (1'h0); (forvar4890 < (1'h0)); forvar4890 = (forvar4890 + (1'h1)))
                    begin
                      reg4891 <= (({(reg3580 - (8'hb2))} + $signed((reg3696 | (8'ha5)))) ?
                          forvar3566 : ($unsigned(reg4850[(4'hb):(1'h0)]) & (&reg4931)));
                      reg4892 <= {((&(forvar4921 ?
                              reg4914 : reg3587)) ~^ ((reg4821 >= forvar4928) ?
                              (reg4938 <<< reg3744) : (!(8'haf))))};
                      reg4893 <= $signed((~|reg3545));
                    end
                  for (forvar4894 = (1'h0); (forvar4894 < (1'h0)); forvar4894 = (forvar4894 + (1'h1)))
                    begin
                      reg4895 <= reg3749;
                      reg4896 <= (reg4792[(2'h3):(2'h2)] <<< (~^forvar3734));
                    end
                  for (forvar4897 = (1'h0); (forvar4897 < (1'h1)); forvar4897 = (forvar4897 + (1'h1)))
                    begin
                      reg4898 <= ((($signed(reg3749) > $signed(forvar3717)) ?
                          $signed($unsigned(forvar4770)) : ($signed(reg4891) ?
                              $unsigned((8'ha9)) : reg3646)) <<< reg3705[(3'h4):(2'h3)]);
                      reg4899 <= reg3625;
                      reg4900 <= reg3557[(4'he):(4'hd)];
                    end
                end
              else
                begin
                  for (forvar4890 = (1'h0); (forvar4890 < (1'h1)); forvar4890 = (forvar4890 + (1'h1)))
                    begin
                      reg4891 <= (~^$unsigned($unsigned((forvar4743 || reg3659))));
                    end
                  for (forvar4892 = (1'h0); (forvar4892 < (2'h3)); forvar4892 = (forvar4892 + (1'h1)))
                    begin
                      reg4893 <= ($signed((~&$signed((8'hb4)))) ?
                          ((^reg4869) ?
                              reg3691[(2'h2):(1'h0)] : forvar3631) : reg4824);
                      reg4894 <= ((reg4874[(3'h4):(3'h4)] ?
                          $signed((^~reg4801)) : reg4936[(2'h2):(1'h1)]) >> reg4823[(3'h5):(2'h2)]);
                      reg4895 <= $unsigned($unsigned($unsigned($unsigned(reg3576))));
                      reg4896 <= forvar3641[(3'h6):(3'h4)];
                    end
                  reg4897 <= reg4768;
                end
              if ((forvar4944 ?
                  reg3741[(3'h5):(1'h0)] : $unsigned($signed((!reg3694)))))
                begin
                  reg4901 <= reg3729;
                  for (forvar4902 = (1'h0); (forvar4902 < (1'h0)); forvar4902 = (forvar4902 + (1'h1)))
                    begin
                      reg4903 <= ($unsigned($unsigned((reg3687 ^ (8'ha8)))) ?
                          forvar3753[(2'h3):(1'h1)] : ($unsigned({(8'ha2)}) ?
                              (!{reg3765}) : $signed($signed(reg4867))));
                    end
                end
              else
                begin
                  for (forvar4901 = (1'h0); (forvar4901 < (1'h0)); forvar4901 = (forvar4901 + (1'h1)))
                    begin
                      reg4902 <= ($signed($signed($unsigned(reg4888))) ?
                          (8'hb3) : $unsigned($unsigned((reg3544 ?
                              forvar4773 : (8'hb2)))));
                      reg4903 <= (^$unsigned((~^reg3632[(3'h4):(3'h4)])));
                      reg4904 <= ((!$unsigned($signed(forvar4866))) + $unsigned((~^$unsigned((8'ha0)))));
                      reg4905 <= reg4904;
                    end
                  for (forvar4906 = (1'h0); (forvar4906 < (2'h2)); forvar4906 = (forvar4906 + (1'h1)))
                    begin
                      reg4907 <= $unsigned($signed(forvar3706));
                      reg4908 <= (!forvar4823[(4'hc):(3'h4)]);
                    end
                  if (({reg3720[(2'h2):(1'h0)]} ?
                      ($signed($signed(forvar4855)) ?
                          reg4743 : $signed((~|reg3575))) : (^~reg4962[(1'h1):(1'h0)])))
                    begin
                      reg4909 <= (((~(forvar3739 ?
                              reg3612 : forvar4911)) + $signed({reg3736})) ?
                          ((~|$unsigned(reg3737)) - $unsigned($signed(reg4844))) : $signed(({reg3551} ?
                              (reg3758 ?
                                  (8'ha3) : (8'hb4)) : reg3662[(2'h3):(1'h1)])));
                      reg4910 <= {$unsigned($signed(reg3639))};
                    end
                  else
                    begin
                      reg4909 <= reg4750[(4'hc):(2'h2)];
                    end
                end
            end
          else
            begin
              if ((({(reg3629 ? reg3555 : (8'hb0))} >= reg4759) ?
                  $unsigned($signed(reg3693)) : ($signed(((8'hb2) | reg3630)) ?
                      reg4747 : ($signed((8'haf)) | (|reg4802)))))
                begin
                  if (($unsigned((&(|(8'hb1)))) ?
                      (reg3656 ?
                          {$signed(reg3678)} : (forvar3641 <= {(8'haa)})) : (((forvar3745 | reg3644) ?
                          $signed(forvar4940) : reg4788) == reg4773)))
                    begin
                      reg4878 <= ({{$unsigned(reg3752)}} * (((forvar4879 ?
                          reg3756 : reg4798) << ((8'ha3) ?
                          reg3645 : reg4822)) <= ((forvar3645 ?
                          wire3540 : reg3689) * (~|reg4806))));
                      reg4879 <= $signed({(|(^reg3687))});
                      reg4880 <= (~{reg3583});
                      reg4881 <= $signed(reg4734[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4878 <= $unsigned($signed({reg3642[(2'h3):(1'h1)]}));
                      reg4879 <= $unsigned(((|(forvar4738 ?
                          reg4758 : reg4767)) | {(^forvar4758)}));
                      reg4880 <= (^(8'hb6));
                      reg4881 <= reg4933;
                    end
                  if ($unsigned((forvar4826[(2'h2):(1'h0)] ?
                      ((reg4913 + reg4802) ?
                          $signed(forvar3660) : (reg3764 ?
                              forvar4822 : reg4962)) : forvar3547)))
                    begin
                      reg4882 <= (((8'hb3) ?
                          ({reg4892} ?
                              $unsigned((8'hb4)) : reg4837) : (!(~&reg4803))) ^ (reg4790[(3'h4):(1'h0)] ?
                          $unsigned(reg3553) : forvar3641));
                      reg4883 <= forvar4753;
                      reg4884 <= {(({forvar4878} || (reg3564 >= wire4864)) && (&reg4883[(2'h3):(1'h0)]))};
                      reg4885 <= {reg3667};
                    end
                  else
                    begin
                      reg4882 <= reg3597;
                      reg4883 <= $unsigned(forvar3734[(3'h5):(3'h4)]);
                      reg4884 <= (8'hb8);
                    end
                end
              else
                begin
                  reg4878 <= $signed((^~(+reg3695)));
                  if (((~|(~^((8'ha2) ? forvar4797 : forvar4911))) ?
                      ((^~$signed(reg4860)) >= (forvar4949[(3'h4):(1'h1)] ?
                          (reg4800 ^ reg3635) : reg4750[(1'h1):(1'h0)])) : (reg3620[(5'h10):(1'h0)] <= ($unsigned(forvar3740) & $signed(reg4888)))))
                    begin
                      reg4879 <= reg3671;
                      reg4880 <= forvar3734[(5'h10):(5'h10)];
                    end
                  else
                    begin
                      reg4879 <= ((8'h9e) ?
                          forvar4752[(4'ha):(3'h4)] : forvar4824);
                      reg4880 <= (reg3696 & ((((8'hb9) ?
                          reg4769 : (8'ha6)) >= (reg4963 ?
                          reg4814 : reg3757)) <= ($signed(forvar4959) ?
                          (-reg3569) : {(8'hb7)})));
                      reg4881 <= (8'ha8);
                      reg4882 <= ($signed(reg3588) >>> (~forvar3626[(1'h0):(1'h0)]));
                    end
                  reg4883 <= (~&$unsigned({$signed((8'hb6))}));
                end
              if (reg4838[(3'h5):(2'h3)])
                begin
                  if ((+(8'had)))
                    begin
                      reg4886 <= (^reg3712);
                      reg4887 <= (((~|(8'hb0)) ?
                              ((^~forvar4896) ?
                                  reg3700[(1'h1):(1'h1)] : {reg4777}) : $unsigned(reg3619[(2'h2):(2'h2)])) ?
                          $signed((~(reg4886 ?
                              reg3674 : reg4870))) : $unsigned((forvar4834 ?
                              (reg4811 ?
                                  (8'hb7) : forvar4746) : (reg4931 + forvar3559))));
                      reg4888 <= reg3553;
                      reg4889 <= $signed((^~reg4780));
                    end
                  else
                    begin
                      reg4886 <= ($signed(reg3614) ?
                          forvar3669 : reg4828[(3'h6):(1'h0)]);
                      reg4887 <= (reg4804[(3'h4):(1'h0)] & reg3707);
                      reg4888 <= reg3587[(4'hb):(4'h8)];
                    end
                  if ((^~(reg4736[(4'he):(4'hc)] ?
                      ({reg4952} >>> (reg3627 ?
                          reg4847 : (8'ha2))) : (+(~|(8'hb4))))))
                    begin
                      reg4890 <= {(~forvar4826)};
                      reg4891 <= ($unsigned((reg3600[(3'h5):(3'h4)] ?
                          forvar4886 : forvar3740)) ~^ reg4779);
                    end
                  else
                    begin
                      reg4890 <= ({$unsigned($signed(reg4919))} == ($unsigned(reg3731[(3'h5):(1'h1)]) + forvar4944));
                      reg4891 <= $unsigned(($signed((forvar4866 ?
                              (8'h9f) : (8'ha8))) ?
                          reg3718[(1'h0):(1'h0)] : (reg4799[(2'h3):(2'h2)] >= (reg4890 ?
                              reg3617 : reg3723))));
                      reg4892 <= $unsigned((($unsigned(reg3696) ?
                          reg3604 : (+wire3540)) ^ $signed((reg4741 ?
                          forvar4906 : (8'hac)))));
                    end
                end
              else
                begin
                  for (forvar4886 = (1'h0); (forvar4886 < (2'h3)); forvar4886 = (forvar4886 + (1'h1)))
                    begin
                      reg4887 <= reg3671[(3'h5):(3'h5)];
                    end
                  reg4888 <= (reg3691[(3'h5):(1'h1)] && {(-reg4781[(1'h1):(1'h1)])});
                  for (forvar4889 = (1'h0); (forvar4889 < (1'h1)); forvar4889 = (forvar4889 + (1'h1)))
                    begin
                      reg4890 <= reg3649;
                    end
                  for (forvar4891 = (1'h0); (forvar4891 < (2'h2)); forvar4891 = (forvar4891 + (1'h1)))
                    begin
                      reg4892 <= (~$signed(forvar3686));
                      reg4893 <= {(reg4797[(1'h0):(1'h0)] ?
                              ({forvar3654} >= reg3730[(2'h2):(2'h2)]) : ((reg4785 == reg3723) << {(8'h9d)}))};
                      reg4894 <= $signed($unsigned(forvar3549[(3'h7):(1'h0)]));
                    end
                end
              for (forvar4895 = (1'h0); (forvar4895 < (2'h3)); forvar4895 = (forvar4895 + (1'h1)))
                begin
                  if (reg3550)
                    begin
                      reg4896 <= ($signed($signed((wire4793 ?
                              (8'ha7) : reg3548))) ?
                          $signed(forvar3654) : forvar4928[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4896 <= $signed((reg3628 << $unsigned(forvar3549)));
                    end
                  if (forvar3742)
                    begin
                      reg4897 <= {$signed({$unsigned(reg3673)})};
                      reg4898 <= forvar4777;
                    end
                  else
                    begin
                      reg4897 <= reg4842;
                      reg4898 <= (reg4803 ?
                          ($signed($signed(forvar4743)) < $unsigned((8'had))) : (forvar4911 ?
                              forvar4852 : {reg3562[(1'h1):(1'h0)]}));
                      reg4899 <= (&{forvar4921[(3'h7):(3'h5)]});
                    end
                end
            end
        end
    end
  assign wire4964 = {(~{reg4950[(3'h7):(3'h5)]})};
  assign wire4965 = (((8'h9c) || forvar4822) | (((forvar4896 ?
                        forvar4822 : reg3603) & {reg4846}) & {(reg3760 ?
                            reg4832 : reg3596)}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1032  (y, clk, wire1037, wire1036, wire1035, wire1034, wire1033);
  output wire [(32'h99):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire1037;
  input wire [(4'hb):(1'h0)] wire1036;
  input wire signed [(3'h5):(1'h0)] wire1035;
  input wire [(4'hd):(1'h0)] wire1034;
  input wire [(5'h10):(1'h0)] wire1033;
  wire signed [(4'hc):(1'h0)] wire3535;
  wire [(2'h3):(1'h0)] wire3534;
  wire signed [(4'he):(1'h0)] wire3532;
  wire [(5'h10):(1'h0)] wire1751;
  wire [(3'h7):(1'h0)] wire1750;
  wire [(2'h3):(1'h0)] wire1749;
  wire [(4'hd):(1'h0)] wire1748;
  wire [(4'ha):(1'h0)] wire1747;
  wire [(3'h6):(1'h0)] wire1746;
  wire signed [(4'hc):(1'h0)] wire1745;
  wire signed [(3'h7):(1'h0)] wire1744;
  wire signed [(4'hf):(1'h0)] wire1742;
  wire [(3'h4):(1'h0)] wire1040;
  wire [(4'he):(1'h0)] wire1039;
  wire [(5'h10):(1'h0)] wire1038;
  assign y = {wire3535,
                 wire3534,
                 wire3532,
                 wire1751,
                 wire1750,
                 wire1749,
                 wire1748,
                 wire1747,
                 wire1746,
                 wire1745,
                 wire1744,
                 wire1742,
                 wire1040,
                 wire1039,
                 wire1038,
                 (1'h0)};
  assign wire1038 = $signed((^~(~^(wire1035 ? wire1035 : wire1034))));
  assign wire1039 = $signed((~&wire1035[(2'h2):(1'h0)]));
  assign wire1040 = $unsigned(wire1038[(2'h2):(1'h1)]);
  module1041 modinst1743 (.wire1045(wire1040), .y(wire1742), .wire1043(wire1035), .wire1042(wire1034), .wire1044(wire1038), .clk(clk));
  assign wire1744 = $signed(wire1034[(1'h1):(1'h0)]);
  assign wire1745 = {{(^~$signed(wire1035))}};
  assign wire1746 = {$signed(((wire1033 >>> wire1039) ?
                            (~^wire1038) : wire1034))};
  assign wire1747 = (&wire1034);
  assign wire1748 = wire1039;
  assign wire1749 = wire1040[(1'h0):(1'h0)];
  assign wire1750 = $signed($unsigned(wire1748[(1'h0):(1'h0)]));
  assign wire1751 = wire1748;
  module1752 modinst3533 (.y(wire3532), .wire1756(wire1748), .wire1755(wire1035), .clk(clk), .wire1753(wire1038), .wire1754(wire1744));
  assign wire3534 = (|(((wire1036 & wire1037) >> $unsigned(wire1033)) > $signed($signed(wire1745))));
  assign wire3535 = $signed(wire1749);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1752  (y, clk, wire1756, wire1755, wire1754, wire1753);
  output wire [(32'h19a8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire1756;
  input wire [(3'h4):(1'h0)] wire1755;
  input wire signed [(3'h7):(1'h0)] wire1754;
  input wire signed [(4'ha):(1'h0)] wire1753;
  wire [(4'hf):(1'h0)] wire3531;
  wire [(3'h7):(1'h0)] wire3035;
  wire [(4'h8):(1'h0)] wire2360;
  wire signed [(4'hf):(1'h0)] wire2359;
  wire [(3'h6):(1'h0)] wire2358;
  wire [(4'ha):(1'h0)] wire2357;
  wire signed [(4'hd):(1'h0)] wire2356;
  wire signed [(4'hc):(1'h0)] wire2355;
  wire signed [(4'hf):(1'h0)] wire2354;
  reg [(5'h10):(1'h0)] reg2353 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2352 = (1'h0);
  reg [(4'hf):(1'h0)] reg2342 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2341 = (1'h0);
  reg [(3'h5):(1'h0)] reg2339 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2336 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2351 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2350 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2349 = (1'h0);
  reg [(4'ha):(1'h0)] reg2348 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2347 = (1'h0);
  reg [(2'h2):(1'h0)] reg2346 = (1'h0);
  reg [(2'h2):(1'h0)] reg2345 = (1'h0);
  reg [(3'h5):(1'h0)] reg2344 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2343 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2342 = (1'h0);
  reg [(4'ha):(1'h0)] reg2341 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2340 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2339 = (1'h0);
  reg [(4'h8):(1'h0)] reg2338 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2337 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2336 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2335 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2334 = (1'h0);
  reg [(4'hd):(1'h0)] reg2333 = (1'h0);
  reg [(4'h8):(1'h0)] reg2332 = (1'h0);
  reg [(3'h7):(1'h0)] reg2331 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2329 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2328 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2327 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2326 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2325 = (1'h0);
  reg [(4'ha):(1'h0)] reg2324 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2323 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2322 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2321 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2320 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2319 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2318 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2317 = (1'h0);
  reg [(3'h4):(1'h0)] reg2316 = (1'h0);
  reg [(4'h8):(1'h0)] reg2315 = (1'h0);
  reg [(4'ha):(1'h0)] reg2314 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2313 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2312 = (1'h0);
  reg [(3'h7):(1'h0)] reg2311 = (1'h0);
  reg [(5'h10):(1'h0)] reg2310 = (1'h0);
  reg [(4'hf):(1'h0)] reg2309 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2307 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2301 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2289 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2288 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2291 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2290 = (1'h0);
  reg [(2'h3):(1'h0)] reg2287 = (1'h0);
  reg [(4'ha):(1'h0)] reg2308 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2307 = (1'h0);
  reg [(3'h7):(1'h0)] reg2305 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2306 = (1'h0);
  reg [(4'he):(1'h0)] forvar2305 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2304 = (1'h0);
  reg [(2'h3):(1'h0)] reg2303 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2302 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2301 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2300 = (1'h0);
  reg [(2'h2):(1'h0)] reg2299 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2298 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2297 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2296 = (1'h0);
  reg [(4'hc):(1'h0)] reg2295 = (1'h0);
  reg [(4'ha):(1'h0)] reg2294 = (1'h0);
  reg [(4'ha):(1'h0)] reg2293 = (1'h0);
  reg [(3'h5):(1'h0)] reg2292 = (1'h0);
  reg [(4'h8):(1'h0)] reg2291 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2290 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2289 = (1'h0);
  reg [(4'hc):(1'h0)] reg2288 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2287 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2232 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2230 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2227 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2225 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2220 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2216 = (1'h0);
  reg [(4'h9):(1'h0)] reg2209 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2208 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2207 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2202 = (1'h0);
  reg [(4'hb):(1'h0)] reg2203 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2201 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2200 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2195 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2187 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2188 = (1'h0);
  reg [(3'h7):(1'h0)] reg2185 = (1'h0);
  reg [(4'he):(1'h0)] forvar2183 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2173 = (1'h0);
  reg [(4'h9):(1'h0)] reg2180 = (1'h0);
  reg [(3'h7):(1'h0)] reg2179 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2177 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2170 = (1'h0);
  reg [(3'h6):(1'h0)] reg2168 = (1'h0);
  reg [(3'h6):(1'h0)] reg2286 = (1'h0);
  reg [(2'h3):(1'h0)] reg2285 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2284 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2283 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2282 = (1'h0);
  reg [(4'hc):(1'h0)] reg2281 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2280 = (1'h0);
  reg [(3'h6):(1'h0)] reg2279 = (1'h0);
  reg [(5'h10):(1'h0)] reg2278 = (1'h0);
  reg [(5'h10):(1'h0)] reg2277 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2276 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2275 = (1'h0);
  reg [(3'h7):(1'h0)] reg2269 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2268 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2265 = (1'h0);
  reg [(2'h3):(1'h0)] reg2264 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2263 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2262 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2255 = (1'h0);
  reg [(3'h4):(1'h0)] reg2256 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2252 = (1'h0);
  reg [(4'he):(1'h0)] reg2248 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2247 = (1'h0);
  reg [(5'h10):(1'h0)] reg2274 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2273 = (1'h0);
  reg [(5'h10):(1'h0)] reg2272 = (1'h0);
  reg [(2'h2):(1'h0)] reg2271 = (1'h0);
  reg [(3'h4):(1'h0)] reg2270 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2269 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2268 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2267 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2266 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2265 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2264 = (1'h0);
  reg [(4'h9):(1'h0)] reg2263 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2262 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2261 = (1'h0);
  reg [(2'h2):(1'h0)] reg2260 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2259 = (1'h0);
  reg [(4'hd):(1'h0)] reg2258 = (1'h0);
  reg [(4'he):(1'h0)] reg2257 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2256 = (1'h0);
  reg [(2'h2):(1'h0)] reg2255 = (1'h0);
  reg [(4'h8):(1'h0)] reg2254 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2253 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2252 = (1'h0);
  reg [(3'h7):(1'h0)] reg2243 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2242 = (1'h0);
  reg [(4'he):(1'h0)] reg2241 = (1'h0);
  reg [(3'h6):(1'h0)] reg2251 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2250 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2249 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2248 = (1'h0);
  reg [(4'hf):(1'h0)] reg2247 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2246 = (1'h0);
  reg [(4'ha):(1'h0)] reg2245 = (1'h0);
  reg [(2'h2):(1'h0)] reg2244 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2243 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2242 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2241 = (1'h0);
  reg [(4'h9):(1'h0)] reg2240 = (1'h0);
  reg [(3'h4):(1'h0)] reg2239 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2238 = (1'h0);
  reg [(4'ha):(1'h0)] reg2237 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2236 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2235 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2234 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2233 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2232 = (1'h0);
  reg [(4'ha):(1'h0)] reg2231 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2230 = (1'h0);
  reg [(4'hc):(1'h0)] reg2229 = (1'h0);
  reg [(4'he):(1'h0)] reg2228 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2227 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2226 = (1'h0);
  reg [(4'he):(1'h0)] reg2225 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2224 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2221 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2223 = (1'h0);
  reg [(4'hd):(1'h0)] reg2222 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2221 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2220 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2219 = (1'h0);
  reg [(2'h3):(1'h0)] reg2218 = (1'h0);
  reg [(2'h2):(1'h0)] reg2217 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2214 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2216 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2215 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2214 = (1'h0);
  reg [(4'h9):(1'h0)] reg2211 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2213 = (1'h0);
  reg [(4'he):(1'h0)] reg2212 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2211 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2210 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2209 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2208 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2175 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2169 = (1'h0);
  reg [(3'h5):(1'h0)] reg2207 = (1'h0);
  reg [(5'h10):(1'h0)] reg2206 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2205 = (1'h0);
  reg [(3'h7):(1'h0)] reg2204 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2203 = (1'h0);
  reg [(4'h8):(1'h0)] reg2202 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2201 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2200 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2199 = (1'h0);
  reg [(4'ha):(1'h0)] reg2198 = (1'h0);
  reg [(4'h8):(1'h0)] reg2197 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2196 = (1'h0);
  reg [(3'h6):(1'h0)] reg2191 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2190 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2195 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2194 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2193 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2192 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2191 = (1'h0);
  reg [(4'hc):(1'h0)] reg2190 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2189 = (1'h0);
  reg [(4'ha):(1'h0)] reg2188 = (1'h0);
  reg [(4'h8):(1'h0)] reg2187 = (1'h0);
  reg [(4'he):(1'h0)] reg2186 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2185 = (1'h0);
  reg [(4'h8):(1'h0)] reg2184 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2183 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2182 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2181 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2180 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2179 = (1'h0);
  reg [(4'hc):(1'h0)] reg2178 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2177 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2176 = (1'h0);
  reg [(4'ha):(1'h0)] reg2175 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2174 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2173 = (1'h0);
  reg [(4'hc):(1'h0)] reg2172 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2171 = (1'h0);
  reg [(3'h4):(1'h0)] reg2170 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2169 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2168 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2135 = (1'h0);
  reg [(4'he):(1'h0)] reg2131 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2130 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2124 = (1'h0);
  reg [(3'h5):(1'h0)] reg2121 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2119 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2117 = (1'h0);
  reg [(2'h3):(1'h0)] reg2113 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2112 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2111 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2109 = (1'h0);
  reg [(4'hb):(1'h0)] reg2167 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2166 = (1'h0);
  reg [(3'h4):(1'h0)] reg2165 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2164 = (1'h0);
  reg [(4'hc):(1'h0)] reg2163 = (1'h0);
  reg [(4'hd):(1'h0)] reg2162 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2161 = (1'h0);
  reg [(4'hd):(1'h0)] reg2160 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2159 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2158 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2157 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2156 = (1'h0);
  reg [(5'h10):(1'h0)] reg2150 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2148 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2143 = (1'h0);
  reg [(3'h4):(1'h0)] reg2155 = (1'h0);
  reg [(3'h4):(1'h0)] reg2154 = (1'h0);
  reg [(4'h9):(1'h0)] reg2153 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2152 = (1'h0);
  reg [(3'h7):(1'h0)] reg2151 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2150 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2149 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2148 = (1'h0);
  reg [(4'hf):(1'h0)] reg2147 = (1'h0);
  reg [(3'h5):(1'h0)] reg2146 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2145 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2144 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2143 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2142 = (1'h0);
  reg [(4'h8):(1'h0)] reg2141 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2140 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2139 = (1'h0);
  reg [(3'h7):(1'h0)] reg2138 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2137 = (1'h0);
  reg [(4'h9):(1'h0)] reg2136 = (1'h0);
  reg [(4'he):(1'h0)] reg2135 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2134 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2133 = (1'h0);
  reg [(4'he):(1'h0)] reg2132 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2131 = (1'h0);
  reg [(2'h3):(1'h0)] reg2130 = (1'h0);
  reg [(4'hb):(1'h0)] reg2129 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2128 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2127 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2126 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2125 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2124 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2123 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2122 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2121 = (1'h0);
  reg [(5'h10):(1'h0)] reg2120 = (1'h0);
  reg [(3'h7):(1'h0)] reg2119 = (1'h0);
  reg [(4'h9):(1'h0)] reg2118 = (1'h0);
  reg [(4'ha):(1'h0)] reg2117 = (1'h0);
  reg [(4'hb):(1'h0)] reg2116 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2115 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2114 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2113 = (1'h0);
  reg [(2'h3):(1'h0)] reg2112 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2111 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2110 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2109 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2087 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2108 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2107 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2106 = (1'h0);
  reg [(2'h3):(1'h0)] reg2105 = (1'h0);
  reg [(3'h4):(1'h0)] reg2104 = (1'h0);
  reg [(4'ha):(1'h0)] reg2102 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2096 = (1'h0);
  reg [(2'h2):(1'h0)] reg2103 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2102 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2101 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2100 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2099 = (1'h0);
  reg [(2'h3):(1'h0)] reg2098 = (1'h0);
  reg [(3'h7):(1'h0)] reg2097 = (1'h0);
  reg [(4'hf):(1'h0)] reg2096 = (1'h0);
  reg [(5'h10):(1'h0)] reg2093 = (1'h0);
  reg [(5'h10):(1'h0)] reg2095 = (1'h0);
  reg [(4'ha):(1'h0)] reg2094 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2093 = (1'h0);
  reg [(4'hd):(1'h0)] reg2092 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2091 = (1'h0);
  reg [(4'hf):(1'h0)] reg2090 = (1'h0);
  reg [(4'h9):(1'h0)] reg2089 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2088 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2087 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2086 = (1'h0);
  reg [(3'h4):(1'h0)] reg2066 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2058 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2056 = (1'h0);
  reg [(4'he):(1'h0)] reg2055 = (1'h0);
  reg [(4'hd):(1'h0)] reg2085 = (1'h0);
  reg [(3'h6):(1'h0)] reg2084 = (1'h0);
  reg [(4'he):(1'h0)] reg2083 = (1'h0);
  reg [(5'h10):(1'h0)] reg2082 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2081 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2078 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2077 = (1'h0);
  reg [(4'hf):(1'h0)] reg2075 = (1'h0);
  reg [(4'hf):(1'h0)] reg2080 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2079 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2078 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2077 = (1'h0);
  reg [(4'hd):(1'h0)] reg2076 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2075 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2074 = (1'h0);
  reg [(3'h4):(1'h0)] reg2073 = (1'h0);
  reg [(4'ha):(1'h0)] reg2072 = (1'h0);
  reg [(4'ha):(1'h0)] reg2071 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2070 = (1'h0);
  reg [(4'hf):(1'h0)] reg2069 = (1'h0);
  reg [(4'he):(1'h0)] forvar2068 = (1'h0);
  reg [(2'h2):(1'h0)] reg2067 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2066 = (1'h0);
  reg [(2'h2):(1'h0)] reg2065 = (1'h0);
  reg [(3'h5):(1'h0)] reg2064 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2063 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2062 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2061 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2060 = (1'h0);
  reg [(4'ha):(1'h0)] reg2059 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2058 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2057 = (1'h0);
  reg [(4'h9):(1'h0)] reg2056 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2055 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2054 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2053 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2052 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2051 = (1'h0);
  reg [(4'hc):(1'h0)] reg2050 = (1'h0);
  reg [(4'ha):(1'h0)] reg2049 = (1'h0);
  reg [(4'hc):(1'h0)] reg2047 = (1'h0);
  reg [(4'h8):(1'h0)] reg2048 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2047 = (1'h0);
  reg [(4'hd):(1'h0)] reg2046 = (1'h0);
  reg [(3'h5):(1'h0)] reg2045 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2044 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2043 = (1'h0);
  reg [(2'h3):(1'h0)] reg2042 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2041 = (1'h0);
  reg [(3'h4):(1'h0)] reg2040 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2039 = (1'h0);
  reg [(4'hd):(1'h0)] reg2038 = (1'h0);
  reg [(2'h2):(1'h0)] reg2037 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2036 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2035 = (1'h0);
  reg [(5'h10):(1'h0)] reg2034 = (1'h0);
  reg [(4'h9):(1'h0)] reg2033 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2030 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2028 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2023 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2017 = (1'h0);
  reg [(4'he):(1'h0)] reg2032 = (1'h0);
  reg [(4'hf):(1'h0)] reg2031 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2030 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2029 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2024 = (1'h0);
  reg [(3'h5):(1'h0)] reg2022 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2021 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2028 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2027 = (1'h0);
  reg [(4'hc):(1'h0)] reg2026 = (1'h0);
  reg [(4'ha):(1'h0)] reg2025 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2024 = (1'h0);
  reg [(4'hc):(1'h0)] reg2023 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2022 = (1'h0);
  reg [(4'ha):(1'h0)] reg2021 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2020 = (1'h0);
  reg [(4'hf):(1'h0)] reg2019 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2015 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2009 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2018 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2014 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2010 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2017 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2016 = (1'h0);
  reg [(4'ha):(1'h0)] reg2015 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2014 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2013 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2012 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2011 = (1'h0);
  reg [(4'h8):(1'h0)] reg2010 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2009 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2008 = (1'h0);
  wire [(2'h2):(1'h0)] wire2007;
  reg signed [(3'h4):(1'h0)] reg2006 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2005 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2004 = (1'h0);
  reg [(3'h7):(1'h0)] reg2003 = (1'h0);
  reg [(4'ha):(1'h0)] reg2002 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2001 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2000 = (1'h0);
  reg [(4'hf):(1'h0)] reg1999 = (1'h0);
  reg [(4'hc):(1'h0)] reg1998 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1997 = (1'h0);
  reg [(4'ha):(1'h0)] reg1996 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1995 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1994 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1993 = (1'h0);
  reg [(3'h7):(1'h0)] reg1992 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1991 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1990 = (1'h0);
  reg [(3'h5):(1'h0)] reg1989 = (1'h0);
  reg [(3'h6):(1'h0)] reg1988 = (1'h0);
  reg [(4'hd):(1'h0)] reg1987 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1986 = (1'h0);
  reg [(3'h5):(1'h0)] reg1985 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1984 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1983 = (1'h0);
  reg [(4'h8):(1'h0)] reg1982 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1981 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1980 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1979 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1978 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1977 = (1'h0);
  reg [(4'hb):(1'h0)] reg1976 = (1'h0);
  reg [(5'h10):(1'h0)] reg1975 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1974 = (1'h0);
  reg [(3'h5):(1'h0)] reg1973 = (1'h0);
  reg [(4'h9):(1'h0)] reg1972 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1971 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1964 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1970 = (1'h0);
  reg [(5'h10):(1'h0)] reg1969 = (1'h0);
  reg [(3'h6):(1'h0)] reg1968 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1967 = (1'h0);
  reg [(2'h3):(1'h0)] reg1966 = (1'h0);
  reg [(4'hc):(1'h0)] reg1965 = (1'h0);
  reg [(3'h4):(1'h0)] reg1964 = (1'h0);
  reg [(4'he):(1'h0)] forvar1963 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1962 = (1'h0);
  reg [(4'hf):(1'h0)] reg1961 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1960 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1959 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1958 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1957 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1956 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1955 = (1'h0);
  reg [(4'hb):(1'h0)] reg1954 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1953 = (1'h0);
  reg [(4'hb):(1'h0)] reg1952 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1951 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1950 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1949 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1948 = (1'h0);
  reg [(5'h10):(1'h0)] reg1947 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1946 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1945 = (1'h0);
  reg [(3'h6):(1'h0)] reg1944 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1943 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1942 = (1'h0);
  reg [(5'h10):(1'h0)] reg1941 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1940 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1939 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1939 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1938 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1937 = (1'h0);
  reg [(2'h3):(1'h0)] reg1936 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1935 = (1'h0);
  reg [(3'h4):(1'h0)] reg1934 = (1'h0);
  reg [(3'h5):(1'h0)] reg1933 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1932 = (1'h0);
  reg [(4'hd):(1'h0)] reg1931 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1930 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1929 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1928 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1927 = (1'h0);
  reg [(3'h7):(1'h0)] reg1926 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1925 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1924 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1923 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1922 = (1'h0);
  reg [(3'h5):(1'h0)] reg1905 = (1'h0);
  reg [(4'hf):(1'h0)] reg1904 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1914 = (1'h0);
  reg [(4'hc):(1'h0)] reg1921 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1920 = (1'h0);
  reg [(3'h7):(1'h0)] reg1919 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1918 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1917 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1916 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1915 = (1'h0);
  reg [(2'h3):(1'h0)] reg1914 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1913 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1912 = (1'h0);
  reg [(3'h5):(1'h0)] reg1911 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1910 = (1'h0);
  reg [(5'h10):(1'h0)] reg1909 = (1'h0);
  reg [(4'h9):(1'h0)] reg1908 = (1'h0);
  reg [(4'h9):(1'h0)] reg1907 = (1'h0);
  reg [(3'h5):(1'h0)] reg1906 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1905 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1904 = (1'h0);
  reg [(3'h4):(1'h0)] reg1903 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1902 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1901 = (1'h0);
  reg [(4'hc):(1'h0)] reg1900 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1899 = (1'h0);
  reg [(4'h8):(1'h0)] reg1898 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1897 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1896 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1894 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1891 = (1'h0);
  reg [(4'hf):(1'h0)] reg1895 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1894 = (1'h0);
  reg [(3'h4):(1'h0)] reg1893 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1892 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1891 = (1'h0);
  reg [(2'h3):(1'h0)] reg1880 = (1'h0);
  reg [(4'h9):(1'h0)] reg1890 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1889 = (1'h0);
  reg [(3'h6):(1'h0)] reg1888 = (1'h0);
  reg [(3'h7):(1'h0)] reg1887 = (1'h0);
  reg [(4'hc):(1'h0)] reg1886 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1885 = (1'h0);
  reg [(3'h5):(1'h0)] reg1884 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1883 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1882 = (1'h0);
  reg [(4'hc):(1'h0)] reg1881 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1880 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1879 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1878 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1877 = (1'h0);
  reg [(4'hf):(1'h0)] reg1876 = (1'h0);
  reg [(4'he):(1'h0)] forvar1875 = (1'h0);
  reg [(3'h4):(1'h0)] reg1874 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1873 = (1'h0);
  reg [(2'h2):(1'h0)] reg1872 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1871 = (1'h0);
  reg [(4'he):(1'h0)] reg1870 = (1'h0);
  reg [(3'h7):(1'h0)] reg1869 = (1'h0);
  reg [(2'h2):(1'h0)] reg1868 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1867 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1866 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1865 = (1'h0);
  reg [(4'he):(1'h0)] reg1864 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1863 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1862 = (1'h0);
  reg [(3'h5):(1'h0)] reg1861 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1860 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1859 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1858 = (1'h0);
  reg [(4'hc):(1'h0)] reg1856 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1850 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1857 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1856 = (1'h0);
  reg [(2'h2):(1'h0)] reg1855 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1854 = (1'h0);
  reg [(5'h10):(1'h0)] reg1853 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1852 = (1'h0);
  reg [(2'h3):(1'h0)] reg1851 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1850 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1849 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1845 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1844 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1840 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1836 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1848 = (1'h0);
  reg [(2'h3):(1'h0)] reg1847 = (1'h0);
  reg [(4'hd):(1'h0)] reg1846 = (1'h0);
  reg [(5'h10):(1'h0)] reg1845 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1844 = (1'h0);
  reg [(3'h6):(1'h0)] reg1843 = (1'h0);
  reg [(3'h6):(1'h0)] reg1842 = (1'h0);
  reg [(2'h2):(1'h0)] reg1841 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1840 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1839 = (1'h0);
  reg [(5'h10):(1'h0)] reg1838 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1837 = (1'h0);
  reg [(4'hb):(1'h0)] reg1836 = (1'h0);
  reg [(3'h7):(1'h0)] reg1835 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1834 = (1'h0);
  reg [(4'h8):(1'h0)] reg1833 = (1'h0);
  reg [(3'h5):(1'h0)] reg1832 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1831 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1830 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1829 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1828 = (1'h0);
  reg [(4'hc):(1'h0)] reg1827 = (1'h0);
  reg [(4'h9):(1'h0)] reg1820 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1826 = (1'h0);
  reg [(4'hc):(1'h0)] reg1825 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1823 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1821 = (1'h0);
  reg [(4'hc):(1'h0)] reg1824 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1823 = (1'h0);
  reg [(3'h4):(1'h0)] reg1822 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1821 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1820 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1819 = (1'h0);
  reg [(4'hc):(1'h0)] reg1818 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1817 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1816 = (1'h0);
  reg [(4'hf):(1'h0)] reg1815 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1814 = (1'h0);
  reg [(4'hb):(1'h0)] reg1813 = (1'h0);
  reg [(4'h9):(1'h0)] reg1812 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1811 = (1'h0);
  reg [(4'hf):(1'h0)] reg1810 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1809 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1808 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1803 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1801 = (1'h0);
  reg [(3'h6):(1'h0)] reg1800 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1798 = (1'h0);
  reg [(3'h5):(1'h0)] reg1807 = (1'h0);
  reg [(3'h7):(1'h0)] reg1806 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1805 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1804 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1803 = (1'h0);
  reg [(4'hf):(1'h0)] reg1802 = (1'h0);
  reg [(4'hf):(1'h0)] reg1801 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1800 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1799 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1798 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1797 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1796 = (1'h0);
  reg [(2'h2):(1'h0)] reg1795 = (1'h0);
  reg [(4'hc):(1'h0)] reg1794 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1793 = (1'h0);
  reg [(2'h3):(1'h0)] reg1792 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1791 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1790 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1789 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1788 = (1'h0);
  reg [(3'h5):(1'h0)] reg1787 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1786 = (1'h0);
  reg [(3'h4):(1'h0)] reg1785 = (1'h0);
  reg [(4'hb):(1'h0)] reg1784 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1783 = (1'h0);
  reg [(3'h5):(1'h0)] reg1782 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1781 = (1'h0);
  reg [(3'h6):(1'h0)] reg1780 = (1'h0);
  reg [(2'h2):(1'h0)] reg1776 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1775 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1773 = (1'h0);
  reg [(2'h3):(1'h0)] reg1779 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1778 = (1'h0);
  reg [(2'h2):(1'h0)] reg1777 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1776 = (1'h0);
  reg [(3'h6):(1'h0)] reg1775 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1774 = (1'h0);
  reg [(3'h6):(1'h0)] reg1773 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1772 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1771 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1770 = (1'h0);
  reg [(3'h5):(1'h0)] reg1769 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1768 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1767 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1766 = (1'h0);
  reg [(4'he):(1'h0)] reg1765 = (1'h0);
  reg [(2'h2):(1'h0)] reg1764 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1763 = (1'h0);
  reg [(3'h4):(1'h0)] reg1762 = (1'h0);
  reg [(5'h10):(1'h0)] reg1761 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1760 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1759 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1758 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1757 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire3037;
  wire signed [(4'hd):(1'h0)] wire3038;
  wire signed [(4'hf):(1'h0)] wire3529;
  assign y = {wire3531,
                 wire3035,
                 wire2360,
                 wire2359,
                 wire2358,
                 wire2357,
                 wire2356,
                 wire2355,
                 wire2354,
                 reg2353,
                 reg2352,
                 reg2342,
                 forvar2341,
                 reg2339,
                 forvar2336,
                 reg2351,
                 reg2350,
                 reg2349,
                 reg2348,
                 forvar2347,
                 reg2346,
                 reg2345,
                 reg2344,
                 reg2343,
                 forvar2342,
                 reg2341,
                 reg2340,
                 forvar2339,
                 reg2338,
                 reg2337,
                 reg2336,
                 reg2335,
                 forvar2334,
                 reg2333,
                 reg2332,
                 reg2331,
                 reg2330,
                 reg2329,
                 reg2328,
                 forvar2327,
                 reg2326,
                 reg2325,
                 reg2324,
                 reg2323,
                 forvar2322,
                 forvar2321,
                 forvar2320,
                 reg2319,
                 reg2318,
                 forvar2317,
                 reg2316,
                 reg2315,
                 reg2314,
                 reg2313,
                 forvar2312,
                 reg2311,
                 reg2310,
                 reg2309,
                 reg2307,
                 forvar2301,
                 forvar2289,
                 forvar2288,
                 forvar2291,
                 reg2290,
                 reg2287,
                 reg2308,
                 forvar2307,
                 reg2305,
                 reg2306,
                 forvar2305,
                 reg2304,
                 reg2303,
                 forvar2302,
                 reg2301,
                 forvar2300,
                 reg2299,
                 reg2298,
                 reg2297,
                 reg2296,
                 reg2295,
                 reg2294,
                 reg2293,
                 reg2292,
                 reg2291,
                 forvar2290,
                 reg2289,
                 reg2288,
                 forvar2287,
                 reg2232,
                 forvar2230,
                 reg2227,
                 forvar2225,
                 forvar2220,
                 forvar2216,
                 reg2209,
                 forvar2208,
                 forvar2207,
                 forvar2202,
                 reg2203,
                 forvar2201,
                 reg2200,
                 forvar2195,
                 forvar2187,
                 forvar2188,
                 reg2185,
                 forvar2183,
                 forvar2173,
                 reg2180,
                 reg2179,
                 reg2177,
                 forvar2170,
                 reg2168,
                 reg2286,
                 reg2285,
                 reg2284,
                 forvar2283,
                 reg2282,
                 reg2281,
                 reg2280,
                 reg2279,
                 reg2278,
                 reg2277,
                 forvar2276,
                 forvar2275,
                 reg2269,
                 forvar2268,
                 reg2265,
                 reg2264,
                 forvar2263,
                 forvar2262,
                 forvar2255,
                 reg2256,
                 reg2252,
                 reg2248,
                 forvar2247,
                 reg2274,
                 reg2273,
                 reg2272,
                 reg2271,
                 reg2270,
                 forvar2269,
                 reg2268,
                 reg2267,
                 reg2266,
                 forvar2265,
                 forvar2264,
                 reg2263,
                 reg2262,
                 reg2261,
                 reg2260,
                 reg2259,
                 reg2258,
                 reg2257,
                 forvar2256,
                 reg2255,
                 reg2254,
                 reg2253,
                 forvar2252,
                 reg2243,
                 forvar2242,
                 reg2241,
                 reg2251,
                 reg2250,
                 reg2249,
                 forvar2248,
                 reg2247,
                 reg2246,
                 reg2245,
                 reg2244,
                 forvar2243,
                 reg2242,
                 forvar2241,
                 reg2240,
                 reg2239,
                 reg2238,
                 reg2237,
                 forvar2236,
                 reg2235,
                 reg2234,
                 reg2233,
                 forvar2232,
                 reg2231,
                 reg2230,
                 reg2229,
                 reg2228,
                 forvar2227,
                 reg2226,
                 reg2225,
                 reg2224,
                 forvar2221,
                 reg2223,
                 reg2222,
                 reg2221,
                 reg2220,
                 reg2219,
                 reg2218,
                 reg2217,
                 reg2214,
                 reg2216,
                 reg2215,
                 forvar2214,
                 reg2211,
                 reg2213,
                 reg2212,
                 forvar2211,
                 reg2210,
                 forvar2209,
                 reg2208,
                 forvar2175,
                 reg2169,
                 reg2207,
                 reg2206,
                 reg2205,
                 reg2204,
                 forvar2203,
                 reg2202,
                 reg2201,
                 forvar2200,
                 reg2199,
                 reg2198,
                 reg2197,
                 forvar2196,
                 reg2191,
                 forvar2190,
                 reg2195,
                 reg2194,
                 reg2193,
                 reg2192,
                 forvar2191,
                 reg2190,
                 reg2189,
                 reg2188,
                 reg2187,
                 reg2186,
                 forvar2185,
                 reg2184,
                 reg2183,
                 reg2182,
                 reg2181,
                 forvar2180,
                 forvar2179,
                 reg2178,
                 forvar2177,
                 reg2176,
                 reg2175,
                 reg2174,
                 reg2173,
                 reg2172,
                 reg2171,
                 reg2170,
                 forvar2169,
                 forvar2168,
                 forvar2135,
                 reg2131,
                 forvar2130,
                 reg2124,
                 reg2121,
                 forvar2119,
                 forvar2117,
                 reg2113,
                 forvar2112,
                 forvar2111,
                 reg2109,
                 reg2167,
                 reg2166,
                 reg2165,
                 reg2164,
                 reg2163,
                 reg2162,
                 forvar2161,
                 reg2160,
                 reg2159,
                 reg2158,
                 forvar2157,
                 forvar2156,
                 reg2150,
                 reg2148,
                 reg2143,
                 reg2155,
                 reg2154,
                 reg2153,
                 forvar2152,
                 reg2151,
                 forvar2150,
                 reg2149,
                 forvar2148,
                 reg2147,
                 reg2146,
                 reg2145,
                 reg2144,
                 forvar2143,
                 forvar2142,
                 reg2141,
                 forvar2140,
                 reg2139,
                 reg2138,
                 reg2137,
                 reg2136,
                 reg2135,
                 reg2134,
                 reg2133,
                 reg2132,
                 forvar2131,
                 reg2130,
                 reg2129,
                 reg2128,
                 forvar2127,
                 reg2126,
                 reg2125,
                 forvar2124,
                 forvar2123,
                 reg2122,
                 forvar2121,
                 reg2120,
                 reg2119,
                 reg2118,
                 reg2117,
                 reg2116,
                 reg2115,
                 reg2114,
                 forvar2113,
                 reg2112,
                 reg2111,
                 forvar2110,
                 forvar2109,
                 reg2087,
                 reg2108,
                 reg2107,
                 reg2106,
                 reg2105,
                 reg2104,
                 reg2102,
                 forvar2096,
                 reg2103,
                 forvar2102,
                 reg2101,
                 reg2100,
                 reg2099,
                 reg2098,
                 reg2097,
                 reg2096,
                 reg2093,
                 reg2095,
                 reg2094,
                 forvar2093,
                 reg2092,
                 reg2091,
                 reg2090,
                 reg2089,
                 forvar2088,
                 forvar2087,
                 forvar2086,
                 reg2066,
                 reg2058,
                 forvar2056,
                 reg2055,
                 reg2085,
                 reg2084,
                 reg2083,
                 reg2082,
                 forvar2081,
                 reg2078,
                 forvar2077,
                 reg2075,
                 reg2080,
                 reg2079,
                 forvar2078,
                 reg2077,
                 reg2076,
                 forvar2075,
                 reg2074,
                 reg2073,
                 reg2072,
                 reg2071,
                 reg2070,
                 reg2069,
                 forvar2068,
                 reg2067,
                 forvar2066,
                 reg2065,
                 reg2064,
                 forvar2063,
                 reg2062,
                 reg2061,
                 reg2060,
                 reg2059,
                 forvar2058,
                 reg2057,
                 reg2056,
                 forvar2055,
                 forvar2054,
                 reg2053,
                 reg2052,
                 forvar2051,
                 reg2050,
                 reg2049,
                 reg2047,
                 reg2048,
                 forvar2047,
                 reg2046,
                 reg2045,
                 forvar2044,
                 reg2043,
                 reg2042,
                 reg2041,
                 reg2040,
                 reg2039,
                 reg2038,
                 reg2037,
                 forvar2036,
                 forvar2035,
                 reg2034,
                 reg2033,
                 reg2030,
                 forvar2028,
                 forvar2023,
                 forvar2017,
                 reg2032,
                 reg2031,
                 forvar2030,
                 reg2029,
                 reg2024,
                 reg2022,
                 forvar2021,
                 reg2028,
                 reg2027,
                 reg2026,
                 reg2025,
                 forvar2024,
                 reg2023,
                 forvar2022,
                 reg2021,
                 reg2020,
                 reg2019,
                 forvar2015,
                 reg2009,
                 reg2018,
                 reg2014,
                 forvar2010,
                 reg2017,
                 reg2016,
                 reg2015,
                 forvar2014,
                 reg2013,
                 reg2012,
                 reg2011,
                 reg2010,
                 forvar2009,
                 reg2008,
                 wire2007,
                 reg2006,
                 reg2005,
                 reg2004,
                 reg2003,
                 reg2002,
                 reg2001,
                 reg2000,
                 reg1999,
                 reg1998,
                 forvar1997,
                 reg1996,
                 reg1995,
                 forvar1994,
                 forvar1993,
                 reg1992,
                 reg1991,
                 reg1990,
                 reg1989,
                 reg1988,
                 reg1987,
                 forvar1986,
                 reg1985,
                 forvar1984,
                 forvar1983,
                 reg1982,
                 reg1981,
                 reg1980,
                 reg1979,
                 reg1978,
                 forvar1977,
                 reg1976,
                 reg1975,
                 forvar1974,
                 reg1973,
                 reg1972,
                 reg1971,
                 forvar1964,
                 reg1970,
                 reg1969,
                 reg1968,
                 reg1967,
                 reg1966,
                 reg1965,
                 reg1964,
                 forvar1963,
                 reg1962,
                 reg1961,
                 reg1960,
                 reg1959,
                 forvar1958,
                 reg1957,
                 reg1956,
                 forvar1955,
                 reg1954,
                 reg1953,
                 reg1952,
                 forvar1951,
                 forvar1950,
                 reg1949,
                 reg1948,
                 reg1947,
                 forvar1946,
                 forvar1945,
                 reg1944,
                 reg1943,
                 forvar1942,
                 reg1941,
                 forvar1940,
                 forvar1939,
                 reg1939,
                 reg1938,
                 reg1937,
                 reg1936,
                 reg1935,
                 reg1934,
                 reg1933,
                 reg1932,
                 reg1931,
                 reg1930,
                 reg1929,
                 reg1928,
                 reg1927,
                 reg1926,
                 forvar1925,
                 forvar1924,
                 forvar1923,
                 forvar1922,
                 reg1905,
                 reg1904,
                 forvar1914,
                 reg1921,
                 forvar1920,
                 reg1919,
                 reg1918,
                 reg1917,
                 reg1916,
                 reg1915,
                 reg1914,
                 reg1913,
                 reg1912,
                 reg1911,
                 reg1910,
                 reg1909,
                 reg1908,
                 reg1907,
                 reg1906,
                 forvar1905,
                 forvar1904,
                 reg1903,
                 forvar1902,
                 forvar1901,
                 reg1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 forvar1896,
                 forvar1894,
                 forvar1891,
                 reg1895,
                 reg1894,
                 reg1893,
                 reg1892,
                 reg1891,
                 reg1880,
                 reg1890,
                 forvar1889,
                 reg1888,
                 reg1887,
                 reg1886,
                 forvar1885,
                 reg1884,
                 reg1883,
                 reg1882,
                 reg1881,
                 forvar1880,
                 forvar1879,
                 forvar1878,
                 reg1877,
                 reg1876,
                 forvar1875,
                 reg1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 reg1870,
                 reg1869,
                 reg1868,
                 forvar1867,
                 reg1866,
                 forvar1865,
                 reg1864,
                 forvar1863,
                 reg1862,
                 reg1861,
                 reg1860,
                 reg1859,
                 forvar1858,
                 reg1856,
                 forvar1850,
                 reg1857,
                 forvar1856,
                 reg1855,
                 forvar1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 reg1850,
                 reg1849,
                 forvar1845,
                 reg1844,
                 forvar1840,
                 forvar1836,
                 reg1848,
                 reg1847,
                 reg1846,
                 reg1845,
                 forvar1844,
                 reg1843,
                 reg1842,
                 reg1841,
                 reg1840,
                 reg1839,
                 reg1838,
                 reg1837,
                 reg1836,
                 reg1835,
                 forvar1834,
                 reg1833,
                 reg1832,
                 reg1831,
                 reg1830,
                 reg1829,
                 forvar1828,
                 reg1827,
                 reg1820,
                 reg1826,
                 reg1825,
                 reg1823,
                 reg1821,
                 reg1824,
                 forvar1823,
                 reg1822,
                 forvar1821,
                 forvar1820,
                 reg1819,
                 reg1818,
                 forvar1817,
                 reg1816,
                 reg1815,
                 reg1814,
                 reg1813,
                 reg1812,
                 reg1811,
                 reg1810,
                 forvar1809,
                 forvar1808,
                 forvar1803,
                 forvar1801,
                 reg1800,
                 forvar1798,
                 reg1807,
                 reg1806,
                 reg1805,
                 reg1804,
                 reg1803,
                 reg1802,
                 reg1801,
                 forvar1800,
                 forvar1799,
                 reg1798,
                 forvar1797,
                 reg1796,
                 reg1795,
                 reg1794,
                 reg1793,
                 reg1792,
                 reg1791,
                 forvar1790,
                 reg1789,
                 forvar1788,
                 reg1787,
                 forvar1786,
                 reg1785,
                 reg1784,
                 reg1783,
                 reg1782,
                 forvar1781,
                 reg1780,
                 reg1776,
                 forvar1775,
                 forvar1773,
                 reg1779,
                 reg1778,
                 reg1777,
                 forvar1776,
                 reg1775,
                 reg1774,
                 reg1773,
                 reg1772,
                 reg1771,
                 reg1770,
                 reg1769,
                 forvar1768,
                 reg1767,
                 reg1766,
                 reg1765,
                 reg1764,
                 reg1763,
                 reg1762,
                 reg1761,
                 forvar1760,
                 forvar1759,
                 forvar1758,
                 forvar1757,
                 wire3037,
                 wire3038,
                 wire3529,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1757 = (1'h0); (forvar1757 < (2'h3)); forvar1757 = (forvar1757 + (1'h1)))
        begin
          for (forvar1758 = (1'h0); (forvar1758 < (1'h0)); forvar1758 = (forvar1758 + (1'h1)))
            begin
              for (forvar1759 = (1'h0); (forvar1759 < (2'h3)); forvar1759 = (forvar1759 + (1'h1)))
                begin
                  for (forvar1760 = (1'h0); (forvar1760 < (2'h3)); forvar1760 = (forvar1760 + (1'h1)))
                    begin
                      reg1761 <= {forvar1758[(2'h2):(2'h2)]};
                      reg1762 <= $signed({forvar1757});
                      reg1763 <= wire1753[(4'h8):(1'h1)];
                      reg1764 <= ($unsigned(reg1761) ?
                          forvar1759 : (-(forvar1760 ?
                              (reg1763 ? forvar1757 : forvar1760) : (8'hb9))));
                    end
                  if ((|$signed(($signed(wire1754) ?
                      (forvar1758 ?
                          wire1754 : forvar1759) : wire1753[(3'h4):(2'h3)]))))
                    begin
                      reg1765 <= forvar1757[(4'h9):(3'h5)];
                      reg1766 <= (~&wire1755[(2'h3):(1'h1)]);
                      reg1767 <= (wire1754[(3'h5):(3'h5)] >= ({(|(8'hb2))} ~^ ({(8'had)} ^~ $unsigned(wire1753))));
                    end
                  else
                    begin
                      reg1765 <= $unsigned(reg1767[(4'ha):(3'h5)]);
                      reg1766 <= ((forvar1758[(1'h0):(1'h0)] ?
                              (&(-wire1754)) : reg1762) ?
                          wire1756[(2'h2):(1'h0)] : $unsigned(wire1755));
                      reg1767 <= ((reg1763[(1'h0):(1'h0)] ^~ ($unsigned(forvar1760) ?
                              (reg1762 != wire1755) : reg1761)) ?
                          reg1766 : wire1755);
                    end
                  for (forvar1768 = (1'h0); (forvar1768 < (1'h0)); forvar1768 = (forvar1768 + (1'h1)))
                    begin
                      reg1769 <= (((8'hb3) <= reg1766[(2'h2):(2'h2)]) ?
                          ((~$unsigned(reg1764)) ?
                              $unsigned($unsigned(forvar1757)) : $signed((!reg1764))) : forvar1760[(2'h3):(2'h2)]);
                      reg1770 <= ($signed((~$unsigned((8'ha3)))) == forvar1760[(1'h0):(1'h0)]);
                      reg1771 <= (^($signed($signed(forvar1757)) != reg1767[(4'hc):(4'h9)]));
                    end
                end
              reg1772 <= (reg1761[(2'h3):(2'h3)] ^~ $unsigned($signed((8'hba))));
              if ($unsigned(reg1769))
                begin
                  if (reg1770)
                    begin
                      reg1773 <= $signed(((~&(reg1769 >= wire1756)) ?
                          ((^~wire1755) <<< reg1770[(3'h7):(3'h7)]) : reg1771[(2'h3):(2'h2)]));
                      reg1774 <= reg1761[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg1773 <= reg1769[(1'h1):(1'h0)];
                      reg1774 <= forvar1768;
                      reg1775 <= reg1763;
                    end
                  for (forvar1776 = (1'h0); (forvar1776 < (2'h3)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 <= {$signed(wire1754)};
                      reg1778 <= reg1761[(2'h2):(1'h0)];
                      reg1779 <= ((~^((~|reg1762) ?
                              $signed(wire1755) : (-wire1754))) ?
                          ((&$signed(wire1755)) & {$signed(reg1763)}) : forvar1757);
                    end
                end
              else
                begin
                  for (forvar1773 = (1'h0); (forvar1773 < (1'h1)); forvar1773 = (forvar1773 + (1'h1)))
                    begin
                      reg1774 <= ($signed($signed(wire1753[(1'h1):(1'h1)])) >> {((forvar1773 ?
                              reg1766 : (8'hb4)) ^ (reg1770 ?
                              reg1764 : reg1765))});
                    end
                  for (forvar1775 = (1'h0); (forvar1775 < (2'h3)); forvar1775 = (forvar1775 + (1'h1)))
                    begin
                      reg1776 <= reg1765;
                      reg1777 <= reg1779[(2'h2):(2'h2)];
                      reg1778 <= reg1771;
                      reg1779 <= ((($unsigned(reg1769) == (wire1753 ?
                              reg1763 : forvar1776)) ?
                          $signed((reg1771 || reg1776)) : (reg1769[(2'h3):(2'h2)] ?
                              $unsigned(wire1756) : ((8'hb4) | forvar1758))) | {(reg1767[(3'h7):(3'h4)] ?
                              $unsigned(forvar1759) : (reg1769 ^~ (8'ha6)))});
                    end
                  reg1780 <= $unsigned({$unsigned((8'had))});
                end
              for (forvar1781 = (1'h0); (forvar1781 < (1'h1)); forvar1781 = (forvar1781 + (1'h1)))
                begin
                  if ($unsigned(reg1764))
                    begin
                      reg1782 <= (8'haf);
                      reg1783 <= wire1755[(2'h3):(1'h1)];
                      reg1784 <= $signed($unsigned($unsigned($signed(wire1753))));
                      reg1785 <= $signed((~$unsigned($unsigned(reg1761))));
                    end
                  else
                    begin
                      reg1782 <= ((~^((reg1782 - reg1779) ?
                              $signed(reg1771) : $signed(wire1756))) ?
                          (reg1776[(2'h2):(2'h2)] <= {reg1761}) : $signed((&((8'ha5) ~^ forvar1768))));
                      reg1783 <= ($signed($signed((reg1762 > reg1776))) ?
                          ({{(8'hb2)}} >>> $signed((^~forvar1759))) : reg1780[(2'h2):(2'h2)]);
                      reg1784 <= $signed($signed($signed((!reg1774))));
                      reg1785 <= forvar1757[(3'h7):(3'h5)];
                    end
                  for (forvar1786 = (1'h0); (forvar1786 < (1'h1)); forvar1786 = (forvar1786 + (1'h1)))
                    begin
                      reg1787 <= $signed({(+wire1753)});
                    end
                end
            end
          for (forvar1788 = (1'h0); (forvar1788 < (1'h1)); forvar1788 = (forvar1788 + (1'h1)))
            begin
              reg1789 <= ($unsigned((~|{reg1761})) < $unsigned(((~^(8'ha6)) ^ (~^wire1754))));
              for (forvar1790 = (1'h0); (forvar1790 < (2'h2)); forvar1790 = (forvar1790 + (1'h1)))
                begin
                  if ((^~forvar1776))
                    begin
                      reg1791 <= {(!reg1770)};
                    end
                  else
                    begin
                      reg1791 <= $signed(forvar1758);
                      reg1792 <= (-($signed((reg1763 <<< reg1779)) + ($unsigned(forvar1760) && {reg1783})));
                      reg1793 <= $signed((+(8'ha6)));
                      reg1794 <= ((($signed(forvar1790) ?
                              $signed(forvar1768) : ((8'ha4) ?
                                  forvar1788 : wire1753)) | forvar1773) ?
                          $signed($signed((+wire1756))) : reg1772);
                    end
                  reg1795 <= (($unsigned(reg1775) && $unsigned((&reg1769))) > ($unsigned(reg1785[(1'h1):(1'h0)]) ?
                      $signed((8'hb6)) : {(forvar1773 * (8'hb9))}));
                end
            end
          reg1796 <= forvar1768[(2'h2):(1'h0)];
        end
      if (reg1794)
        begin
          for (forvar1797 = (1'h0); (forvar1797 < (1'h1)); forvar1797 = (forvar1797 + (1'h1)))
            begin
              reg1798 <= reg1780[(3'h5):(1'h1)];
              for (forvar1799 = (1'h0); (forvar1799 < (1'h0)); forvar1799 = (forvar1799 + (1'h1)))
                begin
                  for (forvar1800 = (1'h0); (forvar1800 < (1'h1)); forvar1800 = (forvar1800 + (1'h1)))
                    begin
                      reg1801 <= ($signed($signed((forvar1790 ?
                          forvar1759 : wire1753))) - $unsigned($unsigned((~&reg1785))));
                      reg1802 <= (reg1761 ?
                          $unsigned(($signed(wire1755) ?
                              (reg1763 ?
                                  reg1764 : (8'ha0)) : (forvar1799 ~^ forvar1797))) : ((~((8'h9d) ?
                                  (8'haf) : forvar1775)) ?
                              wire1756 : $signed((|reg1787))));
                      reg1803 <= ({(~&$signed(reg1791))} ?
                          $signed((forvar1781 - (reg1795 || (8'h9e)))) : {$unsigned($unsigned((8'hb2)))});
                    end
                  if ($unsigned(reg1789[(3'h5):(3'h5)]))
                    begin
                      reg1804 <= wire1754;
                      reg1805 <= (reg1782 >= (~((^~reg1796) << (+reg1764))));
                    end
                  else
                    begin
                      reg1804 <= (-($unsigned($unsigned(reg1773)) ?
                          ($signed((8'h9c)) & $signed(reg1774)) : (^~wire1753)));
                      reg1805 <= ((forvar1757[(2'h3):(2'h2)] ?
                          forvar1800[(4'hc):(1'h0)] : $signed($signed((8'h9c)))) - (($signed(reg1764) & reg1804) ?
                          $unsigned((reg1801 ?
                              forvar1773 : forvar1790)) : (~{forvar1800})));
                      reg1806 <= (~^{(~^(wire1756 ? reg1774 : wire1753))});
                      reg1807 <= $signed($signed(reg1767));
                    end
                end
            end
        end
      else
        begin
          for (forvar1797 = (1'h0); (forvar1797 < (2'h3)); forvar1797 = (forvar1797 + (1'h1)))
            begin
              for (forvar1798 = (1'h0); (forvar1798 < (2'h2)); forvar1798 = (forvar1798 + (1'h1)))
                begin
                  for (forvar1799 = (1'h0); (forvar1799 < (2'h3)); forvar1799 = (forvar1799 + (1'h1)))
                    begin
                      reg1800 <= forvar1788;
                    end
                  for (forvar1801 = (1'h0); (forvar1801 < (2'h2)); forvar1801 = (forvar1801 + (1'h1)))
                    begin
                      reg1802 <= $signed(forvar1797);
                    end
                  for (forvar1803 = (1'h0); (forvar1803 < (2'h2)); forvar1803 = (forvar1803 + (1'h1)))
                    begin
                      reg1804 <= $unsigned($unsigned(forvar1776));
                    end
                  if ((8'ha1))
                    begin
                      reg1805 <= forvar1786;
                      reg1806 <= reg1794[(3'h5):(2'h3)];
                      reg1807 <= {(forvar1797[(3'h7):(3'h7)] ?
                              (~$unsigned(forvar1800)) : reg1796[(2'h2):(1'h0)])};
                    end
                  else
                    begin
                      reg1805 <= $signed((|reg1802[(4'hf):(1'h1)]));
                    end
                end
            end
          for (forvar1808 = (1'h0); (forvar1808 < (2'h3)); forvar1808 = (forvar1808 + (1'h1)))
            begin
              for (forvar1809 = (1'h0); (forvar1809 < (1'h0)); forvar1809 = (forvar1809 + (1'h1)))
                begin
                  if ((|((^(~&reg1801)) ?
                      forvar1776[(3'h6):(3'h5)] : $signed((reg1798 ?
                          forvar1781 : reg1782)))))
                    begin
                      reg1810 <= forvar1808[(1'h1):(1'h0)];
                      reg1811 <= (-(8'ha9));
                      reg1812 <= (forvar1800 ?
                          $signed(($signed(wire1756) * (reg1762 && reg1776))) : ((~|(reg1770 ?
                                  (8'hba) : reg1785)) ?
                              ((reg1804 - forvar1757) & (forvar1788 ?
                                  forvar1760 : forvar1799)) : (~^(~^reg1793))));
                    end
                  else
                    begin
                      reg1810 <= forvar1799[(1'h1):(1'h1)];
                      reg1811 <= reg1765;
                      reg1812 <= $signed({(!$unsigned(reg1782))});
                    end
                  if ((8'hb4))
                    begin
                      reg1813 <= $signed(forvar1786[(1'h0):(1'h0)]);
                      reg1814 <= reg1761;
                      reg1815 <= reg1806[(2'h3):(2'h3)];
                      reg1816 <= reg1796[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1813 <= reg1764[(1'h1):(1'h0)];
                      reg1814 <= (((reg1773[(3'h6):(3'h4)] ?
                          (forvar1775 ?
                              reg1770 : (8'hb7)) : (wire1756 != forvar1801)) >> $unsigned($unsigned(reg1766))) > ($unsigned($unsigned(reg1761)) ?
                          reg1771[(4'hc):(4'ha)] : $unsigned(reg1772)));
                      reg1815 <= {({(reg1762 >>> reg1816)} < (reg1810[(3'h7):(3'h5)] >= $signed(reg1787)))};
                      reg1816 <= ($signed(reg1770) | reg1771[(1'h1):(1'h0)]);
                    end
                end
            end
          for (forvar1817 = (1'h0); (forvar1817 < (2'h2)); forvar1817 = (forvar1817 + (1'h1)))
            begin
              reg1818 <= (|{{reg1766[(3'h7):(3'h6)]}});
              reg1819 <= (({$signed((8'ha7))} ? reg1811 : reg1806) ?
                  (($unsigned((8'hb5)) ? forvar1800 : (reg1784 > (8'hb4))) ?
                      $unsigned(reg1794[(4'ha):(1'h1)]) : forvar1773[(3'h5):(3'h5)]) : forvar1775[(3'h7):(3'h5)]);
            end
          if (reg1807)
            begin
              for (forvar1820 = (1'h0); (forvar1820 < (1'h0)); forvar1820 = (forvar1820 + (1'h1)))
                begin
                  for (forvar1821 = (1'h0); (forvar1821 < (1'h1)); forvar1821 = (forvar1821 + (1'h1)))
                    begin
                      reg1822 <= reg1771;
                    end
                end
              for (forvar1823 = (1'h0); (forvar1823 < (2'h3)); forvar1823 = (forvar1823 + (1'h1)))
                begin
                  if (((&(reg1784[(4'hb):(3'h6)] >= reg1777)) ?
                      (+{$unsigned(forvar1768)}) : $signed(forvar1820[(3'h5):(2'h3)])))
                    begin
                      reg1824 <= (|$unsigned(reg1762[(2'h3):(2'h2)]));
                    end
                  else
                    begin
                      reg1824 <= (wire1754 ?
                          $signed($unsigned(reg1791[(3'h5):(1'h0)])) : {$unsigned(reg1802[(2'h3):(1'h0)])});
                    end
                end
            end
          else
            begin
              if ((({$signed((8'hb0))} ?
                      ((forvar1821 ? reg1776 : (8'hae)) ?
                          (reg1775 == reg1764) : reg1767) : ((forvar1809 + forvar1775) ?
                          $unsigned(forvar1809) : (reg1818 ?
                              forvar1817 : forvar1821))) ?
                  {{$signed((8'ha0))}} : {{(^~forvar1757)}}))
                begin
                  for (forvar1820 = (1'h0); (forvar1820 < (2'h2)); forvar1820 = (forvar1820 + (1'h1)))
                    begin
                      reg1821 <= ((~|forvar1757[(4'h8):(2'h3)]) ?
                          (reg1804[(2'h3):(2'h2)] ^~ (~&forvar1758)) : $unsigned((8'had)));
                      reg1822 <= (~&reg1778[(3'h4):(1'h1)]);
                      reg1823 <= ($signed(reg1816[(3'h5):(2'h2)]) ?
                          $unsigned(reg1785[(2'h3):(1'h0)]) : forvar1801[(2'h3):(1'h0)]);
                      reg1824 <= $unsigned((forvar1773[(3'h4):(2'h2)] ?
                          reg1785 : $signed(forvar1776)));
                    end
                  reg1825 <= (&forvar1808);
                  reg1826 <= ($unsigned(forvar1821) ?
                      (~&$unsigned($unsigned(forvar1800))) : (reg1782[(2'h2):(1'h1)] ?
                          {(forvar1797 ?
                                  reg1805 : forvar1801)} : (&(reg1770 - reg1769))));
                end
              else
                begin
                  if (($signed($signed($unsigned(reg1766))) == reg1800[(2'h3):(1'h1)]))
                    begin
                      reg1820 <= $signed({(((8'hac) ?
                              (8'hb2) : wire1755) <= (^~forvar1798))});
                      reg1821 <= (reg1807[(1'h0):(1'h0)] ?
                          reg1784[(2'h3):(2'h2)] : reg1804);
                      reg1822 <= $unsigned((8'had));
                      reg1823 <= (((-(!reg1778)) ?
                              $signed(reg1803) : ((~&(8'h9c)) >= forvar1759)) ?
                          reg1815[(4'h8):(3'h7)] : $signed($signed((~forvar1759))));
                    end
                  else
                    begin
                      reg1820 <= ((|reg1820) ? reg1807 : {$unsigned(reg1776)});
                      reg1821 <= $signed({$signed(reg1782[(1'h0):(1'h0)])});
                    end
                  if ((forvar1760[(2'h2):(1'h0)] ?
                      (+{reg1792}) : ((!$signed(reg1763)) ?
                          (&(forvar1768 ?
                              forvar1823 : reg1798)) : ((forvar1820 ?
                              forvar1797 : (8'ha7)) | (&reg1787)))))
                    begin
                      reg1824 <= reg1795;
                      reg1825 <= (~$unsigned(reg1796[(1'h1):(1'h1)]));
                      reg1826 <= $unsigned($unsigned(reg1770[(4'ha):(3'h4)]));
                      reg1827 <= (wire1753[(2'h3):(2'h2)] <= $signed(({reg1811} ?
                          $unsigned((8'hb0)) : {forvar1817})));
                    end
                  else
                    begin
                      reg1824 <= ((|forvar1775) <<< ($unsigned($unsigned(forvar1781)) ?
                          (~$signed(wire1753)) : $unsigned((reg1784 ?
                              (8'ha2) : reg1824))));
                      reg1825 <= (^~(({forvar1776} >= (reg1818 && reg1818)) ^~ ((reg1801 || reg1818) ?
                          $signed(reg1794) : $signed(reg1761))));
                      reg1826 <= $unsigned(forvar1768);
                      reg1827 <= reg1792;
                    end
                end
              for (forvar1828 = (1'h0); (forvar1828 < (1'h0)); forvar1828 = (forvar1828 + (1'h1)))
                begin
                  reg1829 <= $signed((^~{(~forvar1823)}));
                  if (reg1794[(3'h5):(1'h0)])
                    begin
                      reg1830 <= ({($signed(wire1753) && $unsigned(reg1796))} ?
                          $unsigned(((forvar1760 ? (8'h9d) : (8'ha5)) ?
                              (reg1774 ?
                                  reg1767 : wire1754) : {forvar1808})) : $unsigned($unsigned({(8'ha6)})));
                      reg1831 <= ((((reg1824 ?
                                  reg1782 : (8'ha1)) == $unsigned(forvar1808)) ?
                              {reg1823} : $signed(reg1780[(2'h2):(1'h1)])) ?
                          (~&$unsigned(forvar1757[(2'h2):(1'h1)])) : reg1826);
                      reg1832 <= $unsigned(forvar1797);
                      reg1833 <= $unsigned($signed((~^forvar1800)));
                    end
                  else
                    begin
                      reg1830 <= forvar1797[(3'h7):(1'h1)];
                      reg1831 <= reg1778;
                      reg1832 <= $signed(((^$signed(forvar1821)) - reg1805[(4'h8):(1'h0)]));
                      reg1833 <= $signed((~(forvar1773 ?
                          {forvar1798} : $signed(forvar1817))));
                    end
                end
              if ((reg1782 < $unsigned($signed((!(8'ha7))))))
                begin
                  for (forvar1834 = (1'h0); (forvar1834 < (2'h2)); forvar1834 = (forvar1834 + (1'h1)))
                    begin
                      reg1835 <= reg1819[(2'h3):(2'h3)];
                      reg1836 <= (($signed((|reg1824)) ?
                              (-(~|reg1792)) : reg1804) ?
                          (-(-$signed(forvar1821))) : $unsigned($signed((reg1805 ?
                              reg1772 : reg1821))));
                    end
                  if ({$unsigned(forvar1786[(2'h2):(1'h0)])})
                    begin
                      reg1837 <= reg1787;
                    end
                  else
                    begin
                      reg1837 <= $unsigned((reg1830 ?
                          reg1766 : reg1822[(2'h2):(2'h2)]));
                      reg1838 <= $unsigned(((~(~^forvar1759)) ?
                          (reg1793 || $unsigned(reg1802)) : ($signed(reg1830) ?
                              (!(8'ha7)) : $signed(forvar1798))));
                      reg1839 <= {(($signed((8'hb3)) ?
                              $unsigned(reg1820) : $signed(forvar1809)) > $unsigned($unsigned(forvar1797)))};
                    end
                  if (({reg1793[(4'h8):(3'h5)]} ?
                      {(reg1764[(2'h2):(1'h0)] ?
                              reg1798[(1'h1):(1'h1)] : (|reg1764))} : (reg1826[(2'h3):(1'h0)] ?
                          ($unsigned((8'haa)) ?
                              (reg1785 ?
                                  wire1754 : forvar1760) : {reg1806}) : $signed((8'ha3)))))
                    begin
                      reg1840 <= reg1769[(3'h5):(1'h1)];
                      reg1841 <= (reg1838[(1'h0):(1'h0)] ~^ (reg1823 ?
                          wire1754 : {(forvar1759 ? (8'ha0) : reg1840)}));
                      reg1842 <= (((~&$unsigned(reg1816)) ^ $signed($signed(reg1829))) - ($unsigned(reg1806) + $signed(((8'hb5) ?
                          reg1800 : (8'hba)))));
                      reg1843 <= (~^(^$unsigned(reg1796[(3'h6):(1'h0)])));
                    end
                  else
                    begin
                      reg1840 <= {reg1801[(3'h5):(1'h0)]};
                      reg1841 <= (~^((^forvar1799[(4'h9):(2'h3)]) ?
                          ($unsigned(reg1839) * reg1806[(3'h7):(3'h7)]) : $signed((forvar1821 <= reg1815))));
                    end
                  for (forvar1844 = (1'h0); (forvar1844 < (1'h0)); forvar1844 = (forvar1844 + (1'h1)))
                    begin
                      reg1845 <= forvar1801;
                      reg1846 <= (~|reg1810[(3'h6):(3'h6)]);
                      reg1847 <= $signed((($unsigned((8'haf)) > {reg1796}) ^~ {{forvar1803}}));
                      reg1848 <= reg1806;
                    end
                end
              else
                begin
                  for (forvar1834 = (1'h0); (forvar1834 < (1'h0)); forvar1834 = (forvar1834 + (1'h1)))
                    begin
                      reg1835 <= $signed(reg1824[(4'ha):(1'h1)]);
                    end
                  for (forvar1836 = (1'h0); (forvar1836 < (1'h0)); forvar1836 = (forvar1836 + (1'h1)))
                    begin
                      reg1837 <= ({{$signed(reg1785)}} ?
                          forvar1820 : $signed(((forvar1759 ?
                              (8'h9e) : forvar1808) + $signed(reg1839))));
                      reg1838 <= (~&$unsigned($signed(reg1827)));
                      reg1839 <= (($signed(reg1816) >= reg1838[(4'hc):(4'h8)]) ?
                          $unsigned($signed(((8'hb2) == reg1764))) : reg1816[(3'h5):(1'h0)]);
                    end
                  for (forvar1840 = (1'h0); (forvar1840 < (2'h2)); forvar1840 = (forvar1840 + (1'h1)))
                    begin
                      reg1841 <= {($unsigned(reg1843) && reg1819)};
                      reg1842 <= $signed(((&{reg1815}) ?
                          (forvar1790 ?
                              (reg1770 << (8'hba)) : (~|reg1805)) : ($unsigned(reg1835) ?
                              $unsigned(reg1761) : {reg1847})));
                      reg1843 <= reg1798[(3'h7):(1'h1)];
                      reg1844 <= forvar1817;
                    end
                  for (forvar1845 = (1'h0); (forvar1845 < (2'h3)); forvar1845 = (forvar1845 + (1'h1)))
                    begin
                      reg1846 <= (reg1795[(1'h0):(1'h0)] && (reg1829 | $unsigned((~^reg1770))));
                      reg1847 <= reg1793[(3'h6):(3'h5)];
                      reg1848 <= $unsigned(reg1835[(3'h4):(1'h0)]);
                      reg1849 <= $unsigned((~($signed(forvar1790) ?
                          $signed(forvar1798) : $signed((8'ha6)))));
                    end
                end
              if (($unsigned($unsigned((forvar1758 ?
                  reg1820 : reg1823))) == forvar1836))
                begin
                  reg1850 <= $unsigned($signed(($unsigned(forvar1845) ?
                      (reg1795 ? reg1818 : reg1773) : (reg1830 > reg1796))));
                  if (forvar1776[(1'h0):(1'h0)])
                    begin
                      reg1851 <= $signed((($unsigned(wire1756) >= $signed(reg1827)) ?
                          reg1837[(2'h3):(1'h1)] : (~$signed((8'hb2)))));
                      reg1852 <= (forvar1799[(3'h7):(3'h5)] ?
                          {reg1779[(1'h1):(1'h0)]} : reg1846);
                    end
                  else
                    begin
                      reg1851 <= (reg1787 ^~ {(8'ha9)});
                      reg1852 <= (forvar1817 | (reg1764 ?
                          $unsigned(reg1822) : forvar1834));
                      reg1853 <= (~((+$unsigned(forvar1760)) ?
                          (-((8'ha8) ? forvar1823 : reg1826)) : forvar1788));
                    end
                  for (forvar1854 = (1'h0); (forvar1854 < (1'h0)); forvar1854 = (forvar1854 + (1'h1)))
                    begin
                      reg1855 <= $signed((({wire1755} + (reg1842 ?
                              reg1848 : reg1832)) ?
                          ((reg1777 ? (8'hab) : (8'ha7)) ?
                              reg1829[(1'h1):(1'h0)] : forvar1828[(4'hc):(1'h0)]) : reg1849[(3'h7):(3'h5)]));
                    end
                  for (forvar1856 = (1'h0); (forvar1856 < (2'h3)); forvar1856 = (forvar1856 + (1'h1)))
                    begin
                      reg1857 <= forvar1800;
                    end
                end
              else
                begin
                  for (forvar1850 = (1'h0); (forvar1850 < (2'h3)); forvar1850 = (forvar1850 + (1'h1)))
                    begin
                      reg1851 <= (~&{forvar1801});
                      reg1852 <= reg1857;
                      reg1853 <= ((($signed(reg1822) <<< ((8'haf) + reg1773)) ?
                              (-forvar1840[(3'h5):(1'h1)]) : forvar1768[(1'h0):(1'h0)]) ?
                          $unsigned(reg1777) : reg1811);
                    end
                  for (forvar1854 = (1'h0); (forvar1854 < (1'h0)); forvar1854 = (forvar1854 + (1'h1)))
                    begin
                      reg1855 <= $unsigned((~((~reg1814) * (~^reg1830))));
                      reg1856 <= ($unsigned((^~reg1802[(1'h0):(1'h0)])) ?
                          ($unsigned((reg1855 ?
                              (8'ha8) : reg1801)) >> reg1800[(2'h2):(1'h1)]) : ((~&(|(8'haa))) && (8'hb1)));
                      reg1857 <= reg1763;
                    end
                  for (forvar1858 = (1'h0); (forvar1858 < (1'h0)); forvar1858 = (forvar1858 + (1'h1)))
                    begin
                      reg1859 <= ((~{$signed(reg1806)}) - $unsigned((8'hac)));
                      reg1860 <= ($signed(reg1764[(2'h2):(1'h1)]) ?
                          $signed(reg1792) : reg1822[(1'h1):(1'h0)]);
                      reg1861 <= $unsigned($signed(reg1832));
                      reg1862 <= (+{((reg1771 ~^ reg1787) == (8'hba))});
                    end
                end
            end
        end
      for (forvar1863 = (1'h0); (forvar1863 < (1'h0)); forvar1863 = (forvar1863 + (1'h1)))
        begin
          reg1864 <= (^~(^~forvar1863[(4'he):(4'hd)]));
        end
    end
  always
    @(posedge clk) begin
      for (forvar1865 = (1'h0); (forvar1865 < (1'h0)); forvar1865 = (forvar1865 + (1'h1)))
        begin
          reg1866 <= reg1792;
          for (forvar1867 = (1'h0); (forvar1867 < (1'h0)); forvar1867 = (forvar1867 + (1'h1)))
            begin
              if (reg1784[(2'h3):(2'h2)])
                begin
                  if ($unsigned((((~&reg1770) >= (forvar1863 < (8'hb0))) ?
                      $unsigned((~|reg1856)) : reg1846[(4'h8):(2'h2)])))
                    begin
                      reg1868 <= forvar1768[(3'h5):(3'h5)];
                      reg1869 <= $unsigned($signed(((~^reg1818) == (forvar1865 ?
                          forvar1760 : reg1833))));
                      reg1870 <= $unsigned($signed(reg1774));
                    end
                  else
                    begin
                      reg1868 <= reg1769[(2'h3):(1'h1)];
                    end
                  if ((((8'hb3) << $signed((reg1836 && reg1775))) && reg1777[(2'h2):(1'h0)]))
                    begin
                      reg1871 <= $signed(reg1851);
                      reg1872 <= $signed(($unsigned((reg1775 >> (8'ha0))) ?
                          ({(8'ha7)} ?
                              $signed(reg1816) : forvar1865) : reg1770));
                      reg1873 <= $signed($unsigned(($unsigned(reg1811) * forvar1840)));
                      reg1874 <= (~^$signed($signed((8'ha4))));
                    end
                  else
                    begin
                      reg1871 <= (+(((~^reg1847) ?
                              (|forvar1809) : reg1847[(2'h2):(1'h1)]) ?
                          forvar1809 : forvar1786[(3'h6):(2'h3)]));
                      reg1872 <= {(|((~&forvar1788) ?
                              (~(8'ha4)) : $signed(reg1824)))};
                      reg1873 <= reg1845[(4'h9):(3'h5)];
                      reg1874 <= ($signed(reg1853[(4'ha):(1'h1)]) >>> reg1869[(1'h1):(1'h1)]);
                    end
                  for (forvar1875 = (1'h0); (forvar1875 < (2'h2)); forvar1875 = (forvar1875 + (1'h1)))
                    begin
                      reg1876 <= $unsigned(forvar1790);
                      reg1877 <= reg1873;
                    end
                end
              else
                begin
                  reg1868 <= $signed(reg1783);
                end
            end
        end
      for (forvar1878 = (1'h0); (forvar1878 < (2'h3)); forvar1878 = (forvar1878 + (1'h1)))
        begin
          for (forvar1879 = (1'h0); (forvar1879 < (1'h0)); forvar1879 = (forvar1879 + (1'h1)))
            begin
              if ($unsigned((reg1855 >> (reg1813 <<< (~reg1853)))))
                begin
                  for (forvar1880 = (1'h0); (forvar1880 < (2'h2)); forvar1880 = (forvar1880 + (1'h1)))
                    begin
                      reg1881 <= {reg1819};
                    end
                  if (forvar1801)
                    begin
                      reg1882 <= (~^({(+reg1870)} ?
                          $unsigned(reg1866) : $unsigned($signed(reg1774))));
                      reg1883 <= (reg1843[(2'h3):(1'h0)] == (reg1877[(3'h6):(2'h3)] <<< ($unsigned(forvar1768) ?
                          (^~reg1789) : $signed(reg1794))));
                      reg1884 <= (forvar1821[(2'h2):(1'h1)] ?
                          reg1791[(3'h6):(3'h6)] : {(^~reg1785)});
                    end
                  else
                    begin
                      reg1882 <= (^reg1766);
                      reg1883 <= {($unsigned((^reg1803)) < (~|reg1884))};
                      reg1884 <= reg1772[(1'h0):(1'h0)];
                    end
                  for (forvar1885 = (1'h0); (forvar1885 < (2'h2)); forvar1885 = (forvar1885 + (1'h1)))
                    begin
                      reg1886 <= $signed((+(!(reg1836 == wire1756))));
                      reg1887 <= $unsigned($signed($unsigned(forvar1856[(4'hb):(1'h1)])));
                      reg1888 <= (!((reg1850[(2'h2):(1'h0)] - $unsigned(reg1826)) ?
                          forvar1854[(3'h5):(1'h0)] : reg1796));
                    end
                  for (forvar1889 = (1'h0); (forvar1889 < (2'h2)); forvar1889 = (forvar1889 + (1'h1)))
                    begin
                      reg1890 <= reg1829[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  reg1880 <= (~&$signed($unsigned((+forvar1844))));
                end
            end
          if (($unsigned(reg1762[(2'h2):(2'h2)]) ^~ (({forvar1758} ?
              ((8'hb0) * (8'hba)) : (^forvar1845)) & $signed((~forvar1786)))))
            begin
              if ((forvar1885 ?
                  (^~{(reg1819 >= reg1876)}) : (~$signed((reg1804 ?
                      reg1826 : forvar1875)))))
                begin
                  if ({(~&((|reg1859) > reg1888[(3'h6):(1'h0)]))})
                    begin
                      reg1891 <= reg1773;
                      reg1892 <= (reg1856[(3'h5):(1'h0)] == $unsigned($signed(forvar1820[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg1891 <= (&(^((reg1870 > forvar1775) + (forvar1885 ~^ (8'hab)))));
                      reg1892 <= $unsigned((($unsigned(forvar1799) ?
                              reg1884[(2'h3):(1'h1)] : $signed(reg1857)) ?
                          ($signed(reg1843) + $unsigned(reg1787)) : $signed((reg1859 <= forvar1836))));
                      reg1893 <= (((8'ha5) ?
                              (((8'hb4) != forvar1798) << (reg1827 ~^ reg1884)) : $signed(reg1820)) ?
                          forvar1875[(1'h1):(1'h0)] : $unsigned(((reg1829 && reg1795) * forvar1758)));
                      reg1894 <= ((&$signed((reg1835 ?
                          reg1844 : (8'hb4)))) & $unsigned(reg1822[(3'h4):(2'h3)]));
                    end
                  reg1895 <= {$signed($signed(forvar1788))};
                end
              else
                begin
                  for (forvar1891 = (1'h0); (forvar1891 < (1'h0)); forvar1891 = (forvar1891 + (1'h1)))
                    begin
                      reg1892 <= reg1785[(2'h2):(2'h2)];
                    end
                end
            end
          else
            begin
              for (forvar1891 = (1'h0); (forvar1891 < (2'h3)); forvar1891 = (forvar1891 + (1'h1)))
                begin
                  if (($signed($signed($unsigned(forvar1797))) << reg1792))
                    begin
                      reg1892 <= (^~reg1829[(1'h1):(1'h1)]);
                      reg1893 <= reg1829;
                    end
                  else
                    begin
                      reg1892 <= forvar1775[(3'h4):(2'h2)];
                    end
                  for (forvar1894 = (1'h0); (forvar1894 < (1'h1)); forvar1894 = (forvar1894 + (1'h1)))
                    begin
                      reg1895 <= $unsigned(forvar1880[(3'h7):(3'h6)]);
                    end
                  for (forvar1896 = (1'h0); (forvar1896 < (1'h0)); forvar1896 = (forvar1896 + (1'h1)))
                    begin
                      reg1897 <= $signed($signed((reg1862 ?
                          $unsigned((8'ha8)) : (reg1847 || reg1780))));
                      reg1898 <= (+reg1820[(3'h5):(2'h3)]);
                      reg1899 <= {($unsigned(forvar1889) ?
                              (~reg1782[(1'h1):(1'h0)]) : $signed((!(8'ha2))))};
                      reg1900 <= forvar1823;
                    end
                end
            end
        end
      for (forvar1901 = (1'h0); (forvar1901 < (1'h1)); forvar1901 = (forvar1901 + (1'h1)))
        begin
          if (reg1890[(2'h2):(1'h0)])
            begin
              for (forvar1902 = (1'h0); (forvar1902 < (2'h2)); forvar1902 = (forvar1902 + (1'h1)))
                begin
                  reg1903 <= (8'ha6);
                end
              for (forvar1904 = (1'h0); (forvar1904 < (2'h3)); forvar1904 = (forvar1904 + (1'h1)))
                begin
                  for (forvar1905 = (1'h0); (forvar1905 < (1'h0)); forvar1905 = (forvar1905 + (1'h1)))
                    begin
                      reg1906 <= (((&reg1829) + reg1868[(1'h0):(1'h0)]) * (|$signed((-reg1871))));
                      reg1907 <= $unsigned((-{(reg1866 ? reg1844 : reg1850)}));
                      reg1908 <= $signed((!$signed((reg1766 - reg1877))));
                      reg1909 <= reg1877[(3'h4):(2'h3)];
                    end
                  if ({$unsigned((-{reg1825}))})
                    begin
                      reg1910 <= $signed($unsigned(reg1784));
                    end
                  else
                    begin
                      reg1910 <= reg1846;
                      reg1911 <= ((~&{reg1877}) && reg1824[(3'h5):(3'h5)]);
                    end
                end
              if (((+$unsigned((reg1831 ? reg1761 : (8'hb6)))) ^~ ((forvar1850 ?
                  $signed(forvar1880) : $unsigned(reg1832)) ^~ ($unsigned(reg1866) & reg1812[(4'h8):(3'h7)]))))
                begin
                  if ($signed(forvar1902[(2'h2):(1'h0)]))
                    begin
                      reg1912 <= ($signed({((8'ha2) ? reg1803 : reg1861)}) ?
                          (($signed(reg1791) ^ $signed(forvar1867)) ?
                              (!(reg1801 || reg1770)) : $unsigned($unsigned(reg1894))) : $signed(($unsigned(reg1853) ?
                              (~|reg1900) : forvar1799[(4'hc):(2'h3)])));
                      reg1913 <= wire1755;
                      reg1914 <= (reg1847[(1'h1):(1'h1)] ^ reg1764);
                      reg1915 <= ({$unsigned((~|reg1911))} ?
                          $unsigned(reg1843[(1'h1):(1'h0)]) : $unsigned(reg1864));
                    end
                  else
                    begin
                      reg1912 <= $unsigned($signed($unsigned(((8'hb9) ?
                          reg1803 : forvar1896))));
                      reg1913 <= $unsigned({(((8'hb3) ?
                              reg1835 : (8'hab)) ~^ $unsigned((8'h9c)))});
                      reg1914 <= ((($signed(forvar1823) ?
                                  $unsigned(reg1883) : $signed(reg1800)) ?
                              (8'ha8) : ($signed(reg1856) ?
                                  (reg1891 * forvar1863) : {reg1880})) ?
                          ($signed((~|reg1831)) ^ ({forvar1875} ?
                              (reg1892 ?
                                  reg1880 : reg1764) : $signed(reg1869))) : $signed(forvar1798[(2'h3):(1'h1)]));
                    end
                  if (reg1825)
                    begin
                      reg1916 <= $unsigned(reg1841);
                    end
                  else
                    begin
                      reg1916 <= $signed(reg1850[(4'hd):(3'h4)]);
                      reg1917 <= reg1852[(3'h7):(3'h7)];
                      reg1918 <= (~^(+reg1818[(2'h2):(1'h1)]));
                      reg1919 <= ((reg1807 <= $unsigned((!(8'had)))) || reg1774);
                    end
                  for (forvar1920 = (1'h0); (forvar1920 < (2'h2)); forvar1920 = (forvar1920 + (1'h1)))
                    begin
                      reg1921 <= forvar1856[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  if ((8'hb2))
                    begin
                      reg1912 <= ((~(8'hb5)) ?
                          ((reg1892 ?
                                  reg1886[(4'h8):(1'h0)] : $unsigned(reg1826)) ?
                              $signed((forvar1781 - reg1836)) : (forvar1865 ?
                                  $unsigned(forvar1757) : $unsigned(reg1886))) : ({$unsigned(forvar1809)} ?
                              forvar1879[(4'h8):(3'h7)] : reg1880[(2'h2):(1'h1)]));
                      reg1913 <= (reg1824 != $unsigned(((forvar1905 || reg1783) ?
                          (forvar1820 ? reg1822 : reg1777) : (^reg1819))));
                    end
                  else
                    begin
                      reg1912 <= ({(8'ha6)} ?
                          $signed(((reg1888 ? forvar1817 : reg1914) ?
                              reg1787[(3'h4):(2'h3)] : {reg1869})) : reg1886);
                      reg1913 <= ((&reg1765[(3'h4):(1'h1)]) & ($signed($signed(forvar1854)) ?
                          $signed((|reg1918)) : {((8'hb5) ?
                                  forvar1840 : reg1827)}));
                    end
                  for (forvar1914 = (1'h0); (forvar1914 < (2'h2)); forvar1914 = (forvar1914 + (1'h1)))
                    begin
                      reg1915 <= forvar1878;
                      reg1916 <= (8'had);
                      reg1917 <= ($unsigned($signed({forvar1790})) ?
                          $signed(reg1816[(1'h0):(1'h0)]) : ((((8'hb4) ?
                              forvar1800 : reg1793) ^~ forvar1828[(3'h7):(3'h4)]) + reg1892[(4'hc):(3'h6)]));
                    end
                end
            end
          else
            begin
              for (forvar1902 = (1'h0); (forvar1902 < (2'h3)); forvar1902 = (forvar1902 + (1'h1)))
                begin
                  if ({forvar1863[(2'h2):(1'h0)]})
                    begin
                      reg1903 <= $unsigned($unsigned($signed(reg1811[(3'h6):(2'h2)])));
                      reg1904 <= reg1765;
                    end
                  else
                    begin
                      reg1903 <= {{forvar1905}};
                      reg1904 <= {$signed($unsigned($unsigned(reg1777)))};
                      reg1905 <= (8'ha4);
                    end
                  reg1906 <= reg1913;
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1922 = (1'h0); (forvar1922 < (1'h0)); forvar1922 = (forvar1922 + (1'h1)))
        begin
          for (forvar1923 = (1'h0); (forvar1923 < (2'h3)); forvar1923 = (forvar1923 + (1'h1)))
            begin
              for (forvar1924 = (1'h0); (forvar1924 < (1'h0)); forvar1924 = (forvar1924 + (1'h1)))
                begin
                  for (forvar1925 = (1'h0); (forvar1925 < (2'h2)); forvar1925 = (forvar1925 + (1'h1)))
                    begin
                      reg1926 <= $unsigned((^reg1862));
                      reg1927 <= $unsigned(reg1798[(1'h1):(1'h0)]);
                      reg1928 <= (((!(reg1910 ?
                          reg1898 : reg1811)) >> ({reg1839} ?
                          $unsigned(reg1777) : (&reg1908))) >> (((^~forvar1775) ~^ (-reg1839)) >> ((^~reg1831) ?
                          (|reg1918) : (forvar1803 | reg1818))));
                      reg1929 <= (+$unsigned((8'hb1)));
                    end
                  if ({$unsigned(($unsigned(reg1824) ~^ {reg1770}))})
                    begin
                      reg1930 <= forvar1879;
                      reg1931 <= ({$unsigned($unsigned(forvar1856))} ?
                          {(~|reg1899[(3'h5):(3'h5)])} : (-forvar1896));
                    end
                  else
                    begin
                      reg1930 <= $unsigned($unsigned($unsigned((reg1897 ?
                          wire1756 : reg1816))));
                      reg1931 <= $unsigned(($unsigned($signed(reg1842)) * (~|(reg1800 ?
                          reg1800 : reg1778))));
                      reg1932 <= forvar1776[(1'h0):(1'h0)];
                    end
                  if ($signed($unsigned((^~(^~(8'hb5))))))
                    begin
                      reg1933 <= $unsigned((reg1887[(2'h2):(1'h1)] ?
                          ((^~(8'hab)) ?
                              reg1908 : (~(8'ha2))) : ({forvar1809} * forvar1817)));
                      reg1934 <= $signed(reg1774[(3'h4):(1'h1)]);
                      reg1935 <= $signed(reg1771);
                      reg1936 <= ($unsigned(reg1812) <= {({reg1805} - forvar1820[(2'h2):(1'h1)])});
                    end
                  else
                    begin
                      reg1933 <= (forvar1879 ?
                          reg1779[(2'h3):(2'h2)] : (8'hb0));
                    end
                  if ((((~^(reg1852 >>> forvar1758)) >> reg1914) ?
                      $signed($signed({reg1815})) : forvar1799[(4'hd):(4'h9)]))
                    begin
                      reg1937 <= (reg1830 <<< $unsigned(({forvar1924} || (|forvar1850))));
                    end
                  else
                    begin
                      reg1937 <= $signed(forvar1798[(1'h0):(1'h0)]);
                      reg1938 <= $signed((((reg1935 ? reg1853 : (8'hb7)) ?
                              (forvar1885 ?
                                  (8'haf) : reg1891) : $signed(reg1887)) ?
                          $signed(wire1754) : reg1850[(3'h7):(3'h7)]));
                    end
                end
            end
          if (forvar1865)
            begin
              reg1939 <= (forvar1865[(1'h0):(1'h0)] ?
                  reg1840 : $signed($unsigned(reg1780)));
            end
          else
            begin
              for (forvar1939 = (1'h0); (forvar1939 < (2'h3)); forvar1939 = (forvar1939 + (1'h1)))
                begin
                  for (forvar1940 = (1'h0); (forvar1940 < (2'h3)); forvar1940 = (forvar1940 + (1'h1)))
                    begin
                      reg1941 <= reg1779[(2'h2):(1'h0)];
                    end
                  for (forvar1942 = (1'h0); (forvar1942 < (2'h3)); forvar1942 = (forvar1942 + (1'h1)))
                    begin
                      reg1943 <= (($unsigned((reg1869 & reg1807)) ?
                          (!$signed((8'hb9))) : $signed($signed(reg1866))) > ($signed(forvar1905) ?
                          forvar1803[(4'hd):(4'h9)] : $unsigned($unsigned(reg1846))));
                      reg1944 <= {reg1846};
                    end
                end
              for (forvar1945 = (1'h0); (forvar1945 < (2'h3)); forvar1945 = (forvar1945 + (1'h1)))
                begin
                  for (forvar1946 = (1'h0); (forvar1946 < (2'h3)); forvar1946 = (forvar1946 + (1'h1)))
                    begin
                      reg1947 <= reg1847[(2'h3):(2'h3)];
                      reg1948 <= (-(reg1849 ?
                          forvar1880 : reg1792[(2'h3):(2'h2)]));
                      reg1949 <= $unsigned(reg1824[(3'h6):(3'h6)]);
                    end
                end
              for (forvar1950 = (1'h0); (forvar1950 < (2'h3)); forvar1950 = (forvar1950 + (1'h1)))
                begin
                  for (forvar1951 = (1'h0); (forvar1951 < (2'h3)); forvar1951 = (forvar1951 + (1'h1)))
                    begin
                      reg1952 <= reg1919;
                      reg1953 <= forvar1880;
                      reg1954 <= (~(~|reg1852));
                    end
                  for (forvar1955 = (1'h0); (forvar1955 < (2'h2)); forvar1955 = (forvar1955 + (1'h1)))
                    begin
                      reg1956 <= $signed($signed($unsigned($signed(reg1895))));
                      reg1957 <= reg1784[(4'h9):(1'h1)];
                    end
                  for (forvar1958 = (1'h0); (forvar1958 < (1'h0)); forvar1958 = (forvar1958 + (1'h1)))
                    begin
                      reg1959 <= $unsigned($unsigned(reg1918[(2'h3):(1'h0)]));
                      reg1960 <= ((forvar1901[(2'h3):(1'h0)] ?
                          {(forvar1797 >> (8'ha5))} : $unsigned(forvar1801[(2'h3):(2'h2)])) > (reg1816[(2'h2):(1'h0)] ?
                          (~&(^reg1887)) : ((^~reg1868) != reg1933)));
                    end
                  if (reg1900)
                    begin
                      reg1961 <= $unsigned($signed({(8'ha5)}));
                    end
                  else
                    begin
                      reg1961 <= $unsigned(((^~((8'haf) ? reg1913 : reg1915)) ?
                          $signed((^~(8'hb3))) : {(reg1804 >= forvar1946)}));
                      reg1962 <= $unsigned($unsigned($signed($signed(reg1778))));
                    end
                end
            end
          for (forvar1963 = (1'h0); (forvar1963 < (2'h2)); forvar1963 = (forvar1963 + (1'h1)))
            begin
              if ($signed($signed($unsigned($signed((8'ha7))))))
                begin
                  if (reg1843[(1'h0):(1'h0)])
                    begin
                      reg1964 <= ((-reg1813) ?
                          reg1937 : (+$unsigned((reg1853 ?
                              reg1877 : forvar1939))));
                      reg1965 <= reg1791;
                    end
                  else
                    begin
                      reg1964 <= $signed($unsigned(((~|forvar1821) & reg1904)));
                      reg1965 <= ($signed(reg1900) ?
                          (forvar1922[(1'h0):(1'h0)] + forvar1799[(4'h8):(1'h0)]) : reg1770);
                      reg1966 <= forvar1828;
                    end
                  if (forvar1828[(2'h3):(1'h0)])
                    begin
                      reg1967 <= reg1933[(2'h2):(1'h0)];
                      reg1968 <= reg1956[(1'h0):(1'h0)];
                      reg1969 <= (($unsigned($signed((8'ha2))) <<< reg1947[(3'h4):(3'h4)]) | forvar1760[(2'h3):(2'h2)]);
                      reg1970 <= $signed(reg1803[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg1967 <= reg1791[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar1964 = (1'h0); (forvar1964 < (1'h1)); forvar1964 = (forvar1964 + (1'h1)))
                    begin
                      reg1965 <= (|$signed((~|(forvar1963 && forvar1809))));
                      reg1966 <= forvar1942;
                      reg1967 <= $unsigned(reg1814);
                      reg1968 <= $unsigned($unsigned({(forvar1879 ?
                              reg1935 : reg1791)}));
                    end
                  if (((($signed(reg1793) ?
                          $signed(reg1897) : {reg1930}) >= ((~(8'ha4)) ?
                          reg1763[(1'h0):(1'h0)] : {reg1810})) ?
                      (-$unsigned($unsigned(reg1801))) : (~(~|$signed(reg1866)))))
                    begin
                      reg1969 <= $unsigned(reg1841);
                      reg1970 <= reg1773;
                      reg1971 <= ($unsigned($unsigned($unsigned(reg1831))) ?
                          (8'ha6) : reg1785);
                      reg1972 <= reg1856;
                    end
                  else
                    begin
                      reg1969 <= ((reg1931 ?
                          $signed(forvar1768[(3'h5):(2'h3)]) : $unsigned((forvar1922 - reg1807))) + (^~reg1780));
                      reg1970 <= (($unsigned(reg1918[(1'h1):(1'h0)]) ?
                              $unsigned((~^reg1836)) : (+(reg1936 >>> reg1853))) ?
                          $unsigned(reg1795) : (forvar1834[(2'h2):(1'h0)] << (~|{reg1778})));
                    end
                  reg1973 <= reg1800;
                  for (forvar1974 = (1'h0); (forvar1974 < (1'h1)); forvar1974 = (forvar1974 + (1'h1)))
                    begin
                      reg1975 <= ({$unsigned({forvar1786})} < {reg1915});
                      reg1976 <= ((~^($signed(reg1944) ~^ $unsigned(reg1973))) ?
                          reg1830 : (reg1851[(2'h3):(1'h1)] >>> $unsigned((!forvar1790))));
                    end
                end
              for (forvar1977 = (1'h0); (forvar1977 < (1'h0)); forvar1977 = (forvar1977 + (1'h1)))
                begin
                  if ($signed($unsigned(reg1928)))
                    begin
                      reg1978 <= reg1860[(2'h2):(1'h0)];
                      reg1979 <= ($unsigned((forvar1834[(2'h2):(1'h1)] ?
                          forvar1951[(1'h0):(1'h0)] : (forvar1820 != (8'hb8)))) || reg1838);
                      reg1980 <= ((&$signed({forvar1955})) * $unsigned($signed($signed(reg1812))));
                    end
                  else
                    begin
                      reg1978 <= {$unsigned(forvar1798)};
                      reg1979 <= $signed((((reg1772 << forvar1798) == (reg1943 * (8'hac))) ~^ ((forvar1844 >>> forvar1885) ?
                          (reg1907 ? reg1766 : reg1826) : (reg1972 ?
                              reg1804 : reg1818))));
                      reg1980 <= (reg1943 <<< forvar1759[(3'h5):(3'h4)]);
                      reg1981 <= ((8'hb1) ?
                          $unsigned($unsigned((reg1956 >>> forvar1963))) : ({(reg1838 ?
                                  reg1962 : reg1869)} == reg1978));
                    end
                  reg1982 <= forvar1799[(3'h4):(3'h4)];
                end
              for (forvar1983 = (1'h0); (forvar1983 < (1'h1)); forvar1983 = (forvar1983 + (1'h1)))
                begin
                  for (forvar1984 = (1'h0); (forvar1984 < (2'h2)); forvar1984 = (forvar1984 + (1'h1)))
                    begin
                      reg1985 <= (reg1772[(4'hc):(2'h2)] ?
                          ((forvar1865[(3'h4):(2'h2)] <<< {forvar1904}) - $unsigned((~|(8'ha4)))) : ((8'ha7) ?
                              (^~$signed(reg1787)) : $signed(reg1853[(4'hb):(1'h1)])));
                    end
                  for (forvar1986 = (1'h0); (forvar1986 < (2'h3)); forvar1986 = (forvar1986 + (1'h1)))
                    begin
                      reg1987 <= ($unsigned(($signed(reg1883) ?
                              (~^(8'ha1)) : $unsigned(reg1793))) ?
                          $signed(({wire1755} ?
                              (~&reg1764) : $unsigned(reg1800))) : {reg1962[(1'h1):(1'h1)]});
                    end
                  if ($signed((~^($unsigned(reg1835) ~^ (reg1793 ?
                      (8'ha8) : (8'h9f))))))
                    begin
                      reg1988 <= (reg1826[(4'h9):(4'h8)] << reg1917);
                    end
                  else
                    begin
                      reg1988 <= {(($unsigned(reg1918) << ((8'hb6) ?
                                  reg1778 : reg1934)) ?
                              (~|((8'ha2) ?
                                  reg1957 : reg1965)) : (~$unsigned(reg1985)))};
                      reg1989 <= $signed(reg1774[(3'h4):(2'h2)]);
                      reg1990 <= $signed(reg1895[(4'he):(3'h4)]);
                    end
                  if ($signed($signed((^(forvar1924 != (8'ha4))))))
                    begin
                      reg1991 <= $signed(reg1990);
                      reg1992 <= $unsigned((~&((reg1872 ?
                          reg1903 : forvar1757) <<< (forvar1977 ?
                          (8'ha2) : reg1860))));
                    end
                  else
                    begin
                      reg1991 <= (&$signed((&reg1978)));
                      reg1992 <= ((reg1988[(1'h0):(1'h0)] > (^~(!forvar1845))) ^ (8'hb3));
                    end
                end
              for (forvar1993 = (1'h0); (forvar1993 < (2'h3)); forvar1993 = (forvar1993 + (1'h1)))
                begin
                  for (forvar1994 = (1'h0); (forvar1994 < (2'h2)); forvar1994 = (forvar1994 + (1'h1)))
                    begin
                      reg1995 <= ($signed(reg1990) ?
                          (($unsigned((8'ha0)) >= (^~forvar1768)) ?
                              (~(reg1880 != (8'ha2))) : reg1802[(4'h8):(3'h6)]) : (~^forvar1950));
                      reg1996 <= forvar1964[(3'h5):(1'h1)];
                    end
                  for (forvar1997 = (1'h0); (forvar1997 < (2'h2)); forvar1997 = (forvar1997 + (1'h1)))
                    begin
                      reg1998 <= reg1929;
                    end
                  if ((&reg1787))
                    begin
                      reg1999 <= reg1825[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg1999 <= (8'had);
                      reg2000 <= (forvar1879 != $signed((reg1869[(3'h4):(2'h3)] ?
                          (reg1792 & reg1905) : $unsigned(reg1773))));
                      reg2001 <= ({reg1829} >>> reg1996[(4'ha):(3'h6)]);
                      reg2002 <= ((~^$signed({forvar1844})) ?
                          $unsigned(($signed(reg1764) ?
                              reg1839 : reg1961[(1'h0):(1'h0)])) : (reg1802 ?
                              {reg1985[(2'h3):(1'h1)]} : (reg1830 <<< ((8'ha5) ?
                                  reg1961 : forvar1951))));
                    end
                  if (reg1871[(4'hc):(4'h9)])
                    begin
                      reg2003 <= (forvar1891[(3'h6):(2'h2)] ?
                          reg1775[(2'h2):(2'h2)] : $unsigned(((-forvar1821) >>> reg1991)));
                      reg2004 <= reg1874;
                    end
                  else
                    begin
                      reg2003 <= ((((-reg1849) ?
                          $signed(reg1928) : (forvar1891 ?
                              reg1763 : forvar1977)) | (8'h9c)) > reg1793[(1'h0):(1'h0)]);
                      reg2004 <= $unsigned({$unsigned((forvar1902 ?
                              reg1961 : reg1971))});
                      reg2005 <= (&((reg1796 ?
                              (reg1847 ? reg1935 : reg1929) : (^~reg1852)) ?
                          $signed($unsigned(forvar1950)) : $unsigned((8'haa))));
                    end
                end
            end
          reg2006 <= wire1755[(2'h3):(2'h2)];
        end
    end
  assign wire2007 = reg1996[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg2008 <= ($unsigned($signed($unsigned(forvar1950))) ?
          ((reg1801[(3'h5):(1'h0)] ?
                  $signed(reg1919) : (reg1999 || forvar1955)) ?
              forvar1946[(2'h2):(2'h2)] : ((forvar1786 ?
                  reg1976 : forvar1854) >>> (~reg1962))) : forvar1776[(1'h1):(1'h1)]);
      if (reg1874)
        begin
          if (reg1975)
            begin
              if (reg2008[(1'h0):(1'h0)])
                begin
                  for (forvar2009 = (1'h0); (forvar2009 < (2'h2)); forvar2009 = (forvar2009 + (1'h1)))
                    begin
                      reg2010 <= $unsigned(reg1874[(2'h2):(1'h1)]);
                      reg2011 <= {$unsigned(($unsigned((8'hb7)) ?
                              {reg1992} : ((8'h9d) > reg1891)))};
                      reg2012 <= (&reg1956[(2'h3):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar2009 = (1'h0); (forvar2009 < (2'h2)); forvar2009 = (forvar2009 + (1'h1)))
                    begin
                      reg2010 <= reg1944;
                      reg2011 <= forvar1925;
                      reg2012 <= ($unsigned(reg1928[(4'hb):(2'h3)]) << reg1973);
                      reg2013 <= reg1908[(2'h3):(1'h1)];
                    end
                  for (forvar2014 = (1'h0); (forvar2014 < (2'h2)); forvar2014 = (forvar2014 + (1'h1)))
                    begin
                      reg2015 <= (&(reg1931 | ((reg2003 ?
                          (8'haa) : (8'hb7)) || $unsigned(reg1853))));
                      reg2016 <= (reg1969 < (!($unsigned(wire1754) * forvar1759[(3'h4):(2'h2)])));
                      reg2017 <= ((({(8'ha5)} >> reg1939) ?
                          reg1935 : $signed((&forvar1878))) <<< forvar1963);
                    end
                end
            end
          else
            begin
              for (forvar2009 = (1'h0); (forvar2009 < (1'h1)); forvar2009 = (forvar2009 + (1'h1)))
                begin
                  for (forvar2010 = (1'h0); (forvar2010 < (1'h1)); forvar2010 = (forvar2010 + (1'h1)))
                    begin
                      reg2011 <= ((~&{(reg1783 ^~ reg1992)}) ?
                          ((reg1835[(3'h4):(2'h3)] ?
                                  (forvar1920 << reg1835) : reg1829) ?
                              ($signed(forvar1878) ?
                                  reg1770 : $signed(reg1762)) : reg1980) : ($signed($unsigned(reg1981)) >= reg1784[(1'h0):(1'h0)]));
                      reg2012 <= $signed($signed($signed($unsigned(reg1968))));
                      reg2013 <= (&(8'hb7));
                    end
                  if (reg1887[(3'h6):(2'h3)])
                    begin
                      reg2014 <= $signed((^~reg1985[(2'h3):(1'h1)]));
                    end
                  else
                    begin
                      reg2014 <= (~($signed(reg1813[(2'h3):(2'h2)]) ~^ reg2011[(5'h10):(3'h6)]));
                      reg2015 <= ((|reg1793) || (-((^reg1908) < $unsigned(reg1850))));
                      reg2016 <= (^reg1987);
                      reg2017 <= ((~|(&forvar1776[(3'h7):(2'h2)])) <= (~|((reg1789 || forvar1773) >> (reg1915 ?
                          reg1776 : forvar1894))));
                    end
                end
              reg2018 <= ({forvar1901[(3'h4):(1'h0)]} <<< reg1909[(3'h6):(1'h0)]);
            end
        end
      else
        begin
          reg2009 <= reg1798;
          if (($signed($signed(forvar1801[(3'h5):(1'h0)])) ^ (8'ha6)))
            begin
              if (($signed(reg2014[(3'h7):(3'h4)]) ^ reg1912[(2'h2):(1'h1)]))
                begin
                  reg2010 <= (reg1938[(1'h1):(1'h1)] - (8'hba));
                end
              else
                begin
                  for (forvar2010 = (1'h0); (forvar2010 < (1'h0)); forvar2010 = (forvar2010 + (1'h1)))
                    begin
                      reg2011 <= reg1859;
                      reg2012 <= $unsigned(reg1906);
                      reg2013 <= reg1806[(2'h3):(1'h1)];
                      reg2014 <= (reg1818 ?
                          (-$signed($signed(forvar1836))) : reg1789);
                    end
                  for (forvar2015 = (1'h0); (forvar2015 < (2'h2)); forvar2015 = (forvar2015 + (1'h1)))
                    begin
                      reg2016 <= $signed(reg1847);
                    end
                  if ($unsigned($signed(({reg1771} >= ((8'h9e) ?
                      (8'ha5) : reg1827)))))
                    begin
                      reg2017 <= (reg1969[(1'h0):(1'h0)] - $unsigned({$signed((8'h9e))}));
                      reg2018 <= ($signed(reg1855) ?
                          $unsigned($unsigned(((8'ha7) >= (8'ha1)))) : ($signed($signed(reg1876)) ?
                              ((8'haa) && (~^(8'hac))) : (+$unsigned(forvar1923))));
                    end
                  else
                    begin
                      reg2017 <= ($signed(($signed((8'hb6)) << (~&reg1782))) != (^((reg2003 ?
                              reg1883 : reg1835) ?
                          reg1964 : (forvar1786 && reg1881))));
                      reg2018 <= reg1893[(2'h3):(1'h0)];
                      reg2019 <= $unsigned($unsigned({reg1976[(4'hb):(4'ha)]}));
                      reg2020 <= $unsigned((reg1967 | forvar1797));
                    end
                end
              if (reg1913[(1'h0):(1'h0)])
                begin
                  reg2021 <= (($unsigned(forvar1786[(3'h4):(1'h0)]) ~^ (!$signed((8'hb6)))) ?
                      (^~$unsigned((^reg1980))) : (reg1904 << $unsigned({reg2010})));
                  for (forvar2022 = (1'h0); (forvar2022 < (1'h0)); forvar2022 = (forvar2022 + (1'h1)))
                    begin
                      reg2023 <= (forvar1768 << {$unsigned((8'hb6))});
                    end
                  for (forvar2024 = (1'h0); (forvar2024 < (1'h1)); forvar2024 = (forvar2024 + (1'h1)))
                    begin
                      reg2025 <= reg1780;
                      reg2026 <= reg1775[(2'h3):(1'h1)];
                      reg2027 <= $signed((((forvar1867 && forvar1863) ?
                              forvar1801 : $unsigned(forvar1939)) ?
                          $signed(reg1972) : ($signed((8'hb8)) + forvar1939[(2'h3):(1'h1)])));
                      reg2028 <= {$unsigned(reg2011)};
                    end
                end
              else
                begin
                  for (forvar2021 = (1'h0); (forvar2021 < (1'h1)); forvar2021 = (forvar2021 + (1'h1)))
                    begin
                      reg2022 <= $signed((reg1825 ?
                          ((reg1823 ?
                              forvar1923 : forvar1781) >>> {reg1899}) : reg2004[(4'hb):(3'h6)]));
                      reg2023 <= {(8'haf)};
                      reg2024 <= reg1836;
                      reg2025 <= (^~{reg1841});
                    end
                  if ((reg1861 <= reg1810[(2'h2):(2'h2)]))
                    begin
                      reg2026 <= forvar1798;
                      reg2027 <= (+$unsigned(forvar1790[(4'h8):(2'h3)]));
                      reg2028 <= $signed(reg1824[(4'ha):(1'h1)]);
                    end
                  else
                    begin
                      reg2026 <= (8'hb1);
                    end
                  reg2029 <= (~&((^reg1856) > $signed($unsigned(reg1939))));
                  for (forvar2030 = (1'h0); (forvar2030 < (1'h1)); forvar2030 = (forvar2030 + (1'h1)))
                    begin
                      reg2031 <= $signed((forvar1798[(3'h6):(1'h0)] << {reg1935[(2'h3):(2'h2)]}));
                    end
                end
              reg2032 <= (forvar1854 > reg1944[(2'h2):(1'h1)]);
            end
          else
            begin
              if (($signed(reg1932[(5'h10):(2'h3)]) ?
                  ((~((8'hb4) | (8'hb2))) ?
                      reg1825[(3'h7):(3'h6)] : ((reg1846 ?
                          reg1990 : (8'hb2)) - $signed(forvar2021))) : ($signed((reg1782 <= reg1844)) + $unsigned({(8'ha7)}))))
                begin
                  for (forvar2010 = (1'h0); (forvar2010 < (2'h2)); forvar2010 = (forvar2010 + (1'h1)))
                    begin
                      reg2011 <= forvar1867[(3'h6):(3'h6)];
                      reg2012 <= $signed((reg1870 ^ ($unsigned(reg1916) ?
                          (reg1862 ?
                              reg1941 : (8'h9d)) : reg1891[(2'h2):(1'h0)])));
                      reg2013 <= ($unsigned(reg1948[(4'ha):(3'h6)]) ?
                          $unsigned(($unsigned(reg1990) ?
                              (^reg1887) : reg1954)) : {($signed(forvar1974) > (forvar1845 <<< reg1812))});
                      reg2014 <= reg1779;
                    end
                  reg2015 <= (~^(^~$signed((reg1777 != reg1916))));
                  reg2016 <= reg1988;
                end
              else
                begin
                  for (forvar2010 = (1'h0); (forvar2010 < (1'h1)); forvar2010 = (forvar2010 + (1'h1)))
                    begin
                      reg2011 <= ($unsigned($unsigned((~^reg1814))) & reg1835);
                      reg2012 <= $signed($signed(({(8'ha1)} ?
                          (reg1936 ?
                              forvar1828 : forvar1946) : $unsigned((8'ha6)))));
                      reg2013 <= reg1839;
                      reg2014 <= ($unsigned(($unsigned(reg1897) ?
                          ((8'hb9) & reg1917) : reg2024[(2'h2):(1'h1)])) ~^ (8'h9e));
                    end
                end
              for (forvar2017 = (1'h0); (forvar2017 < (2'h3)); forvar2017 = (forvar2017 + (1'h1)))
                begin
                  reg2018 <= $unsigned({reg2011[(3'h6):(1'h0)]});
                  if (((((reg1782 + reg1927) == {reg1903}) ^~ $unsigned(forvar1854[(2'h2):(2'h2)])) << ((~reg2031) - $unsigned((reg2024 ?
                      forvar1845 : forvar1773)))))
                    begin
                      reg2019 <= $signed(reg1800);
                      reg2020 <= $signed((|$signed($signed((8'hba)))));
                    end
                  else
                    begin
                      reg2019 <= (({$unsigned(reg1839)} ?
                              $signed((+reg1787)) : reg1908[(2'h3):(1'h0)]) ?
                          reg2002[(4'h9):(2'h2)] : $unsigned($signed($unsigned(reg2000))));
                      reg2020 <= (8'hae);
                      reg2021 <= forvar1914;
                    end
                  reg2022 <= {$signed(((~^reg1985) ~^ $unsigned(reg1890)))};
                end
              for (forvar2023 = (1'h0); (forvar2023 < (2'h2)); forvar2023 = (forvar2023 + (1'h1)))
                begin
                  for (forvar2024 = (1'h0); (forvar2024 < (2'h3)); forvar2024 = (forvar2024 + (1'h1)))
                    begin
                      reg2025 <= (reg1771[(4'he):(4'hb)] != reg1971[(1'h0):(1'h0)]);
                      reg2026 <= (((|((8'haf) ?
                              reg1953 : (8'hb0))) ~^ {$signed(forvar1993)}) ?
                          $signed((^~$signed(reg1967))) : reg1860[(3'h4):(2'h2)]);
                      reg2027 <= reg2020;
                    end
                  for (forvar2028 = (1'h0); (forvar2028 < (1'h0)); forvar2028 = (forvar2028 + (1'h1)))
                    begin
                      reg2029 <= (reg1876 * reg1839);
                      reg2030 <= forvar1875;
                      reg2031 <= {$signed($signed((reg1962 ?
                              reg1774 : forvar1955)))};
                    end
                  if (forvar1940[(2'h3):(2'h3)])
                    begin
                      reg2032 <= reg1842[(1'h0):(1'h0)];
                      reg2033 <= ((8'h9c) + reg2019[(4'hf):(4'hd)]);
                      reg2034 <= reg1970[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg2032 <= $unsigned($unsigned($unsigned((forvar2030 - reg1815))));
                      reg2033 <= $unsigned($unsigned(forvar1801[(1'h0):(1'h0)]));
                    end
                end
              for (forvar2035 = (1'h0); (forvar2035 < (1'h0)); forvar2035 = (forvar2035 + (1'h1)))
                begin
                  for (forvar2036 = (1'h0); (forvar2036 < (1'h0)); forvar2036 = (forvar2036 + (1'h1)))
                    begin
                      reg2037 <= $signed(({(^~reg1767)} ?
                          (~^$signed(reg1998)) : reg1991[(1'h0):(1'h0)]));
                      reg2038 <= (reg1957 ?
                          (8'hba) : (({reg1810} ? reg1880 : reg1960) ?
                              ((8'hba) ~^ reg1938) : ((^~(8'ha6)) ?
                                  $signed(reg1894) : (+wire2007))));
                      reg2039 <= (8'hac);
                    end
                  if (($signed(reg1883) ?
                      (reg1956[(1'h0):(1'h0)] * reg1766) : ((reg1765[(4'h9):(1'h0)] << $signed((8'hb5))) <<< {$unsigned((8'hba))})))
                    begin
                      reg2040 <= $unsigned((((8'hb3) && (reg1832 ?
                          reg2014 : forvar1986)) <= $signed($signed(reg1825))));
                      reg2041 <= ($unsigned((~^$signed(reg1992))) ?
                          $unsigned(forvar1797) : $unsigned((&(8'hb6))));
                      reg2042 <= $unsigned($signed(reg1952));
                      reg2043 <= (reg1782[(1'h1):(1'h1)] ?
                          $unsigned((^~$signed(reg1811))) : ((8'hb1) ^ ({reg2004} ?
                              (forvar1942 ?
                                  reg1771 : forvar1786) : $signed(forvar1800))));
                    end
                  else
                    begin
                      reg2040 <= ((reg2031 ?
                          reg1935[(1'h0):(1'h0)] : (8'ha1)) > (+$unsigned(reg1856[(4'h8):(4'h8)])));
                      reg2041 <= (^(reg1998[(3'h7):(3'h4)] > $unsigned(reg1873)));
                    end
                end
            end
          for (forvar2044 = (1'h0); (forvar2044 < (1'h1)); forvar2044 = (forvar2044 + (1'h1)))
            begin
              reg2045 <= (|reg1873[(3'h5):(3'h5)]);
              reg2046 <= {forvar1984[(3'h5):(1'h1)]};
              if ((8'h9f))
                begin
                  for (forvar2047 = (1'h0); (forvar2047 < (1'h0)); forvar2047 = (forvar2047 + (1'h1)))
                    begin
                      reg2048 <= (~^forvar1878[(3'h4):(1'h0)]);
                    end
                end
              else
                begin
                  if (((&(reg1980 - $unsigned(reg2041))) ?
                      (~&$signed((reg1956 ?
                          reg1975 : reg1763))) : {(reg1890[(3'h4):(2'h3)] >>> (reg1883 > (8'hb2)))}))
                    begin
                      reg2047 <= ($unsigned(wire2007) <= $unsigned($signed({reg1776})));
                      reg2048 <= {{reg1910}};
                      reg2049 <= $signed(((&(^forvar1834)) ?
                          reg1927[(4'ha):(3'h7)] : forvar1951));
                    end
                  else
                    begin
                      reg2047 <= $unsigned((^($signed(reg1762) ?
                          $unsigned(reg1830) : reg2033[(3'h5):(1'h1)])));
                      reg2048 <= reg1970[(1'h1):(1'h0)];
                      reg2049 <= $signed(({(reg1964 ? (8'hab) : reg1947)} ?
                          (((8'ha0) ? reg1899 : reg2004) ?
                              reg1947 : $signed(forvar1894)) : $unsigned((reg1949 ~^ reg1972))));
                      reg2050 <= (($signed($signed(reg1949)) >>> $unsigned((+forvar1940))) * reg1857);
                    end
                  for (forvar2051 = (1'h0); (forvar2051 < (2'h3)); forvar2051 = (forvar2051 + (1'h1)))
                    begin
                      reg2052 <= ((reg2014 + $signed((+forvar1994))) & ($unsigned(reg1804) ?
                          ((forvar1891 ? forvar1942 : (8'hb7)) ?
                              $unsigned(forvar2022) : $signed(reg1820)) : $signed((^reg1949))));
                      reg2053 <= $unsigned(($unsigned(reg1928[(2'h3):(2'h2)]) ?
                          ((8'ha4) ?
                              reg1936[(1'h0):(1'h0)] : (^~(8'ha5))) : (~(reg1777 >= reg1975))));
                    end
                end
            end
          if ({$signed(reg2042[(1'h1):(1'h1)])})
            begin
              for (forvar2054 = (1'h0); (forvar2054 < (2'h2)); forvar2054 = (forvar2054 + (1'h1)))
                begin
                  for (forvar2055 = (1'h0); (forvar2055 < (2'h2)); forvar2055 = (forvar2055 + (1'h1)))
                    begin
                      reg2056 <= (((reg1792 ? {reg1969} : $signed(reg1823)) ?
                          $signed((forvar2023 > reg1980)) : (forvar1821[(1'h1):(1'h1)] >= (reg1938 ?
                              (8'hac) : forvar2035))) | {reg2010});
                      reg2057 <= reg1979;
                    end
                  for (forvar2058 = (1'h0); (forvar2058 < (1'h0)); forvar2058 = (forvar2058 + (1'h1)))
                    begin
                      reg2059 <= reg1931;
                      reg2060 <= (^$unsigned(reg1890));
                      reg2061 <= reg1991[(4'ha):(1'h0)];
                      reg2062 <= (reg1934 && (~|$unsigned((reg1910 >> forvar1905))));
                    end
                  for (forvar2063 = (1'h0); (forvar2063 < (2'h2)); forvar2063 = (forvar2063 + (1'h1)))
                    begin
                      reg2064 <= $unsigned($signed($unsigned(reg1815[(2'h2):(1'h0)])));
                      reg2065 <= reg1825[(3'h7):(3'h4)];
                    end
                  for (forvar2066 = (1'h0); (forvar2066 < (1'h0)); forvar2066 = (forvar2066 + (1'h1)))
                    begin
                      reg2067 <= reg1847[(2'h3):(2'h2)];
                    end
                end
              for (forvar2068 = (1'h0); (forvar2068 < (1'h0)); forvar2068 = (forvar2068 + (1'h1)))
                begin
                  if ((((reg1789[(3'h6):(1'h1)] >> {(8'hac)}) | reg1816[(4'h8):(2'h3)]) ?
                      (($unsigned(reg1859) ~^ wire1754[(2'h2):(1'h1)]) && (&$signed((8'had)))) : reg1770[(3'h7):(3'h4)]))
                    begin
                      reg2069 <= $unsigned($signed($unsigned((-reg1822))));
                    end
                  else
                    begin
                      reg2069 <= forvar1786[(3'h7):(2'h3)];
                      reg2070 <= $unsigned($signed({((8'hb3) * (8'hb0))}));
                      reg2071 <= ((((8'ha0) - {reg1992}) ?
                              $signed($unsigned(forvar1863)) : (~^reg1970)) ?
                          $unsigned(forvar1800[(4'h8):(3'h7)]) : (forvar1836 >= reg1810[(4'hb):(3'h5)]));
                      reg2072 <= (~|$unsigned($signed((reg2020 ?
                          reg1803 : reg1884))));
                    end
                  reg2073 <= {(reg2000 ?
                          $signed((forvar2035 ? reg2027 : reg1973)) : reg1832)};
                  reg2074 <= reg1763;
                end
              if ((~|$unsigned(($signed(reg1943) ?
                  (reg1778 == forvar1914) : (forvar2009 ? reg1959 : reg1820)))))
                begin
                  for (forvar2075 = (1'h0); (forvar2075 < (1'h0)); forvar2075 = (forvar2075 + (1'h1)))
                    begin
                      reg2076 <= $signed(($unsigned($signed(reg2002)) ?
                          $signed(reg1949[(2'h3):(2'h3)]) : $unsigned((reg1941 ?
                              forvar1904 : (8'hac)))));
                    end
                  reg2077 <= reg1943[(3'h6):(2'h2)];
                  for (forvar2078 = (1'h0); (forvar2078 < (2'h2)); forvar2078 = (forvar2078 + (1'h1)))
                    begin
                      reg2079 <= $signed((~^$signed((!reg1943))));
                      reg2080 <= $unsigned((^$signed((reg1882 < reg1891))));
                    end
                end
              else
                begin
                  if (((((forvar1920 ?
                      reg2080 : reg1906) * (-reg1802)) == $unsigned({forvar2021})) << reg2077))
                    begin
                      reg2075 <= (~^reg1787);
                      reg2076 <= (($unsigned($signed((8'ha5))) ?
                              $signed(forvar1776[(3'h7):(1'h1)]) : (8'h9d)) ?
                          ((~|(8'ha2)) ^ (8'haf)) : reg2017);
                    end
                  else
                    begin
                      reg2075 <= reg1789;
                      reg2076 <= ($unsigned({(reg2070 <= forvar1867)}) ?
                          {(~(!reg2015))} : ($signed((reg2076 ?
                              (8'ha8) : reg1823)) < (~|(forvar2009 ?
                              reg1890 : forvar1939))));
                    end
                  for (forvar2077 = (1'h0); (forvar2077 < (1'h1)); forvar2077 = (forvar2077 + (1'h1)))
                    begin
                      reg2078 <= (~|$unsigned(reg1845));
                      reg2079 <= (forvar1993 ?
                          (8'haa) : $unsigned((|(~|(8'ha2)))));
                      reg2080 <= $unsigned({(~^(forvar1865 ^~ (8'ha3)))});
                    end
                  for (forvar2081 = (1'h0); (forvar2081 < (2'h2)); forvar2081 = (forvar2081 + (1'h1)))
                    begin
                      reg2082 <= (((((8'hb5) ?
                          (8'h9f) : reg2079) < reg2003[(2'h2):(1'h0)]) <= $signed(reg1882[(2'h2):(1'h1)])) >>> $signed($signed(forvar1817)));
                      reg2083 <= (forvar1759 ?
                          reg2041 : $signed(((reg2014 >> reg1892) ?
                              $unsigned((8'hb3)) : reg1789)));
                      reg2084 <= $signed(forvar2017);
                    end
                end
              reg2085 <= (^(!(-(reg1985 == (8'hb3)))));
            end
          else
            begin
              if ($unsigned(reg1775[(1'h1):(1'h1)]))
                begin
                  for (forvar2054 = (1'h0); (forvar2054 < (2'h2)); forvar2054 = (forvar2054 + (1'h1)))
                    begin
                      reg2055 <= ((|forvar1840) ?
                          (8'hb9) : (~{forvar2081[(4'h8):(4'h8)]}));
                    end
                  for (forvar2056 = (1'h0); (forvar2056 < (1'h0)); forvar2056 = (forvar2056 + (1'h1)))
                    begin
                      reg2057 <= reg1826;
                      reg2058 <= $signed((-{reg1933}));
                    end
                end
              else
                begin
                  for (forvar2054 = (1'h0); (forvar2054 < (1'h0)); forvar2054 = (forvar2054 + (1'h1)))
                    begin
                      reg2055 <= ((&(~|(forvar1775 ?
                          reg2073 : forvar1854))) ^~ reg1792[(2'h3):(2'h2)]);
                    end
                  if (((~&($signed(reg1829) ?
                      reg1962 : (8'haf))) != $signed(forvar1946)))
                    begin
                      reg2056 <= ($signed(($signed(forvar1823) <<< (reg1840 > reg1990))) ?
                          $unsigned(reg2010[(3'h7):(3'h7)]) : $unsigned((~^reg1794[(3'h6):(2'h2)])));
                      reg2057 <= ((forvar1776 ?
                          ($unsigned((8'h9f)) <= {forvar1768}) : $unsigned(reg1982[(2'h2):(1'h0)])) ~^ ($unsigned(forvar2021[(4'h9):(4'h8)]) ?
                          reg1837[(1'h1):(1'h1)] : (^(!reg1908))));
                    end
                  else
                    begin
                      reg2056 <= ((forvar1984[(4'h8):(3'h7)] <= $signed((^~reg1832))) >= (~^$unsigned($signed(reg1859))));
                    end
                  for (forvar2058 = (1'h0); (forvar2058 < (1'h0)); forvar2058 = (forvar2058 + (1'h1)))
                    begin
                      reg2059 <= $unsigned({($unsigned(reg1982) == (reg1884 ?
                              reg2040 : reg1935))});
                      reg2060 <= (reg2000[(1'h1):(1'h1)] ?
                          (~^((reg1988 >= reg2065) ^~ (~|reg2014))) : $unsigned(reg1872));
                      reg2061 <= (reg1793[(2'h2):(2'h2)] < ((^(reg1787 ?
                              forvar1889 : forvar2051)) ?
                          ((~|reg2055) ~^ $signed(wire2007)) : $unsigned($signed((8'ha2)))));
                      reg2062 <= forvar2047;
                    end
                  for (forvar2063 = (1'h0); (forvar2063 < (1'h1)); forvar2063 = (forvar2063 + (1'h1)))
                    begin
                      reg2064 <= reg2027;
                      reg2065 <= $unsigned(reg1824);
                      reg2066 <= ($unsigned($signed((reg1988 ?
                          reg2073 : reg1916))) ^ (reg1934[(3'h4):(1'h1)] ^ forvar1867));
                    end
                end
            end
        end
      if ($signed({(reg2027 | (reg2040 ? reg1959 : reg2024))}))
        begin
          for (forvar2086 = (1'h0); (forvar2086 < (2'h2)); forvar2086 = (forvar2086 + (1'h1)))
            begin
              for (forvar2087 = (1'h0); (forvar2087 < (1'h0)); forvar2087 = (forvar2087 + (1'h1)))
                begin
                  for (forvar2088 = (1'h0); (forvar2088 < (2'h3)); forvar2088 = (forvar2088 + (1'h1)))
                    begin
                      reg2089 <= reg1880[(2'h3):(1'h1)];
                      reg2090 <= {{reg1877[(1'h0):(1'h0)]}};
                    end
                  reg2091 <= {$signed((reg1886[(4'ha):(1'h1)] ?
                          forvar1801[(2'h3):(2'h3)] : (reg2001 ?
                              reg1769 : forvar1905)))};
                  reg2092 <= reg2034;
                end
              if (($unsigned($unsigned(reg1934[(1'h0):(1'h0)])) ?
                  $unsigned(((reg1780 ? reg1841 : reg1893) ?
                      {forvar1828} : ((8'ha6) ?
                          reg1909 : forvar2086))) : reg1933[(1'h1):(1'h1)]))
                begin
                  for (forvar2093 = (1'h0); (forvar2093 < (2'h3)); forvar2093 = (forvar2093 + (1'h1)))
                    begin
                      reg2094 <= ($unsigned((~$signed(reg1826))) ?
                          $signed(forvar2066) : {(~|$unsigned(forvar2066))});
                    end
                  reg2095 <= (!$signed($signed((reg1776 ^ forvar2077))));
                end
              else
                begin
                  reg2093 <= (^((forvar1986 | forvar1914) ?
                      $signed($signed(reg2082)) : reg1792[(2'h2):(2'h2)]));
                end
              if (forvar1775[(2'h3):(2'h3)])
                begin
                  reg2096 <= ((+$signed((reg1876 ? reg1771 : (8'hba)))) ?
                      (((forvar1997 != reg1832) ?
                              {forvar1850} : $unsigned(forvar1840)) ?
                          $signed($signed(forvar2093)) : ((forvar1986 ~^ reg1765) ~^ reg2024)) : forvar1836[(1'h1):(1'h0)]);
                  if (reg1778)
                    begin
                      reg2097 <= (8'ha2);
                      reg2098 <= reg1929[(1'h1):(1'h0)];
                      reg2099 <= ((~|(8'hba)) ^ (~^forvar2081));
                      reg2100 <= {$signed($signed({reg2024}))};
                    end
                  else
                    begin
                      reg2097 <= $signed({$signed(reg1773)});
                      reg2098 <= (reg1894 + reg2074[(1'h1):(1'h1)]);
                      reg2099 <= {{reg2050}};
                      reg2100 <= (({$unsigned(forvar2017)} & $unsigned({reg1819})) - reg1995[(3'h4):(2'h2)]);
                    end
                  if ($unsigned($unsigned(($signed(reg1835) != reg2024))))
                    begin
                      reg2101 <= $signed($signed(forvar1885[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg2101 <= ({reg1988[(1'h0):(1'h0)]} > reg2089[(3'h4):(2'h3)]);
                    end
                  for (forvar2102 = (1'h0); (forvar2102 < (1'h0)); forvar2102 = (forvar2102 + (1'h1)))
                    begin
                      reg2103 <= (~$unsigned($signed((reg2066 || forvar2068))));
                    end
                end
              else
                begin
                  for (forvar2096 = (1'h0); (forvar2096 < (2'h3)); forvar2096 = (forvar2096 + (1'h1)))
                    begin
                      reg2097 <= ({(+(reg1965 <= forvar2047))} - (8'hb6));
                      reg2098 <= reg2089[(4'h8):(2'h2)];
                    end
                  reg2099 <= (!$unsigned(((reg1793 || reg2064) ?
                      (~|(8'hb9)) : (forvar2022 ? reg1991 : forvar1817))));
                  if (forvar2075[(2'h2):(1'h0)])
                    begin
                      reg2100 <= forvar1945[(4'he):(4'hc)];
                      reg2101 <= reg1765[(1'h1):(1'h0)];
                      reg2102 <= $unsigned(($signed(((8'ha4) > reg2084)) <= $signed((reg1767 + reg2042))));
                      reg2103 <= forvar1891[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg2100 <= ((+{$unsigned(reg1778)}) ?
                          reg2079[(3'h5):(1'h0)] : $unsigned(forvar1809[(3'h5):(3'h4)]));
                    end
                  if ((((~^(forvar1844 && reg1783)) ?
                      (-((8'hb7) && (8'haf))) : $unsigned(((8'h9c) - forvar1823))) >> {(reg1916[(1'h1):(1'h0)] >>> $unsigned(reg1938))}))
                    begin
                      reg2104 <= reg1911;
                      reg2105 <= (reg2072[(4'ha):(4'ha)] != {(((8'hb2) ?
                              (8'hb4) : reg1787) <= $signed((8'hb5)))});
                      reg2106 <= ((($signed(reg2002) ?
                          forvar2088 : {(8'haf)}) & (~&{reg2012})) < reg2050);
                    end
                  else
                    begin
                      reg2104 <= ((((&reg1999) ?
                              ((8'hb5) >>> reg1775) : $signed(reg2043)) ?
                          ($unsigned(reg2106) ?
                              (wire2007 - forvar1775) : (reg2010 ^~ reg1884)) : $unsigned((~(8'hb9)))) ^~ reg2021[(4'h9):(1'h1)]);
                      reg2105 <= ((&(8'ha3)) >= $signed(reg1947[(4'ha):(4'h9)]));
                      reg2106 <= $signed(reg2089);
                      reg2107 <= reg1798;
                    end
                end
            end
          reg2108 <= (forvar2024[(1'h1):(1'h0)] <= reg1835[(3'h4):(1'h1)]);
        end
      else
        begin
          for (forvar2086 = (1'h0); (forvar2086 < (2'h3)); forvar2086 = (forvar2086 + (1'h1)))
            begin
              reg2087 <= (+reg1837);
              for (forvar2088 = (1'h0); (forvar2088 < (2'h2)); forvar2088 = (forvar2088 + (1'h1)))
                begin
                  reg2089 <= (($signed($signed(forvar2063)) == ($unsigned(forvar1799) ?
                      (reg1821 ?
                          reg1765 : wire1754) : ((8'hb5) ~^ reg1914))) == $unsigned($unsigned((~&forvar1828))));
                  if ({(({reg2012} + reg1919) ?
                          {$unsigned(forvar1781)} : (forvar1950 ?
                              (!reg1845) : (!(8'ha1))))})
                    begin
                      reg2090 <= reg1990[(3'h5):(2'h2)];
                      reg2091 <= (($signed((reg2028 >= (8'hba))) * $signed(reg1851[(1'h0):(1'h0)])) ?
                          reg1772[(4'hc):(2'h2)] : reg2072[(4'h8):(2'h3)]);
                      reg2092 <= $signed((+$signed((reg1848 && reg1991))));
                    end
                  else
                    begin
                      reg2090 <= $signed(($signed(reg1796) ?
                          ((|reg2020) >> forvar1920[(4'ha):(3'h6)]) : reg2061[(3'h4):(2'h3)]));
                      reg2091 <= reg1830;
                      reg2092 <= $unsigned($unsigned($unsigned((forvar2066 ?
                          reg1787 : (8'ha3)))));
                      reg2093 <= ((8'hae) <<< ((+((8'h9c) ?
                              reg2004 : forvar1923)) ?
                          reg1791 : $unsigned((!reg2061))));
                    end
                  if ($unsigned($signed(((forvar1945 ? reg2080 : reg2108) ?
                      (^~forvar2075) : reg1930))))
                    begin
                      reg2094 <= forvar1924[(2'h3):(1'h1)];
                      reg2095 <= ($signed((^(reg2078 ? (8'ha4) : reg1930))) ?
                          (!{reg2025[(2'h3):(1'h0)]}) : reg2047);
                      reg2096 <= {$unsigned((~$signed(reg1833)))};
                      reg2097 <= (~reg1813);
                    end
                  else
                    begin
                      reg2094 <= {reg2014[(2'h2):(1'h1)]};
                    end
                end
              reg2098 <= $signed(reg1964[(3'h4):(1'h1)]);
            end
          reg2099 <= {(reg1926 ?
                  (reg2096[(4'ha):(2'h3)] ?
                      reg1934 : (reg1917 ?
                          reg1947 : reg2084)) : (reg1767 | (8'haa)))};
        end
      if (reg1776[(1'h1):(1'h0)])
        begin
          for (forvar2109 = (1'h0); (forvar2109 < (2'h3)); forvar2109 = (forvar2109 + (1'h1)))
            begin
              for (forvar2110 = (1'h0); (forvar2110 < (1'h1)); forvar2110 = (forvar2110 + (1'h1)))
                begin
                  if ($signed({(~|{reg1992})}))
                    begin
                      reg2111 <= (reg1943[(2'h3):(1'h0)] >>> ($unsigned($unsigned(reg2101)) <<< $signed($signed((8'hb3)))));
                      reg2112 <= (forvar1836[(2'h2):(1'h0)] + $signed(reg1916));
                    end
                  else
                    begin
                      reg2111 <= ((reg1807[(3'h5):(3'h5)] || reg1767[(2'h2):(1'h1)]) < (!$unsigned((&forvar1786))));
                    end
                  for (forvar2113 = (1'h0); (forvar2113 < (1'h0)); forvar2113 = (forvar2113 + (1'h1)))
                    begin
                      reg2114 <= reg1821[(3'h4):(2'h2)];
                      reg2115 <= (8'hb3);
                      reg2116 <= ((reg2040 && $signed(reg1953)) ?
                          forvar1854 : reg1861[(2'h3):(2'h3)]);
                    end
                  if (forvar2066[(2'h3):(1'h0)])
                    begin
                      reg2117 <= ((~^wire1756[(3'h5):(2'h3)]) < reg1927);
                      reg2118 <= ({$signed($unsigned((8'h9e)))} | (~|$unsigned((8'ha2))));
                      reg2119 <= (|$unsigned(reg2034[(1'h1):(1'h0)]));
                      reg2120 <= $unsigned($unsigned((!reg1886[(2'h3):(1'h1)])));
                    end
                  else
                    begin
                      reg2117 <= (forvar2068 ?
                          ({reg1855[(1'h1):(1'h0)]} <<< (^~{reg2064})) : ({(reg2033 ?
                                      forvar1798 : reg1840)} ?
                              $signed((reg2042 <= reg2062)) : (-reg1853)));
                      reg2118 <= (-reg1917[(4'h9):(3'h5)]);
                      reg2119 <= (reg1903[(2'h2):(1'h0)] < {reg2111[(1'h0):(1'h0)]});
                    end
                end
            end
          for (forvar2121 = (1'h0); (forvar2121 < (1'h0)); forvar2121 = (forvar2121 + (1'h1)))
            begin
              reg2122 <= $unsigned(reg1964);
              for (forvar2123 = (1'h0); (forvar2123 < (1'h1)); forvar2123 = (forvar2123 + (1'h1)))
                begin
                  for (forvar2124 = (1'h0); (forvar2124 < (2'h3)); forvar2124 = (forvar2124 + (1'h1)))
                    begin
                      reg2125 <= {(&(^(^~(8'hba))))};
                      reg2126 <= {reg2016};
                    end
                  for (forvar2127 = (1'h0); (forvar2127 < (2'h2)); forvar2127 = (forvar2127 + (1'h1)))
                    begin
                      reg2128 <= reg2030[(3'h6):(1'h1)];
                    end
                  if ((reg2065 >>> $signed(reg1991)))
                    begin
                      reg2129 <= reg1972;
                      reg2130 <= reg1826;
                    end
                  else
                    begin
                      reg2129 <= {$unsigned($signed((~^forvar1809)))};
                      reg2130 <= (reg1971[(2'h3):(1'h1)] ?
                          ($unsigned((8'hab)) ?
                              ($unsigned(forvar1768) ?
                                  reg2026 : $signed((8'ha9))) : $signed((reg1776 ?
                                  reg1805 : forvar1891))) : ($unsigned(reg1805) ?
                              reg1793[(3'h6):(1'h1)] : $unsigned($unsigned(forvar2077))));
                    end
                  for (forvar2131 = (1'h0); (forvar2131 < (2'h2)); forvar2131 = (forvar2131 + (1'h1)))
                    begin
                      reg2132 <= (reg1913 << $unsigned($signed((reg1846 ?
                          reg1833 : (8'ha2)))));
                      reg2133 <= reg2106[(2'h2):(1'h0)];
                      reg2134 <= $signed($signed($unsigned($signed((8'hb4)))));
                    end
                end
              if ($signed((-(~|{reg2031}))))
                begin
                  if ($unsigned(({(forvar1867 <<< (8'hb4))} <= ({reg2125} ^~ (reg2087 * reg2120)))))
                    begin
                      reg2135 <= ((&({forvar1858} == (8'ha6))) ?
                          reg1824 : reg1859[(1'h1):(1'h0)]);
                      reg2136 <= $unsigned(reg2064);
                      reg2137 <= forvar2030;
                      reg2138 <= (((|forvar2102[(3'h5):(2'h2)]) || ({reg1975} * $unsigned(reg1836))) ?
                          reg1898 : {reg1912});
                    end
                  else
                    begin
                      reg2135 <= forvar2036;
                      reg2136 <= (!reg2018);
                      reg2137 <= $signed((^~$unsigned((reg1991 ?
                          reg2085 : reg1829))));
                    end
                  reg2139 <= ($signed((&$signed(forvar1880))) ?
                      (reg1948[(1'h0):(1'h0)] <<< {(~^reg1971)}) : ({$signed(reg2016)} ?
                          ((|reg1821) <= $signed(reg1866)) : $unsigned({reg1827})));
                end
              else
                begin
                  reg2135 <= $unsigned(forvar1757);
                end
              for (forvar2140 = (1'h0); (forvar2140 < (2'h2)); forvar2140 = (forvar2140 + (1'h1)))
                begin
                  reg2141 <= (~^$unsigned((8'hb2)));
                end
            end
          for (forvar2142 = (1'h0); (forvar2142 < (1'h1)); forvar2142 = (forvar2142 + (1'h1)))
            begin
              if (((~|((reg1807 << reg2050) ?
                  reg1952 : $unsigned(reg2023))) & (8'hae)))
                begin
                  for (forvar2143 = (1'h0); (forvar2143 < (1'h0)); forvar2143 = (forvar2143 + (1'h1)))
                    begin
                      reg2144 <= $signed($unsigned({reg1779[(2'h3):(1'h0)]}));
                      reg2145 <= $signed(forvar1896);
                      reg2146 <= ((((reg2065 ?
                              reg1766 : reg1771) >>> $signed(forvar1845)) >>> $unsigned($unsigned(reg1931))) ?
                          ({forvar1945[(4'hc):(3'h5)]} >> ($signed((8'h9f)) * reg1785)) : (((forvar2058 > (8'h9c)) > $signed(reg1794)) ?
                              $unsigned(reg2004) : $signed((|reg1784))));
                      reg2147 <= ((((forvar2093 ? reg1926 : (8'hae)) ?
                              reg1815[(4'h8):(1'h1)] : forvar2123[(4'hb):(4'h8)]) >= reg2090) ?
                          {$signed($signed(reg1915))} : ($unsigned(reg1847[(1'h1):(1'h0)]) ?
                              ($unsigned(reg1898) ?
                                  $unsigned(forvar1905) : (forvar1986 <<< reg2129)) : {(&forvar1759)}));
                    end
                  for (forvar2148 = (1'h0); (forvar2148 < (2'h2)); forvar2148 = (forvar2148 + (1'h1)))
                    begin
                      reg2149 <= (forvar2068[(2'h2):(2'h2)] ?
                          reg1842 : ($unsigned((reg1844 << reg1767)) <<< (^(reg2132 + forvar2081))));
                    end
                  for (forvar2150 = (1'h0); (forvar2150 < (1'h1)); forvar2150 = (forvar2150 + (1'h1)))
                    begin
                      reg2151 <= forvar1984[(4'ha):(3'h6)];
                    end
                  for (forvar2152 = (1'h0); (forvar2152 < (1'h1)); forvar2152 = (forvar2152 + (1'h1)))
                    begin
                      reg2153 <= forvar1858[(1'h1):(1'h0)];
                      reg2154 <= {($signed((reg1764 <= reg2017)) ?
                              $signed((reg2024 ?
                                  reg2019 : reg1780)) : {reg2001[(3'h5):(3'h4)]})};
                      reg2155 <= ($unsigned(({reg2073} ?
                              $signed(forvar2086) : $unsigned(forvar2143))) ?
                          $unsigned((((8'hb5) > reg2003) == (forvar1955 && reg2111))) : forvar1875[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  if ($signed((reg1987 ~^ ($signed(reg1836) ?
                      $signed(forvar1885) : $signed(forvar1993)))))
                    begin
                      reg2143 <= $unsigned((((reg1947 >= reg1767) > (reg2104 && (8'hb3))) != $signed($unsigned(forvar1856))));
                      reg2144 <= (&reg1792);
                      reg2145 <= reg2059;
                    end
                  else
                    begin
                      reg2143 <= ({(reg1836 ^~ (reg2141 * reg1968))} ?
                          (reg2017 != (!(reg2149 ?
                              (8'ha7) : forvar2142))) : reg2022);
                      reg2144 <= forvar1924;
                      reg2145 <= reg2139;
                      reg2146 <= ({{reg1954[(4'h9):(3'h5)]}} & reg1767[(3'h7):(3'h7)]);
                    end
                  if ((reg1904 ^ {$unsigned($unsigned(forvar1845))}))
                    begin
                      reg2147 <= ($unsigned($unsigned($unsigned(reg2045))) ?
                          (8'ha4) : (8'ha4));
                      reg2148 <= {reg1824[(3'h5):(1'h1)]};
                      reg2149 <= (((^(|forvar1904)) < reg2058) + (^~$signed(((8'ha7) ?
                          reg2019 : forvar1964))));
                    end
                  else
                    begin
                      reg2147 <= {reg2145};
                      reg2148 <= ((|forvar2123) ?
                          $unsigned(($unsigned((8'ha0)) >= $signed((8'had)))) : (&{(reg2139 ?
                                  reg1976 : reg2032)}));
                      reg2149 <= $unsigned(reg1909[(4'h8):(1'h1)]);
                      reg2150 <= (reg1827 >>> $signed({(reg1769 * reg1943)}));
                    end
                end
              for (forvar2156 = (1'h0); (forvar2156 < (2'h2)); forvar2156 = (forvar2156 + (1'h1)))
                begin
                  for (forvar2157 = (1'h0); (forvar2157 < (1'h0)); forvar2157 = (forvar2157 + (1'h1)))
                    begin
                      reg2158 <= reg2155;
                      reg2159 <= $signed(reg2042);
                      reg2160 <= $unsigned(($unsigned({reg1862}) ?
                          (reg1770[(4'hd):(3'h5)] && (reg1827 | reg2118)) : $unsigned(reg2011)));
                    end
                  for (forvar2161 = (1'h0); (forvar2161 < (1'h1)); forvar2161 = (forvar2161 + (1'h1)))
                    begin
                      reg2162 <= reg1835;
                      reg2163 <= $signed((reg2037 ~^ reg1874[(2'h3):(2'h2)]));
                      reg2164 <= (((reg1818 ?
                              (reg1918 ?
                                  reg1941 : reg1883) : (reg1855 ~^ reg2069)) ?
                          reg2143[(3'h5):(1'h1)] : reg2008[(3'h4):(2'h2)]) >= (((reg1941 * reg1864) ?
                          $unsigned(reg1930) : (reg1860 >>> reg1787)) == ((reg2146 ?
                          forvar2051 : reg2085) || (+reg1796))));
                    end
                  if (forvar2110[(3'h5):(1'h0)])
                    begin
                      reg2165 <= $unsigned($signed((8'hb9)));
                      reg2166 <= forvar1809[(1'h1):(1'h1)];
                      reg2167 <= reg1953[(4'h8):(4'h8)];
                    end
                  else
                    begin
                      reg2165 <= forvar1891[(3'h7):(3'h7)];
                    end
                end
            end
        end
      else
        begin
          reg2109 <= {(reg2039[(1'h0):(1'h0)] ?
                  (((8'hb0) * reg2039) >= forvar2093) : (~|$unsigned(reg1967)))};
          for (forvar2110 = (1'h0); (forvar2110 < (2'h2)); forvar2110 = (forvar2110 + (1'h1)))
            begin
              for (forvar2111 = (1'h0); (forvar2111 < (2'h2)); forvar2111 = (forvar2111 + (1'h1)))
                begin
                  for (forvar2112 = (1'h0); (forvar2112 < (1'h1)); forvar2112 = (forvar2112 + (1'h1)))
                    begin
                      reg2113 <= reg2070[(4'hd):(4'hd)];
                      reg2114 <= forvar2143;
                      reg2115 <= reg1789;
                      reg2116 <= reg1826;
                    end
                end
              for (forvar2117 = (1'h0); (forvar2117 < (1'h1)); forvar2117 = (forvar2117 + (1'h1)))
                begin
                  reg2118 <= ($unsigned({$signed(forvar1790)}) != $signed($unsigned($signed(reg1777))));
                  for (forvar2119 = (1'h0); (forvar2119 < (1'h1)); forvar2119 = (forvar2119 + (1'h1)))
                    begin
                      reg2120 <= $signed($signed((8'hb3)));
                      reg2121 <= {(|reg2023)};
                      reg2122 <= $signed({((reg2114 ? reg1919 : reg1769) ?
                              ((8'hb2) > (8'h9e)) : $signed(forvar2124))});
                    end
                  for (forvar2123 = (1'h0); (forvar2123 < (1'h0)); forvar2123 = (forvar2123 + (1'h1)))
                    begin
                      reg2124 <= ((+reg2087) << (reg2058 < ((|forvar2036) ^ (~&reg1883))));
                      reg2125 <= reg1872;
                    end
                  reg2126 <= reg1892[(2'h3):(1'h0)];
                end
              for (forvar2127 = (1'h0); (forvar2127 < (1'h1)); forvar2127 = (forvar2127 + (1'h1)))
                begin
                  if (reg1772[(3'h6):(1'h1)])
                    begin
                      reg2128 <= $signed($unsigned(($signed(reg1779) >> (forvar1885 != reg2062))));
                    end
                  else
                    begin
                      reg2128 <= $signed(($unsigned(forvar1891[(2'h2):(1'h0)]) ^ ($signed(reg2100) ?
                          (8'hae) : $unsigned(reg1872))));
                      reg2129 <= (!(+$signed((reg2160 ^~ reg1987))));
                    end
                  for (forvar2130 = (1'h0); (forvar2130 < (2'h2)); forvar2130 = (forvar2130 + (1'h1)))
                    begin
                      reg2131 <= $signed((^~$unsigned(reg1825)));
                      reg2132 <= {$signed(reg1953)};
                      reg2133 <= (~|reg2141[(3'h7):(3'h7)]);
                      reg2134 <= reg1869[(1'h0):(1'h0)];
                    end
                  for (forvar2135 = (1'h0); (forvar2135 < (1'h1)); forvar2135 = (forvar2135 + (1'h1)))
                    begin
                      reg2136 <= ((-((~forvar1858) ?
                          (reg1852 | reg1766) : (reg1813 ~^ reg2145))) >> (|{(forvar1942 >> reg2132)}));
                      reg2137 <= reg1893;
                    end
                  reg2138 <= (8'hb9);
                end
            end
          reg2139 <= (!{$unsigned((|reg1857))});
        end
    end
  always
    @(posedge clk) begin
      if ({$unsigned({reg1787[(2'h3):(2'h2)]})})
        begin
          if ((!(-reg1912)))
            begin
              for (forvar2168 = (1'h0); (forvar2168 < (1'h1)); forvar2168 = (forvar2168 + (1'h1)))
                begin
                  for (forvar2169 = (1'h0); (forvar2169 < (1'h0)); forvar2169 = (forvar2169 + (1'h1)))
                    begin
                      reg2170 <= ((reg2039[(3'h4):(1'h0)] ?
                          ({reg1833} == $unsigned(forvar2081)) : $signed({reg1837})) != (($signed(reg1981) ?
                              (^~reg2023) : (forvar1775 ^~ forvar2148)) ?
                          ((reg1859 << (8'hab)) > (reg1968 + (8'hb4))) : {(reg1864 ?
                                  (8'h9f) : (8'hac))}));
                      reg2171 <= $signed(forvar1878);
                      reg2172 <= $signed((^reg1917[(4'h9):(3'h6)]));
                      reg2173 <= (8'hb4);
                    end
                  reg2174 <= reg2136[(1'h0):(1'h0)];
                  if (reg2097[(2'h2):(1'h1)])
                    begin
                      reg2175 <= (($unsigned({wire1754}) + reg2124[(2'h2):(2'h2)]) ^~ (reg2003 > {(~^reg1887)}));
                      reg2176 <= reg2046[(4'h9):(3'h5)];
                    end
                  else
                    begin
                      reg2175 <= reg2030[(2'h3):(2'h2)];
                      reg2176 <= ($unsigned(reg1929) ?
                          ((~(&(8'ha2))) + reg2175) : (($signed(forvar1760) ?
                              (forvar1788 ?
                                  (8'h9f) : reg1935) : $signed(reg2022)) ^ reg2074));
                    end
                  for (forvar2177 = (1'h0); (forvar2177 < (2'h2)); forvar2177 = (forvar2177 + (1'h1)))
                    begin
                      reg2178 <= reg1970[(1'h0):(1'h0)];
                    end
                end
              for (forvar2179 = (1'h0); (forvar2179 < (2'h3)); forvar2179 = (forvar2179 + (1'h1)))
                begin
                  for (forvar2180 = (1'h0); (forvar2180 < (2'h3)); forvar2180 = (forvar2180 + (1'h1)))
                    begin
                      reg2181 <= $unsigned(reg2029);
                      reg2182 <= $unsigned(reg1926);
                      reg2183 <= $unsigned(forvar1889[(2'h3):(2'h2)]);
                    end
                  reg2184 <= ((8'haa) ? (8'haf) : {$unsigned((8'hb0))});
                  for (forvar2185 = (1'h0); (forvar2185 < (1'h1)); forvar2185 = (forvar2185 + (1'h1)))
                    begin
                      reg2186 <= reg2047[(4'ha):(4'h9)];
                      reg2187 <= $signed({(!reg2065[(1'h0):(1'h0)])});
                      reg2188 <= $signed(reg1787);
                      reg2189 <= (reg2117 ? reg1928 : reg1898[(3'h7):(3'h7)]);
                    end
                end
              if ({$unsigned((~|(reg1956 + reg1840)))})
                begin
                  reg2190 <= ($signed(({forvar2063} ?
                          reg2074[(2'h3):(1'h1)] : forvar2148[(4'ha):(4'ha)])) ?
                      (($unsigned((8'hb9)) != ((8'hb6) ?
                          reg2108 : reg1953)) | {(reg2031 ~^ forvar1940)}) : (~|(^$unsigned((8'ha7)))));
                  for (forvar2191 = (1'h0); (forvar2191 < (2'h3)); forvar2191 = (forvar2191 + (1'h1)))
                    begin
                      reg2192 <= ((forvar1901 ?
                          (~|(reg2069 & reg2039)) : reg2090[(4'hf):(1'h0)]) | $unsigned($unsigned($unsigned(forvar2112))));
                      reg2193 <= (reg1869[(1'h1):(1'h1)] ?
                          forvar2063 : $signed((8'hb4)));
                      reg2194 <= reg1845[(4'hb):(3'h4)];
                      reg2195 <= (~^((((8'ha6) == reg2117) ?
                          $unsigned(reg1762) : (reg1776 ?
                              (8'h9f) : reg2042)) ^ ((~(8'ha3)) ?
                          $signed(reg1884) : (forvar1986 ?
                              reg1833 : reg1965))));
                    end
                end
              else
                begin
                  for (forvar2190 = (1'h0); (forvar2190 < (2'h3)); forvar2190 = (forvar2190 + (1'h1)))
                    begin
                      reg2191 <= {($unsigned((reg2116 ? (8'ha7) : reg1848)) ?
                              reg1856[(2'h2):(2'h2)] : (((8'h9f) ?
                                  reg1982 : reg2077) ^~ (reg1771 * reg1798)))};
                      reg2192 <= $signed($signed(((8'ha5) << forvar2088)));
                    end
                  reg2193 <= reg2074;
                end
              for (forvar2196 = (1'h0); (forvar2196 < (1'h0)); forvar2196 = (forvar2196 + (1'h1)))
                begin
                  if ((~|forvar1809))
                    begin
                      reg2197 <= reg1778;
                    end
                  else
                    begin
                      reg2197 <= reg2003[(3'h5):(2'h2)];
                      reg2198 <= $unsigned((-(reg2033[(4'h8):(1'h1)] ?
                          $signed(reg1792) : (reg1829 ? reg2005 : reg2038))));
                      reg2199 <= reg1816[(2'h2):(1'h1)];
                    end
                  for (forvar2200 = (1'h0); (forvar2200 < (1'h0)); forvar2200 = (forvar2200 + (1'h1)))
                    begin
                      reg2201 <= forvar1820;
                      reg2202 <= (^~reg2018);
                    end
                  for (forvar2203 = (1'h0); (forvar2203 < (1'h0)); forvar2203 = (forvar2203 + (1'h1)))
                    begin
                      reg2204 <= (forvar2112 && forvar1845[(4'h9):(1'h1)]);
                      reg2205 <= reg1947;
                      reg2206 <= {$unsigned(forvar1808[(2'h3):(1'h1)])};
                    end
                  reg2207 <= reg1784[(4'hb):(3'h6)];
                end
            end
          else
            begin
              for (forvar2168 = (1'h0); (forvar2168 < (2'h3)); forvar2168 = (forvar2168 + (1'h1)))
                begin
                  if (reg2207[(2'h3):(1'h0)])
                    begin
                      reg2169 <= (reg1980[(3'h7):(1'h1)] - (!((-(8'hae)) ?
                          reg1991[(2'h2):(2'h2)] : (!(8'ha1)))));
                      reg2170 <= {(reg1904[(4'ha):(2'h2)] != forvar2068[(4'ha):(1'h1)])};
                    end
                  else
                    begin
                      reg2169 <= (forvar1863 <= reg2172);
                    end
                  if ($signed(reg2012[(3'h4):(2'h2)]))
                    begin
                      reg2171 <= reg1998[(2'h3):(1'h0)];
                      reg2172 <= ((!forvar1923[(2'h2):(2'h2)]) ?
                          {(8'hb3)} : ({$unsigned(reg2172)} ?
                              (+((8'h9d) ?
                                  reg2126 : forvar1803)) : {$signed(reg2039)}));
                      reg2173 <= (8'ha2);
                      reg2174 <= (reg2017[(4'h9):(3'h7)] < ($signed(forvar2131) && (forvar2113 + forvar1759[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg2171 <= reg2058[(2'h2):(1'h0)];
                    end
                  for (forvar2175 = (1'h0); (forvar2175 < (2'h2)); forvar2175 = (forvar2175 + (1'h1)))
                    begin
                      reg2176 <= (reg2080 ?
                          $signed(reg1777) : ($unsigned(reg1957[(1'h0):(1'h0)]) ?
                              ((~&reg1787) != (^~reg2128)) : $signed((reg1919 == (8'haa)))));
                    end
                end
            end
          reg2208 <= forvar1836[(2'h3):(1'h0)];
          for (forvar2209 = (1'h0); (forvar2209 < (2'h2)); forvar2209 = (forvar2209 + (1'h1)))
            begin
              if ($unsigned($unsigned((&reg1953[(3'h7):(2'h2)]))))
                begin
                  reg2210 <= ((~|reg1874[(2'h3):(1'h0)]) ?
                      (^$signed(((8'ha8) >>> reg1762))) : $unsigned(reg2097));
                  for (forvar2211 = (1'h0); (forvar2211 < (2'h3)); forvar2211 = (forvar2211 + (1'h1)))
                    begin
                      reg2212 <= (~&(&{(reg1877 >= (8'hae))}));
                      reg2213 <= {($signed((~|forvar2047)) ?
                              (~(^reg2004)) : reg1921[(4'hb):(3'h5)])};
                    end
                end
              else
                begin
                  if ((((~|{forvar1856}) >> ($unsigned(reg1913) ?
                          $signed((8'hba)) : $unsigned(reg2018))) ?
                      reg1886 : reg2169))
                    begin
                      reg2210 <= (~^((^~(8'hb3)) - reg1948[(1'h0):(1'h0)]));
                      reg2211 <= (({$signed(reg1965)} ?
                          $signed((~forvar1997)) : reg1881[(3'h4):(3'h4)]) + reg2023);
                    end
                  else
                    begin
                      reg2210 <= (&(((8'hba) ?
                          $unsigned(reg2023) : (reg1959 ?
                              reg1908 : reg1992)) && (^~forvar2017[(2'h2):(1'h0)])));
                      reg2211 <= $signed(reg2020);
                      reg2212 <= $unsigned($unsigned({(~&reg2205)}));
                      reg2213 <= reg1802[(4'hc):(4'h8)];
                    end
                end
              if ($signed((reg2109 ?
                  reg1827[(3'h7):(2'h3)] : ((forvar2066 ?
                      (8'ha8) : reg1871) ~^ ((8'ha4) ^~ reg2163)))))
                begin
                  for (forvar2214 = (1'h0); (forvar2214 < (1'h1)); forvar2214 = (forvar2214 + (1'h1)))
                    begin
                      reg2215 <= (|reg1861);
                    end
                  if ((forvar1984[(4'hb):(1'h1)] ?
                      reg1887 : $unsigned(forvar2124)))
                    begin
                      reg2216 <= (8'hba);
                    end
                  else
                    begin
                      reg2216 <= (reg1810[(4'hb):(3'h5)] + reg1883);
                    end
                end
              else
                begin
                  if (($signed(($signed(reg2197) ?
                          $unsigned(reg1811) : {forvar1760})) ?
                      {{(reg2092 ?
                                  forvar2110 : (8'hab))}} : $unsigned(($unsigned(reg2107) || (reg1843 <<< reg2189)))))
                    begin
                      reg2214 <= (&$signed((forvar2015[(4'h8):(4'h8)] >> {reg2025})));
                    end
                  else
                    begin
                      reg2214 <= forvar2148;
                      reg2215 <= $unsigned((+(forvar2203 - forvar1914[(4'h8):(3'h5)])));
                      reg2216 <= reg2070[(4'hc):(4'ha)];
                    end
                  if ($unsigned(((|(+(8'ha7))) == (^~(reg1792 > reg1829)))))
                    begin
                      reg2217 <= $unsigned(({$unsigned(reg1891)} >> ($unsigned(reg1933) - (reg1877 ?
                          (8'hac) : forvar2142))));
                      reg2218 <= $unsigned($unsigned($unsigned((reg2095 >> forvar1788))));
                      reg2219 <= $unsigned(($unsigned((^(8'h9f))) - $signed((reg2195 + (8'hae)))));
                      reg2220 <= {({(reg2116 <<< forvar1923)} ^ (forvar1808 ?
                              reg2124[(4'ha):(3'h7)] : $unsigned(forvar1942)))};
                    end
                  else
                    begin
                      reg2217 <= (reg2164 ?
                          (^{$signed(reg1947)}) : (reg2111 ?
                              {(reg1919 ?
                                      forvar2143 : reg1910)} : {{reg1970}}));
                      reg2218 <= (reg1823 >>> ({$unsigned(forvar2063)} ?
                          $unsigned((forvar1803 ?
                              reg1874 : forvar1803)) : ($signed(reg1800) > reg2169[(3'h5):(3'h5)])));
                    end
                end
              if (($unsigned(((reg1990 ? reg2211 : reg2191) ?
                  (~|reg2197) : $signed(reg1784))) || (+{$signed(reg1850)})))
                begin
                  if ((~|(((|forvar2175) << $unsigned((8'ha1))) ?
                      $signed(reg2126) : $signed((8'hb2)))))
                    begin
                      reg2221 <= (reg1981[(2'h2):(2'h2)] || reg2208);
                      reg2222 <= $unsigned(reg2113);
                      reg2223 <= (~((~reg2053[(2'h3):(1'h1)]) + (reg1842 != (^~(8'h9e)))));
                    end
                  else
                    begin
                      reg2221 <= $unsigned($signed(({reg2144} * (-forvar1867))));
                    end
                end
              else
                begin
                  for (forvar2221 = (1'h0); (forvar2221 < (1'h0)); forvar2221 = (forvar2221 + (1'h1)))
                    begin
                      reg2222 <= $unsigned((&($signed(reg2052) <<< reg1794[(2'h2):(2'h2)])));
                    end
                  if ($signed(($unsigned((reg2165 << reg2186)) + (^~(|forvar2123)))))
                    begin
                      reg2223 <= reg1853[(4'hd):(3'h5)];
                      reg2224 <= reg1851;
                      reg2225 <= (reg1780[(2'h3):(1'h1)] ?
                          $unsigned(((reg2184 == reg1837) ?
                              $unsigned(forvar2131) : $signed(reg1845))) : (8'hb6));
                    end
                  else
                    begin
                      reg2223 <= ($unsigned((|forvar1863)) - ({forvar1904} ?
                          forvar1905 : ((8'had) ? (+forvar2150) : (&reg2145))));
                      reg2224 <= (+$signed((+$unsigned(reg1771))));
                      reg2225 <= ($unsigned((~&reg2112)) ?
                          reg1905[(3'h5):(1'h0)] : $signed((reg2182 ?
                              $unsigned(reg1876) : (reg2024 < reg1791))));
                      reg2226 <= (^((~^reg2201[(2'h3):(2'h3)]) ?
                          {reg1840[(4'ha):(4'h9)]} : $unsigned($unsigned((8'hb1)))));
                    end
                  for (forvar2227 = (1'h0); (forvar2227 < (2'h3)); forvar2227 = (forvar2227 + (1'h1)))
                    begin
                      reg2228 <= (({reg1827} ?
                          reg2033[(4'h8):(2'h2)] : $signed($signed(reg1982))) | $unsigned(reg2215[(1'h1):(1'h0)]));
                      reg2229 <= $signed((-reg1943[(4'h8):(3'h6)]));
                      reg2230 <= ((^~(~&$unsigned(reg2070))) * (-(reg2201[(3'h6):(3'h4)] ?
                          reg1987[(2'h2):(2'h2)] : $unsigned(forvar2177))));
                      reg2231 <= $signed({(reg1996 ?
                              $unsigned(reg2023) : $unsigned(forvar1920))});
                    end
                end
              for (forvar2232 = (1'h0); (forvar2232 < (1'h1)); forvar2232 = (forvar2232 + (1'h1)))
                begin
                  if (reg2001)
                    begin
                      reg2233 <= $signed($unsigned(forvar2024));
                      reg2234 <= $unsigned({{forvar2063}});
                    end
                  else
                    begin
                      reg2233 <= (~&(^(~^(reg2183 ? forvar2168 : reg2125))));
                      reg2234 <= reg2182;
                      reg2235 <= $unsigned(((reg2080 > $unsigned(reg2060)) ?
                          (^~(reg2118 ?
                              forvar1820 : reg1936)) : (|(^reg2037))));
                    end
                  for (forvar2236 = (1'h0); (forvar2236 < (1'h1)); forvar2236 = (forvar2236 + (1'h1)))
                    begin
                      reg2237 <= (forvar2009[(1'h0):(1'h0)] ?
                          forvar2203 : reg2000[(1'h0):(1'h0)]);
                      reg2238 <= $signed((~reg2146));
                      reg2239 <= {((&{forvar1920}) ?
                              $signed((reg2059 ?
                                  reg1873 : reg1792)) : $unsigned(reg1881))};
                      reg2240 <= ((|((reg1978 ?
                              reg1980 : (8'hb3)) < $signed(forvar2030))) ?
                          {((reg2141 ? reg2173 : reg2141) ?
                                  {forvar1786} : reg2235[(4'hd):(4'hd)])} : $signed(($unsigned((8'ha0)) >>> {reg2193})));
                    end
                end
            end
          if ((~reg1991[(2'h3):(2'h2)]))
            begin
              if (reg1857)
                begin
                  for (forvar2241 = (1'h0); (forvar2241 < (2'h3)); forvar2241 = (forvar2241 + (1'h1)))
                    begin
                      reg2242 <= forvar1760[(2'h2):(1'h1)];
                    end
                  for (forvar2243 = (1'h0); (forvar2243 < (1'h0)); forvar2243 = (forvar2243 + (1'h1)))
                    begin
                      reg2244 <= reg1967[(4'hb):(2'h3)];
                      reg2245 <= reg1802[(4'hd):(1'h0)];
                      reg2246 <= $signed(reg1971);
                      reg2247 <= reg2189;
                    end
                  for (forvar2248 = (1'h0); (forvar2248 < (1'h0)); forvar2248 = (forvar2248 + (1'h1)))
                    begin
                      reg2249 <= $signed(forvar2009);
                      reg2250 <= (-((|((8'hb7) & (8'hb7))) ?
                          {(reg1996 | forvar1798)} : ((^~(8'hb2)) ?
                              $unsigned(reg2005) : (reg2214 <<< reg2080))));
                      reg2251 <= ({(+{(8'hab)})} ?
                          reg2076[(2'h2):(1'h1)] : reg1976[(2'h3):(1'h0)]);
                    end
                end
              else
                begin
                  reg2241 <= forvar1836;
                  for (forvar2242 = (1'h0); (forvar2242 < (1'h1)); forvar2242 = (forvar2242 + (1'h1)))
                    begin
                      reg2243 <= $unsigned($unsigned(((forvar1891 || reg2235) < forvar2248[(2'h3):(2'h2)])));
                      reg2244 <= $signed(($signed($unsigned(reg1823)) <<< $signed((~|reg1897))));
                      reg2245 <= reg1917[(3'h5):(2'h2)];
                    end
                end
              for (forvar2252 = (1'h0); (forvar2252 < (1'h0)); forvar2252 = (forvar2252 + (1'h1)))
                begin
                  if ($signed($unsigned($signed((reg2242 ?
                      (8'ha5) : (8'haa))))))
                    begin
                      reg2253 <= $unsigned((reg2144 ?
                          reg1990[(4'hb):(4'h9)] : $signed($signed(reg2150))));
                    end
                  else
                    begin
                      reg2253 <= {({$signed(reg2046)} & $unsigned(reg2182))};
                      reg2254 <= reg2090;
                      reg2255 <= forvar2086[(2'h2):(1'h0)];
                    end
                  for (forvar2256 = (1'h0); (forvar2256 < (1'h0)); forvar2256 = (forvar2256 + (1'h1)))
                    begin
                      reg2257 <= {{((forvar2096 ? reg2158 : (8'h9d)) ?
                                  $unsigned(forvar1920) : {reg2229})}};
                      reg2258 <= ((~{forvar1891[(2'h2):(2'h2)]}) != (reg2024 ?
                          (reg2215[(4'h9):(3'h5)] * (8'hb8)) : $unsigned($unsigned(forvar1781))));
                      reg2259 <= $signed($signed(((reg1915 ?
                          reg2175 : reg2233) + forvar1844[(2'h2):(1'h0)])));
                    end
                  if ((+reg2002))
                    begin
                      reg2260 <= ($unsigned((~|((8'hb9) ?
                              reg2225 : forvar1905))) ?
                          ($signed((reg1956 ^~ (8'ha1))) ?
                              reg1904[(4'hd):(2'h3)] : $signed((|(8'h9e)))) : ((((8'ha5) <= forvar1896) ?
                                  (!reg2042) : $unsigned(reg2122)) ?
                              (-(~|forvar1878)) : forvar1924[(3'h7):(2'h2)]));
                      reg2261 <= $unsigned($unsigned({$signed(forvar2221)}));
                      reg2262 <= reg1948[(1'h1):(1'h0)];
                      reg2263 <= reg2100[(4'h8):(2'h2)];
                    end
                  else
                    begin
                      reg2260 <= (reg1919[(2'h3):(1'h1)] ?
                          {{forvar1977}} : ($signed($unsigned(reg1789)) ?
                              ((reg2111 ?
                                  reg1909 : forvar2232) << forvar1942[(3'h6):(3'h4)]) : forvar2030));
                      reg2261 <= $unsigned($unsigned(($unsigned(reg1836) ?
                          $signed(reg2250) : (~(8'hb1)))));
                    end
                end
              for (forvar2264 = (1'h0); (forvar2264 < (2'h3)); forvar2264 = (forvar2264 + (1'h1)))
                begin
                  for (forvar2265 = (1'h0); (forvar2265 < (1'h0)); forvar2265 = (forvar2265 + (1'h1)))
                    begin
                      reg2266 <= $signed((((reg2224 ?
                              forvar2203 : reg2095) ~^ $signed((8'ha4))) ?
                          ((-forvar2177) ?
                              (reg1823 & reg1829) : reg1880) : reg2075));
                      reg2267 <= (~&$unsigned((8'h9e)));
                      reg2268 <= $signed(reg1900[(1'h1):(1'h1)]);
                    end
                  for (forvar2269 = (1'h0); (forvar2269 < (2'h3)); forvar2269 = (forvar2269 + (1'h1)))
                    begin
                      reg2270 <= $unsigned((^($signed(reg2176) ?
                          (reg1964 ? reg1935 : reg2025) : $unsigned((8'had)))));
                      reg2271 <= $unsigned($signed(forvar1844[(1'h1):(1'h1)]));
                    end
                  if ((($unsigned((forvar2179 != reg2235)) != (^(|reg2221))) ?
                      ((!(&reg2181)) < (&{reg2122})) : ($unsigned($unsigned(reg2254)) ?
                          (forvar2156[(3'h5):(1'h1)] ?
                              (^~forvar2009) : {reg1870}) : $signed((forvar2093 >= forvar1808)))))
                    begin
                      reg2272 <= $unsigned(reg1959[(3'h4):(2'h3)]);
                      reg2273 <= $signed(reg1811);
                    end
                  else
                    begin
                      reg2272 <= $unsigned(((reg2027[(3'h4):(3'h4)] ?
                              reg2145 : (forvar2081 ^ (8'hab))) ?
                          (reg2220 != reg2181[(3'h4):(1'h0)]) : ((^~(8'hb8)) * (~&(8'h9e)))));
                    end
                end
              reg2274 <= (^$unsigned((reg2084 <= {forvar2256})));
            end
          else
            begin
              for (forvar2241 = (1'h0); (forvar2241 < (2'h3)); forvar2241 = (forvar2241 + (1'h1)))
                begin
                  for (forvar2242 = (1'h0); (forvar2242 < (2'h3)); forvar2242 = (forvar2242 + (1'h1)))
                    begin
                      reg2243 <= reg1904[(1'h0):(1'h0)];
                      reg2244 <= reg1870;
                      reg2245 <= (^$unsigned(((forvar2150 ?
                              forvar2130 : reg1943) ?
                          forvar2066 : reg2240)));
                      reg2246 <= {((~|(reg2151 ?
                              (8'hb0) : reg1937)) >= (reg1912[(1'h1):(1'h1)] ?
                              (reg2250 || reg1952) : (forvar2200 * forvar1757)))};
                    end
                  for (forvar2247 = (1'h0); (forvar2247 < (1'h0)); forvar2247 = (forvar2247 + (1'h1)))
                    begin
                      reg2248 <= forvar2232[(1'h0):(1'h0)];
                      reg2249 <= (~&(+$signed((reg1876 ? reg1913 : reg2204))));
                      reg2250 <= forvar1817;
                    end
                  if ($signed(($unsigned((reg2220 ? forvar1951 : reg2014)) ?
                      ($unsigned((8'ha6)) ?
                          reg2120 : ((8'hb3) ^~ reg1921)) : (reg2097[(1'h0):(1'h0)] + $unsigned(reg2189)))))
                    begin
                      reg2251 <= $unsigned({{reg1820}});
                      reg2252 <= reg2107[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2251 <= $signed(((((8'h9d) >= (8'hae)) >> (forvar2148 ?
                              reg1835 : reg1823)) ?
                          reg1842[(3'h5):(2'h2)] : $signed(reg1953)));
                      reg2252 <= ($unsigned((-reg1859[(1'h1):(1'h0)])) << $signed($signed(reg2188)));
                      reg2253 <= $signed((forvar1891 ?
                          ($signed(reg2113) ?
                              $unsigned(forvar2264) : (reg2077 > reg2254)) : {(reg2079 ?
                                  (8'ha4) : forvar1840)}));
                      reg2254 <= $unsigned((($unsigned(reg1962) >> (~^reg1991)) ?
                          ({reg1765} - (^~(8'haf))) : (8'hac)));
                    end
                end
              if (((&{(reg2074 | reg1852)}) ?
                  reg2220[(1'h1):(1'h0)] : reg2083[(4'he):(4'hc)]))
                begin
                  reg2255 <= {$signed($unsigned((!reg2042)))};
                  if ($unsigned($signed($signed($unsigned(reg2124)))))
                    begin
                      reg2256 <= (+reg2202);
                      reg2257 <= ($signed(((reg1990 ?
                              (8'hae) : reg1880) >= {forvar1844})) ?
                          $signed($signed((forvar1858 ~^ reg2105))) : ((8'ha6) ?
                              ($unsigned(reg2005) <= forvar2140[(1'h0):(1'h0)]) : (reg2040 ^~ $unsigned(reg2028))));
                      reg2258 <= wire2007;
                      reg2259 <= (-(~&forvar1865[(4'h8):(3'h7)]));
                    end
                  else
                    begin
                      reg2256 <= $unsigned((8'hb1));
                      reg2257 <= {$signed($signed((forvar2180 - reg2084)))};
                    end
                  if (((!$signed(forvar2078)) && (&{$unsigned(forvar2185)})))
                    begin
                      reg2260 <= ((!$signed((~^(8'hb8)))) ?
                          $unsigned(($unsigned(reg1894) ?
                              reg2250 : (reg2129 << forvar2214))) : reg2017[(4'he):(1'h1)]);
                    end
                  else
                    begin
                      reg2260 <= reg2210[(3'h7):(3'h5)];
                    end
                  reg2261 <= (8'ha2);
                end
              else
                begin
                  for (forvar2255 = (1'h0); (forvar2255 < (2'h2)); forvar2255 = (forvar2255 + (1'h1)))
                    begin
                      reg2256 <= (~reg2050);
                      reg2257 <= ((~{$unsigned((8'hb3))}) - {$unsigned({reg2160})});
                      reg2258 <= $signed($unsigned(reg2189));
                      reg2259 <= ($signed(forvar2156[(4'h8):(3'h4)]) ?
                          (+$signed(((8'h9f) ?
                              reg1795 : reg1778))) : (!{(8'hb4)}));
                    end
                end
              for (forvar2262 = (1'h0); (forvar2262 < (2'h3)); forvar2262 = (forvar2262 + (1'h1)))
                begin
                  for (forvar2263 = (1'h0); (forvar2263 < (1'h1)); forvar2263 = (forvar2263 + (1'h1)))
                    begin
                      reg2264 <= {((~^$unsigned(reg1844)) == $signed((reg2189 ?
                              forvar1955 : reg1884)))};
                      reg2265 <= reg1802[(4'h9):(4'h8)];
                      reg2266 <= reg2026;
                      reg2267 <= reg2055;
                    end
                  for (forvar2268 = (1'h0); (forvar2268 < (2'h2)); forvar2268 = (forvar2268 + (1'h1)))
                    begin
                      reg2269 <= $signed($signed($signed(forvar2140[(1'h0):(1'h0)])));
                      reg2270 <= {($unsigned($signed(forvar2264)) || $unsigned(forvar1790[(3'h5):(3'h5)]))};
                      reg2271 <= (~&(((~^forvar1983) ^ (forvar2111 != reg2011)) & {$signed(forvar2055)}));
                    end
                  if ((reg2111[(4'h9):(4'h9)] ?
                      ((reg2151[(3'h5):(1'h1)] + (forvar2086 | reg1821)) >= ((forvar2262 ?
                          reg2034 : (8'ha9)) >>> (&reg1957))) : ({{reg1824}} | forvar2015)))
                    begin
                      reg2272 <= $signed($signed((+$unsigned(reg2015))));
                      reg2273 <= reg2223;
                    end
                  else
                    begin
                      reg2272 <= reg1988;
                      reg2273 <= {{((reg2250 >>> reg2089) ^ (forvar2023 ?
                                  reg2167 : wire1755))}};
                      reg2274 <= reg1857;
                    end
                end
              for (forvar2275 = (1'h0); (forvar2275 < (1'h0)); forvar2275 = (forvar2275 + (1'h1)))
                begin
                  for (forvar2276 = (1'h0); (forvar2276 < (2'h3)); forvar2276 = (forvar2276 + (1'h1)))
                    begin
                      reg2277 <= ((($signed(reg2045) || $signed(forvar2209)) ?
                              reg2031[(4'ha):(3'h7)] : (((8'hb1) ?
                                  reg1973 : (8'ha6)) < $signed(reg1926))) ?
                          $signed({reg2053}) : (((reg1971 & reg1981) > (reg2228 && forvar1905)) ?
                              (reg2187 > ((8'h9e) ?
                                  forvar2123 : wire1756)) : (-(reg2091 ~^ reg1850))));
                      reg2278 <= $signed(reg1936[(1'h0):(1'h0)]);
                    end
                  if ($unsigned((((^~reg1866) ?
                      ((8'hb5) & reg1840) : {forvar1901}) < (reg1829 <<< forvar2117[(1'h1):(1'h0)]))))
                    begin
                      reg2279 <= $unsigned((reg1903 > (+forvar1803[(3'h4):(3'h4)])));
                      reg2280 <= reg2060[(3'h6):(1'h0)];
                      reg2281 <= (-reg2134[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2279 <= $signed($unsigned(reg2119[(1'h1):(1'h0)]));
                      reg2280 <= $unsigned(forvar1865[(1'h0):(1'h0)]);
                      reg2281 <= $unsigned((8'had));
                      reg2282 <= (|(8'hb5));
                    end
                  for (forvar2283 = (1'h0); (forvar2283 < (2'h3)); forvar2283 = (forvar2283 + (1'h1)))
                    begin
                      reg2284 <= ($unsigned($signed({forvar1808})) ?
                          ((^((8'ha3) ? reg2128 : reg2064)) <<< (-(reg2183 ?
                              reg2173 : reg2070))) : {(!$unsigned(reg2245))});
                      reg2285 <= forvar2009[(4'hc):(4'hb)];
                      reg2286 <= reg2017;
                    end
                end
            end
        end
      else
        begin
          reg2168 <= (|reg1913[(3'h4):(2'h2)]);
          if (({(+reg1844[(2'h2):(1'h1)])} ?
              reg2137[(1'h0):(1'h0)] : $unsigned(((reg1900 ?
                      reg2147 : (8'h9d)) ?
                  forvar2276[(1'h0):(1'h0)] : ((8'hb3) & reg2248)))))
            begin
              for (forvar2169 = (1'h0); (forvar2169 < (1'h1)); forvar2169 = (forvar2169 + (1'h1)))
                begin
                  for (forvar2170 = (1'h0); (forvar2170 < (1'h0)); forvar2170 = (forvar2170 + (1'h1)))
                    begin
                      reg2171 <= $signed(reg2147[(4'he):(4'h8)]);
                      reg2172 <= ((8'h9c) << {$signed($signed(reg1852))});
                      reg2173 <= forvar1800;
                      reg2174 <= $unsigned($signed(($signed(forvar2036) ?
                          $signed(reg2247) : reg1851)));
                    end
                  for (forvar2175 = (1'h0); (forvar2175 < (1'h1)); forvar2175 = (forvar2175 + (1'h1)))
                    begin
                      reg2176 <= ($unsigned($signed((~reg2178))) | $signed((+{reg2273})));
                      reg2177 <= reg2055[(3'h7):(3'h4)];
                      reg2178 <= (~((~$unsigned(reg2103)) ?
                          $signed($signed(reg1832)) : {(reg1822 != forvar1858)}));
                      reg2179 <= reg2034[(4'h9):(3'h7)];
                    end
                end
              reg2180 <= (~^reg1887);
            end
          else
            begin
              if ((~^(~|$signed($unsigned(reg2175)))))
                begin
                  for (forvar2169 = (1'h0); (forvar2169 < (2'h3)); forvar2169 = (forvar2169 + (1'h1)))
                    begin
                      reg2170 <= {(^~((~&reg2014) > $unsigned(reg1909)))};
                      reg2171 <= {(&reg2201)};
                      reg2172 <= forvar1983;
                      reg2173 <= (|((forvar2117[(2'h3):(1'h1)] * $signed(reg1931)) || $signed((reg2013 << reg2016))));
                    end
                  reg2174 <= (reg2003[(1'h0):(1'h0)] ?
                      reg1990[(3'h5):(3'h4)] : (8'haa));
                  for (forvar2175 = (1'h0); (forvar2175 < (1'h0)); forvar2175 = (forvar2175 + (1'h1)))
                    begin
                      reg2176 <= reg1847[(1'h0):(1'h0)];
                      reg2177 <= reg1992[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar2169 = (1'h0); (forvar2169 < (2'h3)); forvar2169 = (forvar2169 + (1'h1)))
                    begin
                      reg2170 <= reg1776;
                      reg2171 <= $unsigned(($unsigned((forvar1836 * reg1807)) ?
                          $unsigned(reg2116) : (8'hab)));
                      reg2172 <= forvar2169[(3'h4):(1'h0)];
                    end
                  for (forvar2173 = (1'h0); (forvar2173 < (1'h1)); forvar2173 = (forvar2173 + (1'h1)))
                    begin
                      reg2174 <= ((reg2057[(1'h1):(1'h0)] && ((reg2139 ?
                          (8'had) : reg2083) <<< {reg1980})) <<< $unsigned((~^(reg2149 ?
                          reg1936 : reg2178))));
                      reg2175 <= $unsigned(reg1807[(1'h1):(1'h0)]);
                      reg2176 <= $unsigned($unsigned(reg2198));
                      reg2177 <= ($signed(((~^(8'ha7)) ?
                          $unsigned(reg1912) : forvar2161)) >>> reg1825);
                    end
                  if ((~($signed($unsigned(reg2132)) ?
                      (~|$unsigned(reg2249)) : ((~^reg2018) ?
                          {reg2114} : reg2122[(2'h2):(1'h0)]))))
                    begin
                      reg2178 <= reg2270;
                      reg2179 <= ({(^(^~reg1988))} * (8'ha8));
                      reg2180 <= $signed((reg2052[(2'h2):(1'h0)] ?
                          (reg2155[(2'h3):(2'h2)] * $signed(reg1769)) : $unsigned($unsigned(reg2102))));
                      reg2181 <= ((((reg2117 ?
                              reg1952 : (8'hb2)) ^~ $signed(reg2268)) > $signed(((8'had) ?
                              reg2125 : (8'hb0)))) ?
                          (forvar1974 ~^ reg1861[(1'h0):(1'h0)]) : reg2096);
                    end
                  else
                    begin
                      reg2178 <= $signed(reg2109[(4'h9):(2'h3)]);
                      reg2179 <= reg1787;
                    end
                  reg2182 <= $unsigned((~|(reg2103[(2'h2):(1'h1)] >>> $signed(forvar2088))));
                end
              if ($unsigned({{$signed(forvar1950)}}))
                begin
                  for (forvar2183 = (1'h0); (forvar2183 < (2'h3)); forvar2183 = (forvar2183 + (1'h1)))
                    begin
                      reg2184 <= $signed(reg2198);
                      reg2185 <= (({$signed(reg2262)} ?
                              (|$unsigned((8'hb3))) : {$unsigned((8'had))}) ?
                          {((&(8'hb9)) ?
                                  forvar1799[(4'hc):(3'h4)] : forvar2152)} : forvar2191[(1'h1):(1'h0)]);
                      reg2186 <= ((^~forvar1939[(3'h4):(3'h4)]) ?
                          $signed((~&$signed((8'h9e)))) : reg1842[(1'h0):(1'h0)]);
                      reg2187 <= (((|$unsigned((8'hae))) != forvar2168[(4'h9):(3'h4)]) ?
                          (8'h9f) : reg1887);
                    end
                  for (forvar2188 = (1'h0); (forvar2188 < (1'h1)); forvar2188 = (forvar2188 + (1'h1)))
                    begin
                      reg2189 <= $unsigned((((~&forvar2066) ?
                          $signed((8'ha9)) : (reg1872 << reg2181)) <<< {(reg1782 ?
                              reg1990 : reg1849)}));
                    end
                  if ($unsigned((~|{(reg2238 >= forvar1788)})))
                    begin
                      reg2190 <= (~^$signed($unsigned(reg2019)));
                      reg2191 <= (((!(forvar1889 ? forvar1955 : reg2083)) ?
                          forvar1939[(3'h5):(2'h3)] : $signed(forvar2183[(4'h9):(4'h9)])) != ($signed((~&reg1881)) <<< $unsigned((reg2216 ?
                          (8'ha0) : reg2131))));
                    end
                  else
                    begin
                      reg2190 <= {($signed($unsigned(reg2267)) ?
                              forvar1799 : $unsigned(forvar1902[(1'h1):(1'h0)]))};
                    end
                end
              else
                begin
                  if (($signed((8'hb4)) ?
                      (-$unsigned($unsigned(reg2045))) : (^~{(~&(8'hb9))})))
                    begin
                      reg2183 <= reg2183;
                      reg2184 <= reg2163[(3'h4):(1'h1)];
                      reg2185 <= ($unsigned($unsigned((reg1880 ?
                          reg1873 : (8'hb2)))) && {reg2067});
                      reg2186 <= reg1821;
                    end
                  else
                    begin
                      reg2183 <= ($signed($signed((8'ha2))) & $signed(forvar1760[(2'h3):(1'h0)]));
                    end
                  for (forvar2187 = (1'h0); (forvar2187 < (2'h3)); forvar2187 = (forvar2187 + (1'h1)))
                    begin
                      reg2188 <= (^(+reg2269[(3'h5):(2'h3)]));
                      reg2189 <= $signed($unsigned($unsigned((~reg1846))));
                    end
                  if ({$unsigned((reg2176[(4'h9):(1'h0)] ?
                          $signed((8'had)) : forvar2131))})
                    begin
                      reg2190 <= $unsigned((~&({forvar1902} ?
                          (reg2005 < reg2090) : (reg2240 ?
                              reg2279 : (8'ha4)))));
                    end
                  else
                    begin
                      reg2190 <= forvar2023[(1'h1):(1'h0)];
                      reg2191 <= $signed($unsigned($unsigned((~|reg1964))));
                      reg2192 <= $signed(($signed((^~reg2136)) ^ reg2141[(3'h4):(1'h1)]));
                      reg2193 <= reg2037;
                    end
                  reg2194 <= (reg2228 ?
                      $unsigned((reg2251[(3'h6):(1'h0)] ?
                          (8'ha0) : reg1852[(3'h7):(2'h3)])) : forvar2009);
                end
              for (forvar2195 = (1'h0); (forvar2195 < (2'h2)); forvar2195 = (forvar2195 + (1'h1)))
                begin
                  for (forvar2196 = (1'h0); (forvar2196 < (1'h1)); forvar2196 = (forvar2196 + (1'h1)))
                    begin
                      reg2197 <= $unsigned((8'ha2));
                    end
                end
              if ((($unsigned((forvar1863 << forvar2123)) ?
                      (-reg1776[(1'h0):(1'h0)]) : ((!reg1823) * (-reg2010))) ?
                  $unsigned(reg2126[(4'hc):(1'h0)]) : {$signed((^reg1820))}))
                begin
                  if (((!(&$signed(reg2066))) ^~ (8'hb1)))
                    begin
                      reg2198 <= (!$signed(($signed(reg2065) != $unsigned(reg1864))));
                      reg2199 <= ($signed((8'hae)) ?
                          $unsigned((forvar2075[(3'h6):(1'h1)] ?
                              $signed(reg2052) : (reg2277 ?
                                  reg1976 : (8'h9d)))) : reg1769);
                      reg2200 <= (|reg1845);
                    end
                  else
                    begin
                      reg2198 <= reg1761[(1'h1):(1'h0)];
                      reg2199 <= reg1996;
                      reg2200 <= ((&$unsigned((^~reg2060))) * reg1921);
                    end
                  for (forvar2201 = (1'h0); (forvar2201 < (1'h0)); forvar2201 = (forvar2201 + (1'h1)))
                    begin
                      reg2202 <= (^~(+(~&(reg2233 != reg2001))));
                      reg2203 <= {$signed($unsigned(reg2092))};
                    end
                  if ($signed($unsigned($unsigned((forvar2140 < reg2117)))))
                    begin
                      reg2204 <= forvar2221;
                      reg2205 <= (($unsigned(forvar1840[(1'h0):(1'h0)]) ?
                          (reg2149 && (-reg2150)) : ((~^reg2067) > $signed(forvar1880))) ~^ (forvar1896 ^~ $unsigned(((8'hb2) ?
                          forvar2017 : (8'hab)))));
                      reg2206 <= forvar2110;
                    end
                  else
                    begin
                      reg2204 <= {reg1969};
                      reg2205 <= $unsigned(($signed($unsigned(reg2092)) ?
                          $unsigned((reg2118 <= reg2184)) : {(reg1776 << (8'haa))}));
                      reg2206 <= forvar1983[(4'h9):(2'h3)];
                    end
                end
              else
                begin
                  if ((+reg2018))
                    begin
                      reg2198 <= {$unsigned($unsigned(forvar2130))};
                      reg2199 <= {((!$signed(reg2135)) != forvar1997)};
                      reg2200 <= forvar2209;
                      reg2201 <= $unsigned(($unsigned((forvar2248 ?
                          forvar2180 : (8'hb5))) >> $unsigned(reg2045)));
                    end
                  else
                    begin
                      reg2198 <= $unsigned($signed(($signed(reg1829) << ((8'ha8) - reg1827))));
                      reg2199 <= ({(((8'hab) ?
                              reg2144 : forvar2169) <= $signed((8'hb8)))} ~^ reg2191);
                    end
                  for (forvar2202 = (1'h0); (forvar2202 < (2'h2)); forvar2202 = (forvar2202 + (1'h1)))
                    begin
                      reg2203 <= (forvar2150 ?
                          (((^~reg2248) ?
                                  (reg2030 >= forvar1896) : (reg1976 ?
                                      reg2244 : reg2234)) ?
                              forvar1773[(2'h2):(2'h2)] : forvar2077[(4'h8):(3'h6)]) : reg2200[(3'h6):(3'h5)]);
                      reg2204 <= reg2169;
                      reg2205 <= ({$unsigned($unsigned(reg1849))} ?
                          (^{reg2141}) : $unsigned((((8'ha9) ^~ forvar1773) * $signed(forvar2087))));
                      reg2206 <= $unsigned((forvar1878[(1'h0):(1'h0)] ^~ $signed(forvar1994)));
                    end
                end
            end
          for (forvar2207 = (1'h0); (forvar2207 < (2'h2)); forvar2207 = (forvar2207 + (1'h1)))
            begin
              if ({$signed($unsigned((~reg2013)))})
                begin
                  for (forvar2208 = (1'h0); (forvar2208 < (1'h0)); forvar2208 = (forvar2208 + (1'h1)))
                    begin
                      reg2209 <= ($unsigned($signed({reg2082})) ?
                          (((!wire1753) ^ {reg1933}) & $signed((!reg1811))) : $signed($unsigned(reg1767[(4'h9):(4'h9)])));
                      reg2210 <= ($signed({(!forvar2179)}) - (-forvar2169));
                      reg2211 <= (^~((8'ha2) >>> forvar2236));
                      reg2212 <= $signed($unsigned($signed(((8'hb2) == reg2246))));
                    end
                  if (($unsigned((8'ha9)) ?
                      (^~(((8'h9e) >= reg1893) * reg2006)) : $signed(reg1766[(4'hc):(3'h4)])))
                    begin
                      reg2213 <= {(8'ha1)};
                      reg2214 <= (reg2094[(2'h3):(2'h3)] ^~ {((~&reg2264) ?
                              (reg2250 ? reg1769 : reg1956) : (~|reg2224))});
                      reg2215 <= reg2220;
                    end
                  else
                    begin
                      reg2213 <= $unsigned({$signed(reg1991[(1'h0):(1'h0)])});
                      reg2214 <= (reg1982[(2'h2):(1'h0)] ?
                          reg1931[(4'hd):(1'h0)] : (($unsigned(reg2198) != (^reg1930)) ?
                              $unsigned(reg2222) : reg2091));
                      reg2215 <= (((-forvar2088[(3'h5):(1'h0)]) ?
                          forvar2236 : reg2246) ~^ ($unsigned(reg1764[(2'h2):(2'h2)]) < (^~forvar2044)));
                    end
                end
              else
                begin
                  for (forvar2208 = (1'h0); (forvar2208 < (2'h3)); forvar2208 = (forvar2208 + (1'h1)))
                    begin
                      reg2209 <= ($unsigned((&(reg1846 ?
                              reg2268 : forvar1950))) ?
                          reg1771 : $signed($unsigned($signed(reg1831))));
                      reg2210 <= $unsigned(($unsigned(reg2103[(2'h2):(2'h2)]) ^~ forvar2117[(3'h7):(3'h6)]));
                      reg2211 <= $signed((&reg2079));
                    end
                  reg2212 <= $unsigned({(~^$signed(reg1821))});
                  if ((8'hba))
                    begin
                      reg2213 <= forvar2161;
                    end
                  else
                    begin
                      reg2213 <= (reg2183[(1'h1):(1'h0)] & {$signed($signed(reg2005))});
                      reg2214 <= ((forvar1983[(4'hd):(1'h1)] ?
                          $signed(reg2195) : (forvar2275[(3'h5):(3'h4)] ?
                              wire1756[(2'h3):(2'h3)] : (reg2224 ?
                                  reg2267 : forvar2180))) < (reg2024[(2'h2):(1'h0)] ?
                          $signed((8'hb9)) : (!(reg2278 ? reg2099 : (8'h9d)))));
                      reg2215 <= ((forvar2208 ?
                              reg1981[(3'h5):(3'h5)] : $unsigned($signed(reg2160))) ?
                          $signed(reg2189[(2'h3):(2'h3)]) : $signed((~$signed(reg1979))));
                    end
                end
              if ((forvar2183 ? (reg1844 >> $unsigned({forvar2243})) : (8'hb5)))
                begin
                  for (forvar2216 = (1'h0); (forvar2216 < (2'h2)); forvar2216 = (forvar2216 + (1'h1)))
                    begin
                      reg2217 <= (reg1861[(2'h3):(1'h0)] ?
                          $unsigned(($unsigned(forvar2056) ?
                              $unsigned(reg2235) : (reg1880 ^~ (8'hab)))) : $signed(($unsigned(reg2103) ?
                              (|forvar2262) : ((8'ha6) << forvar2056))));
                      reg2218 <= {($signed((reg2186 ^~ reg2071)) ?
                              $signed((reg2138 ?
                                  reg1981 : forvar1889)) : ((~reg1872) ?
                                  (8'ha7) : (+forvar1854)))};
                      reg2219 <= ($signed($unsigned((~^(8'hba)))) < (reg2284[(2'h2):(1'h1)] <<< reg2126[(4'ha):(4'ha)]));
                    end
                  for (forvar2220 = (1'h0); (forvar2220 < (2'h2)); forvar2220 = (forvar2220 + (1'h1)))
                    begin
                      reg2221 <= {$signed(((^reg1853) ?
                              (reg2164 ^~ reg1932) : ((8'hb6) >= reg2282)))};
                      reg2222 <= {$unsigned(((reg2171 && reg1839) == $signed(reg1855)))};
                      reg2223 <= (~^(reg1765 ?
                          {(forvar1798 & forvar1878)} : $signed(forvar2190[(3'h4):(2'h2)])));
                      reg2224 <= (-($signed(reg1961[(2'h2):(2'h2)]) ?
                          $signed((reg2022 && reg2145)) : reg1798[(1'h1):(1'h1)]));
                    end
                  for (forvar2225 = (1'h0); (forvar2225 < (1'h0)); forvar2225 = (forvar2225 + (1'h1)))
                    begin
                      reg2226 <= {{forvar2225[(3'h4):(2'h3)]}};
                      reg2227 <= $unsigned(($signed({reg1841}) ?
                          ((forvar1836 >>> forvar1939) < forvar2068[(3'h4):(1'h0)]) : reg2223[(3'h6):(2'h2)]));
                      reg2228 <= reg1892[(4'hb):(4'hb)];
                      reg2229 <= reg2139;
                    end
                  for (forvar2230 = (1'h0); (forvar2230 < (1'h0)); forvar2230 = (forvar2230 + (1'h1)))
                    begin
                      reg2231 <= ($signed((!$signed(reg1898))) ?
                          (|reg2249) : (reg2116 ?
                              reg2267 : (!$signed((8'hb7)))));
                      reg2232 <= (reg1835[(3'h7):(3'h5)] ?
                          (^$signed($signed(reg1789))) : ({forvar1863} >= (~^reg2285)));
                    end
                end
              else
                begin
                  for (forvar2216 = (1'h0); (forvar2216 < (1'h0)); forvar2216 = (forvar2216 + (1'h1)))
                    begin
                      reg2217 <= reg1919;
                      reg2218 <= (-reg2153[(3'h6):(2'h2)]);
                      reg2219 <= (8'hb9);
                      reg2220 <= $unsigned($unsigned(reg2093[(4'hd):(4'ha)]));
                    end
                end
            end
        end
      if (((({reg1886} << reg2163[(1'h1):(1'h1)]) ?
          $signed(reg1935[(2'h3):(1'h1)]) : $signed($unsigned(reg2237))) && (reg2023 ~^ $signed(reg1918))))
        begin
          if ({$signed(((forvar1963 ?
                  reg1776 : reg1895) == (reg1998 ^ (8'ha6))))})
            begin
              for (forvar2287 = (1'h0); (forvar2287 < (1'h1)); forvar2287 = (forvar2287 + (1'h1)))
                begin
                  if ($signed((!forvar1983[(4'h8):(3'h6)])))
                    begin
                      reg2288 <= reg2001[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2288 <= (&{((8'ha2) <<< reg1849)});
                      reg2289 <= forvar1786[(3'h5):(2'h2)];
                    end
                  for (forvar2290 = (1'h0); (forvar2290 < (1'h1)); forvar2290 = (forvar2290 + (1'h1)))
                    begin
                      reg2291 <= reg1851;
                      reg2292 <= ($unsigned($signed(reg2291[(1'h0):(1'h0)])) != (((reg2254 == (8'hb2)) ?
                              (forvar2256 ? reg2039 : reg2282) : (~reg1793)) ?
                          reg2197 : $signed((forvar1946 == reg1887))));
                      reg2293 <= reg2207[(2'h2):(1'h1)];
                      reg2294 <= (~&{$signed($signed(forvar2230))});
                    end
                  if ((+(reg2075[(1'h1):(1'h0)] - $signed((reg2237 & forvar2030)))))
                    begin
                      reg2295 <= (~&$unsigned($signed($signed(forvar2179))));
                      reg2296 <= $unsigned(reg1766);
                    end
                  else
                    begin
                      reg2295 <= reg1791;
                    end
                  if ($unsigned($unsigned($signed(reg1964[(1'h0):(1'h0)]))))
                    begin
                      reg2297 <= (~^((~&$signed(reg2095)) != forvar2161));
                      reg2298 <= {($unsigned((reg2034 ?
                              reg2166 : forvar1942)) & $signed($signed(forvar2263)))};
                    end
                  else
                    begin
                      reg2297 <= $signed(reg2120[(4'ha):(4'ha)]);
                      reg2298 <= reg2281;
                      reg2299 <= $signed(((&(reg1841 >= reg1769)) != $signed($signed(reg1821))));
                    end
                end
              for (forvar2300 = (1'h0); (forvar2300 < (2'h3)); forvar2300 = (forvar2300 + (1'h1)))
                begin
                  reg2301 <= reg1976[(4'h9):(1'h0)];
                  for (forvar2302 = (1'h0); (forvar2302 < (2'h2)); forvar2302 = (forvar2302 + (1'h1)))
                    begin
                      reg2303 <= $unsigned(forvar2179[(4'hb):(1'h0)]);
                      reg2304 <= (!{forvar1865[(2'h2):(1'h1)]});
                    end
                end
              if (reg2165)
                begin
                  for (forvar2305 = (1'h0); (forvar2305 < (2'h2)); forvar2305 = (forvar2305 + (1'h1)))
                    begin
                      reg2306 <= (8'hae);
                    end
                end
              else
                begin
                  if (reg1964[(1'h0):(1'h0)])
                    begin
                      reg2305 <= $unsigned(forvar1817);
                      reg2306 <= (8'haf);
                    end
                  else
                    begin
                      reg2305 <= ($signed(((^~reg2148) & (~^reg1853))) ?
                          (&$unsigned({reg1821})) : (8'h9d));
                    end
                end
              for (forvar2307 = (1'h0); (forvar2307 < (2'h3)); forvar2307 = (forvar2307 + (1'h1)))
                begin
                  reg2308 <= reg2225[(4'hb):(1'h0)];
                end
            end
          else
            begin
              reg2287 <= $unsigned($unsigned(forvar2117));
              if (reg1978)
                begin
                  if ((reg2271[(1'h1):(1'h1)] | {$unsigned((8'had))}))
                    begin
                      reg2288 <= {$unsigned($unsigned(reg1910[(4'hd):(3'h7)]))};
                      reg2289 <= reg2160[(4'h8):(1'h0)];
                      reg2290 <= $unsigned({reg2229[(3'h5):(1'h0)]});
                    end
                  else
                    begin
                      reg2288 <= $signed($unsigned($unsigned($signed(forvar2030))));
                      reg2289 <= {(forvar2191[(4'hb):(4'ha)] ?
                              $unsigned($signed((8'h9c))) : reg1794)};
                    end
                  for (forvar2291 = (1'h0); (forvar2291 < (2'h2)); forvar2291 = (forvar2291 + (1'h1)))
                    begin
                      reg2292 <= ((({reg1825} >> $unsigned(reg1970)) | (forvar1845 * (wire1753 ?
                          reg2020 : (8'hb0)))) | (-(8'h9f)));
                      reg2293 <= (~^$unsigned($signed($signed(forvar2209))));
                      reg2294 <= ((^~reg1959[(4'ha):(1'h1)]) >> $unsigned($signed($signed(reg2143))));
                    end
                end
              else
                begin
                  if ({($unsigned((reg1851 == reg1961)) & reg2104[(2'h2):(1'h1)])})
                    begin
                      reg2288 <= (&reg2192[(1'h1):(1'h1)]);
                      reg2289 <= $unsigned((forvar2230[(4'he):(4'h8)] ?
                          $signed(reg1779) : reg1776[(1'h1):(1'h1)]));
                      reg2290 <= (reg2201 & $unsigned(forvar2119));
                      reg2291 <= reg1990[(4'hd):(3'h7)];
                    end
                  else
                    begin
                      reg2288 <= ((forvar1984 ?
                          {$signed(wire1756)} : forvar1845[(4'ha):(1'h0)]) <= ({reg2108} >= reg2141));
                      reg2289 <= {($unsigned(((8'ha7) <<< forvar1993)) ?
                              forvar2081 : $signed((8'hb3)))};
                      reg2290 <= $unsigned(((8'hb7) ^~ (^~reg1864)));
                      reg2291 <= $signed(reg2180[(3'h7):(3'h4)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar2287 = (1'h0); (forvar2287 < (1'h1)); forvar2287 = (forvar2287 + (1'h1)))
            begin
              for (forvar2288 = (1'h0); (forvar2288 < (2'h2)); forvar2288 = (forvar2288 + (1'h1)))
                begin
                  for (forvar2289 = (1'h0); (forvar2289 < (1'h0)); forvar2289 = (forvar2289 + (1'h1)))
                    begin
                      reg2290 <= ((~|(reg1900 + $signed(reg2017))) && reg1807[(1'h0):(1'h0)]);
                    end
                  for (forvar2291 = (1'h0); (forvar2291 < (1'h1)); forvar2291 = (forvar2291 + (1'h1)))
                    begin
                      reg2292 <= reg1793;
                      reg2293 <= (&$unsigned(({forvar1786} <<< (reg1861 <<< reg2070))));
                      reg2294 <= ((~|(-(forvar2202 ^ reg1772))) << (((forvar1845 ?
                              (8'hae) : reg2147) ?
                          reg2019[(4'he):(3'h4)] : (~(8'h9d))) <<< ($unsigned((8'ha1)) ^ {forvar2117})));
                      reg2295 <= ($unsigned($unsigned((&forvar2170))) ^ ($unsigned(((8'haf) ?
                          forvar1889 : reg1792)) || reg2268[(1'h0):(1'h0)]));
                    end
                  if ({(~(~&(^~reg2041)))})
                    begin
                      reg2296 <= reg2212[(3'h5):(3'h5)];
                      reg2297 <= $unsigned($unsigned(($unsigned(reg2288) ?
                          reg1943 : ((8'hb4) ? (8'hb4) : (8'hae)))));
                      reg2298 <= {{((-(8'hba)) >> (|reg1857))}};
                    end
                  else
                    begin
                      reg2296 <= ((((-(8'haa)) ?
                              $unsigned((8'ha0)) : $unsigned(reg1787)) ?
                          ((~&reg2082) <= {forvar1759}) : ({reg2186} ?
                              {reg1852} : reg2173)) | $unsigned(((reg2083 & reg2281) >>> (+(8'h9c)))));
                      reg2297 <= reg1787[(3'h4):(2'h2)];
                      reg2298 <= reg1891[(3'h4):(2'h2)];
                      reg2299 <= {$signed($unsigned({reg1803}))};
                    end
                end
            end
          for (forvar2300 = (1'h0); (forvar2300 < (2'h2)); forvar2300 = (forvar2300 + (1'h1)))
            begin
              for (forvar2301 = (1'h0); (forvar2301 < (2'h3)); forvar2301 = (forvar2301 + (1'h1)))
                begin
                  for (forvar2302 = (1'h0); (forvar2302 < (2'h2)); forvar2302 = (forvar2302 + (1'h1)))
                    begin
                      reg2303 <= reg2299[(1'h1):(1'h1)];
                      reg2304 <= {$unsigned({reg2059[(4'h9):(3'h7)]})};
                    end
                end
              for (forvar2305 = (1'h0); (forvar2305 < (2'h2)); forvar2305 = (forvar2305 + (1'h1)))
                begin
                  reg2306 <= $unsigned(reg1821[(3'h6):(3'h6)]);
                  if (reg2208)
                    begin
                      reg2307 <= (~^$signed({{reg2046}}));
                      reg2308 <= {(&$unsigned(reg1898))};
                      reg2309 <= (-$signed((forvar1963 ?
                          (reg1876 ?
                              reg2242 : forvar1997) : $unsigned(reg2079))));
                      reg2310 <= reg1821[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2307 <= forvar2268;
                      reg2308 <= (-({(reg1949 ~^ reg2128)} ?
                          $signed(reg2266) : reg1910[(3'h4):(2'h2)]));
                    end
                  reg2311 <= reg1892[(1'h1):(1'h0)];
                  for (forvar2312 = (1'h0); (forvar2312 < (1'h1)); forvar2312 = (forvar2312 + (1'h1)))
                    begin
                      reg2313 <= (($unsigned(reg1917) - forvar2287[(3'h7):(3'h7)]) ?
                          $signed((reg2264 <<< (reg2050 ?
                              reg2280 : reg2164))) : $unsigned(({reg1941} | (8'ha2))));
                      reg2314 <= ((~&reg1894) ?
                          $signed(((forvar2252 ?
                              reg2186 : forvar2175) + (~^reg1763))) : reg2211[(4'h9):(3'h6)]);
                      reg2315 <= reg2065;
                      reg2316 <= $unsigned({forvar1759});
                    end
                end
              for (forvar2317 = (1'h0); (forvar2317 < (2'h2)); forvar2317 = (forvar2317 + (1'h1)))
                begin
                  if (reg2188)
                    begin
                      reg2318 <= $unsigned((reg2240[(1'h1):(1'h1)] ?
                          $signed((forvar1879 ? reg1911 : (8'hae))) : reg2193));
                      reg2319 <= $signed(($unsigned((8'ha7)) * $unsigned($unsigned(reg1952))));
                    end
                  else
                    begin
                      reg2318 <= ((8'hb1) ?
                          reg2307[(4'ha):(3'h5)] : $unsigned(({reg2124} ?
                              reg1859[(1'h1):(1'h0)] : (reg2053 ?
                                  forvar1854 : reg1939))));
                    end
                end
            end
        end
      for (forvar2320 = (1'h0); (forvar2320 < (2'h3)); forvar2320 = (forvar2320 + (1'h1)))
        begin
          for (forvar2321 = (1'h0); (forvar2321 < (1'h1)); forvar2321 = (forvar2321 + (1'h1)))
            begin
              for (forvar2322 = (1'h0); (forvar2322 < (1'h1)); forvar2322 = (forvar2322 + (1'h1)))
                begin
                  if (reg1794)
                    begin
                      reg2323 <= (reg2194 ?
                          ($unsigned($unsigned(reg2135)) << (~^reg2173)) : reg2080[(3'h6):(2'h3)]);
                      reg2324 <= $signed((^~(+reg2207[(2'h2):(1'h0)])));
                      reg2325 <= reg1819[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg2323 <= $unsigned(reg2006[(3'h4):(2'h3)]);
                      reg2324 <= (~&$unsigned($signed((!forvar2288))));
                      reg2325 <= reg2279[(2'h3):(2'h2)];
                      reg2326 <= ((^reg1911) && (wire1753 ?
                          (!(reg2126 ?
                              forvar2111 : reg1868)) : (forvar2241[(2'h2):(1'h0)] ?
                              (reg1899 >> (8'hab)) : (forvar2170 ?
                                  reg2164 : reg2065))));
                    end
                  for (forvar2327 = (1'h0); (forvar2327 < (1'h0)); forvar2327 = (forvar2327 + (1'h1)))
                    begin
                      reg2328 <= (forvar2320 && $unsigned($unsigned($unsigned(reg2194))));
                      reg2329 <= reg1778[(2'h2):(1'h1)];
                      reg2330 <= (forvar2320 >>> reg1972);
                      reg2331 <= reg2039[(1'h1):(1'h1)];
                    end
                  if (($signed($unsigned((reg2033 <= (8'hb9)))) ?
                      ($unsigned((^~reg2304)) ?
                          $signed(forvar2256) : reg1952[(2'h2):(1'h1)]) : ($unsigned(reg1909) + reg1813)))
                    begin
                      reg2332 <= (reg2078 ? (^~{{wire1756}}) : (8'hae));
                    end
                  else
                    begin
                      reg2332 <= (forvar1878 ?
                          $signed($signed($signed(reg2028))) : ({(!reg2022)} ?
                              (reg2135[(4'h8):(3'h4)] << (~reg1967)) : $signed($signed(reg1888))));
                      reg2333 <= ($signed(reg2194) ?
                          $unsigned((^((8'ha0) - reg2289))) : $unsigned($signed({forvar1951})));
                    end
                end
              if (((!(~^(reg2313 + reg1857))) ?
                  $unsigned($unsigned($signed(reg2022))) : {reg2092}))
                begin
                  for (forvar2334 = (1'h0); (forvar2334 < (1'h1)); forvar2334 = (forvar2334 + (1'h1)))
                    begin
                      reg2335 <= ({($unsigned(reg2177) ?
                              (^reg2303) : $unsigned((8'ha3)))} * (~(-$signed(reg2177))));
                      reg2336 <= (8'ha1);
                      reg2337 <= (~|(8'ha1));
                      reg2338 <= reg2241;
                    end
                  for (forvar2339 = (1'h0); (forvar2339 < (2'h2)); forvar2339 = (forvar2339 + (1'h1)))
                    begin
                      reg2340 <= forvar1875;
                      reg2341 <= {reg2225};
                    end
                  for (forvar2342 = (1'h0); (forvar2342 < (2'h3)); forvar2342 = (forvar2342 + (1'h1)))
                    begin
                      reg2343 <= $unsigned($unsigned({(~(8'h9e))}));
                      reg2344 <= $signed({reg2112});
                      reg2345 <= (~$unsigned((8'ha6)));
                      reg2346 <= ((~forvar1891[(2'h2):(1'h0)]) && ((+(forvar2169 ?
                              reg2229 : reg1815)) ?
                          ({forvar2150} != (^~reg2061)) : {$signed(forvar2017)}));
                    end
                  for (forvar2347 = (1'h0); (forvar2347 < (2'h3)); forvar2347 = (forvar2347 + (1'h1)))
                    begin
                      reg2348 <= reg2306;
                      reg2349 <= $signed($unsigned($signed(forvar1920)));
                      reg2350 <= (+({reg2003[(1'h1):(1'h1)]} ?
                          $signed(reg2078) : forvar1994));
                      reg2351 <= $signed(reg2225);
                    end
                end
              else
                begin
                  for (forvar2334 = (1'h0); (forvar2334 < (2'h3)); forvar2334 = (forvar2334 + (1'h1)))
                    begin
                      reg2335 <= ((reg2102 && $unsigned((~&reg2351))) <<< reg1898);
                    end
                  for (forvar2336 = (1'h0); (forvar2336 < (1'h0)); forvar2336 = (forvar2336 + (1'h1)))
                    begin
                      reg2337 <= ($unsigned($signed((reg2323 ?
                          (8'hb1) : reg2049))) | (!($signed(forvar2290) ?
                          {reg2009} : $signed(reg2145))));
                      reg2338 <= reg2138;
                      reg2339 <= (~|{$signed(reg2048[(2'h2):(1'h1)])});
                    end
                  reg2340 <= ($signed((((8'hb8) ? forvar1790 : forvar2113) ?
                          $signed(reg2266) : $signed(reg2017))) ?
                      (8'ha0) : (&($unsigned(reg1981) ? {reg1880} : (8'haa))));
                  for (forvar2341 = (1'h0); (forvar2341 < (2'h2)); forvar2341 = (forvar2341 + (1'h1)))
                    begin
                      reg2342 <= $unsigned(((reg1962 ?
                          (-reg2234) : (forvar2119 * reg2013)) + ((forvar2124 & reg2173) ?
                          ((8'h9e) ?
                              forvar1836 : reg1804) : $unsigned((8'haa)))));
                      reg2343 <= (((8'h9d) == forvar2265[(2'h2):(1'h0)]) ?
                          $unsigned((|reg1921)) : reg2314);
                      reg2344 <= {(-$signed($signed(forvar2255)))};
                      reg2345 <= $unsigned({($signed(reg2033) ?
                              ((8'ha3) == reg1927) : (reg2169 ?
                                  forvar1955 : reg2337))});
                    end
                end
              reg2352 <= reg2102;
              reg2353 <= $signed((^$signed($signed((8'ha6)))));
            end
        end
    end
  assign wire2354 = ((($signed(reg2003) - forvar1923) > {(forvar1905 ?
                                reg2252 : forvar2225)}) ?
                        {((^~reg1947) ?
                                (reg2008 ?
                                    (8'hb8) : reg2132) : (reg1771 == forvar2142))} : (reg2108[(2'h2):(1'h1)] ?
                            $signed((&forvar2301)) : (~^reg1872)));
  assign wire2355 = (~$unsigned(($unsigned(reg1806) ?
                        (reg2132 <<< reg2059) : {reg2037})));
  assign wire2356 = reg1927[(3'h6):(3'h5)];
  assign wire2357 = {$signed($unsigned(forvar2175))};
  assign wire2358 = $unsigned({(forvar2268[(4'h8):(4'h8)] ?
                            reg1771 : ((8'hb9) * reg2135))});
  assign wire2359 = reg1847[(2'h3):(1'h0)];
  assign wire2360 = (+reg1936);
  module2361 modinst3036 (.clk(clk), .wire2365(forvar2014), .wire2363(reg2129), .wire2366(reg2203), .wire2364(reg1928), .y(wire3035), .wire2362(forvar1809));
  assign wire3037 = $unsigned((~(^~reg1804)));
  assign wire3038 = forvar2196[(4'h8):(3'h5)];
  module3039 modinst3530 (.y(wire3529), .clk(clk), .wire3043(reg2258), .wire3041(forvar1809), .wire3044(forvar2030), .wire3040(reg2307), .wire3042(reg1761));
  assign wire3531 = $unsigned(reg2183[(4'h8):(3'h7)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1041
#( parameter param1741 = (^((((8'hb0) ? (8'hab) : (8'ha8)) ? (8'hb6) : ((8'ha1) == (8'hb0))) - (((8'hb9) + (8'hb9)) ? {(8'ha8)} : ((8'hb8) | (8'hb5))))) )
(y, clk, wire1045, wire1044, wire1043, wire1042);
  output wire [(32'h15a8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire1045;
  input wire signed [(5'h10):(1'h0)] wire1044;
  input wire [(3'h5):(1'h0)] wire1043;
  input wire [(4'hd):(1'h0)] wire1042;
  wire signed [(3'h6):(1'h0)] wire1739;
  reg [(4'hf):(1'h0)] reg1531 = (1'h0);
  wire [(3'h5):(1'h0)] wire1530;
  reg [(3'h6):(1'h0)] forvar1510 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1504 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1503 = (1'h0);
  reg [(3'h4):(1'h0)] reg1502 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1529 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1528 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1527 = (1'h0);
  reg [(5'h10):(1'h0)] reg1526 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1525 = (1'h0);
  reg [(4'hc):(1'h0)] reg1524 = (1'h0);
  reg [(4'hc):(1'h0)] reg1523 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1522 = (1'h0);
  reg [(4'he):(1'h0)] reg1521 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1520 = (1'h0);
  reg [(5'h10):(1'h0)] reg1519 = (1'h0);
  reg [(3'h6):(1'h0)] reg1518 = (1'h0);
  reg [(2'h2):(1'h0)] reg1517 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1516 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1515 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1509 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1514 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1513 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1512 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1511 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1510 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1509 = (1'h0);
  reg [(3'h4):(1'h0)] reg1508 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1507 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1506 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1505 = (1'h0);
  reg [(3'h5):(1'h0)] reg1504 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1503 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1502 = (1'h0);
  reg [(4'h9):(1'h0)] reg1501 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1500 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1499 = (1'h0);
  reg [(4'hb):(1'h0)] reg1498 = (1'h0);
  reg [(2'h2):(1'h0)] reg1497 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1495 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1492 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1491 = (1'h0);
  reg [(3'h6):(1'h0)] reg1484 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1482 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1481 = (1'h0);
  reg [(3'h7):(1'h0)] reg1496 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1495 = (1'h0);
  reg [(3'h6):(1'h0)] reg1494 = (1'h0);
  reg [(2'h3):(1'h0)] reg1493 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1492 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1491 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1490 = (1'h0);
  reg [(5'h10):(1'h0)] reg1489 = (1'h0);
  reg [(4'hc):(1'h0)] reg1488 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1487 = (1'h0);
  reg [(3'h7):(1'h0)] reg1486 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1485 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1484 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1479 = (1'h0);
  reg [(5'h10):(1'h0)] reg1483 = (1'h0);
  reg [(4'hd):(1'h0)] reg1482 = (1'h0);
  reg [(3'h5):(1'h0)] reg1481 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1480 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1479 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1478 = (1'h0);
  reg [(3'h7):(1'h0)] reg1477 = (1'h0);
  reg [(2'h3):(1'h0)] reg1476 = (1'h0);
  reg [(4'he):(1'h0)] reg1475 = (1'h0);
  reg [(3'h6):(1'h0)] reg1474 = (1'h0);
  reg [(3'h5):(1'h0)] reg1473 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1472 = (1'h0);
  reg [(4'hd):(1'h0)] reg1471 = (1'h0);
  reg [(4'he):(1'h0)] reg1470 = (1'h0);
  reg [(4'hb):(1'h0)] reg1469 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1468 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1461 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1460 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1457 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1467 = (1'h0);
  reg [(4'h8):(1'h0)] reg1466 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1465 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1464 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1463 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1462 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1461 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1460 = (1'h0);
  reg [(5'h10):(1'h0)] reg1459 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1458 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1457 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1456 = (1'h0);
  reg [(4'hb):(1'h0)] reg1455 = (1'h0);
  reg [(3'h6):(1'h0)] reg1453 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1449 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1448 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1447 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1446 = (1'h0);
  reg [(4'hc):(1'h0)] reg1440 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1439 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1437 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1436 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1429 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1454 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1453 = (1'h0);
  reg [(4'hb):(1'h0)] reg1452 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1451 = (1'h0);
  reg [(4'h8):(1'h0)] reg1450 = (1'h0);
  reg [(5'h10):(1'h0)] reg1449 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1448 = (1'h0);
  reg [(2'h2):(1'h0)] reg1447 = (1'h0);
  reg [(3'h7):(1'h0)] reg1446 = (1'h0);
  reg [(2'h3):(1'h0)] reg1445 = (1'h0);
  reg [(4'hc):(1'h0)] reg1444 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1443 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1442 = (1'h0);
  reg [(4'ha):(1'h0)] reg1441 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1440 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1439 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1438 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1437 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1436 = (1'h0);
  reg [(4'ha):(1'h0)] reg1435 = (1'h0);
  reg [(4'hf):(1'h0)] reg1434 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1433 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1426 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1433 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1432 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1431 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1430 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1429 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1428 = (1'h0);
  reg [(4'hc):(1'h0)] reg1427 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1426 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1425 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1424 = (1'h0);
  wire [(3'h4):(1'h0)] wire1423;
  reg [(3'h7):(1'h0)] reg1415 = (1'h0);
  reg [(4'hc):(1'h0)] reg1412 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1422 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1421 = (1'h0);
  reg [(4'h8):(1'h0)] reg1420 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1419 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1418 = (1'h0);
  reg [(4'he):(1'h0)] reg1417 = (1'h0);
  reg [(4'ha):(1'h0)] reg1416 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1415 = (1'h0);
  reg [(3'h5):(1'h0)] reg1414 = (1'h0);
  reg [(4'hb):(1'h0)] reg1413 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1412 = (1'h0);
  reg [(5'h10):(1'h0)] reg1407 = (1'h0);
  reg [(4'ha):(1'h0)] reg1411 = (1'h0);
  reg [(4'ha):(1'h0)] reg1410 = (1'h0);
  reg [(4'ha):(1'h0)] reg1409 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1407 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1406 = (1'h0);
  reg [(3'h7):(1'h0)] reg1405 = (1'h0);
  reg [(3'h4):(1'h0)] reg1404 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1397 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1396 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1403 = (1'h0);
  reg [(4'hd):(1'h0)] reg1402 = (1'h0);
  reg [(4'hc):(1'h0)] reg1401 = (1'h0);
  reg [(3'h7):(1'h0)] reg1400 = (1'h0);
  reg [(4'hc):(1'h0)] reg1399 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1398 = (1'h0);
  reg [(4'h9):(1'h0)] reg1397 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1396 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1395 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1394 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1393 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1392 = (1'h0);
  reg [(4'hf):(1'h0)] reg1391 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1390 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1389 = (1'h0);
  reg [(4'hd):(1'h0)] reg1388 = (1'h0);
  reg [(4'hd):(1'h0)] reg1387 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1386 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1385 = (1'h0);
  reg [(4'hc):(1'h0)] reg1384 = (1'h0);
  reg [(4'ha):(1'h0)] reg1383 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1382 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1381 = (1'h0);
  reg [(4'hc):(1'h0)] reg1380 = (1'h0);
  reg [(4'hd):(1'h0)] reg1379 = (1'h0);
  reg [(5'h10):(1'h0)] reg1378 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1377 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1376 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1375 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1374 = (1'h0);
  reg [(3'h7):(1'h0)] reg1373 = (1'h0);
  reg [(2'h2):(1'h0)] reg1372 = (1'h0);
  reg [(4'h9):(1'h0)] reg1371 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1370 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1369 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1368 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1367 = (1'h0);
  reg [(3'h5):(1'h0)] reg1340 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1336 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1366 = (1'h0);
  reg [(3'h4):(1'h0)] reg1365 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1364 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1363 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1362 = (1'h0);
  reg [(4'h9):(1'h0)] reg1361 = (1'h0);
  reg [(3'h7):(1'h0)] reg1360 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1359 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1358 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1357 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1356 = (1'h0);
  reg [(3'h6):(1'h0)] reg1355 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1354 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1353 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1352 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1344 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1351 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1350 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1349 = (1'h0);
  reg [(4'hc):(1'h0)] reg1348 = (1'h0);
  reg [(3'h7):(1'h0)] reg1347 = (1'h0);
  reg [(5'h10):(1'h0)] reg1346 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1345 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1344 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1343 = (1'h0);
  reg [(4'hc):(1'h0)] reg1342 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1341 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1340 = (1'h0);
  reg [(5'h10):(1'h0)] reg1335 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1339 = (1'h0);
  reg [(5'h10):(1'h0)] reg1338 = (1'h0);
  reg [(3'h6):(1'h0)] reg1337 = (1'h0);
  reg [(4'hc):(1'h0)] reg1336 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1335 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1334 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1333 = (1'h0);
  reg [(4'hd):(1'h0)] reg1332 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1331 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1330 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1329 = (1'h0);
  reg [(4'hc):(1'h0)] reg1328 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1327 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1326 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1325 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1323 = (1'h0);
  reg [(5'h10):(1'h0)] reg1322 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1324 = (1'h0);
  reg [(4'he):(1'h0)] reg1323 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1322 = (1'h0);
  reg [(2'h3):(1'h0)] reg1321 = (1'h0);
  reg [(4'he):(1'h0)] forvar1320 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1319 = (1'h0);
  reg [(3'h5):(1'h0)] reg1318 = (1'h0);
  reg [(4'hc):(1'h0)] reg1317 = (1'h0);
  reg [(2'h2):(1'h0)] reg1316 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1315 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1314 = (1'h0);
  reg [(4'h9):(1'h0)] reg1313 = (1'h0);
  reg [(4'hf):(1'h0)] reg1312 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1311 = (1'h0);
  reg [(4'hd):(1'h0)] reg1310 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1309 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1296 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1292 = (1'h0);
  reg [(2'h3):(1'h0)] reg1291 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1290 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1287 = (1'h0);
  reg [(3'h5):(1'h0)] reg1288 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1306 = (1'h0);
  reg [(4'hb):(1'h0)] reg1308 = (1'h0);
  reg [(3'h4):(1'h0)] reg1307 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1306 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1305 = (1'h0);
  reg [(4'h9):(1'h0)] reg1304 = (1'h0);
  reg [(4'hd):(1'h0)] reg1303 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1302 = (1'h0);
  reg [(5'h10):(1'h0)] reg1301 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1300 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1299 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1298 = (1'h0);
  reg [(4'h9):(1'h0)] reg1297 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1296 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1295 = (1'h0);
  reg [(3'h7):(1'h0)] reg1294 = (1'h0);
  reg [(3'h7):(1'h0)] reg1293 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1292 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1291 = (1'h0);
  reg [(3'h4):(1'h0)] reg1290 = (1'h0);
  reg [(2'h2):(1'h0)] reg1289 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1288 = (1'h0);
  reg [(4'ha):(1'h0)] reg1287 = (1'h0);
  reg [(4'h9):(1'h0)] reg1269 = (1'h0);
  reg [(4'hc):(1'h0)] reg1286 = (1'h0);
  reg [(2'h2):(1'h0)] reg1285 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1284 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1283 = (1'h0);
  reg [(2'h2):(1'h0)] reg1282 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1280 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1277 = (1'h0);
  reg [(3'h6):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1275 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1273 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1271 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1260 = (1'h0);
  reg [(4'hb):(1'h0)] reg1281 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1264 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1263 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1261 = (1'h0);
  reg [(4'h8):(1'h0)] reg1259 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1280 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1279 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1278 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1277 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1276 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1275 = (1'h0);
  reg [(4'h9):(1'h0)] reg1274 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1266 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1273 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1272 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1271 = (1'h0);
  reg [(2'h3):(1'h0)] reg1270 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1269 = (1'h0);
  reg [(2'h2):(1'h0)] reg1268 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1267 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1266 = (1'h0);
  reg [(5'h10):(1'h0)] reg1265 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1264 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1263 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1262 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1261 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1260 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1259 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1258 = (1'h0);
  reg [(2'h3):(1'h0)] reg1257 = (1'h0);
  reg [(5'h10):(1'h0)] reg1256 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1255 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1254 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1253 = (1'h0);
  reg [(4'he):(1'h0)] reg1250 = (1'h0);
  reg [(5'h10):(1'h0)] reg1248 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1246 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1244 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1235 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1238 = (1'h0);
  reg [(2'h2):(1'h0)] reg1252 = (1'h0);
  reg [(4'he):(1'h0)] reg1251 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1250 = (1'h0);
  reg [(4'hf):(1'h0)] reg1249 = (1'h0);
  reg [(4'he):(1'h0)] forvar1248 = (1'h0);
  reg [(2'h3):(1'h0)] reg1247 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1246 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1245 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1244 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1243 = (1'h0);
  reg [(4'h9):(1'h0)] reg1242 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1241 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1240 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1239 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1238 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1237 = (1'h0);
  reg [(4'hb):(1'h0)] reg1233 = (1'h0);
  reg [(3'h4):(1'h0)] reg1236 = (1'h0);
  reg [(4'h8):(1'h0)] reg1235 = (1'h0);
  reg [(4'ha):(1'h0)] reg1234 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1233 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1232 = (1'h0);
  reg [(4'he):(1'h0)] reg1231 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1230 = (1'h0);
  reg [(4'ha):(1'h0)] reg1229 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1228 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1227 = (1'h0);
  reg [(3'h4):(1'h0)] reg1226 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1225 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1224 = (1'h0);
  reg [(2'h3):(1'h0)] reg1223 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1222 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1221 = (1'h0);
  reg [(3'h6):(1'h0)] reg1220 = (1'h0);
  reg [(3'h4):(1'h0)] reg1219 = (1'h0);
  reg [(2'h3):(1'h0)] reg1218 = (1'h0);
  reg [(4'h8):(1'h0)] reg1217 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1216 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1212 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1204 = (1'h0);
  reg [(3'h6):(1'h0)] reg1203 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1202 = (1'h0);
  reg [(4'hf):(1'h0)] reg1215 = (1'h0);
  reg [(4'h8):(1'h0)] reg1214 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1213 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1211 = (1'h0);
  reg [(4'h8):(1'h0)] reg1208 = (1'h0);
  reg [(4'hd):(1'h0)] reg1212 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1211 = (1'h0);
  reg [(4'hf):(1'h0)] reg1210 = (1'h0);
  reg [(3'h4):(1'h0)] reg1209 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1208 = (1'h0);
  reg [(4'ha):(1'h0)] reg1207 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1206 = (1'h0);
  reg [(4'ha):(1'h0)] reg1205 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1204 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1203 = (1'h0);
  reg [(4'h9):(1'h0)] reg1202 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1188 = (1'h0);
  reg [(4'hf):(1'h0)] reg1201 = (1'h0);
  reg [(5'h10):(1'h0)] reg1200 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1199 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1198 = (1'h0);
  reg [(4'he):(1'h0)] reg1197 = (1'h0);
  reg [(3'h6):(1'h0)] reg1196 = (1'h0);
  reg [(2'h3):(1'h0)] reg1195 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1194 = (1'h0);
  reg [(3'h7):(1'h0)] reg1193 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1192 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1191 = (1'h0);
  reg [(2'h3):(1'h0)] reg1190 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1189 = (1'h0);
  reg [(4'h8):(1'h0)] reg1188 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1187 = (1'h0);
  reg [(4'he):(1'h0)] reg1186 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1183 = (1'h0);
  reg [(2'h2):(1'h0)] reg1185 = (1'h0);
  reg [(3'h5):(1'h0)] reg1184 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1183 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1181 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1177 = (1'h0);
  reg [(4'h9):(1'h0)] reg1175 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1174 = (1'h0);
  reg [(4'hc):(1'h0)] reg1182 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1181 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1180 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1179 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1178 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1177 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1176 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1175 = (1'h0);
  reg [(3'h4):(1'h0)] reg1174 = (1'h0);
  reg [(4'he):(1'h0)] forvar1173 = (1'h0);
  reg [(4'h9):(1'h0)] reg1172 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1165 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1171 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1170 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1169 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1168 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1160 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1156 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1170 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1169 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1168 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1167 = (1'h0);
  reg [(4'hf):(1'h0)] reg1166 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1165 = (1'h0);
  reg [(5'h10):(1'h0)] reg1164 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1163 = (1'h0);
  reg [(4'hb):(1'h0)] reg1159 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1158 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1154 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1162 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1160 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1159 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1158 = (1'h0);
  reg [(3'h4):(1'h0)] reg1155 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1157 = (1'h0);
  reg [(4'h8):(1'h0)] reg1156 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1155 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1154 = (1'h0);
  reg [(4'hb):(1'h0)] reg1153 = (1'h0);
  reg [(4'hf):(1'h0)] reg1152 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1151 = (1'h0);
  reg [(4'hd):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1149 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1148 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1147 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1146 = (1'h0);
  reg [(3'h7):(1'h0)] reg1145 = (1'h0);
  reg [(4'he):(1'h0)] reg1144 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1143 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1142 = (1'h0);
  reg [(4'hf):(1'h0)] reg1141 = (1'h0);
  reg [(5'h10):(1'h0)] reg1140 = (1'h0);
  reg [(4'hf):(1'h0)] reg1130 = (1'h0);
  reg [(2'h3):(1'h0)] reg1129 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1128 = (1'h0);
  reg [(4'h8):(1'h0)] reg1126 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1123 = (1'h0);
  reg [(5'h10):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1120 = (1'h0);
  reg [(4'ha):(1'h0)] reg1119 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1117 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1114 = (1'h0);
  reg [(4'hc):(1'h0)] reg1139 = (1'h0);
  reg [(3'h6):(1'h0)] reg1138 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1137 = (1'h0);
  reg [(4'hd):(1'h0)] reg1136 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1135 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1134 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1133 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1132 = (1'h0);
  reg [(4'hd):(1'h0)] reg1131 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1130 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1129 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1128 = (1'h0);
  reg [(3'h4):(1'h0)] reg1127 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1126 = (1'h0);
  reg [(4'hb):(1'h0)] reg1125 = (1'h0);
  reg [(4'h9):(1'h0)] reg1124 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1123 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1122 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1121 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1120 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1119 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1118 = (1'h0);
  reg [(4'h9):(1'h0)] reg1117 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1116 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1115 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1114 = (1'h0);
  reg [(5'h10):(1'h0)] reg1113 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1112 = (1'h0);
  reg [(4'h9):(1'h0)] reg1111 = (1'h0);
  reg [(4'he):(1'h0)] reg1110 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1109 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1108 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1107 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1106 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1105 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1104 = (1'h0);
  reg [(4'ha):(1'h0)] reg1103 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1102 = (1'h0);
  reg [(4'hd):(1'h0)] reg1101 = (1'h0);
  reg [(4'hc):(1'h0)] reg1100 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1099 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1098 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1097 = (1'h0);
  reg [(4'hb):(1'h0)] reg1096 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1095 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1094 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1085 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1083 = (1'h0);
  reg [(4'he):(1'h0)] reg1093 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1092 = (1'h0);
  reg [(2'h3):(1'h0)] reg1091 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1090 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1089 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1088 = (1'h0);
  reg [(4'he):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1086 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1085 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1084 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1083 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1082 = (1'h0);
  reg [(4'ha):(1'h0)] reg1081 = (1'h0);
  reg [(5'h10):(1'h0)] reg1080 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1079 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1078 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1077 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1076 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1075 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1074 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1065 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1061 = (1'h0);
  reg [(4'hc):(1'h0)] reg1073 = (1'h0);
  reg [(4'h9):(1'h0)] reg1072 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1071 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1070 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1069 = (1'h0);
  reg [(4'hc):(1'h0)] reg1068 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1067 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1066 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1065 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1064 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1063 = (1'h0);
  reg [(4'h8):(1'h0)] reg1062 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1061 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1060 = (1'h0);
  reg [(4'h9):(1'h0)] reg1059 = (1'h0);
  reg [(5'h10):(1'h0)] reg1058 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1057 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1056 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1055 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1054 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1053 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1052 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1051 = (1'h0);
  reg [(4'he):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1049 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1048 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1047 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire1046;
  assign y = {wire1739,
                 reg1531,
                 wire1530,
                 forvar1510,
                 forvar1504,
                 reg1503,
                 reg1502,
                 reg1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 forvar1525,
                 reg1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 forvar1520,
                 reg1519,
                 reg1518,
                 reg1517,
                 forvar1516,
                 forvar1515,
                 forvar1509,
                 reg1514,
                 reg1513,
                 reg1512,
                 reg1511,
                 reg1510,
                 reg1509,
                 reg1508,
                 reg1507,
                 reg1506,
                 reg1505,
                 reg1504,
                 forvar1503,
                 forvar1502,
                 reg1501,
                 reg1500,
                 forvar1499,
                 reg1498,
                 reg1497,
                 reg1495,
                 forvar1492,
                 reg1491,
                 reg1484,
                 forvar1482,
                 forvar1481,
                 reg1496,
                 forvar1495,
                 reg1494,
                 reg1493,
                 reg1492,
                 forvar1491,
                 reg1490,
                 reg1489,
                 reg1488,
                 reg1487,
                 reg1486,
                 reg1485,
                 forvar1484,
                 reg1479,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1480,
                 forvar1479,
                 forvar1478,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1471,
                 reg1470,
                 reg1469,
                 forvar1468,
                 reg1461,
                 forvar1460,
                 reg1457,
                 reg1467,
                 reg1466,
                 forvar1465,
                 reg1464,
                 reg1463,
                 reg1462,
                 forvar1461,
                 reg1460,
                 reg1459,
                 reg1458,
                 forvar1457,
                 forvar1456,
                 reg1455,
                 reg1453,
                 forvar1449,
                 reg1448,
                 forvar1447,
                 forvar1446,
                 reg1440,
                 reg1439,
                 forvar1437,
                 forvar1436,
                 forvar1429,
                 reg1454,
                 forvar1453,
                 reg1452,
                 reg1451,
                 reg1450,
                 reg1449,
                 forvar1448,
                 reg1447,
                 reg1446,
                 reg1445,
                 reg1444,
                 forvar1443,
                 reg1442,
                 reg1441,
                 forvar1440,
                 forvar1439,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1434,
                 forvar1433,
                 reg1426,
                 reg1433,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 forvar1426,
                 forvar1425,
                 reg1424,
                 wire1423,
                 reg1415,
                 reg1412,
                 reg1422,
                 forvar1421,
                 reg1420,
                 forvar1419,
                 reg1418,
                 reg1417,
                 reg1416,
                 forvar1415,
                 reg1414,
                 reg1413,
                 forvar1412,
                 reg1407,
                 reg1411,
                 reg1410,
                 reg1409,
                 reg1408,
                 forvar1407,
                 reg1406,
                 reg1405,
                 reg1404,
                 forvar1397,
                 reg1396,
                 reg1403,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1399,
                 reg1398,
                 reg1397,
                 forvar1396,
                 forvar1395,
                 reg1394,
                 reg1393,
                 forvar1392,
                 reg1391,
                 forvar1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 forvar1386,
                 forvar1385,
                 reg1384,
                 reg1383,
                 reg1382,
                 reg1381,
                 reg1380,
                 reg1379,
                 reg1378,
                 reg1377,
                 reg1376,
                 forvar1375,
                 reg1374,
                 reg1373,
                 reg1372,
                 reg1371,
                 forvar1370,
                 forvar1369,
                 forvar1368,
                 forvar1367,
                 reg1340,
                 forvar1336,
                 reg1366,
                 reg1365,
                 reg1364,
                 reg1363,
                 forvar1362,
                 reg1361,
                 reg1360,
                 forvar1359,
                 reg1358,
                 reg1357,
                 forvar1356,
                 reg1355,
                 reg1354,
                 forvar1353,
                 reg1352,
                 reg1344,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 reg1347,
                 reg1346,
                 reg1345,
                 forvar1344,
                 reg1343,
                 reg1342,
                 reg1341,
                 forvar1340,
                 reg1335,
                 reg1339,
                 reg1338,
                 reg1337,
                 reg1336,
                 forvar1335,
                 forvar1334,
                 reg1333,
                 reg1332,
                 reg1331,
                 reg1330,
                 forvar1329,
                 reg1328,
                 forvar1327,
                 reg1326,
                 reg1325,
                 forvar1323,
                 reg1322,
                 reg1324,
                 reg1323,
                 forvar1322,
                 reg1321,
                 forvar1320,
                 forvar1319,
                 reg1318,
                 reg1317,
                 reg1316,
                 forvar1315,
                 reg1314,
                 reg1313,
                 reg1312,
                 reg1311,
                 reg1310,
                 forvar1309,
                 reg1296,
                 reg1292,
                 reg1291,
                 forvar1290,
                 forvar1287,
                 reg1288,
                 reg1306,
                 reg1308,
                 reg1307,
                 forvar1306,
                 reg1305,
                 reg1304,
                 reg1303,
                 reg1302,
                 reg1301,
                 reg1300,
                 reg1299,
                 reg1298,
                 reg1297,
                 forvar1296,
                 reg1295,
                 reg1294,
                 reg1293,
                 forvar1292,
                 forvar1291,
                 reg1290,
                 reg1289,
                 forvar1288,
                 reg1287,
                 reg1269,
                 reg1286,
                 reg1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 forvar1280,
                 forvar1277,
                 reg1276,
                 reg1275,
                 forvar1273,
                 forvar1271,
                 reg1260,
                 reg1281,
                 reg1264,
                 forvar1263,
                 forvar1261,
                 reg1259,
                 reg1280,
                 reg1279,
                 reg1278,
                 reg1277,
                 forvar1276,
                 forvar1275,
                 reg1274,
                 reg1266,
                 reg1273,
                 reg1272,
                 reg1271,
                 reg1270,
                 forvar1269,
                 reg1268,
                 reg1267,
                 forvar1266,
                 reg1265,
                 forvar1264,
                 reg1263,
                 reg1262,
                 reg1261,
                 forvar1260,
                 forvar1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 reg1255,
                 forvar1254,
                 reg1253,
                 reg1250,
                 reg1248,
                 reg1246,
                 forvar1244,
                 forvar1235,
                 forvar1238,
                 reg1252,
                 reg1251,
                 forvar1250,
                 reg1249,
                 forvar1248,
                 reg1247,
                 forvar1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 reg1241,
                 reg1240,
                 reg1239,
                 reg1238,
                 reg1237,
                 reg1233,
                 reg1236,
                 reg1235,
                 reg1234,
                 forvar1233,
                 reg1232,
                 reg1231,
                 reg1230,
                 reg1229,
                 forvar1228,
                 reg1227,
                 reg1226,
                 reg1225,
                 forvar1224,
                 reg1223,
                 reg1222,
                 forvar1221,
                 reg1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 forvar1216,
                 forvar1212,
                 reg1204,
                 reg1203,
                 forvar1202,
                 reg1215,
                 reg1214,
                 reg1213,
                 forvar1211,
                 reg1208,
                 reg1212,
                 reg1211,
                 reg1210,
                 reg1209,
                 forvar1208,
                 reg1207,
                 forvar1206,
                 reg1205,
                 forvar1204,
                 forvar1203,
                 reg1202,
                 forvar1188,
                 reg1201,
                 reg1200,
                 reg1199,
                 reg1198,
                 reg1197,
                 reg1196,
                 reg1195,
                 reg1194,
                 reg1193,
                 reg1192,
                 reg1191,
                 reg1190,
                 reg1189,
                 reg1188,
                 reg1187,
                 reg1186,
                 forvar1183,
                 reg1185,
                 reg1184,
                 reg1183,
                 forvar1181,
                 forvar1177,
                 reg1175,
                 forvar1174,
                 reg1182,
                 reg1181,
                 reg1180,
                 reg1179,
                 reg1178,
                 reg1177,
                 reg1176,
                 forvar1175,
                 reg1174,
                 forvar1173,
                 reg1172,
                 forvar1165,
                 reg1171,
                 forvar1170,
                 reg1169,
                 reg1168,
                 forvar1160,
                 forvar1156,
                 reg1170,
                 forvar1169,
                 forvar1168,
                 reg1167,
                 reg1166,
                 reg1165,
                 reg1164,
                 forvar1163,
                 reg1159,
                 forvar1158,
                 reg1154,
                 reg1162,
                 reg1161,
                 reg1160,
                 forvar1159,
                 reg1158,
                 reg1155,
                 reg1157,
                 reg1156,
                 forvar1155,
                 forvar1154,
                 reg1153,
                 reg1152,
                 forvar1151,
                 reg1150,
                 reg1149,
                 reg1148,
                 forvar1147,
                 forvar1146,
                 reg1145,
                 reg1144,
                 reg1143,
                 forvar1142,
                 reg1141,
                 reg1140,
                 reg1130,
                 reg1129,
                 forvar1128,
                 reg1126,
                 reg1123,
                 reg1109,
                 reg1120,
                 reg1119,
                 forvar1117,
                 reg1114,
                 reg1139,
                 reg1138,
                 forvar1137,
                 reg1136,
                 reg1135,
                 reg1134,
                 reg1133,
                 reg1132,
                 reg1131,
                 forvar1130,
                 forvar1129,
                 reg1128,
                 reg1127,
                 forvar1126,
                 reg1125,
                 reg1124,
                 forvar1123,
                 reg1122,
                 reg1121,
                 forvar1120,
                 forvar1119,
                 reg1118,
                 reg1117,
                 reg1116,
                 reg1115,
                 forvar1114,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1110,
                 forvar1109,
                 reg1108,
                 reg1107,
                 forvar1106,
                 reg1105,
                 reg1104,
                 reg1103,
                 forvar1102,
                 reg1101,
                 reg1100,
                 reg1099,
                 forvar1098,
                 reg1097,
                 reg1096,
                 forvar1095,
                 forvar1094,
                 forvar1085,
                 reg1083,
                 reg1093,
                 reg1092,
                 reg1091,
                 reg1090,
                 reg1089,
                 forvar1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 reg1084,
                 forvar1083,
                 reg1082,
                 reg1081,
                 reg1080,
                 forvar1079,
                 reg1078,
                 forvar1077,
                 reg1076,
                 forvar1075,
                 forvar1074,
                 reg1065,
                 reg1061,
                 reg1073,
                 reg1072,
                 reg1071,
                 reg1070,
                 reg1069,
                 reg1068,
                 reg1067,
                 reg1066,
                 forvar1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 forvar1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1057,
                 reg1056,
                 reg1055,
                 forvar1054,
                 reg1053,
                 reg1052,
                 reg1051,
                 reg1050,
                 forvar1049,
                 forvar1048,
                 forvar1047,
                 wire1046,
                 (1'h0)};
  assign wire1046 = (8'hb3);
  always
    @(posedge clk) begin
      for (forvar1047 = (1'h0); (forvar1047 < (1'h1)); forvar1047 = (forvar1047 + (1'h1)))
        begin
          for (forvar1048 = (1'h0); (forvar1048 < (1'h1)); forvar1048 = (forvar1048 + (1'h1)))
            begin
              for (forvar1049 = (1'h0); (forvar1049 < (2'h3)); forvar1049 = (forvar1049 + (1'h1)))
                begin
                  if ((|forvar1047[(3'h4):(3'h4)]))
                    begin
                      reg1050 <= ((forvar1047[(3'h5):(3'h4)] != (!$signed(forvar1047))) & forvar1049);
                    end
                  else
                    begin
                      reg1050 <= ($unsigned(reg1050[(4'he):(4'ha)]) && {forvar1049[(3'h4):(1'h0)]});
                      reg1051 <= $signed($unsigned(((^forvar1049) ?
                          reg1050[(2'h3):(1'h0)] : (~&forvar1049))));
                    end
                  if ($unsigned(wire1046[(4'hc):(3'h6)]))
                    begin
                      reg1052 <= (wire1042 <<< reg1050);
                    end
                  else
                    begin
                      reg1052 <= (((((8'haa) ? wire1045 : reg1051) ?
                              reg1050[(4'hd):(3'h4)] : (wire1043 | wire1045)) ?
                          reg1051[(5'h10):(3'h7)] : wire1043) && wire1044);
                      reg1053 <= ((^~wire1046[(1'h0):(1'h0)]) <= (^~{(^~wire1044)}));
                    end
                  for (forvar1054 = (1'h0); (forvar1054 < (2'h2)); forvar1054 = (forvar1054 + (1'h1)))
                    begin
                      reg1055 <= ((+$signed($unsigned(forvar1047))) ?
                          wire1046 : (reg1050 > {$signed(reg1052)}));
                      reg1056 <= ($unsigned(({wire1044} > {wire1044})) == $signed(($unsigned(wire1043) >>> wire1042[(3'h5):(3'h4)])));
                    end
                  if (reg1050[(4'hd):(3'h5)])
                    begin
                      reg1057 <= $unsigned($signed(wire1044));
                      reg1058 <= (~^(8'h9e));
                      reg1059 <= wire1044[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg1057 <= (^(((^~(8'hb8)) != reg1056) == ($unsigned(reg1053) & (8'ha3))));
                    end
                end
              if ((forvar1049[(2'h2):(1'h0)] - (reg1053 | wire1043)))
                begin
                  reg1060 <= $unsigned(forvar1049);
                  for (forvar1061 = (1'h0); (forvar1061 < (2'h2)); forvar1061 = (forvar1061 + (1'h1)))
                    begin
                      reg1062 <= (8'hb7);
                      reg1063 <= $unsigned((wire1043 ?
                          forvar1061[(4'h8):(2'h2)] : ($signed(reg1051) <<< (reg1059 ?
                              (8'hb5) : reg1050))));
                      reg1064 <= ((~^$signed(forvar1054)) ?
                          (~^wire1044) : (($signed(reg1058) <<< $unsigned(wire1042)) ?
                              reg1059 : reg1062[(2'h2):(1'h0)]));
                    end
                  for (forvar1065 = (1'h0); (forvar1065 < (2'h2)); forvar1065 = (forvar1065 + (1'h1)))
                    begin
                      reg1066 <= (forvar1048[(4'h8):(1'h0)] && (reg1064 ~^ reg1050));
                      reg1067 <= reg1064;
                      reg1068 <= $unsigned(reg1053[(4'h8):(2'h3)]);
                      reg1069 <= (reg1068[(2'h3):(1'h0)] ^ (reg1057[(3'h5):(1'h1)] ?
                          $signed(reg1066[(1'h1):(1'h1)]) : {reg1055}));
                    end
                  if ($unsigned($signed($signed($unsigned(wire1045)))))
                    begin
                      reg1070 <= reg1057[(3'h7):(1'h1)];
                      reg1071 <= wire1042[(4'ha):(1'h1)];
                      reg1072 <= $unsigned(reg1053);
                      reg1073 <= ((~&reg1058[(3'h6):(1'h0)]) != ($unsigned(((8'hb2) ?
                          (8'hb8) : forvar1047)) ^ ((reg1050 ?
                          reg1067 : reg1068) ^ wire1045[(2'h2):(2'h2)])));
                    end
                  else
                    begin
                      reg1070 <= $signed((~|$signed((-wire1045))));
                      reg1071 <= $unsigned((reg1050 ?
                          {{reg1072}} : $unsigned($signed(reg1060))));
                      reg1072 <= $signed(($unsigned(reg1060[(1'h0):(1'h0)]) ?
                          reg1073 : reg1069));
                    end
                end
              else
                begin
                  if ((~&($signed((~forvar1054)) ?
                      (!(-forvar1065)) : (^(reg1062 >> (8'haf))))))
                    begin
                      reg1060 <= (reg1073 >>> (forvar1054 + wire1046[(4'hb):(3'h6)]));
                    end
                  else
                    begin
                      reg1060 <= (~$signed(reg1053));
                      reg1061 <= (-reg1051);
                    end
                  if (reg1073[(1'h1):(1'h1)])
                    begin
                      reg1062 <= reg1069[(3'h5):(1'h0)];
                      reg1063 <= {wire1046[(4'h8):(1'h1)]};
                      reg1064 <= {$signed({(^~(8'hba))})};
                      reg1065 <= $signed((&(&forvar1065[(3'h6):(1'h0)])));
                    end
                  else
                    begin
                      reg1062 <= ((8'hb6) <<< $unsigned((&(forvar1048 < (8'ha9)))));
                      reg1063 <= ((forvar1065[(2'h3):(2'h2)] <= $unsigned((reg1060 ?
                              reg1065 : (8'ha1)))) ?
                          (^~(~&(wire1043 ~^ wire1045))) : reg1072);
                      reg1064 <= $unsigned((8'hb4));
                      reg1065 <= (8'h9f);
                    end
                  if (reg1057)
                    begin
                      reg1066 <= (|$signed(reg1051));
                    end
                  else
                    begin
                      reg1066 <= forvar1065;
                      reg1067 <= ({$signed(forvar1048[(1'h1):(1'h1)])} < (+$signed(reg1063[(3'h7):(3'h4)])));
                      reg1068 <= $unsigned($signed($unsigned((~wire1043))));
                      reg1069 <= reg1073;
                    end
                end
              for (forvar1074 = (1'h0); (forvar1074 < (1'h0)); forvar1074 = (forvar1074 + (1'h1)))
                begin
                  for (forvar1075 = (1'h0); (forvar1075 < (2'h3)); forvar1075 = (forvar1075 + (1'h1)))
                    begin
                      reg1076 <= (((^$unsigned(reg1070)) < $unsigned(reg1060[(1'h0):(1'h0)])) ?
                          (!$unsigned(wire1046[(4'he):(2'h2)])) : (^~(-((8'had) ?
                              reg1062 : reg1070))));
                    end
                end
              for (forvar1077 = (1'h0); (forvar1077 < (2'h3)); forvar1077 = (forvar1077 + (1'h1)))
                begin
                  reg1078 <= (-reg1050[(4'he):(4'hd)]);
                  for (forvar1079 = (1'h0); (forvar1079 < (2'h2)); forvar1079 = (forvar1079 + (1'h1)))
                    begin
                      reg1080 <= (+(reg1078[(4'ha):(2'h3)] ?
                          {$unsigned(reg1050)} : reg1064));
                      reg1081 <= (forvar1048[(4'h8):(1'h0)] >= {{reg1059}});
                    end
                end
            end
          if (($signed(reg1061[(4'hb):(2'h2)]) | (((~reg1050) ^~ reg1055) ?
              $signed(reg1073) : ((^reg1070) ?
                  $signed(reg1078) : (forvar1048 << wire1044)))))
            begin
              reg1082 <= (~|reg1064[(1'h0):(1'h0)]);
              for (forvar1083 = (1'h0); (forvar1083 < (2'h3)); forvar1083 = (forvar1083 + (1'h1)))
                begin
                  if (((8'ha8) == (reg1082 * {forvar1065[(3'h5):(3'h5)]})))
                    begin
                      reg1084 <= wire1046[(4'hb):(2'h2)];
                      reg1085 <= ($unsigned(reg1052[(2'h3):(2'h2)]) ?
                          {(~|reg1081)} : (^{{wire1045}}));
                      reg1086 <= $signed(($unsigned((!reg1064)) ^ ((forvar1048 ?
                          (8'ha3) : forvar1047) ^ forvar1054[(1'h0):(1'h0)])));
                      reg1087 <= reg1082;
                    end
                  else
                    begin
                      reg1084 <= {$signed(reg1072)};
                      reg1085 <= forvar1049;
                      reg1086 <= forvar1065;
                      reg1087 <= (reg1062 ?
                          $signed($signed(wire1042)) : reg1059[(3'h4):(1'h1)]);
                    end
                  for (forvar1088 = (1'h0); (forvar1088 < (1'h0)); forvar1088 = (forvar1088 + (1'h1)))
                    begin
                      reg1089 <= $signed(reg1078[(1'h0):(1'h0)]);
                      reg1090 <= (((8'h9f) ^ {(^~reg1060)}) <<< $unsigned({(|reg1071)}));
                      reg1091 <= (reg1061[(1'h0):(1'h0)] ?
                          (^reg1070[(4'hc):(1'h0)]) : $unsigned(reg1082[(2'h3):(1'h1)]));
                      reg1092 <= ($unsigned(((^~(8'ha1)) ~^ reg1069)) ?
                          (reg1090[(2'h2):(1'h1)] ?
                              reg1052[(1'h1):(1'h0)] : (8'h9f)) : (~|((8'had) | $unsigned((8'h9d)))));
                    end
                end
            end
          else
            begin
              reg1082 <= (~forvar1079);
              if ((reg1078[(3'h7):(3'h7)] ^ $unsigned((((8'hb5) ?
                  reg1058 : reg1081) <<< (forvar1079 ? reg1084 : reg1055)))))
                begin
                  for (forvar1083 = (1'h0); (forvar1083 < (2'h2)); forvar1083 = (forvar1083 + (1'h1)))
                    begin
                      reg1084 <= $signed(reg1065[(3'h4):(1'h1)]);
                      reg1085 <= reg1069;
                      reg1086 <= reg1084[(2'h2):(2'h2)];
                      reg1087 <= (8'ha4);
                    end
                  for (forvar1088 = (1'h0); (forvar1088 < (2'h3)); forvar1088 = (forvar1088 + (1'h1)))
                    begin
                      reg1089 <= $unsigned((^~$unsigned((!forvar1065))));
                      reg1090 <= $unsigned((&($signed(forvar1065) ?
                          reg1057[(4'h8):(3'h5)] : ((8'ha0) ?
                              reg1059 : forvar1088))));
                      reg1091 <= $signed($unsigned(((~&reg1051) < $unsigned((8'ha0)))));
                      reg1092 <= (reg1080 ?
                          {wire1043} : $unsigned({{forvar1065}}));
                    end
                  reg1093 <= forvar1049[(3'h4):(2'h3)];
                end
              else
                begin
                  reg1083 <= $unsigned({(~$unsigned(reg1060))});
                  if (wire1046[(4'ha):(3'h6)])
                    begin
                      reg1084 <= reg1069[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1084 <= reg1064[(4'h8):(3'h6)];
                    end
                  for (forvar1085 = (1'h0); (forvar1085 < (1'h0)); forvar1085 = (forvar1085 + (1'h1)))
                    begin
                      reg1086 <= (reg1078 ?
                          (~reg1060) : (((8'hb4) ?
                                  (~&(8'had)) : ((8'hae) <= reg1052)) ?
                              $signed(reg1091[(2'h3):(2'h3)]) : $unsigned((8'hb5))));
                    end
                end
              for (forvar1094 = (1'h0); (forvar1094 < (1'h0)); forvar1094 = (forvar1094 + (1'h1)))
                begin
                  for (forvar1095 = (1'h0); (forvar1095 < (2'h3)); forvar1095 = (forvar1095 + (1'h1)))
                    begin
                      reg1096 <= $unsigned($signed((^reg1050)));
                      reg1097 <= (~|{((~^reg1065) ? (-reg1056) : (^(8'h9f)))});
                    end
                  for (forvar1098 = (1'h0); (forvar1098 < (1'h1)); forvar1098 = (forvar1098 + (1'h1)))
                    begin
                      reg1099 <= ({((8'hb2) ?
                              $signed(reg1078) : (reg1081 ?
                                  wire1043 : reg1081))} ^ reg1056);
                      reg1100 <= reg1065[(3'h4):(1'h0)];
                      reg1101 <= reg1082;
                    end
                  for (forvar1102 = (1'h0); (forvar1102 < (1'h0)); forvar1102 = (forvar1102 + (1'h1)))
                    begin
                      reg1103 <= $unsigned($signed(((!reg1081) ?
                          (~|forvar1075) : (-(8'hae)))));
                      reg1104 <= $unsigned((~&$unsigned($unsigned(forvar1094))));
                      reg1105 <= reg1050[(4'h8):(3'h5)];
                    end
                  for (forvar1106 = (1'h0); (forvar1106 < (1'h0)); forvar1106 = (forvar1106 + (1'h1)))
                    begin
                      reg1107 <= $unsigned(($signed((reg1103 << (8'hb2))) && forvar1079[(1'h1):(1'h1)]));
                      reg1108 <= reg1103;
                    end
                end
            end
        end
      if ({$unsigned($signed(reg1056))})
        begin
          if (reg1096)
            begin
              for (forvar1109 = (1'h0); (forvar1109 < (1'h0)); forvar1109 = (forvar1109 + (1'h1)))
                begin
                  reg1110 <= reg1090;
                  if (wire1046)
                    begin
                      reg1111 <= (-($unsigned(forvar1102[(2'h2):(1'h0)]) >= reg1080[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg1111 <= ($unsigned(forvar1083[(1'h0):(1'h0)]) ?
                          (+((forvar1048 ^~ reg1053) <<< {(8'haa)})) : reg1086);
                      reg1112 <= ((reg1111[(4'h9):(3'h5)] >= reg1111[(2'h2):(1'h0)]) ?
                          $unsigned({(reg1058 <= (8'hb8))}) : ((~^reg1083) ?
                              $signed(reg1100) : {reg1090}));
                    end
                  reg1113 <= (~|$unsigned(reg1071[(1'h0):(1'h0)]));
                  for (forvar1114 = (1'h0); (forvar1114 < (2'h2)); forvar1114 = (forvar1114 + (1'h1)))
                    begin
                      reg1115 <= $unsigned((reg1061 | reg1062));
                      reg1116 <= $unsigned(reg1058[(4'h8):(4'h8)]);
                      reg1117 <= forvar1074[(1'h1):(1'h1)];
                      reg1118 <= ($signed(((~&reg1083) - (forvar1047 ?
                              wire1044 : (8'ha3)))) ?
                          $signed(reg1097) : {reg1064[(2'h3):(2'h2)]});
                    end
                end
              for (forvar1119 = (1'h0); (forvar1119 < (2'h2)); forvar1119 = (forvar1119 + (1'h1)))
                begin
                  for (forvar1120 = (1'h0); (forvar1120 < (2'h3)); forvar1120 = (forvar1120 + (1'h1)))
                    begin
                      reg1121 <= ((reg1087[(4'hc):(1'h1)] | {(8'ha9)}) ~^ $unsigned((8'h9d)));
                      reg1122 <= reg1113;
                    end
                  for (forvar1123 = (1'h0); (forvar1123 < (1'h0)); forvar1123 = (forvar1123 + (1'h1)))
                    begin
                      reg1124 <= (-(((^~(8'ha6)) == (reg1096 ?
                          reg1117 : reg1084)) | forvar1109[(1'h1):(1'h0)]));
                    end
                  if ((8'ha6))
                    begin
                      reg1125 <= $unsigned(($signed($signed(reg1061)) * {(reg1110 ?
                              reg1064 : reg1082)}));
                    end
                  else
                    begin
                      reg1125 <= {reg1085};
                    end
                  for (forvar1126 = (1'h0); (forvar1126 < (2'h3)); forvar1126 = (forvar1126 + (1'h1)))
                    begin
                      reg1127 <= {reg1051};
                      reg1128 <= (!forvar1123[(3'h7):(2'h3)]);
                    end
                end
              for (forvar1129 = (1'h0); (forvar1129 < (2'h2)); forvar1129 = (forvar1129 + (1'h1)))
                begin
                  for (forvar1130 = (1'h0); (forvar1130 < (2'h3)); forvar1130 = (forvar1130 + (1'h1)))
                    begin
                      reg1131 <= ((~^(reg1111[(2'h2):(2'h2)] ?
                              {reg1066} : $unsigned(reg1115))) ?
                          (reg1053 ?
                              reg1087 : ($signed((8'ha1)) ?
                                  $unsigned((8'hb5)) : (reg1056 ^ (8'hb7)))) : (forvar1114[(1'h0):(1'h0)] ?
                              reg1096 : reg1058[(4'ha):(3'h5)]));
                      reg1132 <= $signed(reg1103[(3'h4):(2'h3)]);
                      reg1133 <= (reg1068[(4'h8):(3'h4)] ?
                          reg1104 : $signed($signed((~|reg1090))));
                      reg1134 <= (8'hb2);
                    end
                  if ({(~&reg1082[(2'h2):(1'h1)])})
                    begin
                      reg1135 <= $unsigned($signed((~&reg1100[(3'h4):(1'h1)])));
                      reg1136 <= (((^(&reg1068)) ?
                          reg1117[(3'h6):(1'h1)] : $signed(forvar1098[(1'h0):(1'h0)])) + ((wire1044[(3'h5):(1'h0)] ~^ $unsigned(reg1110)) > (-reg1113[(4'hc):(4'h9)])));
                    end
                  else
                    begin
                      reg1135 <= (forvar1129[(1'h1):(1'h1)] - {reg1050});
                      reg1136 <= reg1073[(2'h3):(2'h3)];
                    end
                  for (forvar1137 = (1'h0); (forvar1137 < (1'h1)); forvar1137 = (forvar1137 + (1'h1)))
                    begin
                      reg1138 <= forvar1102;
                    end
                  reg1139 <= ($unsigned(((forvar1061 >>> reg1068) >>> $unsigned(reg1116))) > reg1108[(2'h3):(1'h0)]);
                end
            end
          else
            begin
              if (reg1091)
                begin
                  for (forvar1109 = (1'h0); (forvar1109 < (2'h2)); forvar1109 = (forvar1109 + (1'h1)))
                    begin
                      reg1110 <= forvar1098[(2'h2):(2'h2)];
                      reg1111 <= reg1125;
                      reg1112 <= $signed($signed($signed(forvar1119[(4'h9):(3'h7)])));
                      reg1113 <= ((reg1059[(2'h3):(1'h0)] ~^ (-(^(8'hac)))) ?
                          {(8'ha6)} : $unsigned(forvar1047[(2'h2):(1'h0)]));
                    end
                  if ((-reg1100))
                    begin
                      reg1114 <= ($unsigned($unsigned(reg1050[(3'h5):(1'h0)])) ?
                          (reg1059 || reg1101[(2'h3):(2'h2)]) : (8'hb2));
                      reg1115 <= (~reg1136);
                      reg1116 <= reg1100[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1114 <= (forvar1061[(3'h6):(2'h3)] >> reg1097[(4'he):(3'h5)]);
                    end
                  for (forvar1117 = (1'h0); (forvar1117 < (1'h1)); forvar1117 = (forvar1117 + (1'h1)))
                    begin
                      reg1118 <= reg1112;
                    end
                  if (forvar1049[(3'h4):(2'h2)])
                    begin
                      reg1119 <= $signed($unsigned((&(~&(8'hb5)))));
                    end
                  else
                    begin
                      reg1119 <= $unsigned(reg1066);
                      reg1120 <= ($signed(wire1042) >>> ($unsigned((forvar1088 * reg1058)) ?
                          $signed($unsigned(reg1097)) : ((reg1112 ~^ wire1043) >> wire1042[(2'h2):(1'h0)])));
                      reg1121 <= reg1103[(3'h5):(3'h4)];
                    end
                end
              else
                begin
                  if ($unsigned((((~reg1125) * (reg1132 ?
                      forvar1137 : reg1113)) > $signed((forvar1095 ?
                      (8'ha1) : reg1052)))))
                    begin
                      reg1109 <= $unsigned((~&($unsigned(reg1136) ?
                          (8'hb3) : (reg1052 <<< forvar1065))));
                      reg1110 <= reg1091;
                      reg1111 <= {forvar1079};
                      reg1112 <= (-$unsigned($unsigned((^~(8'hab)))));
                    end
                  else
                    begin
                      reg1109 <= {$unsigned(reg1103[(3'h4):(2'h2)])};
                      reg1110 <= forvar1098[(2'h2):(1'h1)];
                      reg1111 <= reg1081[(3'h6):(1'h0)];
                    end
                end
              reg1122 <= reg1060[(1'h0):(1'h0)];
              if ($signed(reg1109[(4'hb):(4'hb)]))
                begin
                  if ($unsigned($signed(forvar1130)))
                    begin
                      reg1123 <= {reg1083};
                      reg1124 <= (forvar1117 ~^ (reg1065 ?
                          $unsigned((^reg1063)) : ({forvar1065} << (reg1092 + reg1053))));
                      reg1125 <= (8'hac);
                      reg1126 <= (($unsigned((|(8'h9d))) * $signed((reg1070 != reg1061))) | reg1076[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg1123 <= reg1076;
                      reg1124 <= (((forvar1085 ?
                          (8'hb5) : reg1051[(5'h10):(5'h10)]) > $signed(reg1093)) == reg1108[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  reg1123 <= reg1119[(4'h9):(3'h5)];
                  if (reg1113)
                    begin
                      reg1124 <= ((!(+$signed(forvar1098))) != reg1107);
                      reg1125 <= (!($unsigned(forvar1061) ?
                          reg1073[(1'h1):(1'h0)] : {$unsigned((8'hb2))}));
                      reg1126 <= (~&(((reg1084 ~^ forvar1129) ?
                              (^~reg1124) : reg1093) ?
                          (|reg1114[(2'h3):(1'h0)]) : ((reg1072 ~^ forvar1106) ?
                              (~&reg1112) : $unsigned(forvar1137))));
                      reg1127 <= (!forvar1077);
                    end
                  else
                    begin
                      reg1124 <= $unsigned($signed((&$unsigned(reg1081))));
                      reg1125 <= (&$unsigned((-wire1046[(3'h4):(2'h2)])));
                    end
                  for (forvar1128 = (1'h0); (forvar1128 < (1'h1)); forvar1128 = (forvar1128 + (1'h1)))
                    begin
                      reg1129 <= ((($signed(reg1139) ?
                              (reg1128 >>> reg1121) : reg1065[(3'h5):(2'h2)]) ?
                          (+{reg1107}) : ((reg1072 & reg1103) - ((8'h9f) ~^ reg1050))) || forvar1114[(2'h3):(2'h3)]);
                      reg1130 <= forvar1094;
                      reg1131 <= reg1117;
                      reg1132 <= forvar1083;
                    end
                end
              reg1133 <= (8'ha3);
            end
          if (reg1084)
            begin
              reg1140 <= $unsigned(forvar1061);
            end
          else
            begin
              if ($signed((8'h9d)))
                begin
                  if (($signed(((+forvar1109) ?
                          $unsigned(forvar1130) : reg1126[(1'h0):(1'h0)])) ?
                      $unsigned(reg1116) : (~|reg1089[(3'h6):(1'h1)])))
                    begin
                      reg1140 <= $signed($signed(forvar1109[(3'h7):(3'h6)]));
                      reg1141 <= (+$signed(((reg1140 ?
                          reg1136 : (8'hb8)) >= reg1134[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg1140 <= reg1090;
                    end
                end
              else
                begin
                  reg1140 <= forvar1088[(1'h1):(1'h1)];
                  reg1141 <= ((+(!$signed(forvar1126))) ?
                      $unsigned($unsigned(reg1125)) : reg1111);
                  for (forvar1142 = (1'h0); (forvar1142 < (2'h2)); forvar1142 = (forvar1142 + (1'h1)))
                    begin
                      reg1143 <= reg1050;
                      reg1144 <= $signed((((reg1083 ? reg1111 : reg1089) ?
                              (forvar1126 ? reg1055 : reg1117) : (~^reg1097)) ?
                          reg1072[(1'h1):(1'h0)] : $unsigned($signed(reg1121))));
                      reg1145 <= $unsigned($signed(reg1123[(4'h8):(3'h6)]));
                    end
                end
            end
          for (forvar1146 = (1'h0); (forvar1146 < (1'h1)); forvar1146 = (forvar1146 + (1'h1)))
            begin
              for (forvar1147 = (1'h0); (forvar1147 < (1'h1)); forvar1147 = (forvar1147 + (1'h1)))
                begin
                  reg1148 <= $signed($unsigned(forvar1109));
                  reg1149 <= $unsigned(reg1133[(3'h7):(1'h1)]);
                end
              reg1150 <= ((((reg1148 ? reg1093 : reg1060) ?
                          $unsigned(reg1078) : (reg1104 ? reg1103 : reg1133)) ?
                      $signed((wire1043 ? forvar1137 : reg1065)) : reg1065) ?
                  reg1130 : $unsigned($unsigned((reg1111 == reg1053))));
            end
          for (forvar1151 = (1'h0); (forvar1151 < (2'h3)); forvar1151 = (forvar1151 + (1'h1)))
            begin
              reg1152 <= $unsigned((~|((|reg1113) || (8'ha2))));
              reg1153 <= reg1134;
            end
        end
      else
        begin
          reg1109 <= reg1097;
        end
      if ($signed(($signed(forvar1146) < forvar1147[(1'h0):(1'h0)])))
        begin
          for (forvar1154 = (1'h0); (forvar1154 < (2'h3)); forvar1154 = (forvar1154 + (1'h1)))
            begin
              for (forvar1155 = (1'h0); (forvar1155 < (1'h0)); forvar1155 = (forvar1155 + (1'h1)))
                begin
                  reg1156 <= (~^(^~$signed($signed(forvar1120))));
                end
              reg1157 <= forvar1095;
            end
        end
      else
        begin
          if ($signed($signed({$signed(forvar1155)})))
            begin
              if ((8'ha7))
                begin
                  for (forvar1154 = (1'h0); (forvar1154 < (1'h1)); forvar1154 = (forvar1154 + (1'h1)))
                    begin
                      reg1155 <= reg1127;
                      reg1156 <= reg1057;
                      reg1157 <= (~&((~&$unsigned(reg1125)) | (((8'ha3) ?
                          reg1099 : forvar1120) & $signed(forvar1147))));
                      reg1158 <= (~^$signed($unsigned($signed(reg1118))));
                    end
                  for (forvar1159 = (1'h0); (forvar1159 < (2'h2)); forvar1159 = (forvar1159 + (1'h1)))
                    begin
                      reg1160 <= (8'ha1);
                      reg1161 <= (^~(~reg1116));
                      reg1162 <= (|$signed(($signed((8'ha1)) && reg1122)));
                    end
                end
              else
                begin
                  if ((8'hb3))
                    begin
                      reg1154 <= $unsigned(((~|forvar1088[(4'h9):(3'h5)]) <<< ((reg1111 ?
                              reg1085 : (8'ha7)) ?
                          reg1135 : (~^reg1132))));
                      reg1155 <= $signed($signed(reg1065[(2'h3):(1'h0)]));
                      reg1156 <= reg1086;
                    end
                  else
                    begin
                      reg1154 <= (reg1099[(3'h6):(1'h0)] ?
                          ($signed($unsigned(forvar1155)) ?
                              (^reg1135) : $signed(reg1092)) : ({$unsigned(forvar1147)} ?
                              (~^forvar1120) : $signed($unsigned(reg1069))));
                      reg1155 <= {reg1112[(1'h1):(1'h0)]};
                      reg1156 <= $signed((forvar1079 << $unsigned($signed(reg1100))));
                      reg1157 <= (8'h9f);
                    end
                  for (forvar1158 = (1'h0); (forvar1158 < (2'h3)); forvar1158 = (forvar1158 + (1'h1)))
                    begin
                      reg1159 <= (forvar1049[(2'h3):(2'h2)] - reg1065);
                      reg1160 <= (forvar1129[(4'ha):(3'h4)] != ((+$unsigned((8'hb1))) <= reg1131[(4'h8):(3'h5)]));
                      reg1161 <= $signed(forvar1047[(1'h0):(1'h0)]);
                    end
                end
              for (forvar1163 = (1'h0); (forvar1163 < (1'h1)); forvar1163 = (forvar1163 + (1'h1)))
                begin
                  if ($unsigned(($signed((reg1160 ? reg1091 : reg1157)) ?
                      forvar1126 : (|(reg1122 ? (8'had) : reg1117)))))
                    begin
                      reg1164 <= ({((forvar1079 ?
                                  (8'ha2) : (8'hb0)) ^ ((8'ha6) * forvar1098))} ?
                          $unsigned($unsigned($unsigned((8'hba)))) : (((reg1078 ?
                                  forvar1114 : reg1148) <<< (reg1090 ?
                                  forvar1147 : (8'hba))) ?
                              $signed($unsigned(reg1085)) : {(reg1085 ?
                                      reg1096 : reg1159)}));
                      reg1165 <= reg1066;
                      reg1166 <= (~|(((wire1044 ? reg1139 : forvar1128) ?
                              (forvar1098 || reg1051) : (reg1139 ?
                                  forvar1130 : reg1160)) ?
                          ($signed((8'haf)) ?
                              {reg1148} : $unsigned(reg1099)) : reg1080[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg1164 <= ((8'hb6) + forvar1047[(2'h2):(1'h0)]);
                      reg1165 <= (~|(reg1165[(3'h6):(1'h0)] ?
                          forvar1047[(1'h1):(1'h1)] : reg1112[(2'h2):(1'h0)]));
                      reg1166 <= (8'haf);
                      reg1167 <= $signed($unsigned(($signed(forvar1154) ?
                          $signed(reg1059) : $signed(reg1103))));
                    end
                end
              for (forvar1168 = (1'h0); (forvar1168 < (1'h1)); forvar1168 = (forvar1168 + (1'h1)))
                begin
                  for (forvar1169 = (1'h0); (forvar1169 < (1'h1)); forvar1169 = (forvar1169 + (1'h1)))
                    begin
                      reg1170 <= $unsigned(reg1058);
                    end
                end
            end
          else
            begin
              for (forvar1154 = (1'h0); (forvar1154 < (2'h2)); forvar1154 = (forvar1154 + (1'h1)))
                begin
                  reg1155 <= (^~$signed((reg1105 <= (reg1084 > reg1058))));
                  for (forvar1156 = (1'h0); (forvar1156 < (1'h1)); forvar1156 = (forvar1156 + (1'h1)))
                    begin
                      reg1157 <= $signed((8'h9c));
                      reg1158 <= $signed(($unsigned((reg1138 ^ reg1059)) ^~ {((8'ha5) << reg1073)}));
                      reg1159 <= ($signed({(reg1153 ^~ forvar1088)}) < (reg1112[(1'h0):(1'h0)] ?
                          forvar1079[(2'h2):(2'h2)] : $signed((~&(8'had)))));
                    end
                end
              if ((+$unsigned(reg1143[(4'h9):(3'h4)])))
                begin
                  for (forvar1160 = (1'h0); (forvar1160 < (2'h2)); forvar1160 = (forvar1160 + (1'h1)))
                    begin
                      reg1161 <= forvar1085[(3'h7):(1'h1)];
                      reg1162 <= reg1167;
                    end
                  for (forvar1163 = (1'h0); (forvar1163 < (2'h2)); forvar1163 = (forvar1163 + (1'h1)))
                    begin
                      reg1164 <= $signed(reg1071);
                      reg1165 <= (+$signed(reg1156[(2'h3):(1'h0)]));
                    end
                  if ((~^(8'ha4)))
                    begin
                      reg1166 <= {(~$signed((forvar1094 ? (8'had) : (8'h9f))))};
                      reg1167 <= (reg1141 && reg1132[(3'h7):(1'h1)]);
                      reg1168 <= (reg1141 << $signed(((|reg1085) ^ $unsigned(reg1087))));
                      reg1169 <= {$signed($unsigned((reg1123 <= forvar1095)))};
                    end
                  else
                    begin
                      reg1166 <= forvar1130[(3'h7):(3'h7)];
                      reg1167 <= $unsigned($unsigned((~|forvar1114)));
                    end
                  for (forvar1170 = (1'h0); (forvar1170 < (1'h1)); forvar1170 = (forvar1170 + (1'h1)))
                    begin
                      reg1171 <= $unsigned(forvar1154);
                    end
                end
              else
                begin
                  if ((-(8'ha8)))
                    begin
                      reg1160 <= $signed((reg1117 == reg1141[(1'h0):(1'h0)]));
                      reg1161 <= (forvar1130 >= reg1121);
                    end
                  else
                    begin
                      reg1160 <= reg1168[(2'h3):(1'h0)];
                      reg1161 <= {((reg1112[(2'h2):(2'h2)] ?
                                  $unsigned((8'hb9)) : reg1076[(4'h9):(1'h1)]) ?
                              ($signed(forvar1102) ?
                                  (8'haf) : {(8'hb6)}) : $signed({forvar1158}))};
                      reg1162 <= ($unsigned(wire1042) <= (reg1093 ?
                          $signed(((8'h9f) ?
                              (8'hb1) : forvar1160)) : $unsigned(reg1091[(2'h3):(1'h0)])));
                    end
                  for (forvar1163 = (1'h0); (forvar1163 < (2'h2)); forvar1163 = (forvar1163 + (1'h1)))
                    begin
                      reg1164 <= {reg1111[(2'h3):(1'h1)]};
                    end
                  for (forvar1165 = (1'h0); (forvar1165 < (1'h1)); forvar1165 = (forvar1165 + (1'h1)))
                    begin
                      reg1166 <= {{(^(reg1087 ? reg1100 : forvar1075))}};
                      reg1167 <= $signed($signed(forvar1160[(1'h1):(1'h1)]));
                      reg1168 <= ({({reg1153} ?
                              (&(8'ha4)) : (~&forvar1083))} ~^ (-(+(~&reg1107))));
                      reg1169 <= $unsigned(forvar1047);
                    end
                  for (forvar1170 = (1'h0); (forvar1170 < (1'h1)); forvar1170 = (forvar1170 + (1'h1)))
                    begin
                      reg1171 <= $unsigned(reg1065);
                    end
                end
              reg1172 <= $unsigned(reg1123);
            end
          for (forvar1173 = (1'h0); (forvar1173 < (2'h2)); forvar1173 = (forvar1173 + (1'h1)))
            begin
              if ((^~forvar1128))
                begin
                  reg1174 <= reg1153;
                  for (forvar1175 = (1'h0); (forvar1175 < (2'h3)); forvar1175 = (forvar1175 + (1'h1)))
                    begin
                      reg1176 <= ((((reg1084 ? reg1165 : forvar1074) ?
                          (forvar1074 ? reg1133 : forvar1094) : (reg1080 ?
                              (8'ha5) : reg1082)) <= $signed(reg1114[(4'hf):(4'h8)])) >= $unsigned($unsigned($unsigned(forvar1175))));
                      reg1177 <= ($unsigned($signed(forvar1098[(1'h0):(1'h0)])) ?
                          $unsigned((forvar1175 ?
                              $signed(reg1104) : (reg1144 ?
                                  (8'h9e) : forvar1095))) : $signed(($unsigned(reg1053) ?
                              reg1164 : (|forvar1102))));
                      reg1178 <= (^reg1078);
                    end
                  if (forvar1098)
                    begin
                      reg1179 <= forvar1163;
                      reg1180 <= (reg1069[(2'h2):(2'h2)] || $signed($signed(((8'hb4) ?
                          (8'ha3) : reg1064))));
                    end
                  else
                    begin
                      reg1179 <= (~|reg1081);
                      reg1180 <= $signed(forvar1128[(4'h9):(4'h9)]);
                      reg1181 <= (($signed(reg1109) << {$unsigned(reg1125)}) || reg1170);
                      reg1182 <= ($signed(forvar1137[(1'h0):(1'h0)]) + $signed(({wire1043} << (8'hba))));
                    end
                end
              else
                begin
                  for (forvar1174 = (1'h0); (forvar1174 < (2'h2)); forvar1174 = (forvar1174 + (1'h1)))
                    begin
                      reg1175 <= ((+(8'ha2)) >> $unsigned(wire1046[(4'hc):(4'hc)]));
                      reg1176 <= reg1157;
                    end
                  for (forvar1177 = (1'h0); (forvar1177 < (2'h2)); forvar1177 = (forvar1177 + (1'h1)))
                    begin
                      reg1178 <= reg1155;
                      reg1179 <= reg1078;
                    end
                  reg1180 <= $unsigned((~|(reg1145[(2'h2):(2'h2)] != (forvar1169 ?
                      reg1060 : reg1070))));
                  for (forvar1181 = (1'h0); (forvar1181 < (2'h3)); forvar1181 = (forvar1181 + (1'h1)))
                    begin
                      reg1182 <= (reg1150[(3'h4):(2'h2)] ?
                          (((reg1130 || forvar1106) >>> {reg1055}) & ((8'hb4) ?
                              ((8'ha0) >>> reg1057) : $signed(forvar1181))) : $unsigned($unsigned(reg1092[(2'h2):(1'h1)])));
                    end
                end
              if (($signed(forvar1054) ~^ (({reg1055} ?
                  $signed(forvar1175) : (~|reg1179)) != (reg1169 << reg1128))))
                begin
                  if ((8'h9c))
                    begin
                      reg1183 <= (!reg1153);
                      reg1184 <= {$unsigned((&(forvar1083 == reg1148)))};
                      reg1185 <= forvar1177;
                    end
                  else
                    begin
                      reg1183 <= $signed((reg1175[(2'h3):(1'h0)] >= reg1092));
                    end
                end
              else
                begin
                  for (forvar1183 = (1'h0); (forvar1183 < (1'h1)); forvar1183 = (forvar1183 + (1'h1)))
                    begin
                      reg1184 <= $signed(reg1050[(2'h3):(2'h3)]);
                      reg1185 <= $unsigned(((+(forvar1129 ?
                          reg1097 : reg1161)) >>> $unsigned((~&forvar1083))));
                      reg1186 <= $signed((reg1136 != $unsigned((reg1168 <= reg1109))));
                    end
                end
              if ((($unsigned($unsigned(reg1149)) <<< (forvar1075[(3'h5):(2'h3)] && forvar1117)) << reg1078[(3'h6):(3'h5)]))
                begin
                  if ($unsigned(forvar1061))
                    begin
                      reg1187 <= reg1164[(1'h1):(1'h1)];
                      reg1188 <= (((&(reg1161 ?
                          reg1123 : forvar1126)) && reg1105[(3'h5):(1'h1)]) != $signed(((reg1090 ~^ reg1086) ~^ $unsigned(reg1128))));
                      reg1189 <= forvar1085[(3'h6):(3'h5)];
                      reg1190 <= $signed({$unsigned((reg1155 - (8'ha3)))});
                    end
                  else
                    begin
                      reg1187 <= $unsigned($signed((!$signed(reg1110))));
                      reg1188 <= {$unsigned((((8'hb2) ?
                              (8'h9c) : reg1068) && reg1055[(3'h5):(2'h2)]))};
                    end
                  if ($signed((forvar1177[(3'h4):(3'h4)] <<< forvar1151)))
                    begin
                      reg1191 <= $signed(($signed($unsigned(forvar1106)) >= (&reg1078[(3'h4):(2'h2)])));
                      reg1192 <= reg1157[(3'h4):(2'h3)];
                      reg1193 <= ((forvar1181[(3'h7):(3'h5)] ?
                          $unsigned($unsigned(reg1165)) : reg1105) ~^ ($signed((reg1145 + reg1068)) ^ (~|reg1189[(1'h0):(1'h0)])));
                      reg1194 <= (~^forvar1142[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg1191 <= (+$unsigned(({forvar1123} <<< (reg1156 >>> reg1068))));
                      reg1192 <= (forvar1074 ?
                          forvar1102 : ($signed(reg1099) ?
                              (~|reg1100[(3'h5):(3'h4)]) : $signed($signed((8'hab)))));
                      reg1193 <= ((reg1100 ?
                              (!(reg1122 << reg1165)) : reg1162) ?
                          {(~|(reg1134 == reg1051))} : $unsigned(reg1183[(3'h5):(1'h1)]));
                    end
                  if (($unsigned(($unsigned((8'ha0)) > forvar1117)) != reg1090[(4'ha):(3'h4)]))
                    begin
                      reg1195 <= reg1097;
                      reg1196 <= (~^($signed((~|(8'haa))) ?
                          ((reg1170 + reg1118) ?
                              (forvar1137 == (8'ha0)) : {(8'haf)}) : $signed((~^reg1122))));
                      reg1197 <= (8'h9f);
                    end
                  else
                    begin
                      reg1195 <= (!{reg1193});
                      reg1196 <= (~(forvar1106[(2'h3):(1'h0)] < (^~(reg1180 ?
                          (8'ha6) : wire1046))));
                    end
                  if (reg1182)
                    begin
                      reg1198 <= (^$unsigned($signed((^~reg1155))));
                      reg1199 <= $unsigned((8'hb6));
                      reg1200 <= forvar1094;
                    end
                  else
                    begin
                      reg1198 <= reg1154[(4'h8):(2'h3)];
                      reg1199 <= reg1127[(2'h3):(1'h0)];
                      reg1200 <= forvar1173;
                      reg1201 <= (+$signed({$unsigned(forvar1106)}));
                    end
                end
              else
                begin
                  reg1187 <= ((!reg1117[(4'h9):(1'h1)]) == $signed(forvar1154));
                  for (forvar1188 = (1'h0); (forvar1188 < (1'h0)); forvar1188 = (forvar1188 + (1'h1)))
                    begin
                      reg1189 <= ($signed(reg1105) ?
                          $unsigned($signed(reg1140[(3'h5):(1'h0)])) : (&reg1144[(3'h4):(2'h2)]));
                      reg1190 <= ($signed({(reg1116 ?
                              reg1199 : reg1143)}) >>> $unsigned(reg1115[(4'h9):(3'h7)]));
                      reg1191 <= $unsigned(reg1115);
                    end
                  if (forvar1083[(2'h2):(2'h2)])
                    begin
                      reg1192 <= (^~reg1131);
                      reg1193 <= $signed((reg1195[(1'h0):(1'h0)] ?
                          $unsigned((reg1201 <= reg1128)) : $signed($signed(reg1176))));
                      reg1194 <= {(~&reg1136[(3'h5):(1'h0)])};
                      reg1195 <= (-($unsigned((forvar1173 ?
                              reg1120 : forvar1159)) ?
                          reg1087[(4'h9):(1'h1)] : $unsigned({reg1099})));
                    end
                  else
                    begin
                      reg1192 <= wire1045;
                      reg1193 <= reg1152[(4'hf):(3'h4)];
                    end
                end
            end
          if ({$unsigned((8'hae))})
            begin
              reg1202 <= $signed(reg1062[(3'h4):(1'h0)]);
              for (forvar1203 = (1'h0); (forvar1203 < (1'h1)); forvar1203 = (forvar1203 + (1'h1)))
                begin
                  for (forvar1204 = (1'h0); (forvar1204 < (1'h0)); forvar1204 = (forvar1204 + (1'h1)))
                    begin
                      reg1205 <= $signed(reg1092);
                    end
                end
              if ($signed((forvar1117[(2'h3):(1'h1)] ~^ $unsigned(reg1127))))
                begin
                  for (forvar1206 = (1'h0); (forvar1206 < (1'h1)); forvar1206 = (forvar1206 + (1'h1)))
                    begin
                      reg1207 <= forvar1159;
                    end
                  for (forvar1208 = (1'h0); (forvar1208 < (1'h0)); forvar1208 = (forvar1208 + (1'h1)))
                    begin
                      reg1209 <= (forvar1120[(1'h0):(1'h0)] < $signed(({forvar1154} != $signed(reg1058))));
                      reg1210 <= $signed(reg1202);
                      reg1211 <= $unsigned(($unsigned(forvar1120[(5'h10):(4'he)]) ?
                          reg1066[(4'hc):(3'h4)] : (!reg1159[(3'h5):(1'h1)])));
                      reg1212 <= $unsigned($unsigned(($unsigned(forvar1168) >>> reg1120)));
                    end
                end
              else
                begin
                  for (forvar1206 = (1'h0); (forvar1206 < (1'h1)); forvar1206 = (forvar1206 + (1'h1)))
                    begin
                      reg1207 <= forvar1168[(1'h0):(1'h0)];
                      reg1208 <= reg1133;
                    end
                  if ($unsigned(reg1063[(2'h2):(2'h2)]))
                    begin
                      reg1209 <= forvar1129[(4'hd):(4'hc)];
                      reg1210 <= reg1209;
                    end
                  else
                    begin
                      reg1209 <= {reg1199[(1'h1):(1'h1)]};
                    end
                  for (forvar1211 = (1'h0); (forvar1211 < (1'h1)); forvar1211 = (forvar1211 + (1'h1)))
                    begin
                      reg1212 <= (~|$unsigned((~^reg1169)));
                    end
                  if (reg1134[(2'h2):(1'h1)])
                    begin
                      reg1213 <= $signed($unsigned($signed(reg1153)));
                      reg1214 <= (reg1080[(3'h4):(1'h0)] ~^ (^~$unsigned({forvar1168})));
                    end
                  else
                    begin
                      reg1213 <= forvar1159[(3'h5):(3'h4)];
                      reg1214 <= {{(~$signed(reg1073))}};
                      reg1215 <= reg1168[(3'h5):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar1202 = (1'h0); (forvar1202 < (2'h3)); forvar1202 = (forvar1202 + (1'h1)))
                begin
                  if ({reg1130[(4'he):(2'h3)]})
                    begin
                      reg1203 <= reg1078;
                      reg1204 <= reg1179;
                    end
                  else
                    begin
                      reg1203 <= reg1084;
                      reg1204 <= {$signed($signed(reg1108[(4'h9):(2'h2)]))};
                      reg1205 <= (~|(8'h9d));
                    end
                  for (forvar1206 = (1'h0); (forvar1206 < (1'h1)); forvar1206 = (forvar1206 + (1'h1)))
                    begin
                      reg1207 <= $signed(reg1145);
                      reg1208 <= (~^((~^reg1062) ?
                          ((reg1083 ? reg1177 : reg1212) <= (forvar1154 ?
                              reg1127 : reg1071)) : {$signed(reg1194)}));
                      reg1209 <= (-reg1133);
                    end
                  if ((forvar1165[(2'h3):(1'h0)] ?
                      reg1181 : $unsigned(($unsigned(reg1080) - $unsigned(reg1171)))))
                    begin
                      reg1210 <= $unsigned({$unsigned((|(8'hba)))});
                      reg1211 <= reg1194[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg1210 <= (~^reg1154[(1'h0):(1'h0)]);
                      reg1211 <= $unsigned(($unsigned($unsigned(forvar1211)) ?
                          ((reg1128 ?
                              reg1057 : forvar1137) | forvar1137[(1'h0):(1'h0)]) : (^$signed(reg1160))));
                    end
                end
              for (forvar1212 = (1'h0); (forvar1212 < (2'h2)); forvar1212 = (forvar1212 + (1'h1)))
                begin
                  if (reg1212)
                    begin
                      reg1213 <= (forvar1165 ?
                          reg1091[(2'h3):(2'h3)] : (reg1164 ?
                              ((reg1182 | reg1109) ?
                                  (forvar1079 ?
                                      reg1159 : reg1117) : (8'ha5)) : ($unsigned(forvar1130) >>> $signed(forvar1158))));
                      reg1214 <= forvar1142;
                      reg1215 <= reg1072;
                    end
                  else
                    begin
                      reg1213 <= $signed({{reg1188}});
                      reg1214 <= ((~|(reg1133[(2'h3):(1'h0)] <= (^forvar1109))) ?
                          $signed($unsigned((reg1175 <<< (8'hba)))) : ({(reg1203 ?
                                  forvar1146 : reg1179)} > $unsigned($signed(reg1202))));
                    end
                end
              for (forvar1216 = (1'h0); (forvar1216 < (2'h2)); forvar1216 = (forvar1216 + (1'h1)))
                begin
                  if ({(($signed(reg1105) ? $unsigned(reg1065) : (~&reg1060)) ?
                          reg1119 : {{(8'h9c)}})})
                    begin
                      reg1217 <= forvar1106[(2'h3):(2'h2)];
                      reg1218 <= {$unsigned($unsigned(((8'haa) | reg1110)))};
                      reg1219 <= (!($signed((|reg1195)) ?
                          reg1170[(3'h7):(2'h3)] : ((reg1213 >= forvar1109) ?
                              (forvar1177 ~^ reg1107) : (-reg1114))));
                      reg1220 <= $unsigned(((+(forvar1151 ?
                              reg1174 : reg1208)) ?
                          reg1187 : (~&(reg1164 << reg1060))));
                    end
                  else
                    begin
                      reg1217 <= ((reg1064[(4'hd):(4'hc)] <= ((~&forvar1155) ?
                              forvar1130 : (~|reg1183))) ?
                          ($unsigned(reg1096[(3'h6):(3'h6)]) ?
                              forvar1129 : (reg1156 ^~ (reg1210 * reg1123))) : ((forvar1175[(1'h1):(1'h0)] ?
                                  (~^reg1128) : (!forvar1174)) ?
                              forvar1088 : (forvar1188 ?
                                  $signed(reg1130) : $signed((8'hb7)))));
                      reg1218 <= (8'haa);
                      reg1219 <= ((({forvar1216} && (~(8'haa))) ?
                          $signed((reg1132 ?
                              (8'hac) : reg1208)) : $signed((8'hb4))) != $unsigned($signed(wire1046[(4'ha):(4'h9)])));
                    end
                  for (forvar1221 = (1'h0); (forvar1221 < (2'h2)); forvar1221 = (forvar1221 + (1'h1)))
                    begin
                      reg1222 <= $signed($signed({$unsigned(forvar1065)}));
                    end
                  reg1223 <= $signed(($unsigned($signed(reg1096)) ?
                      $unsigned((reg1086 > reg1191)) : ((|reg1080) ?
                          forvar1074[(1'h1):(1'h0)] : (forvar1126 ?
                              (8'hac) : reg1194))));
                end
              for (forvar1224 = (1'h0); (forvar1224 < (1'h0)); forvar1224 = (forvar1224 + (1'h1)))
                begin
                  if ({({$signed(reg1061)} ? reg1065[(2'h3):(2'h2)] : reg1101)})
                    begin
                      reg1225 <= $unsigned(({(^~reg1195)} ?
                          reg1129 : $signed((&forvar1123))));
                      reg1226 <= (($unsigned({reg1090}) == reg1058) ?
                          reg1103[(3'h5):(1'h1)] : (reg1127 >= wire1043[(2'h2):(2'h2)]));
                      reg1227 <= $signed(reg1153[(4'ha):(3'h4)]);
                    end
                  else
                    begin
                      reg1225 <= (8'hb5);
                      reg1226 <= forvar1170;
                      reg1227 <= $unsigned($unsigned((reg1126[(1'h1):(1'h1)] ?
                          $signed(forvar1077) : $unsigned((8'hb3)))));
                    end
                  for (forvar1228 = (1'h0); (forvar1228 < (1'h0)); forvar1228 = (forvar1228 + (1'h1)))
                    begin
                      reg1229 <= $signed(((-forvar1181) >> reg1129[(1'h0):(1'h0)]));
                      reg1230 <= (^$unsigned((reg1104[(2'h2):(1'h0)] * (forvar1117 ?
                          reg1055 : reg1051))));
                      reg1231 <= forvar1158;
                      reg1232 <= $unsigned(forvar1130[(3'h4):(3'h4)]);
                    end
                end
            end
          if (($signed($signed({reg1097})) ?
              $signed($signed((forvar1169 > (8'ha0)))) : $unsigned($signed((^~forvar1106)))))
            begin
              if ($signed((~&reg1066)))
                begin
                  for (forvar1233 = (1'h0); (forvar1233 < (2'h3)); forvar1233 = (forvar1233 + (1'h1)))
                    begin
                      reg1234 <= (((^reg1150[(4'h9):(3'h4)]) ?
                          (&(reg1110 * forvar1075)) : reg1149[(3'h4):(3'h4)]) ^ (~((8'ha7) ^~ reg1217)));
                      reg1235 <= wire1046[(4'hd):(4'ha)];
                      reg1236 <= forvar1173;
                    end
                end
              else
                begin
                  if ({(({reg1211} ? forvar1065 : (!reg1175)) ?
                          (-(+reg1129)) : reg1232[(4'h8):(3'h5)])})
                    begin
                      reg1233 <= (|$unsigned((8'hab)));
                      reg1234 <= ({{$unsigned((8'hb6))}} ?
                          (~^reg1083) : (~&$signed((reg1199 ?
                              forvar1077 : (8'ha9)))));
                      reg1235 <= {$signed($signed($unsigned(reg1168)))};
                    end
                  else
                    begin
                      reg1233 <= ($signed(reg1197[(2'h3):(2'h3)]) ?
                          {({forvar1158} ?
                                  (8'hb4) : $unsigned(reg1186))} : reg1135[(2'h3):(1'h1)]);
                      reg1234 <= $unsigned(forvar1129);
                      reg1235 <= reg1172[(2'h2):(1'h1)];
                    end
                  reg1236 <= reg1193[(3'h6):(3'h5)];
                  reg1237 <= $unsigned({(forvar1106[(3'h5):(2'h2)] ?
                          (forvar1208 ? reg1060 : reg1174) : (8'hb5))});
                  if (((~^({(8'haa)} & (reg1159 ? wire1043 : forvar1224))) ?
                      $signed($signed(forvar1130[(1'h0):(1'h0)])) : ({reg1089} ?
                          reg1223 : reg1068[(3'h7):(2'h2)])))
                    begin
                      reg1238 <= $unsigned(((forvar1151[(3'h7):(3'h7)] ?
                              (forvar1147 & (8'h9d)) : ((8'ha2) & reg1187)) ?
                          $signed(((8'hac) ?
                              reg1166 : forvar1170)) : ((reg1112 | reg1145) >> (forvar1208 ?
                              forvar1154 : forvar1085))));
                      reg1239 <= reg1227[(4'h8):(1'h0)];
                      reg1240 <= (!reg1167);
                      reg1241 <= {((8'hae) ?
                              {reg1105[(3'h6):(3'h4)]} : forvar1211[(3'h6):(2'h3)])};
                    end
                  else
                    begin
                      reg1238 <= ($unsigned($signed({reg1097})) + $signed((-{reg1072})));
                      reg1239 <= $unsigned($signed(({reg1223} != $unsigned(forvar1088))));
                      reg1240 <= $unsigned(reg1156);
                      reg1241 <= reg1155[(3'h4):(1'h0)];
                    end
                end
              if (((((&forvar1048) > $signed(reg1062)) <= ((reg1213 ?
                          reg1081 : forvar1224) ?
                      (!forvar1126) : forvar1088)) ?
                  {$signed($unsigned(forvar1049))} : (~&$unsigned((reg1205 ?
                      forvar1154 : reg1231)))))
                begin
                  reg1242 <= $unsigned(reg1185[(2'h2):(2'h2)]);
                end
              else
                begin
                  if ($unsigned(reg1238[(3'h6):(1'h1)]))
                    begin
                      reg1242 <= $unsigned((^forvar1233[(1'h0):(1'h0)]));
                      reg1243 <= $signed(reg1180);
                      reg1244 <= $unsigned((^~(reg1124[(4'h8):(1'h0)] > ((8'hb2) & wire1043))));
                      reg1245 <= (-$signed({forvar1147}));
                    end
                  else
                    begin
                      reg1242 <= $unsigned($unsigned((-reg1226)));
                      reg1243 <= $unsigned((reg1103[(3'h4):(1'h0)] ?
                          (!reg1055[(3'h5):(3'h5)]) : {(~reg1187)}));
                      reg1244 <= (reg1136[(4'hb):(1'h1)] ?
                          (reg1152 ?
                              $signed((+reg1118)) : (((8'ha3) == forvar1221) >> $unsigned(reg1090))) : $signed(reg1191[(4'hc):(4'h9)]));
                      reg1245 <= {(^reg1107[(1'h1):(1'h0)])};
                    end
                end
              for (forvar1246 = (1'h0); (forvar1246 < (1'h0)); forvar1246 = (forvar1246 + (1'h1)))
                begin
                  reg1247 <= (reg1066 ?
                      $unsigned(reg1130) : forvar1160[(4'ha):(2'h2)]);
                  for (forvar1248 = (1'h0); (forvar1248 < (1'h1)); forvar1248 = (forvar1248 + (1'h1)))
                    begin
                      reg1249 <= (reg1066 ^ $unsigned(reg1116[(2'h3):(1'h0)]));
                    end
                  for (forvar1250 = (1'h0); (forvar1250 < (1'h1)); forvar1250 = (forvar1250 + (1'h1)))
                    begin
                      reg1251 <= $unsigned(reg1114);
                      reg1252 <= $unsigned($unsigned(((+reg1085) ?
                          reg1133 : $unsigned((8'haf)))));
                    end
                end
            end
          else
            begin
              if ((8'haa))
                begin
                  for (forvar1233 = (1'h0); (forvar1233 < (1'h0)); forvar1233 = (forvar1233 + (1'h1)))
                    begin
                      reg1234 <= reg1180;
                      reg1235 <= reg1050[(4'hb):(4'h9)];
                    end
                  if ($unsigned((~&reg1189)))
                    begin
                      reg1236 <= (~^(!{$unsigned((8'ha3))}));
                    end
                  else
                    begin
                      reg1236 <= $signed((((reg1112 >>> forvar1165) ?
                          (^reg1234) : $unsigned((8'h9e))) >= reg1188[(1'h0):(1'h0)]));
                    end
                  reg1237 <= (~|(~^($unsigned(reg1217) ?
                      (reg1068 >= reg1175) : reg1166[(4'hc):(3'h7)])));
                  for (forvar1238 = (1'h0); (forvar1238 < (1'h1)); forvar1238 = (forvar1238 + (1'h1)))
                    begin
                      reg1239 <= reg1241;
                      reg1240 <= {$unsigned((-(reg1156 ?
                              forvar1102 : forvar1074)))};
                      reg1241 <= $unsigned(($signed($unsigned(forvar1177)) * {$signed(reg1183)}));
                    end
                end
              else
                begin
                  for (forvar1233 = (1'h0); (forvar1233 < (2'h3)); forvar1233 = (forvar1233 + (1'h1)))
                    begin
                      reg1234 <= (reg1160 ?
                          forvar1163 : ((reg1211 != reg1110[(1'h0):(1'h0)]) > ((|reg1168) ?
                              (reg1083 | forvar1202) : reg1057)));
                    end
                  for (forvar1235 = (1'h0); (forvar1235 < (2'h3)); forvar1235 = (forvar1235 + (1'h1)))
                    begin
                      reg1236 <= {($unsigned(((8'ha7) ? reg1105 : wire1044)) ?
                              {reg1158} : $signed((reg1220 ?
                                  reg1144 : reg1210)))};
                      reg1237 <= $unsigned({($unsigned(reg1150) + (~&reg1219))});
                    end
                end
              reg1242 <= ($unsigned($signed(reg1126[(3'h6):(1'h1)])) < (8'ha9));
              reg1243 <= $signed(reg1160[(4'h9):(4'h8)]);
              for (forvar1244 = (1'h0); (forvar1244 < (2'h2)); forvar1244 = (forvar1244 + (1'h1)))
                begin
                  reg1245 <= (-(-$signed($signed((8'hb1)))));
                  if ((~((^$signed(forvar1158)) ?
                      ((reg1092 << reg1214) ?
                          {(8'had)} : forvar1077) : ($unsigned((8'ha8)) ?
                          forvar1047[(2'h2):(1'h1)] : $signed(reg1215)))))
                    begin
                      reg1246 <= {((^~reg1184[(1'h1):(1'h0)]) ?
                              ($unsigned(reg1143) * reg1061[(1'h0):(1'h0)]) : $signed((forvar1228 ?
                                  (8'hb7) : reg1125)))};
                    end
                  else
                    begin
                      reg1246 <= reg1145[(2'h2):(1'h1)];
                      reg1247 <= $signed((((reg1237 >> reg1055) ?
                              (forvar1114 ?
                                  forvar1238 : reg1188) : (reg1201 ^ reg1112)) ?
                          $signed($unsigned(reg1182)) : {(reg1230 >= wire1045)}));
                      reg1248 <= forvar1221;
                      reg1249 <= reg1072;
                    end
                  if ({$unsigned({$unsigned((8'ha5))})})
                    begin
                      reg1250 <= reg1219[(2'h2):(1'h0)];
                      reg1251 <= (reg1087[(4'h8):(4'h8)] ?
                          ((8'hb9) & ({reg1119} >> (reg1066 * forvar1183))) : ((reg1226[(1'h0):(1'h0)] == $signed(reg1208)) >>> reg1133[(3'h4):(1'h1)]));
                      reg1252 <= $unsigned({$signed((|reg1063))});
                      reg1253 <= (($unsigned((forvar1120 * reg1192)) * (+reg1108)) ?
                          ((^~{(8'ha5)}) ?
                              $unsigned($unsigned(reg1092)) : (reg1166 ^~ ((8'hae) < reg1215))) : ($signed((!reg1225)) < (8'ha3)));
                    end
                  else
                    begin
                      reg1250 <= {$unsigned($unsigned($signed(reg1103)))};
                      reg1251 <= reg1097;
                      reg1252 <= forvar1085;
                    end
                  for (forvar1254 = (1'h0); (forvar1254 < (1'h0)); forvar1254 = (forvar1254 + (1'h1)))
                    begin
                      reg1255 <= $unsigned((((~(8'hb9)) ?
                              reg1087 : reg1236[(2'h2):(1'h1)]) ?
                          ($unsigned(reg1104) ~^ wire1042[(3'h5):(1'h1)]) : reg1237));
                      reg1256 <= reg1219;
                      reg1257 <= (~|$unsigned(reg1096));
                      reg1258 <= (reg1126 ?
                          reg1160[(4'hf):(4'hd)] : $signed(reg1129[(2'h3):(1'h0)]));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned($signed((forvar1120 || forvar1188))))
        begin
          if (($signed($unsigned((^reg1212))) ?
              (!($unsigned((8'ha4)) ?
                  (reg1159 > reg1227) : {reg1181})) : $unsigned((8'ha6))))
            begin
              for (forvar1259 = (1'h0); (forvar1259 < (2'h3)); forvar1259 = (forvar1259 + (1'h1)))
                begin
                  for (forvar1260 = (1'h0); (forvar1260 < (2'h2)); forvar1260 = (forvar1260 + (1'h1)))
                    begin
                      reg1261 <= ((^~reg1108) > reg1255[(2'h3):(1'h1)]);
                      reg1262 <= {$signed(reg1186[(2'h3):(1'h0)])};
                    end
                  reg1263 <= (forvar1175[(1'h0):(1'h0)] & (8'ha9));
                  for (forvar1264 = (1'h0); (forvar1264 < (2'h2)); forvar1264 = (forvar1264 + (1'h1)))
                    begin
                      reg1265 <= (reg1143 - ((reg1076[(4'h9):(2'h2)] ?
                              reg1180 : reg1129) ?
                          $unsigned((~^(8'haa))) : $signed({reg1072})));
                    end
                end
              if (reg1130[(1'h1):(1'h1)])
                begin
                  for (forvar1266 = (1'h0); (forvar1266 < (1'h0)); forvar1266 = (forvar1266 + (1'h1)))
                    begin
                      reg1267 <= ($unsigned(reg1249[(3'h5):(1'h0)]) ?
                          (($signed(reg1056) | (reg1178 ^ forvar1211)) + $unsigned(reg1185)) : wire1042[(1'h0):(1'h0)]);
                      reg1268 <= ($unsigned($unsigned(forvar1156)) < (forvar1173[(4'hc):(3'h6)] ?
                          $unsigned($signed((8'h9e))) : $unsigned(forvar1074[(2'h2):(1'h0)])));
                    end
                  for (forvar1269 = (1'h0); (forvar1269 < (2'h2)); forvar1269 = (forvar1269 + (1'h1)))
                    begin
                      reg1270 <= (reg1226 - $unsigned(($unsigned(reg1225) <<< $signed(reg1214))));
                      reg1271 <= ($unsigned(((^forvar1047) + reg1087)) >> (+{forvar1088[(1'h0):(1'h0)]}));
                      reg1272 <= reg1245;
                      reg1273 <= $unsigned($signed(reg1214[(4'h8):(1'h1)]));
                    end
                end
              else
                begin
                  if ($signed(reg1082[(1'h0):(1'h0)]))
                    begin
                      reg1266 <= (reg1211[(2'h2):(1'h0)] + reg1053);
                      reg1267 <= $unsigned(reg1229[(2'h3):(2'h3)]);
                      reg1268 <= {forvar1211};
                    end
                  else
                    begin
                      reg1266 <= {{reg1065[(3'h7):(1'h0)]}};
                    end
                end
              reg1274 <= (reg1149 && $signed($unsigned((^reg1086))));
              for (forvar1275 = (1'h0); (forvar1275 < (1'h1)); forvar1275 = (forvar1275 + (1'h1)))
                begin
                  for (forvar1276 = (1'h0); (forvar1276 < (2'h3)); forvar1276 = (forvar1276 + (1'h1)))
                    begin
                      reg1277 <= $signed((reg1136 ?
                          $unsigned($unsigned(forvar1266)) : $signed(reg1272[(1'h1):(1'h0)])));
                      reg1278 <= $signed(($unsigned((8'ha7)) | (+$unsigned(reg1122))));
                      reg1279 <= forvar1049;
                      reg1280 <= ($unsigned(reg1105[(2'h2):(2'h2)]) - $signed(reg1128));
                    end
                end
            end
          else
            begin
              reg1259 <= $unsigned(((~&forvar1211[(2'h3):(2'h2)]) && (|(~reg1064))));
              for (forvar1260 = (1'h0); (forvar1260 < (1'h0)); forvar1260 = (forvar1260 + (1'h1)))
                begin
                  for (forvar1261 = (1'h0); (forvar1261 < (2'h2)); forvar1261 = (forvar1261 + (1'h1)))
                    begin
                      reg1262 <= (forvar1216 ?
                          $signed(((~reg1087) <<< (reg1237 & (8'hb2)))) : (({reg1073} || {reg1215}) ?
                              $unsigned(forvar1206) : ((forvar1154 ?
                                      (8'hb3) : forvar1129) ?
                                  (reg1166 ~^ reg1140) : (reg1174 == forvar1248))));
                    end
                  for (forvar1263 = (1'h0); (forvar1263 < (1'h0)); forvar1263 = (forvar1263 + (1'h1)))
                    begin
                      reg1264 <= reg1267[(3'h4):(3'h4)];
                      reg1265 <= wire1046;
                      reg1266 <= {$signed((|(reg1273 ? reg1093 : forvar1146)))};
                      reg1267 <= forvar1233[(2'h2):(1'h1)];
                    end
                end
            end
          reg1281 <= $signed((reg1218[(2'h3):(2'h3)] + $unsigned((reg1244 * forvar1151))));
        end
      else
        begin
          if ($signed((~|reg1121)))
            begin
              if ({forvar1211[(3'h6):(3'h6)]})
                begin
                  for (forvar1259 = (1'h0); (forvar1259 < (2'h2)); forvar1259 = (forvar1259 + (1'h1)))
                    begin
                      reg1260 <= {(|$unsigned(((8'hae) ? (8'hb5) : (8'hb9))))};
                      reg1261 <= ((reg1144[(4'hd):(3'h4)] ^~ ((|reg1116) ?
                          (|forvar1146) : (reg1103 ?
                              forvar1098 : reg1169))) ~^ {reg1051});
                    end
                  if ((|reg1081[(3'h7):(3'h7)]))
                    begin
                      reg1262 <= $signed($signed($unsigned(forvar1048)));
                      reg1263 <= ((~($signed((8'ha0)) & reg1255)) ?
                          $unsigned((8'haf)) : $unsigned(($signed((8'haf)) >>> (reg1066 << reg1108))));
                      reg1264 <= $unsigned($unsigned((reg1188 ?
                          (|(8'ha8)) : $unsigned(reg1121))));
                      reg1265 <= (reg1211[(3'h4):(1'h1)] - ({(reg1059 ?
                                  forvar1077 : forvar1130)} ?
                          (~|{reg1063}) : (reg1236[(2'h3):(1'h1)] || (forvar1173 ?
                              (8'hb9) : forvar1088))));
                    end
                  else
                    begin
                      reg1262 <= $signed({$signed(reg1148[(2'h3):(1'h0)])});
                      reg1263 <= {(~|(!(&reg1069)))};
                      reg1264 <= reg1270;
                    end
                  if (reg1062)
                    begin
                      reg1266 <= forvar1054;
                      reg1267 <= $signed((^$unsigned((reg1086 ?
                          reg1232 : (8'ha0)))));
                      reg1268 <= {reg1161[(2'h2):(1'h0)]};
                    end
                  else
                    begin
                      reg1266 <= (-(reg1084[(3'h6):(3'h5)] >>> (forvar1142 ?
                          (reg1222 ? reg1073 : forvar1202) : (reg1069 ?
                              reg1222 : reg1135))));
                      reg1267 <= ((^(~|{forvar1147})) ?
                          reg1281 : (reg1252 ?
                              (reg1136 ?
                                  $unsigned(forvar1246) : forvar1183) : reg1198));
                      reg1268 <= (^forvar1130[(4'h9):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar1259 = (1'h0); (forvar1259 < (1'h0)); forvar1259 = (forvar1259 + (1'h1)))
                    begin
                      reg1260 <= (-(+$unsigned((&reg1155))));
                      reg1261 <= reg1135[(1'h0):(1'h0)];
                      reg1262 <= $unsigned($unsigned((forvar1168[(2'h2):(1'h1)] ~^ reg1059[(2'h3):(1'h0)])));
                      reg1263 <= (forvar1154 ?
                          $unsigned((!(~&reg1233))) : reg1226);
                    end
                  for (forvar1264 = (1'h0); (forvar1264 < (1'h0)); forvar1264 = (forvar1264 + (1'h1)))
                    begin
                      reg1265 <= (~^{((~forvar1203) ?
                              (forvar1211 ?
                                  reg1068 : reg1117) : reg1226[(2'h2):(2'h2)])});
                      reg1266 <= ((+reg1168[(2'h3):(2'h3)]) - (|forvar1168));
                    end
                end
              for (forvar1269 = (1'h0); (forvar1269 < (2'h2)); forvar1269 = (forvar1269 + (1'h1)))
                begin
                  reg1270 <= ({$signed($unsigned((8'haa)))} < $unsigned($unsigned((^forvar1170))));
                  for (forvar1271 = (1'h0); (forvar1271 < (2'h2)); forvar1271 = (forvar1271 + (1'h1)))
                    begin
                      reg1272 <= forvar1048[(3'h4):(2'h3)];
                    end
                end
              if ($unsigned((^((^reg1272) ? reg1119 : reg1164))))
                begin
                  for (forvar1273 = (1'h0); (forvar1273 < (1'h0)); forvar1273 = (forvar1273 + (1'h1)))
                    begin
                      reg1274 <= {(8'haa)};
                      reg1275 <= reg1169;
                      reg1276 <= reg1052;
                      reg1277 <= reg1274;
                    end
                  if (reg1281)
                    begin
                      reg1278 <= $unsigned($signed(forvar1117));
                    end
                  else
                    begin
                      reg1278 <= $unsigned(reg1153);
                    end
                end
              else
                begin
                  for (forvar1273 = (1'h0); (forvar1273 < (1'h0)); forvar1273 = (forvar1273 + (1'h1)))
                    begin
                      reg1274 <= $unsigned({$signed($unsigned(reg1209))});
                      reg1275 <= ((forvar1266[(1'h0):(1'h0)] ~^ $signed(forvar1173[(3'h5):(3'h4)])) != reg1261[(4'hc):(4'hc)]);
                      reg1276 <= forvar1177;
                    end
                  for (forvar1277 = (1'h0); (forvar1277 < (1'h1)); forvar1277 = (forvar1277 + (1'h1)))
                    begin
                      reg1278 <= $signed($signed(reg1176[(3'h7):(3'h7)]));
                      reg1279 <= $unsigned(reg1261);
                    end
                  for (forvar1280 = (1'h0); (forvar1280 < (2'h2)); forvar1280 = (forvar1280 + (1'h1)))
                    begin
                      reg1281 <= reg1117[(3'h4):(1'h0)];
                      reg1282 <= reg1183;
                    end
                  if (reg1266[(1'h1):(1'h0)])
                    begin
                      reg1283 <= $unsigned($signed({(reg1058 ?
                              reg1148 : reg1140)}));
                    end
                  else
                    begin
                      reg1283 <= (^~(+(!forvar1083)));
                      reg1284 <= $unsigned({$signed({wire1044})});
                      reg1285 <= (8'ha8);
                      reg1286 <= reg1222;
                    end
                end
            end
          else
            begin
              reg1259 <= (reg1235[(2'h3):(2'h2)] ?
                  reg1247[(1'h0):(1'h0)] : (8'ha5));
              for (forvar1260 = (1'h0); (forvar1260 < (2'h2)); forvar1260 = (forvar1260 + (1'h1)))
                begin
                  if ((8'hb7))
                    begin
                      reg1261 <= (8'hab);
                      reg1262 <= ($signed(forvar1065) ?
                          (forvar1094[(3'h7):(3'h7)] <<< reg1092[(2'h3):(2'h3)]) : $signed(((^~reg1170) ?
                              (|reg1118) : reg1105[(4'hc):(4'h8)])));
                    end
                  else
                    begin
                      reg1261 <= (reg1183 + ($signed(reg1258) ?
                          ((forvar1147 ^ wire1042) ?
                              forvar1088 : {reg1192}) : (!(reg1279 || forvar1151))));
                      reg1262 <= $unsigned(forvar1156[(3'h7):(1'h0)]);
                      reg1263 <= ((+$signed(forvar1170)) ?
                          (-$unsigned(reg1277)) : (($signed(forvar1048) >>> forvar1077) ?
                              $signed((~^reg1149)) : ($signed(reg1115) ?
                                  (reg1242 ?
                                      (8'ha4) : (8'h9c)) : reg1130[(4'ha):(3'h6)])));
                      reg1264 <= (($unsigned({forvar1130}) != forvar1259[(2'h3):(2'h2)]) ?
                          forvar1169 : {reg1212});
                    end
                  if ((8'had))
                    begin
                      reg1265 <= reg1092[(1'h1):(1'h0)];
                      reg1266 <= ($signed(reg1168) ?
                          ((~|reg1135) ?
                              (((8'hb0) >>> reg1215) == (~^reg1213)) : {((8'haf) >> reg1144)}) : $unsigned($signed(reg1153[(2'h2):(1'h1)])));
                      reg1267 <= {(8'hba)};
                      reg1268 <= reg1239[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg1265 <= ($unsigned(reg1172) ?
                          (^~(forvar1109 << (~^reg1189))) : ((^~((8'hb1) ?
                                  reg1246 : forvar1183)) ?
                              (~$signed(reg1190)) : (8'hb7)));
                      reg1266 <= $unsigned((&$signed((forvar1117 - (8'hb0)))));
                    end
                  if (forvar1119[(3'h4):(1'h0)])
                    begin
                      reg1269 <= {$signed($signed((reg1154 ~^ forvar1088)))};
                      reg1270 <= reg1203;
                    end
                  else
                    begin
                      reg1269 <= reg1181;
                      reg1270 <= {$signed(reg1090)};
                      reg1271 <= (^{({(8'hb2)} == reg1064[(5'h10):(4'h9)])});
                      reg1272 <= {{{(reg1065 << reg1129)}}};
                    end
                  reg1273 <= ((((~^(8'had)) == $unsigned(forvar1128)) >>> $unsigned((|wire1045))) * reg1133[(1'h0):(1'h0)]);
                end
            end
          if ($signed(($signed($signed(forvar1246)) ?
              {$unsigned(reg1057)} : $signed(reg1063))))
            begin
              reg1287 <= reg1236;
              for (forvar1288 = (1'h0); (forvar1288 < (2'h3)); forvar1288 = (forvar1288 + (1'h1)))
                begin
                  if (((~forvar1147[(3'h6):(3'h5)]) ?
                      reg1191[(1'h1):(1'h0)] : ({((8'hb8) ~^ reg1283)} ?
                          forvar1250 : forvar1250[(3'h5):(1'h1)])))
                    begin
                      reg1289 <= {(|reg1271[(2'h2):(1'h1)])};
                    end
                  else
                    begin
                      reg1289 <= reg1179[(4'hc):(1'h1)];
                      reg1290 <= (8'haa);
                    end
                end
              for (forvar1291 = (1'h0); (forvar1291 < (2'h2)); forvar1291 = (forvar1291 + (1'h1)))
                begin
                  for (forvar1292 = (1'h0); (forvar1292 < (1'h0)); forvar1292 = (forvar1292 + (1'h1)))
                    begin
                      reg1293 <= forvar1129;
                      reg1294 <= reg1060;
                      reg1295 <= {$signed($signed(((8'haa) && forvar1095)))};
                    end
                  for (forvar1296 = (1'h0); (forvar1296 < (2'h2)); forvar1296 = (forvar1296 + (1'h1)))
                    begin
                      reg1297 <= (($signed(reg1133[(4'h8):(3'h4)]) ?
                          ($unsigned((8'ha3)) & (|forvar1181)) : reg1287) != (^$unsigned((^reg1171))));
                      reg1298 <= wire1042;
                      reg1299 <= reg1115[(2'h2):(1'h0)];
                      reg1300 <= {(+forvar1088)};
                    end
                  if (reg1231)
                    begin
                      reg1301 <= (forvar1088[(3'h7):(1'h1)] ?
                          $signed((8'h9f)) : reg1225);
                      reg1302 <= reg1078;
                      reg1303 <= (8'ha7);
                      reg1304 <= $signed((^~{reg1070}));
                    end
                  else
                    begin
                      reg1301 <= ($signed(reg1289[(1'h0):(1'h0)]) ?
                          $unsigned((((8'ha7) ?
                              reg1238 : forvar1079) | reg1260[(2'h2):(1'h0)])) : $signed(forvar1263[(3'h5):(1'h0)]));
                    end
                end
              if ($signed((~|{{reg1200}})))
                begin
                  reg1305 <= ((reg1205[(4'h9):(4'h8)] ?
                      $signed((forvar1244 != reg1202)) : (!$signed(reg1255))) - $unsigned($unsigned(reg1212)));
                  for (forvar1306 = (1'h0); (forvar1306 < (2'h2)); forvar1306 = (forvar1306 + (1'h1)))
                    begin
                      reg1307 <= (((~(forvar1169 ?
                              reg1277 : forvar1280)) >= (reg1175 > $signed(reg1113))) ?
                          reg1086[(3'h5):(3'h4)] : $unsigned(($signed(reg1223) ?
                              forvar1077 : reg1113)));
                      reg1308 <= (($signed($signed(reg1262)) | $unsigned($unsigned((8'ha4)))) ?
                          ((((8'ha2) ?
                                  reg1204 : reg1250) >> forvar1170[(3'h4):(1'h1)]) ?
                              reg1152 : (8'hba)) : forvar1158);
                    end
                end
              else
                begin
                  if (((|reg1072) ?
                      (forvar1244 ?
                          forvar1233[(2'h3):(2'h3)] : (&(!forvar1288))) : (({(8'hb6)} == forvar1154[(1'h0):(1'h0)]) ?
                          forvar1280[(3'h6):(3'h4)] : {(reg1091 ?
                                  reg1159 : reg1063)})))
                    begin
                      reg1305 <= $unsigned($signed(reg1214[(3'h6):(3'h6)]));
                    end
                  else
                    begin
                      reg1305 <= (reg1058 ^~ $unsigned({forvar1271[(1'h1):(1'h0)]}));
                      reg1306 <= (~&(~&$signed(reg1263[(1'h1):(1'h0)])));
                    end
                end
            end
          else
            begin
              if ((forvar1269 ?
                  $signed(reg1053[(2'h3):(2'h2)]) : ((~&(|reg1297)) + {(reg1209 ?
                          reg1133 : reg1153)})))
                begin
                  if ((((reg1205[(3'h7):(3'h4)] || (forvar1102 ?
                          reg1298 : (8'hab))) << $signed($unsigned(reg1273))) ?
                      reg1305[(2'h2):(1'h0)] : $unsigned($unsigned(reg1060))))
                    begin
                      reg1287 <= wire1044;
                      reg1288 <= $unsigned((|((reg1278 ?
                          reg1194 : reg1061) || ((8'hb9) >>> reg1192))));
                    end
                  else
                    begin
                      reg1287 <= $signed((reg1211[(2'h2):(2'h2)] ?
                          ((8'h9c) ?
                              reg1275 : (&(8'hb8))) : $signed((-(8'ha5)))));
                    end
                end
              else
                begin
                  for (forvar1287 = (1'h0); (forvar1287 < (2'h3)); forvar1287 = (forvar1287 + (1'h1)))
                    begin
                      reg1288 <= $signed(((reg1285[(1'h0):(1'h0)] ?
                          $unsigned(reg1181) : $signed(forvar1094)) ^ ({forvar1248} ?
                          forvar1206 : ((8'hb3) ? (8'had) : reg1190))));
                      reg1289 <= (!reg1116[(1'h1):(1'h1)]);
                    end
                end
              if (($signed((reg1242[(4'h8):(2'h3)] ?
                  $signed((8'h9d)) : $unsigned(reg1165))) - (!$unsigned(reg1250))))
                begin
                  for (forvar1290 = (1'h0); (forvar1290 < (2'h3)); forvar1290 = (forvar1290 + (1'h1)))
                    begin
                      reg1291 <= reg1060[(2'h3):(1'h1)];
                      reg1292 <= {(($signed(reg1072) ?
                              wire1042 : (^reg1308)) <<< (reg1100 <= (-reg1120)))};
                      reg1293 <= reg1286;
                      reg1294 <= $unsigned({reg1232[(4'h8):(2'h3)]});
                    end
                  if ($signed((|$signed((reg1110 > reg1187)))))
                    begin
                      reg1295 <= {forvar1273};
                      reg1296 <= reg1155;
                      reg1297 <= forvar1266[(2'h3):(2'h2)];
                      reg1298 <= $unsigned({$unsigned((reg1213 >> reg1149))});
                    end
                  else
                    begin
                      reg1295 <= ((reg1258 ^~ (~|(8'ha2))) ?
                          (8'hba) : (^(!$signed(forvar1188))));
                      reg1296 <= ((8'hab) * reg1091[(2'h2):(1'h0)]);
                    end
                end
              else
                begin
                  if ($signed(reg1090))
                    begin
                      reg1290 <= $signed((~^(reg1281[(4'ha):(4'h9)] ?
                          $unsigned(reg1073) : $signed(forvar1075))));
                      reg1291 <= ($signed($unsigned((~&reg1096))) ?
                          $signed(reg1279) : ({$signed(forvar1221)} ?
                              reg1080 : (^~forvar1130[(4'h9):(4'h8)])));
                    end
                  else
                    begin
                      reg1290 <= reg1237[(2'h2):(2'h2)];
                      reg1291 <= $signed(reg1285[(2'h2):(2'h2)]);
                    end
                  for (forvar1292 = (1'h0); (forvar1292 < (1'h1)); forvar1292 = (forvar1292 + (1'h1)))
                    begin
                      reg1293 <= $signed($unsigned($unsigned($unsigned((8'hac)))));
                      reg1294 <= (($unsigned($unsigned(reg1135)) || $unsigned($unsigned(reg1121))) ~^ {reg1188});
                      reg1295 <= (&forvar1163[(2'h3):(2'h2)]);
                    end
                end
            end
          for (forvar1309 = (1'h0); (forvar1309 < (2'h2)); forvar1309 = (forvar1309 + (1'h1)))
            begin
              if (reg1218)
                begin
                  reg1310 <= reg1300;
                  if ($signed((reg1295 ^~ $signed((reg1108 ?
                      forvar1077 : forvar1109)))))
                    begin
                      reg1311 <= reg1149;
                      reg1312 <= $unsigned(reg1108[(1'h1):(1'h0)]);
                      reg1313 <= ((($signed(reg1261) & (forvar1159 ?
                          (8'ha5) : forvar1146)) * ($unsigned(reg1069) ~^ reg1135[(3'h5):(1'h0)])) >= ((((8'ha4) ?
                              (8'ha4) : reg1083) & reg1099[(3'h7):(2'h3)]) ?
                          {reg1096} : ((~reg1118) > $signed(forvar1126))));
                      reg1314 <= $unsigned({(~forvar1130)});
                    end
                  else
                    begin
                      reg1311 <= $unsigned(($unsigned((forvar1109 ?
                          forvar1273 : (8'hb6))) - forvar1233));
                      reg1312 <= reg1107[(1'h1):(1'h0)];
                    end
                  for (forvar1315 = (1'h0); (forvar1315 < (2'h2)); forvar1315 = (forvar1315 + (1'h1)))
                    begin
                      reg1316 <= forvar1106[(4'ha):(3'h5)];
                      reg1317 <= $unsigned($unsigned($unsigned(((8'hb2) ?
                          reg1235 : reg1299))));
                      reg1318 <= reg1053;
                    end
                end
              else
                begin
                  reg1310 <= (reg1055[(4'ha):(3'h5)] ? forvar1277 : reg1096);
                  if ({reg1292[(3'h6):(3'h6)]})
                    begin
                      reg1311 <= {($signed(reg1064[(4'he):(4'h9)]) ?
                              (reg1144 ?
                                  $unsigned(reg1284) : (8'hae)) : {forvar1077})};
                    end
                  else
                    begin
                      reg1311 <= ($signed(reg1178) >>> $unsigned($signed((~^reg1065))));
                    end
                  reg1312 <= $unsigned(reg1062);
                end
              for (forvar1319 = (1'h0); (forvar1319 < (1'h0)); forvar1319 = (forvar1319 + (1'h1)))
                begin
                  for (forvar1320 = (1'h0); (forvar1320 < (2'h2)); forvar1320 = (forvar1320 + (1'h1)))
                    begin
                      reg1321 <= {reg1312[(3'h5):(2'h3)]};
                    end
                end
              if ((reg1083[(4'ha):(3'h6)] ?
                  (!$unsigned((+(8'hb2)))) : $signed((((8'h9e) ?
                      reg1251 : reg1127) < $signed(reg1122)))))
                begin
                  for (forvar1322 = (1'h0); (forvar1322 < (1'h0)); forvar1322 = (forvar1322 + (1'h1)))
                    begin
                      reg1323 <= (reg1107 ^ reg1124);
                    end
                  reg1324 <= forvar1074;
                end
              else
                begin
                  reg1322 <= reg1170[(3'h6):(3'h5)];
                  for (forvar1323 = (1'h0); (forvar1323 < (2'h3)); forvar1323 = (forvar1323 + (1'h1)))
                    begin
                      reg1324 <= (reg1305[(1'h0):(1'h0)] <<< $unsigned((reg1273[(1'h1):(1'h1)] ?
                          $signed(reg1239) : $unsigned(reg1282))));
                      reg1325 <= $signed(reg1293);
                      reg1326 <= (&($signed((|reg1156)) ? (8'hb2) : (8'hb6)));
                    end
                  for (forvar1327 = (1'h0); (forvar1327 < (2'h3)); forvar1327 = (forvar1327 + (1'h1)))
                    begin
                      reg1328 <= reg1072[(3'h6):(1'h1)];
                    end
                end
              for (forvar1329 = (1'h0); (forvar1329 < (1'h0)); forvar1329 = (forvar1329 + (1'h1)))
                begin
                  if ($signed({($signed(forvar1246) ^ reg1122[(4'hc):(4'h8)])}))
                    begin
                      reg1330 <= reg1241[(4'hb):(2'h3)];
                      reg1331 <= $signed({((~^reg1087) ?
                              {(8'hb1)} : $unsigned(forvar1128))});
                      reg1332 <= {(|{reg1271})};
                    end
                  else
                    begin
                      reg1330 <= {(((forvar1079 ~^ reg1194) || (reg1237 * reg1313)) ?
                              reg1284 : {(forvar1075 << reg1230)})};
                      reg1331 <= ((+reg1232[(3'h7):(1'h1)]) >> $unsigned((reg1070[(1'h0):(1'h0)] == forvar1156)));
                      reg1332 <= ((&{reg1288[(3'h5):(1'h1)]}) ?
                          {reg1252} : reg1131);
                      reg1333 <= {((forvar1235[(2'h2):(1'h1)] ?
                                  $signed(reg1301) : reg1301[(5'h10):(5'h10)]) ?
                              $signed(reg1169[(2'h2):(2'h2)]) : $signed((+forvar1074)))};
                    end
                end
            end
        end
      for (forvar1334 = (1'h0); (forvar1334 < (2'h2)); forvar1334 = (forvar1334 + (1'h1)))
        begin
          if ((forvar1273 ?
              reg1255[(2'h2):(1'h0)] : (((~reg1226) ?
                  (reg1330 <<< forvar1296) : {reg1188}) < ((reg1090 <= reg1055) ?
                  $unsigned(reg1274) : (reg1274 ? reg1168 : forvar1165)))))
            begin
              if ((reg1204 ?
                  $signed($unsigned((^reg1326))) : (reg1184[(1'h1):(1'h1)] ?
                      $signed((forvar1137 ?
                          reg1187 : reg1124)) : $signed((forvar1168 ?
                          reg1229 : reg1273)))))
                begin
                  for (forvar1335 = (1'h0); (forvar1335 < (2'h2)); forvar1335 = (forvar1335 + (1'h1)))
                    begin
                      reg1336 <= $signed($signed(($signed((8'hb5)) ~^ $signed((8'hb4)))));
                      reg1337 <= ($unsigned(forvar1224) ?
                          reg1159 : forvar1254[(2'h3):(1'h0)]);
                      reg1338 <= ((((~reg1333) <<< $unsigned(reg1328)) ?
                              (^reg1215[(4'hd):(1'h0)]) : {reg1252[(1'h1):(1'h1)]}) ?
                          reg1086[(4'h9):(3'h7)] : (^~((-reg1186) ?
                              (+forvar1309) : reg1190)));
                      reg1339 <= $signed({({reg1051} ?
                              (reg1154 ?
                                  (8'ha8) : wire1045) : (forvar1049 * (8'ha6)))});
                    end
                end
              else
                begin
                  reg1335 <= forvar1061;
                end
              if (({(reg1176[(3'h7):(1'h1)] > (reg1066 >= forvar1188))} != (reg1104[(1'h0):(1'h0)] & $unsigned(reg1171))))
                begin
                  for (forvar1340 = (1'h0); (forvar1340 < (1'h1)); forvar1340 = (forvar1340 + (1'h1)))
                    begin
                      reg1341 <= $signed(({reg1280} | reg1322));
                      reg1342 <= $signed(($signed((~&reg1267)) ?
                          (forvar1233 ?
                              (wire1043 ?
                                  reg1292 : forvar1163) : (~^reg1101)) : reg1323[(4'he):(3'h4)]));
                      reg1343 <= $unsigned($unsigned(forvar1128[(3'h7):(3'h7)]));
                    end
                  for (forvar1344 = (1'h0); (forvar1344 < (1'h1)); forvar1344 = (forvar1344 + (1'h1)))
                    begin
                      reg1345 <= forvar1334[(2'h2):(1'h1)];
                      reg1346 <= (((reg1136[(3'h4):(2'h3)] == ((8'ha7) >>> reg1128)) ?
                              forvar1083[(2'h2):(1'h1)] : reg1161[(1'h1):(1'h0)]) ?
                          (|((^reg1082) & reg1185[(1'h0):(1'h0)])) : ((8'hb5) ?
                              (^~$signed(reg1204)) : forvar1203));
                    end
                  if (reg1197[(4'hb):(3'h7)])
                    begin
                      reg1347 <= (+reg1087[(4'h8):(3'h7)]);
                    end
                  else
                    begin
                      reg1347 <= reg1346;
                      reg1348 <= (~^forvar1117);
                      reg1349 <= forvar1259;
                    end
                  if ($unsigned((~^reg1271[(2'h2):(1'h1)])))
                    begin
                      reg1350 <= forvar1260[(2'h2):(1'h0)];
                      reg1351 <= ($unsigned(reg1347[(2'h2):(1'h0)]) <= $signed((!reg1240)));
                    end
                  else
                    begin
                      reg1350 <= ({$signed($signed(reg1342))} & $unsigned($signed({reg1116})));
                      reg1351 <= ((reg1067 + $signed(reg1219)) ?
                          reg1073 : $signed($signed({reg1161})));
                    end
                end
              else
                begin
                  for (forvar1340 = (1'h0); (forvar1340 < (2'h3)); forvar1340 = (forvar1340 + (1'h1)))
                    begin
                      reg1341 <= $unsigned((^$unsigned(reg1304)));
                      reg1342 <= ((reg1113[(4'hd):(3'h6)] ?
                              forvar1147 : $signed({forvar1174})) ?
                          $signed(forvar1221) : (~|($unsigned((8'h9d)) ?
                              forvar1174 : (reg1093 ? (8'ha3) : reg1145))));
                      reg1343 <= reg1192[(3'h4):(2'h3)];
                    end
                  if ($signed((($signed(reg1261) ?
                          (~&reg1333) : $signed(wire1045)) ?
                      reg1164 : reg1282)))
                    begin
                      reg1344 <= forvar1142;
                      reg1345 <= reg1096;
                      reg1346 <= reg1124[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg1344 <= $signed((reg1068[(2'h3):(2'h3)] ?
                          $signed($unsigned(reg1276)) : forvar1204[(1'h0):(1'h0)]));
                      reg1345 <= ($unsigned(($unsigned(reg1086) ?
                          {reg1230} : {reg1085})) + $unsigned(reg1187[(2'h3):(1'h1)]));
                      reg1346 <= (((&reg1134[(3'h6):(3'h6)]) ^ $unsigned({wire1045})) ?
                          $signed((reg1252 + forvar1117[(3'h7):(3'h7)])) : ($signed((8'hb8)) ?
                              ((&reg1197) ?
                                  forvar1327[(1'h1):(1'h1)] : reg1130) : $unsigned(reg1223)));
                    end
                end
              reg1352 <= forvar1119[(4'hc):(4'h8)];
              if (forvar1137[(2'h2):(1'h1)])
                begin
                  for (forvar1353 = (1'h0); (forvar1353 < (1'h0)); forvar1353 = (forvar1353 + (1'h1)))
                    begin
                      reg1354 <= $unsigned(reg1214[(3'h7):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar1353 = (1'h0); (forvar1353 < (1'h1)); forvar1353 = (forvar1353 + (1'h1)))
                    begin
                      reg1354 <= $signed($unsigned(forvar1188[(4'hc):(3'h5)]));
                      reg1355 <= (reg1290[(2'h3):(1'h1)] ^ $signed(forvar1102[(1'h1):(1'h1)]));
                    end
                  for (forvar1356 = (1'h0); (forvar1356 < (1'h1)); forvar1356 = (forvar1356 + (1'h1)))
                    begin
                      reg1357 <= ($signed($signed(reg1104[(4'h8):(1'h1)])) ?
                          reg1126 : ((8'hb1) ^~ wire1043[(3'h4):(1'h0)]));
                      reg1358 <= ((reg1066[(3'h4):(2'h3)] ?
                              reg1335 : $signed((reg1080 ^ (8'hb6)))) ?
                          {forvar1287[(1'h0):(1'h0)]} : (~&reg1093));
                    end
                  for (forvar1359 = (1'h0); (forvar1359 < (2'h2)); forvar1359 = (forvar1359 + (1'h1)))
                    begin
                      reg1360 <= forvar1126[(3'h5):(1'h1)];
                      reg1361 <= {$signed((~forvar1315))};
                    end
                  for (forvar1362 = (1'h0); (forvar1362 < (2'h2)); forvar1362 = (forvar1362 + (1'h1)))
                    begin
                      reg1363 <= (~^reg1081);
                      reg1364 <= $signed(reg1143);
                      reg1365 <= forvar1048[(3'h7):(3'h6)];
                      reg1366 <= ($signed({$unsigned(forvar1156)}) | reg1119);
                    end
                end
            end
          else
            begin
              if ($signed({$unsigned(reg1177[(2'h2):(2'h2)])}))
                begin
                  reg1335 <= ($unsigned($unsigned((^~forvar1290))) ?
                      {reg1251} : ($signed($unsigned(forvar1188)) ^ (forvar1188[(2'h3):(1'h0)] | reg1181[(1'h0):(1'h0)])));
                  for (forvar1336 = (1'h0); (forvar1336 < (1'h1)); forvar1336 = (forvar1336 + (1'h1)))
                    begin
                      reg1337 <= ((reg1322[(4'h9):(4'h8)] ?
                              $unsigned($signed((8'ha1))) : $signed((8'ha9))) ?
                          $signed(((~&(8'h9f)) ?
                              ((8'hb8) ?
                                  forvar1216 : forvar1048) : $signed(forvar1109))) : $unsigned(reg1213));
                      reg1338 <= $signed({$unsigned((forvar1173 != forvar1102))});
                    end
                end
              else
                begin
                  for (forvar1335 = (1'h0); (forvar1335 < (1'h1)); forvar1335 = (forvar1335 + (1'h1)))
                    begin
                      reg1336 <= (reg1168 ?
                          reg1128[(5'h10):(4'h8)] : ((~^(reg1181 ?
                                  (8'hb3) : forvar1175)) ?
                              (~$signed((8'h9c))) : (|(^forvar1061))));
                      reg1337 <= $unsigned(reg1253[(3'h5):(3'h4)]);
                    end
                  reg1338 <= {(reg1164 ?
                          ({reg1245} ?
                              $unsigned(reg1057) : reg1128[(2'h3):(1'h1)]) : (^~$signed(forvar1137)))};
                  reg1339 <= reg1209[(2'h3):(2'h3)];
                  if ($unsigned($signed(forvar1329[(2'h2):(1'h1)])))
                    begin
                      reg1340 <= $signed($unsigned(({reg1076} <= $unsigned(reg1092))));
                    end
                  else
                    begin
                      reg1340 <= $signed($signed($unsigned($unsigned((8'ha1)))));
                      reg1341 <= ((^reg1189[(1'h1):(1'h1)]) << ($unsigned({reg1323}) && reg1063));
                      reg1342 <= $unsigned((-reg1168[(2'h2):(1'h1)]));
                    end
                end
            end
        end
      for (forvar1367 = (1'h0); (forvar1367 < (2'h3)); forvar1367 = (forvar1367 + (1'h1)))
        begin
          for (forvar1368 = (1'h0); (forvar1368 < (1'h1)); forvar1368 = (forvar1368 + (1'h1)))
            begin
              for (forvar1369 = (1'h0); (forvar1369 < (1'h1)); forvar1369 = (forvar1369 + (1'h1)))
                begin
                  for (forvar1370 = (1'h0); (forvar1370 < (1'h1)); forvar1370 = (forvar1370 + (1'h1)))
                    begin
                      reg1371 <= $signed(((reg1255[(2'h3):(2'h3)] * forvar1170) >>> $unsigned((|forvar1367))));
                      reg1372 <= ($unsigned($signed((reg1114 ?
                          forvar1159 : (8'hb3)))) * ($unsigned((reg1365 ?
                          forvar1322 : (8'hb8))) < ({forvar1370} << ((8'hb6) ?
                          reg1060 : reg1357))));
                      reg1373 <= $signed($unsigned(($unsigned(reg1357) <= (reg1293 <<< forvar1160))));
                      reg1374 <= ((reg1331 ?
                          $signed($signed(reg1330)) : (^(forvar1146 ?
                              reg1366 : forvar1288))) != ($unsigned(((8'h9e) <= reg1338)) ?
                          (^~$signed(reg1281)) : ((&reg1209) ?
                              $signed(reg1090) : (+reg1078))));
                    end
                  for (forvar1375 = (1'h0); (forvar1375 < (2'h3)); forvar1375 = (forvar1375 + (1'h1)))
                    begin
                      reg1376 <= forvar1208;
                    end
                  if ((reg1311[(3'h5):(2'h2)] ?
                      ({(^reg1139)} ^~ (+$unsigned(reg1301))) : ({reg1113[(4'ha):(4'ha)]} ?
                          ($signed(forvar1275) ^~ reg1317[(3'h6):(1'h0)]) : reg1249)))
                    begin
                      reg1377 <= ((((!reg1225) ? (8'ha3) : $unsigned(reg1124)) ?
                          $signed($signed(reg1234)) : ({forvar1266} ?
                              $signed(forvar1088) : (reg1291 ?
                                  forvar1203 : reg1256))) ^ $unsigned(reg1053[(4'h8):(1'h1)]));
                      reg1378 <= (-reg1287[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1377 <= (~&$signed($signed(reg1283)));
                    end
                end
              if (reg1165[(1'h1):(1'h0)])
                begin
                  reg1379 <= forvar1160[(4'ha):(1'h1)];
                  reg1380 <= {(($signed(reg1119) <= $signed((8'h9e))) ?
                          reg1321 : $unsigned((^(8'hb8))))};
                  if ($signed($unsigned(($signed(forvar1362) ?
                      $signed(forvar1048) : (forvar1287 ?
                          forvar1120 : reg1089)))))
                    begin
                      reg1381 <= reg1212[(2'h3):(2'h2)];
                      reg1382 <= ((~&forvar1292) ?
                          forvar1156 : ((~|forvar1094[(4'h9):(3'h5)]) < (|$signed(reg1196))));
                      reg1383 <= reg1125[(4'h9):(3'h7)];
                    end
                  else
                    begin
                      reg1381 <= (~|forvar1212);
                      reg1382 <= (($signed($unsigned(reg1057)) <<< (^((8'ha4) ?
                              reg1234 : reg1061))) ?
                          $unsigned($unsigned(reg1112[(1'h1):(1'h0)])) : ($unsigned($signed((8'ha8))) * forvar1362));
                      reg1383 <= ($signed(($signed(reg1082) ?
                              forvar1175[(1'h1):(1'h1)] : reg1084)) ?
                          forvar1175 : $unsigned((8'ha0)));
                      reg1384 <= $signed(reg1289);
                    end
                end
              else
                begin
                  if ($unsigned(forvar1146))
                    begin
                      reg1379 <= forvar1296[(4'h9):(4'h8)];
                      reg1380 <= ((~|reg1299) ?
                          forvar1228 : ((|$signed((8'h9e))) | ($unsigned(reg1177) ?
                              forvar1160[(2'h3):(1'h1)] : (reg1236 >> reg1328))));
                    end
                  else
                    begin
                      reg1379 <= ((forvar1098 ?
                          reg1207[(4'h8):(3'h4)] : $unsigned((reg1358 >> reg1239))) ^~ (forvar1154[(2'h2):(1'h0)] && reg1141[(4'hb):(2'h3)]));
                    end
                  reg1381 <= reg1372;
                  reg1382 <= reg1218[(2'h3):(2'h3)];
                end
              for (forvar1385 = (1'h0); (forvar1385 < (1'h0)); forvar1385 = (forvar1385 + (1'h1)))
                begin
                  for (forvar1386 = (1'h0); (forvar1386 < (1'h1)); forvar1386 = (forvar1386 + (1'h1)))
                    begin
                      reg1387 <= ($unsigned(($unsigned(forvar1260) != $unsigned(forvar1259))) || ($signed({reg1230}) ?
                          $signed($signed(reg1291)) : (forvar1367[(2'h3):(1'h1)] >= $signed((8'hb9)))));
                    end
                  if ((reg1215[(3'h6):(1'h0)] <= reg1258))
                    begin
                      reg1388 <= forvar1340;
                      reg1389 <= reg1086[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg1388 <= forvar1129;
                      reg1389 <= reg1295;
                    end
                  for (forvar1390 = (1'h0); (forvar1390 < (2'h3)); forvar1390 = (forvar1390 + (1'h1)))
                    begin
                      reg1391 <= (~|(reg1266 ?
                          {$unsigned(reg1120)} : (&$signed(reg1217))));
                    end
                  for (forvar1392 = (1'h0); (forvar1392 < (1'h1)); forvar1392 = (forvar1392 + (1'h1)))
                    begin
                      reg1393 <= (~^reg1231);
                    end
                end
              reg1394 <= reg1324;
            end
          for (forvar1395 = (1'h0); (forvar1395 < (2'h3)); forvar1395 = (forvar1395 + (1'h1)))
            begin
              if (reg1200[(4'hc):(3'h7)])
                begin
                  for (forvar1396 = (1'h0); (forvar1396 < (2'h2)); forvar1396 = (forvar1396 + (1'h1)))
                    begin
                      reg1397 <= forvar1276[(2'h2):(1'h1)];
                      reg1398 <= ((~|$unsigned((reg1241 ?
                              forvar1368 : reg1354))) ?
                          $unsigned(forvar1165[(4'h8):(1'h0)]) : forvar1174);
                      reg1399 <= (8'ha7);
                    end
                  if (reg1204[(1'h1):(1'h1)])
                    begin
                      reg1400 <= forvar1362[(2'h3):(1'h1)];
                      reg1401 <= (reg1242 & {(+(reg1184 ^~ forvar1098))});
                      reg1402 <= (&$unsigned($signed((~|reg1394))));
                    end
                  else
                    begin
                      reg1400 <= {$unsigned({(+reg1233)})};
                      reg1401 <= (forvar1359[(3'h4):(2'h3)] ?
                          $unsigned(($unsigned((8'hac)) ?
                              (-reg1052) : (~reg1380))) : $signed($signed(reg1350[(4'h8):(3'h4)])));
                      reg1402 <= reg1119[(2'h2):(1'h1)];
                    end
                  reg1403 <= (forvar1228[(4'he):(3'h7)] >> $unsigned(reg1345));
                end
              else
                begin
                  reg1396 <= (~^reg1169);
                  for (forvar1397 = (1'h0); (forvar1397 < (2'h3)); forvar1397 = (forvar1397 + (1'h1)))
                    begin
                      reg1398 <= (^~(|$unsigned((!reg1363))));
                      reg1399 <= (+(reg1398[(1'h0):(1'h0)] <= forvar1048));
                      reg1400 <= reg1312[(4'hd):(4'hb)];
                    end
                  if ($unsigned($signed(((8'hb9) ?
                      $signed(forvar1273) : (forvar1119 ? reg1277 : (8'hb3))))))
                    begin
                      reg1401 <= (forvar1224 ^ $unsigned($signed((~forvar1142))));
                      reg1402 <= (-$signed({(reg1207 ? forvar1235 : reg1233)}));
                      reg1403 <= {(&forvar1336[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg1401 <= reg1220;
                    end
                  if ({reg1081})
                    begin
                      reg1404 <= {{$signed(reg1399)}};
                    end
                  else
                    begin
                      reg1404 <= forvar1170;
                      reg1405 <= ((|$signed({(8'haf)})) ?
                          {(~&(reg1050 <<< reg1245))} : reg1256[(4'hc):(1'h1)]);
                      reg1406 <= $unsigned((~&$unsigned(reg1387[(4'h9):(4'h8)])));
                    end
                end
              if ({$signed(((reg1282 ? reg1091 : reg1132) ?
                      forvar1212[(3'h5):(3'h5)] : (!reg1378)))})
                begin
                  for (forvar1407 = (1'h0); (forvar1407 < (2'h3)); forvar1407 = (forvar1407 + (1'h1)))
                    begin
                      reg1408 <= wire1042;
                      reg1409 <= {(forvar1309 <= (^~reg1396))};
                      reg1410 <= forvar1047;
                    end
                  reg1411 <= reg1396;
                end
              else
                begin
                  reg1407 <= $signed(reg1060[(2'h3):(2'h2)]);
                end
              if ({((+$unsigned(wire1042)) ~^ ((forvar1142 || (8'hab)) ?
                      (reg1138 < reg1264) : (reg1112 ^ reg1136)))})
                begin
                  for (forvar1412 = (1'h0); (forvar1412 < (1'h0)); forvar1412 = (forvar1412 + (1'h1)))
                    begin
                      reg1413 <= ((|{$signed(reg1184)}) ?
                          (^~$signed(forvar1269)) : $unsigned($unsigned($signed(reg1209))));
                      reg1414 <= (forvar1263[(1'h1):(1'h0)] >>> forvar1183);
                    end
                  for (forvar1415 = (1'h0); (forvar1415 < (1'h1)); forvar1415 = (forvar1415 + (1'h1)))
                    begin
                      reg1416 <= (&(^~(8'ha1)));
                      reg1417 <= $unsigned(forvar1170[(1'h0):(1'h0)]);
                      reg1418 <= $signed((8'hb8));
                    end
                  for (forvar1419 = (1'h0); (forvar1419 < (1'h0)); forvar1419 = (forvar1419 + (1'h1)))
                    begin
                      reg1420 <= forvar1329;
                    end
                  for (forvar1421 = (1'h0); (forvar1421 < (2'h2)); forvar1421 = (forvar1421 + (1'h1)))
                    begin
                      reg1422 <= ($unsigned(((reg1303 - reg1226) ?
                          reg1191[(1'h1):(1'h0)] : (reg1135 ?
                              (8'h9f) : reg1134))) < $unsigned(((|reg1382) ?
                          (^~forvar1320) : reg1282[(1'h1):(1'h0)])));
                    end
                end
              else
                begin
                  if ((({(~^reg1241)} ?
                          (reg1287 ^~ reg1314) : ((reg1154 ?
                              reg1201 : reg1171) != reg1131)) ?
                      (+($signed(reg1168) ?
                          $signed(reg1323) : reg1402[(4'hd):(4'hd)])) : (($signed((8'ha6)) ?
                              reg1377 : $signed(reg1055)) ?
                          ((|(8'hb1)) & (^~reg1286)) : reg1101[(4'hb):(1'h0)])))
                    begin
                      reg1412 <= reg1220[(2'h3):(1'h0)];
                      reg1413 <= $signed((~^reg1235[(3'h6):(1'h1)]));
                      reg1414 <= (+($signed((forvar1386 > reg1235)) ?
                          $unsigned(forvar1315) : $signed((reg1188 && reg1091))));
                    end
                  else
                    begin
                      reg1412 <= $unsigned((!reg1412));
                      reg1413 <= ((~^((forvar1079 << reg1177) ?
                          forvar1280[(4'he):(3'h7)] : (reg1121 && (8'ha4)))) & reg1188);
                      reg1414 <= reg1226;
                      reg1415 <= (|($unsigned(reg1133[(4'ha):(4'h8)]) | ($signed(reg1107) ?
                          (-reg1105) : (+reg1227))));
                    end
                end
            end
        end
    end
  assign wire1423 = {{forvar1386[(3'h4):(3'h4)]}};
  always
    @(posedge clk) begin
      reg1424 <= ((8'hb0) >= $signed($unsigned({reg1240})));
      for (forvar1425 = (1'h0); (forvar1425 < (2'h2)); forvar1425 = (forvar1425 + (1'h1)))
        begin
          if ($unsigned(((~|$unsigned(reg1068)) >= reg1062)))
            begin
              if ($signed($signed(((reg1384 ? (8'hb9) : forvar1130) ?
                  reg1057 : $signed((8'ha7))))))
                begin
                  for (forvar1426 = (1'h0); (forvar1426 < (2'h3)); forvar1426 = (forvar1426 + (1'h1)))
                    begin
                      reg1427 <= (-((8'hac) ?
                          (reg1252 >> (~(8'ha0))) : forvar1216));
                      reg1428 <= (&$signed($signed($signed(reg1223))));
                      reg1429 <= ((~&((8'h9c) == {reg1247})) - $unsigned($signed((forvar1169 ?
                          forvar1244 : forvar1415))));
                    end
                  if ({(reg1234[(2'h3):(2'h2)] ~^ forvar1233[(1'h0):(1'h0)])})
                    begin
                      reg1430 <= reg1186[(4'he):(3'h4)];
                      reg1431 <= {$signed($unsigned((forvar1273 < (8'ha2))))};
                      reg1432 <= reg1239;
                      reg1433 <= ({$signed($signed(forvar1085))} ?
                          {(reg1346[(4'hf):(3'h6)] | reg1273)} : reg1318[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg1430 <= ((reg1232[(2'h3):(2'h2)] != (8'ha0)) >>> forvar1233[(4'h8):(1'h0)]);
                      reg1431 <= ($signed($unsigned($signed((8'h9e)))) + reg1223[(2'h2):(2'h2)]);
                    end
                end
              else
                begin
                  if (reg1296[(2'h3):(1'h0)])
                    begin
                      reg1426 <= ((8'ha8) ? reg1085 : reg1145);
                    end
                  else
                    begin
                      reg1426 <= reg1411;
                      reg1427 <= {((+$signed(forvar1340)) ?
                              ((reg1170 <<< (8'ha2)) ?
                                  (reg1183 < reg1230) : forvar1228) : (((8'ha6) ?
                                      (8'haa) : reg1159) ?
                                  $signed((8'ha4)) : ((8'hb3) && reg1384)))};
                    end
                  reg1428 <= (|$signed(((~^(8'hb9)) >> (forvar1306 ?
                      reg1431 : reg1345))));
                  if ({($signed((reg1342 ?
                          reg1402 : forvar1344)) ^~ (&$unsigned(forvar1375)))})
                    begin
                      reg1429 <= $signed(forvar1386);
                      reg1430 <= (~|reg1180[(3'h6):(1'h0)]);
                      reg1431 <= reg1202[(2'h2):(2'h2)];
                      reg1432 <= ((reg1433 << forvar1425) ?
                          $unsigned(reg1060) : (|({reg1138} ?
                              $signed(forvar1320) : $signed(reg1058))));
                    end
                  else
                    begin
                      reg1429 <= forvar1273[(4'he):(4'hb)];
                      reg1430 <= $unsigned(reg1150);
                      reg1431 <= reg1233[(1'h1):(1'h1)];
                    end
                  for (forvar1433 = (1'h0); (forvar1433 < (1'h0)); forvar1433 = (forvar1433 + (1'h1)))
                    begin
                      reg1434 <= $signed(reg1355[(1'h0):(1'h0)]);
                      reg1435 <= ((8'hb6) || (-reg1432[(1'h1):(1'h0)]));
                      reg1436 <= reg1376[(1'h1):(1'h0)];
                      reg1437 <= ($signed(reg1136) >>> forvar1129[(1'h1):(1'h0)]);
                    end
                end
              reg1438 <= (&($unsigned(reg1065[(3'h6):(1'h1)]) ?
                  (~|$unsigned(reg1153)) : (reg1332 && (~|forvar1117))));
              for (forvar1439 = (1'h0); (forvar1439 < (1'h1)); forvar1439 = (forvar1439 + (1'h1)))
                begin
                  for (forvar1440 = (1'h0); (forvar1440 < (1'h1)); forvar1440 = (forvar1440 + (1'h1)))
                    begin
                      reg1441 <= $signed(($unsigned(reg1124) ?
                          (forvar1188 <= forvar1216) : $signed($unsigned(reg1414))));
                      reg1442 <= {(reg1172[(2'h3):(1'h0)] > $unsigned(reg1250[(4'hd):(4'h8)]))};
                    end
                  for (forvar1443 = (1'h0); (forvar1443 < (1'h0)); forvar1443 = (forvar1443 + (1'h1)))
                    begin
                      reg1444 <= (((~$unsigned(reg1291)) ?
                              (~^reg1207[(3'h6):(2'h3)]) : reg1195[(1'h1):(1'h1)]) ?
                          reg1349 : (~|$signed((forvar1159 * forvar1329))));
                      reg1445 <= ((((~reg1251) ?
                              $signed((8'h9f)) : reg1267[(3'h5):(1'h1)]) ^ reg1115) ?
                          ($unsigned($signed(reg1281)) >= {reg1335[(2'h2):(1'h0)]}) : $unsigned({$unsigned(reg1183)}));
                      reg1446 <= reg1212;
                      reg1447 <= forvar1269;
                    end
                  for (forvar1448 = (1'h0); (forvar1448 < (2'h2)); forvar1448 = (forvar1448 + (1'h1)))
                    begin
                      reg1449 <= (reg1442[(3'h4):(1'h1)] ?
                          $signed((reg1398[(3'h6):(1'h1)] >>> reg1377)) : $unsigned((reg1231 & (reg1444 != forvar1169))));
                      reg1450 <= reg1347[(2'h3):(1'h0)];
                      reg1451 <= ($unsigned(reg1092[(4'he):(1'h1)]) + reg1379);
                      reg1452 <= (^reg1213[(2'h2):(1'h1)]);
                    end
                end
              for (forvar1453 = (1'h0); (forvar1453 < (2'h3)); forvar1453 = (forvar1453 + (1'h1)))
                begin
                  reg1454 <= wire1043;
                end
            end
          else
            begin
              if (forvar1061[(4'h9):(2'h3)])
                begin
                  for (forvar1426 = (1'h0); (forvar1426 < (2'h2)); forvar1426 = (forvar1426 + (1'h1)))
                    begin
                      reg1427 <= {reg1124[(4'h8):(1'h1)]};
                      reg1428 <= (($unsigned((&(8'hb7))) ?
                              (reg1417[(3'h5):(1'h1)] ?
                                  (^reg1164) : (~&forvar1147)) : ((|reg1168) && (reg1404 ?
                                  forvar1315 : reg1053))) ?
                          {(^$signed(wire1044))} : $signed($unsigned((wire1042 ?
                              reg1446 : (8'h9d)))));
                    end
                  for (forvar1429 = (1'h0); (forvar1429 < (1'h0)); forvar1429 = (forvar1429 + (1'h1)))
                    begin
                      reg1430 <= ($unsigned((~^$signed(reg1125))) - $unsigned($signed(((8'hb2) << reg1120))));
                      reg1431 <= (+reg1159[(2'h2):(2'h2)]);
                      reg1432 <= ($unsigned($signed($signed(forvar1216))) ?
                          $signed($unsigned(reg1230[(3'h7):(1'h0)])) : (-forvar1233[(2'h3):(2'h2)]));
                    end
                  for (forvar1433 = (1'h0); (forvar1433 < (2'h3)); forvar1433 = (forvar1433 + (1'h1)))
                    begin
                      reg1434 <= $signed((!({forvar1098} ?
                          (-reg1285) : (forvar1439 ? reg1363 : reg1153))));
                      reg1435 <= $signed(((reg1428[(4'h9):(2'h2)] ^~ (forvar1061 < reg1377)) ?
                          $signed($signed((8'h9d))) : {(~^reg1072)}));
                    end
                end
              else
                begin
                  if ((~&({forvar1238} ?
                      ((forvar1114 ?
                          forvar1142 : reg1435) * (forvar1263 >= reg1433)) : $unsigned((reg1444 || reg1255)))))
                    begin
                      reg1426 <= (forvar1181[(4'h9):(1'h0)] - $unsigned(($signed(reg1100) ?
                          $unsigned(forvar1221) : (!reg1323))));
                    end
                  else
                    begin
                      reg1426 <= $signed($signed(((reg1374 >>> forvar1320) ?
                          {(8'ha4)} : forvar1233[(2'h2):(2'h2)])));
                      reg1427 <= (~&$unsigned($unsigned((~^reg1300))));
                    end
                end
              for (forvar1436 = (1'h0); (forvar1436 < (1'h0)); forvar1436 = (forvar1436 + (1'h1)))
                begin
                  for (forvar1437 = (1'h0); (forvar1437 < (1'h1)); forvar1437 = (forvar1437 + (1'h1)))
                    begin
                      reg1438 <= $signed((~reg1280));
                      reg1439 <= {((~(^reg1259)) <= forvar1208[(2'h2):(1'h1)])};
                    end
                  if ($signed(reg1435[(3'h4):(2'h2)]))
                    begin
                      reg1440 <= $unsigned((~^(|$signed(forvar1120))));
                      reg1441 <= {$signed($signed((~|forvar1244)))};
                      reg1442 <= $unsigned($signed((~reg1261[(4'hc):(4'hb)])));
                    end
                  else
                    begin
                      reg1440 <= ($unsigned({$unsigned(reg1265)}) ?
                          reg1424 : (^~(8'hba)));
                      reg1441 <= reg1361[(1'h0):(1'h0)];
                    end
                  for (forvar1443 = (1'h0); (forvar1443 < (1'h1)); forvar1443 = (forvar1443 + (1'h1)))
                    begin
                      reg1444 <= {(8'hb2)};
                    end
                  reg1445 <= {(|$unsigned((reg1436 + reg1215)))};
                end
              for (forvar1446 = (1'h0); (forvar1446 < (1'h1)); forvar1446 = (forvar1446 + (1'h1)))
                begin
                  for (forvar1447 = (1'h0); (forvar1447 < (2'h2)); forvar1447 = (forvar1447 + (1'h1)))
                    begin
                      reg1448 <= ($signed($signed($signed(reg1059))) ?
                          reg1450[(2'h3):(2'h3)] : (reg1251[(3'h4):(2'h3)] == reg1093));
                    end
                  for (forvar1449 = (1'h0); (forvar1449 < (2'h2)); forvar1449 = (forvar1449 + (1'h1)))
                    begin
                      reg1450 <= reg1201[(1'h1):(1'h0)];
                      reg1451 <= $signed($unsigned($signed({reg1322})));
                    end
                  if (((forvar1336 ~^ ((reg1372 ~^ reg1258) ?
                      (reg1192 ?
                          reg1379 : forvar1271) : $unsigned(forvar1079))) >= reg1363))
                    begin
                      reg1452 <= ((forvar1160 == $signed(((8'ha0) == (8'hb5)))) ?
                          ((+reg1373) ?
                              reg1092[(4'hc):(3'h6)] : (^~$signed(forvar1094))) : forvar1259);
                      reg1453 <= (|(reg1212[(1'h0):(1'h0)] ~^ (~reg1322)));
                      reg1454 <= (~&(~&{reg1405}));
                    end
                  else
                    begin
                      reg1452 <= (reg1300 | $signed(($signed(reg1345) > $unsigned(reg1389))));
                      reg1453 <= $signed((~&$unsigned((-forvar1277))));
                      reg1454 <= (!(((~reg1222) < (reg1314 ?
                          reg1352 : reg1157)) != $unsigned(forvar1386)));
                    end
                  reg1455 <= forvar1183[(1'h0):(1'h0)];
                end
            end
          for (forvar1456 = (1'h0); (forvar1456 < (1'h0)); forvar1456 = (forvar1456 + (1'h1)))
            begin
              if ((~&(-(reg1424[(3'h7):(3'h4)] ?
                  $signed(reg1067) : $unsigned((8'ha6))))))
                begin
                  for (forvar1457 = (1'h0); (forvar1457 < (2'h2)); forvar1457 = (forvar1457 + (1'h1)))
                    begin
                      reg1458 <= $unsigned((8'hb2));
                      reg1459 <= ({(reg1255[(4'h8):(3'h4)] ?
                              {reg1342} : $signed(reg1179))} | $signed(reg1160));
                    end
                  reg1460 <= $unsigned(reg1387[(4'ha):(3'h5)]);
                  for (forvar1461 = (1'h0); (forvar1461 < (2'h2)); forvar1461 = (forvar1461 + (1'h1)))
                    begin
                      reg1462 <= (-reg1116);
                      reg1463 <= ((((reg1428 * reg1193) >>> $unsigned(reg1351)) ?
                          (~^{reg1189}) : (((8'hab) ? reg1158 : reg1281) ?
                              (forvar1075 - reg1080) : reg1152)) == forvar1277[(4'hf):(4'he)]);
                      reg1464 <= reg1403;
                    end
                  for (forvar1465 = (1'h0); (forvar1465 < (2'h3)); forvar1465 = (forvar1465 + (1'h1)))
                    begin
                      reg1466 <= ($signed($signed((~^reg1432))) ?
                          (-((reg1167 << (8'ha8)) <<< $unsigned(reg1214))) : ({{reg1104}} + ((|reg1326) ?
                              reg1180[(4'hb):(2'h2)] : $unsigned(forvar1177))));
                      reg1467 <= (~&forvar1368);
                    end
                end
              else
                begin
                  if ($unsigned({reg1289[(2'h2):(1'h1)]}))
                    begin
                      reg1457 <= $unsigned((^~forvar1448));
                    end
                  else
                    begin
                      reg1457 <= $unsigned(reg1160);
                      reg1458 <= (~|({{forvar1276}} ?
                          $signed($unsigned(reg1171)) : ((^~reg1381) | ((8'hab) + reg1405))));
                      reg1459 <= reg1188[(4'h8):(3'h7)];
                    end
                  for (forvar1460 = (1'h0); (forvar1460 < (2'h3)); forvar1460 = (forvar1460 + (1'h1)))
                    begin
                      reg1461 <= forvar1460[(1'h1):(1'h1)];
                      reg1462 <= $signed((reg1460 | reg1417));
                      reg1463 <= $signed($unsigned($unsigned($signed(forvar1175))));
                    end
                end
              if ((8'ha1))
                begin
                  for (forvar1468 = (1'h0); (forvar1468 < (1'h1)); forvar1468 = (forvar1468 + (1'h1)))
                    begin
                      reg1469 <= {$unsigned($signed(reg1203))};
                      reg1470 <= (8'h9c);
                      reg1471 <= $unsigned(($unsigned((reg1195 ?
                          reg1366 : forvar1340)) | ({reg1193} - (reg1270 ^~ reg1133))));
                      reg1472 <= ((^~$unsigned({(8'h9d)})) ?
                          $signed($signed(reg1234)) : (^$signed(reg1400[(1'h1):(1'h0)])));
                    end
                  reg1473 <= (~|forvar1370[(3'h5):(3'h5)]);
                  if (($signed($signed(reg1229)) + $signed($unsigned((reg1165 ?
                      reg1360 : (8'haf))))))
                    begin
                      reg1474 <= (^($unsigned($signed(reg1253)) ?
                          $unsigned({reg1278}) : forvar1259[(1'h0):(1'h0)]));
                      reg1475 <= (($signed((+forvar1156)) ?
                          (!reg1193[(1'h0):(1'h0)]) : (~^((8'ha5) ?
                              reg1174 : reg1454))) >= $signed((^~forvar1174[(3'h4):(2'h3)])));
                    end
                  else
                    begin
                      reg1474 <= reg1076[(3'h7):(3'h5)];
                      reg1475 <= (&($signed(reg1405) << $unsigned({wire1046})));
                      reg1476 <= {forvar1440[(1'h1):(1'h1)]};
                      reg1477 <= {{$signed((reg1377 ? reg1276 : forvar1154))}};
                    end
                end
              else
                begin
                  for (forvar1468 = (1'h0); (forvar1468 < (1'h1)); forvar1468 = (forvar1468 + (1'h1)))
                    begin
                      reg1469 <= ((^(!reg1475)) ?
                          (~|{forvar1159}) : forvar1457[(4'ha):(3'h7)]);
                      reg1470 <= $signed((((|forvar1079) & $unsigned(forvar1340)) ?
                          ($signed(forvar1065) ^~ (!reg1360)) : reg1245));
                    end
                  if (reg1244[(1'h1):(1'h1)])
                    begin
                      reg1471 <= reg1186[(4'hb):(2'h2)];
                      reg1472 <= $unsigned($signed($signed($signed(forvar1244))));
                    end
                  else
                    begin
                      reg1471 <= reg1341[(1'h1):(1'h0)];
                      reg1472 <= ((forvar1271 ?
                              reg1225 : ((reg1073 ? reg1289 : reg1101) ?
                                  $signed(reg1273) : ((8'hb3) ?
                                      reg1464 : reg1239))) ?
                          {forvar1221} : $signed($signed((reg1187 <<< forvar1465))));
                      reg1473 <= ($unsigned((~|(reg1267 >> reg1144))) ?
                          $signed($signed($signed((8'ha4)))) : reg1081);
                    end
                end
            end
        end
      for (forvar1478 = (1'h0); (forvar1478 < (2'h2)); forvar1478 = (forvar1478 + (1'h1)))
        begin
          if (reg1372)
            begin
              if (forvar1320[(4'hb):(3'h6)])
                begin
                  for (forvar1479 = (1'h0); (forvar1479 < (2'h2)); forvar1479 = (forvar1479 + (1'h1)))
                    begin
                      reg1480 <= {reg1172};
                      reg1481 <= $signed((((^reg1441) >>> $signed((8'hb2))) ?
                          ((^~reg1196) ?
                              $unsigned(reg1249) : (~|reg1063)) : $signed($signed(reg1207))));
                      reg1482 <= ({(reg1275 ~^ (-reg1372))} ?
                          ($unsigned(reg1400) ?
                              ((reg1422 >= reg1160) - (reg1432 >> forvar1137)) : reg1411[(1'h1):(1'h1)]) : $signed(((reg1066 ?
                                  forvar1437 : reg1175) ?
                              $signed(reg1103) : (reg1323 ?
                                  reg1164 : reg1279))));
                      reg1483 <= (forvar1266[(1'h0):(1'h0)] * (^((forvar1183 ?
                              forvar1419 : reg1476) ?
                          {reg1060} : forvar1415)));
                    end
                end
              else
                begin
                  reg1479 <= (forvar1296[(4'hd):(4'hb)] >= ($signed({(8'ha1)}) < forvar1109[(4'h9):(3'h7)]));
                end
              for (forvar1484 = (1'h0); (forvar1484 < (1'h1)); forvar1484 = (forvar1484 + (1'h1)))
                begin
                  if ((reg1399 - reg1154[(3'h4):(2'h3)]))
                    begin
                      reg1485 <= $signed(reg1420);
                      reg1486 <= $unsigned((((forvar1246 <= forvar1277) ?
                              $unsigned(forvar1117) : reg1138) ?
                          {(reg1373 ? forvar1461 : reg1292)} : reg1218));
                    end
                  else
                    begin
                      reg1485 <= {(|{(+(8'hb6))})};
                      reg1486 <= forvar1244;
                      reg1487 <= {{((^forvar1386) == $unsigned(forvar1147))}};
                    end
                  if (((~|(^~forvar1147)) < ((~$signed(reg1461)) ?
                      $unsigned(((8'ha0) <<< reg1293)) : reg1232)))
                    begin
                      reg1488 <= $signed($signed({forvar1291[(4'hb):(3'h5)]}));
                      reg1489 <= ((8'hb6) | forvar1412);
                      reg1490 <= $unsigned($unsigned($unsigned((~(8'h9f)))));
                    end
                  else
                    begin
                      reg1488 <= ({$unsigned((!forvar1336))} > reg1236[(2'h3):(2'h2)]);
                      reg1489 <= reg1416[(2'h3):(1'h1)];
                    end
                  for (forvar1491 = (1'h0); (forvar1491 < (1'h0)); forvar1491 = (forvar1491 + (1'h1)))
                    begin
                      reg1492 <= (^~$unsigned($signed((~forvar1260))));
                      reg1493 <= (~^$unsigned(($unsigned(forvar1453) >= (reg1249 >>> (8'ha0)))));
                      reg1494 <= $unsigned({$unsigned(reg1310)});
                    end
                  for (forvar1495 = (1'h0); (forvar1495 < (1'h1)); forvar1495 = (forvar1495 + (1'h1)))
                    begin
                      reg1496 <= $unsigned(reg1093[(3'h5):(2'h3)]);
                    end
                end
            end
          else
            begin
              for (forvar1479 = (1'h0); (forvar1479 < (2'h3)); forvar1479 = (forvar1479 + (1'h1)))
                begin
                  reg1480 <= (^~$unsigned((8'ha3)));
                end
              for (forvar1481 = (1'h0); (forvar1481 < (1'h0)); forvar1481 = (forvar1481 + (1'h1)))
                begin
                  for (forvar1482 = (1'h0); (forvar1482 < (2'h3)); forvar1482 = (forvar1482 + (1'h1)))
                    begin
                      reg1483 <= $signed($unsigned($unsigned((reg1110 >= reg1201))));
                      reg1484 <= forvar1443[(4'h8):(1'h1)];
                      reg1485 <= reg1150[(4'hc):(3'h4)];
                      reg1486 <= reg1292;
                    end
                  if ((~^reg1259))
                    begin
                      reg1487 <= reg1447;
                      reg1488 <= (!(8'hb0));
                      reg1489 <= $unsigned((reg1460 ?
                          ($unsigned(reg1185) ?
                              (~&reg1328) : forvar1126[(2'h2):(1'h1)]) : (~^forvar1478)));
                      reg1490 <= (reg1464 ?
                          ((8'h9c) ?
                              {(reg1260 < reg1182)} : {(&reg1266)}) : $signed({$unsigned(reg1065)}));
                    end
                  else
                    begin
                      reg1487 <= reg1080;
                    end
                  reg1491 <= $signed((^((reg1483 ?
                      reg1396 : (8'ha4)) >>> (~forvar1212))));
                  for (forvar1492 = (1'h0); (forvar1492 < (2'h2)); forvar1492 = (forvar1492 + (1'h1)))
                    begin
                      reg1493 <= (+reg1343);
                      reg1494 <= {$unsigned(forvar1334[(3'h4):(2'h2)])};
                      reg1495 <= reg1062;
                      reg1496 <= reg1415;
                    end
                end
              reg1497 <= (^forvar1291);
              if ({reg1475})
                begin
                  reg1498 <= (~$signed($unsigned(forvar1154)));
                end
              else
                begin
                  reg1498 <= {$unsigned((forvar1425[(3'h5):(1'h1)] ?
                          {reg1354} : (^reg1144)))};
                  for (forvar1499 = (1'h0); (forvar1499 < (1'h1)); forvar1499 = (forvar1499 + (1'h1)))
                    begin
                      reg1500 <= reg1275[(4'ha):(2'h2)];
                    end
                end
            end
          reg1501 <= reg1461[(2'h2):(1'h1)];
          if ((($signed((reg1169 - reg1138)) ?
              $signed($signed(forvar1327)) : $unsigned((!reg1217))) >> (((~|(8'hb6)) ?
              (~^reg1186) : (~&forvar1146)) - {$unsigned(reg1065)})))
            begin
              for (forvar1502 = (1'h0); (forvar1502 < (1'h0)); forvar1502 = (forvar1502 + (1'h1)))
                begin
                  for (forvar1503 = (1'h0); (forvar1503 < (1'h1)); forvar1503 = (forvar1503 + (1'h1)))
                    begin
                      reg1504 <= {(+forvar1395)};
                      reg1505 <= forvar1397[(3'h5):(3'h4)];
                      reg1506 <= reg1130;
                    end
                  reg1507 <= (~^(|forvar1370[(1'h0):(1'h0)]));
                  reg1508 <= reg1126;
                end
              if ((-reg1260))
                begin
                  reg1509 <= (~^$signed(((forvar1094 ? reg1232 : reg1177) ?
                      $signed(forvar1211) : reg1412)));
                  reg1510 <= reg1260;
                  if ($unsigned($signed(reg1396[(4'h8):(2'h2)])))
                    begin
                      reg1511 <= $signed($signed($unsigned((reg1286 ^ reg1463))));
                    end
                  else
                    begin
                      reg1511 <= forvar1291;
                      reg1512 <= wire1044[(4'he):(3'h6)];
                      reg1513 <= ({$signed($signed(reg1304))} != (forvar1119 ?
                          {$unsigned(forvar1048)} : (((8'ha8) <<< (8'ha4)) < {forvar1181})));
                    end
                  reg1514 <= ($signed($signed($signed(reg1473))) > reg1434[(4'h8):(3'h7)]);
                end
              else
                begin
                  for (forvar1509 = (1'h0); (forvar1509 < (1'h1)); forvar1509 = (forvar1509 + (1'h1)))
                    begin
                      reg1510 <= {$signed($signed($signed(reg1328)))};
                    end
                end
              for (forvar1515 = (1'h0); (forvar1515 < (1'h0)); forvar1515 = (forvar1515 + (1'h1)))
                begin
                  for (forvar1516 = (1'h0); (forvar1516 < (1'h0)); forvar1516 = (forvar1516 + (1'h1)))
                    begin
                      reg1517 <= ((|($signed(reg1506) ?
                          (~^reg1246) : $signed(reg1124))) < $unsigned(((reg1417 & reg1219) ?
                          $unsigned(reg1076) : (+forvar1246))));
                      reg1518 <= $signed(((~$unsigned(reg1447)) ?
                          ($signed((8'hb8)) & $signed((8'hb7))) : $unsigned((~^reg1057))));
                      reg1519 <= forvar1356[(1'h1):(1'h1)];
                    end
                  for (forvar1520 = (1'h0); (forvar1520 < (1'h0)); forvar1520 = (forvar1520 + (1'h1)))
                    begin
                      reg1521 <= $signed({$signed($unsigned(reg1131))});
                      reg1522 <= $signed(reg1272);
                      reg1523 <= {$unsigned(({reg1227} ^ (reg1424 ?
                              forvar1509 : reg1301)))};
                      reg1524 <= $signed($signed(forvar1137));
                    end
                  for (forvar1525 = (1'h0); (forvar1525 < (1'h1)); forvar1525 = (forvar1525 + (1'h1)))
                    begin
                      reg1526 <= ((((reg1076 - reg1508) + {reg1332}) ?
                              ($signed(reg1139) ?
                                  reg1413 : forvar1429) : $unsigned((forvar1468 & reg1136))) ?
                          reg1346[(3'h6):(1'h1)] : (reg1394[(2'h2):(1'h1)] ?
                              forvar1395[(4'hc):(4'h9)] : {(reg1056 != reg1513)}));
                    end
                  if ((reg1495[(3'h4):(2'h3)] ?
                      $unsigned($unsigned((reg1346 * reg1066))) : $unsigned((~^$unsigned(forvar1516)))))
                    begin
                      reg1527 <= $unsigned(reg1103[(3'h6):(3'h6)]);
                      reg1528 <= (8'ha2);
                      reg1529 <= (forvar1263 + reg1449[(4'hc):(2'h2)]);
                    end
                  else
                    begin
                      reg1527 <= {$signed(reg1354[(1'h1):(1'h1)])};
                      reg1528 <= reg1435;
                    end
                end
            end
          else
            begin
              if ((|$unsigned({(&reg1135)})))
                begin
                  if ((~&$signed((forvar1271[(1'h0):(1'h0)] <<< (^~reg1277)))))
                    begin
                      reg1502 <= reg1218;
                      reg1503 <= reg1433;
                    end
                  else
                    begin
                      reg1502 <= $unsigned($signed(($unsigned(forvar1491) <<< reg1197[(4'ha):(1'h1)])));
                      reg1503 <= $unsigned((~reg1256));
                      reg1504 <= (reg1155[(2'h2):(1'h0)] ?
                          $unsigned(((|reg1067) ?
                              reg1265[(5'h10):(4'h9)] : $unsigned(reg1399))) : {($signed((8'h9f)) ?
                                  forvar1516[(2'h2):(2'h2)] : (forvar1106 ?
                                      (8'hb2) : reg1357))});
                      reg1505 <= ((~|$signed((~&reg1066))) == ($unsigned((~^reg1383)) ?
                          ($unsigned(reg1411) | {forvar1396}) : $signed($signed(reg1348))));
                    end
                  if (((reg1060 ?
                      reg1416 : {(!(8'ha8))}) + $unsigned(forvar1429[(2'h2):(1'h0)])))
                    begin
                      reg1506 <= $unsigned(((((8'hb4) != (8'ha4)) <= (8'hb5)) ?
                          (forvar1137 ?
                              reg1314[(3'h5):(1'h1)] : $unsigned(forvar1126)) : {((8'h9f) ?
                                  reg1444 : forvar1327)}));
                      reg1507 <= (+$signed($signed((reg1194 ?
                          reg1335 : forvar1188))));
                      reg1508 <= forvar1502;
                      reg1509 <= reg1145[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1506 <= $signed(reg1297);
                      reg1507 <= $signed($unsigned(($unsigned(reg1169) <= reg1279[(1'h1):(1'h0)])));
                    end
                end
              else
                begin
                  if (reg1187[(2'h2):(1'h1)])
                    begin
                      reg1502 <= forvar1224;
                      reg1503 <= reg1290[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg1502 <= forvar1436[(4'h8):(2'h3)];
                      reg1503 <= {{{reg1401}}};
                    end
                  for (forvar1504 = (1'h0); (forvar1504 < (1'h0)); forvar1504 = (forvar1504 + (1'h1)))
                    begin
                      reg1505 <= $unsigned((~|(^reg1457[(4'h9):(3'h5)])));
                      reg1506 <= ((reg1321 << $unsigned(reg1529[(1'h1):(1'h0)])) == reg1143[(3'h5):(1'h1)]);
                    end
                end
              for (forvar1510 = (1'h0); (forvar1510 < (2'h2)); forvar1510 = (forvar1510 + (1'h1)))
                begin
                  if (($signed($unsigned((&forvar1425))) << forvar1495))
                    begin
                      reg1511 <= reg1322;
                    end
                  else
                    begin
                      reg1511 <= $unsigned(forvar1356[(4'ha):(3'h4)]);
                      reg1512 <= reg1414[(2'h3):(1'h0)];
                      reg1513 <= ((reg1354 ?
                              (^((8'hb9) ?
                                  reg1313 : reg1222)) : ($signed((8'ha7)) ~^ (~&forvar1065))) ?
                          reg1250 : (({reg1184} <<< reg1360[(3'h6):(3'h5)]) & (+$unsigned(reg1277))));
                      reg1514 <= (~^reg1452[(2'h3):(1'h0)]);
                    end
                end
            end
        end
    end
  assign wire1530 = reg1125[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      reg1531 <= $unsigned((reg1231 ? (|{reg1219}) : $signed({reg1089})));
    end
  module1532 modinst1740 (wire1739, clk, reg1438, reg1509, reg1072, reg1510);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1532  (y, clk, wire1536, wire1535, wire1534, wire1533);
  output wire [(32'h840):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire1536;
  input wire [(4'hd):(1'h0)] wire1535;
  input wire signed [(4'h9):(1'h0)] wire1534;
  input wire [(4'hf):(1'h0)] wire1533;
  wire [(5'h10):(1'h0)] wire1738;
  wire signed [(3'h5):(1'h0)] wire1737;
  wire signed [(3'h4):(1'h0)] wire1736;
  wire signed [(2'h3):(1'h0)] wire1735;
  wire [(3'h7):(1'h0)] wire1734;
  reg signed [(2'h2):(1'h0)] reg1733 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1732 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1731 = (1'h0);
  reg [(4'hb):(1'h0)] reg1730 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1729 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1728 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1727 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1726 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1718 = (1'h0);
  reg [(4'hd):(1'h0)] reg1725 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1724 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1723 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1722 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1721 = (1'h0);
  reg [(4'hc):(1'h0)] reg1720 = (1'h0);
  reg [(4'hc):(1'h0)] reg1719 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1718 = (1'h0);
  reg [(4'he):(1'h0)] reg1717 = (1'h0);
  reg [(3'h6):(1'h0)] reg1716 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1715 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1714 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1713 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1712 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1711 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1710 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1709 = (1'h0);
  reg [(2'h2):(1'h0)] reg1708 = (1'h0);
  reg [(4'h9):(1'h0)] reg1707 = (1'h0);
  reg [(4'hd):(1'h0)] reg1706 = (1'h0);
  reg [(2'h3):(1'h0)] reg1705 = (1'h0);
  reg [(4'hd):(1'h0)] reg1704 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1703 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1702 = (1'h0);
  reg [(2'h3):(1'h0)] reg1696 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1702 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1701 = (1'h0);
  reg [(3'h6):(1'h0)] reg1700 = (1'h0);
  reg [(2'h2):(1'h0)] reg1699 = (1'h0);
  reg [(4'hc):(1'h0)] reg1698 = (1'h0);
  reg [(2'h3):(1'h0)] reg1697 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1696 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1695 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1694 = (1'h0);
  reg [(3'h6):(1'h0)] reg1693 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1692 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1691 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1690 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1689 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1671 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1670 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1685 = (1'h0);
  reg [(4'he):(1'h0)] forvar1684 = (1'h0);
  reg [(3'h4):(1'h0)] reg1688 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1687 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1686 = (1'h0);
  reg [(4'he):(1'h0)] forvar1685 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1684 = (1'h0);
  reg [(4'he):(1'h0)] reg1683 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1682 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1681 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1680 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1679 = (1'h0);
  reg [(4'ha):(1'h0)] reg1678 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1677 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1676 = (1'h0);
  reg [(4'h8):(1'h0)] reg1675 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1674 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1673 = (1'h0);
  reg [(5'h10):(1'h0)] reg1672 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1671 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1670 = (1'h0);
  reg [(4'hf):(1'h0)] reg1669 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1668 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1659 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1648 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1653 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1639 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1638 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1647 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1644 = (1'h0);
  reg [(2'h2):(1'h0)] reg1649 = (1'h0);
  reg [(3'h6):(1'h0)] reg1646 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1643 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1632 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1629 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1627 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1667 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1666 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1665 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1664 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1663 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1655 = (1'h0);
  reg [(4'h9):(1'h0)] reg1662 = (1'h0);
  reg [(4'ha):(1'h0)] reg1661 = (1'h0);
  reg [(3'h6):(1'h0)] reg1660 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1659 = (1'h0);
  reg [(4'h8):(1'h0)] reg1658 = (1'h0);
  reg [(3'h5):(1'h0)] reg1657 = (1'h0);
  reg [(2'h3):(1'h0)] reg1656 = (1'h0);
  reg [(4'he):(1'h0)] reg1655 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1642 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1637 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1633 = (1'h0);
  reg [(4'h8):(1'h0)] reg1628 = (1'h0);
  reg [(3'h4):(1'h0)] reg1625 = (1'h0);
  reg [(2'h2):(1'h0)] reg1654 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1653 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1652 = (1'h0);
  reg [(4'hf):(1'h0)] reg1651 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1650 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1649 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1648 = (1'h0);
  reg [(4'he):(1'h0)] reg1647 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1646 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1645 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1641 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1644 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1643 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1642 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1641 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1640 = (1'h0);
  reg [(4'hf):(1'h0)] reg1639 = (1'h0);
  reg [(4'h8):(1'h0)] reg1638 = (1'h0);
  reg [(4'he):(1'h0)] reg1637 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1636 = (1'h0);
  reg [(3'h4):(1'h0)] reg1635 = (1'h0);
  reg [(4'hd):(1'h0)] reg1634 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1633 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1632 = (1'h0);
  reg [(3'h7):(1'h0)] reg1631 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1630 = (1'h0);
  reg [(3'h4):(1'h0)] reg1629 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1628 = (1'h0);
  reg [(4'he):(1'h0)] reg1627 = (1'h0);
  reg [(4'hd):(1'h0)] reg1626 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1625 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1624 = (1'h0);
  reg [(2'h3):(1'h0)] reg1623 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1622 = (1'h0);
  reg [(4'h9):(1'h0)] reg1621 = (1'h0);
  reg [(4'hc):(1'h0)] reg1620 = (1'h0);
  reg [(4'hb):(1'h0)] reg1619 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1618 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1617 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1599 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1616 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1615 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1614 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1613 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1612 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1611 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1610 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1609 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1608 = (1'h0);
  reg [(4'he):(1'h0)] reg1607 = (1'h0);
  reg [(4'hc):(1'h0)] reg1606 = (1'h0);
  reg [(4'hd):(1'h0)] reg1605 = (1'h0);
  reg [(4'hf):(1'h0)] reg1604 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1603 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1602 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1601 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1600 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1599 = (1'h0);
  reg [(3'h5):(1'h0)] reg1598 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1597 = (1'h0);
  reg [(3'h6):(1'h0)] reg1596 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1595 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1594 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1593 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1592 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1591 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1590 = (1'h0);
  reg [(3'h6):(1'h0)] reg1589 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1588 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1587 = (1'h0);
  reg [(5'h10):(1'h0)] reg1579 = (1'h0);
  reg [(4'hd):(1'h0)] reg1586 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1585 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1584 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1583 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1582 = (1'h0);
  reg [(4'h8):(1'h0)] reg1581 = (1'h0);
  reg [(4'hd):(1'h0)] reg1580 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1579 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1578 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1577 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1576 = (1'h0);
  reg [(4'hf):(1'h0)] reg1575 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1574 = (1'h0);
  reg [(5'h10):(1'h0)] reg1573 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1572 = (1'h0);
  reg [(2'h3):(1'h0)] reg1571 = (1'h0);
  reg [(4'ha):(1'h0)] reg1570 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1569 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1568 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1560 = (1'h0);
  reg [(4'hb):(1'h0)] reg1567 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1566 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1565 = (1'h0);
  reg [(5'h10):(1'h0)] reg1564 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1563 = (1'h0);
  reg [(4'h9):(1'h0)] reg1562 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1561 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1560 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1559 = (1'h0);
  reg [(5'h10):(1'h0)] reg1558 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1557 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1556 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1555 = (1'h0);
  reg [(3'h7):(1'h0)] reg1554 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1553 = (1'h0);
  reg [(4'h8):(1'h0)] reg1552 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1551 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1550 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1549 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1548 = (1'h0);
  reg [(3'h6):(1'h0)] reg1547 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1546 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1545 = (1'h0);
  reg [(4'he):(1'h0)] reg1544 = (1'h0);
  reg [(3'h4):(1'h0)] reg1542 = (1'h0);
  reg [(4'h8):(1'h0)] reg1543 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1542 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1541 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1540 = (1'h0);
  wire [(4'ha):(1'h0)] wire1539;
  wire signed [(4'he):(1'h0)] wire1538;
  wire [(4'ha):(1'h0)] wire1537;
  assign y = {wire1738,
                 wire1737,
                 wire1736,
                 wire1735,
                 wire1734,
                 reg1733,
                 forvar1732,
                 reg1731,
                 reg1730,
                 reg1729,
                 reg1728,
                 forvar1727,
                 forvar1726,
                 forvar1718,
                 reg1725,
                 reg1724,
                 reg1723,
                 forvar1722,
                 reg1721,
                 reg1720,
                 reg1719,
                 reg1718,
                 reg1717,
                 reg1716,
                 reg1715,
                 forvar1714,
                 forvar1713,
                 reg1712,
                 reg1711,
                 forvar1710,
                 reg1709,
                 reg1708,
                 reg1707,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1703,
                 forvar1702,
                 reg1696,
                 reg1702,
                 reg1701,
                 reg1700,
                 reg1699,
                 reg1698,
                 reg1697,
                 forvar1696,
                 reg1695,
                 reg1694,
                 reg1693,
                 forvar1692,
                 forvar1691,
                 forvar1690,
                 forvar1689,
                 reg1671,
                 reg1670,
                 reg1685,
                 forvar1684,
                 reg1688,
                 reg1687,
                 reg1686,
                 forvar1685,
                 reg1684,
                 reg1683,
                 reg1682,
                 reg1681,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 forvar1674,
                 reg1673,
                 reg1672,
                 forvar1671,
                 forvar1670,
                 reg1669,
                 forvar1668,
                 reg1659,
                 forvar1648,
                 forvar1653,
                 forvar1639,
                 forvar1638,
                 forvar1647,
                 forvar1644,
                 reg1649,
                 reg1646,
                 forvar1643,
                 forvar1632,
                 forvar1629,
                 forvar1627,
                 reg1667,
                 reg1666,
                 reg1665,
                 reg1664,
                 forvar1663,
                 forvar1655,
                 reg1662,
                 reg1661,
                 reg1660,
                 forvar1659,
                 reg1658,
                 reg1657,
                 reg1656,
                 reg1655,
                 forvar1642,
                 forvar1637,
                 reg1633,
                 reg1628,
                 reg1625,
                 reg1654,
                 reg1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 forvar1649,
                 reg1648,
                 reg1647,
                 forvar1646,
                 reg1645,
                 forvar1641,
                 reg1644,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 reg1637,
                 reg1636,
                 reg1635,
                 reg1634,
                 forvar1633,
                 reg1632,
                 reg1631,
                 reg1630,
                 reg1629,
                 forvar1628,
                 reg1627,
                 reg1626,
                 forvar1625,
                 forvar1624,
                 reg1623,
                 forvar1622,
                 reg1621,
                 reg1620,
                 reg1619,
                 forvar1618,
                 forvar1617,
                 reg1599,
                 reg1616,
                 reg1615,
                 reg1614,
                 reg1613,
                 forvar1612,
                 reg1611,
                 reg1610,
                 reg1609,
                 forvar1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1603,
                 reg1602,
                 reg1601,
                 reg1600,
                 forvar1599,
                 reg1598,
                 forvar1597,
                 reg1596,
                 reg1595,
                 reg1594,
                 forvar1593,
                 forvar1592,
                 reg1591,
                 reg1590,
                 reg1589,
                 forvar1588,
                 forvar1587,
                 reg1579,
                 reg1586,
                 reg1585,
                 reg1584,
                 reg1583,
                 forvar1582,
                 reg1581,
                 reg1580,
                 forvar1579,
                 reg1578,
                 reg1577,
                 reg1576,
                 reg1575,
                 forvar1574,
                 reg1573,
                 forvar1572,
                 reg1571,
                 reg1570,
                 reg1569,
                 reg1568,
                 forvar1560,
                 reg1567,
                 forvar1566,
                 reg1565,
                 reg1564,
                 reg1563,
                 reg1562,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1558,
                 forvar1557,
                 reg1556,
                 reg1555,
                 reg1554,
                 forvar1553,
                 reg1552,
                 reg1551,
                 reg1550,
                 reg1549,
                 reg1548,
                 reg1547,
                 forvar1546,
                 reg1545,
                 reg1544,
                 reg1542,
                 reg1543,
                 forvar1542,
                 forvar1541,
                 forvar1540,
                 wire1539,
                 wire1538,
                 wire1537,
                 (1'h0)};
  assign wire1537 = ((wire1536[(3'h4):(2'h3)] ?
                        (^(^(8'hb1))) : (^wire1533[(1'h0):(1'h0)])) || ({wire1534} ?
                        (wire1533[(3'h6):(1'h0)] ?
                            wire1535 : $unsigned(wire1533)) : (^(wire1536 >= (8'haf)))));
  assign wire1538 = wire1534;
  assign wire1539 = $signed((wire1537 && (wire1533 ?
                        $unsigned(wire1534) : (wire1534 ?
                            wire1536 : wire1537))));
  always
    @(posedge clk) begin
      for (forvar1540 = (1'h0); (forvar1540 < (1'h0)); forvar1540 = (forvar1540 + (1'h1)))
        begin
          for (forvar1541 = (1'h0); (forvar1541 < (2'h2)); forvar1541 = (forvar1541 + (1'h1)))
            begin
              if (forvar1540[(1'h0):(1'h0)])
                begin
                  for (forvar1542 = (1'h0); (forvar1542 < (2'h3)); forvar1542 = (forvar1542 + (1'h1)))
                    begin
                      reg1543 <= (wire1534 ^~ $unsigned({forvar1542[(1'h1):(1'h1)]}));
                    end
                end
              else
                begin
                  if (forvar1540)
                    begin
                      reg1542 <= forvar1540;
                      reg1543 <= reg1543[(2'h2):(2'h2)];
                      reg1544 <= forvar1542;
                      reg1545 <= reg1544[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg1542 <= wire1537[(3'h7):(2'h2)];
                    end
                  for (forvar1546 = (1'h0); (forvar1546 < (2'h2)); forvar1546 = (forvar1546 + (1'h1)))
                    begin
                      reg1547 <= {$signed(forvar1542)};
                      reg1548 <= $signed($unsigned(reg1543[(3'h6):(3'h5)]));
                    end
                  if ((wire1534[(3'h5):(3'h4)] ?
                      $unsigned((|reg1544[(1'h0):(1'h0)])) : ((+wire1538) == (~|wire1533[(1'h0):(1'h0)]))))
                    begin
                      reg1549 <= (reg1545[(2'h2):(2'h2)] >= (-({wire1537} * (~|wire1535))));
                      reg1550 <= wire1533;
                      reg1551 <= ($signed(forvar1541) && ((^$signed(wire1534)) ?
                          wire1539 : wire1538));
                    end
                  else
                    begin
                      reg1549 <= {wire1537};
                      reg1550 <= (~$unsigned(wire1538[(4'hc):(4'ha)]));
                      reg1551 <= ($unsigned({(wire1534 - reg1550)}) ?
                          (8'ha8) : $unsigned((8'hb7)));
                      reg1552 <= $unsigned(((8'hb9) ?
                          {forvar1540} : (^(wire1537 != wire1534))));
                    end
                  for (forvar1553 = (1'h0); (forvar1553 < (1'h1)); forvar1553 = (forvar1553 + (1'h1)))
                    begin
                      reg1554 <= ($signed(reg1543[(3'h7):(2'h2)]) ?
                          $unsigned($unsigned(forvar1542[(1'h1):(1'h1)])) : wire1534);
                      reg1555 <= $unsigned(($unsigned($signed(reg1552)) ?
                          reg1552[(3'h4):(3'h4)] : (~&$signed(wire1536))));
                      reg1556 <= ($unsigned((reg1552 ?
                              wire1537[(3'h5):(1'h0)] : (reg1555 ?
                                  wire1537 : wire1534))) ?
                          wire1535[(3'h6):(1'h1)] : (reg1552[(1'h0):(1'h0)] ?
                              wire1537[(3'h5):(1'h0)] : $signed((&wire1536))));
                    end
                end
              for (forvar1557 = (1'h0); (forvar1557 < (1'h0)); forvar1557 = (forvar1557 + (1'h1)))
                begin
                  reg1558 <= ($signed($unsigned({reg1542})) ?
                      {$signed($unsigned(wire1535))} : $unsigned(wire1534));
                end
              reg1559 <= (~(((forvar1541 - reg1551) && $signed((8'ha5))) ?
                  forvar1540[(4'h8):(3'h5)] : (+reg1554)));
              if (wire1538)
                begin
                  reg1560 <= reg1559;
                  if ($signed(reg1542))
                    begin
                      reg1561 <= reg1548[(2'h2):(2'h2)];
                      reg1562 <= (reg1555 ?
                          (~((reg1552 ? reg1555 : (8'ha5)) ?
                              reg1545[(2'h3):(1'h1)] : (reg1545 >= reg1555))) : reg1548);
                      reg1563 <= forvar1546[(5'h10):(4'h9)];
                      reg1564 <= $signed(($signed($signed(reg1555)) >>> ($unsigned(reg1560) ~^ (forvar1546 ?
                          reg1555 : wire1536))));
                    end
                  else
                    begin
                      reg1561 <= {((~|$unsigned(reg1548)) ?
                              {(^~reg1544)} : $signed({reg1548}))};
                      reg1562 <= {reg1556[(2'h2):(1'h0)]};
                    end
                  reg1565 <= {$signed($unsigned($unsigned(reg1545)))};
                  for (forvar1566 = (1'h0); (forvar1566 < (1'h1)); forvar1566 = (forvar1566 + (1'h1)))
                    begin
                      reg1567 <= (^reg1543[(3'h6):(3'h5)]);
                    end
                end
              else
                begin
                  for (forvar1560 = (1'h0); (forvar1560 < (2'h2)); forvar1560 = (forvar1560 + (1'h1)))
                    begin
                      reg1561 <= reg1564;
                      reg1562 <= {reg1564[(3'h7):(1'h0)]};
                    end
                  if (($signed(wire1536[(2'h3):(1'h1)]) ?
                      (-$signed((reg1555 >> reg1555))) : (+$unsigned($unsigned(reg1542)))))
                    begin
                      reg1563 <= (8'had);
                      reg1564 <= reg1549;
                      reg1565 <= $unsigned($unsigned(reg1559[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg1563 <= {(((^~reg1565) & $signed(forvar1541)) != ($unsigned(reg1552) || $signed(forvar1560)))};
                      reg1564 <= $unsigned($unsigned(reg1565[(1'h1):(1'h0)]));
                    end
                  for (forvar1566 = (1'h0); (forvar1566 < (1'h1)); forvar1566 = (forvar1566 + (1'h1)))
                    begin
                      reg1567 <= ($unsigned(forvar1566) ?
                          wire1539 : (reg1549[(1'h0):(1'h0)] ?
                              (8'hab) : ((!(8'ha0)) >= $unsigned(forvar1566))));
                      reg1568 <= ($signed(wire1534[(1'h0):(1'h0)]) * $signed((~&reg1544)));
                      reg1569 <= ($signed((8'hb5)) ?
                          reg1559[(2'h2):(1'h0)] : ($signed((~^reg1549)) >> ((reg1560 && reg1555) * ((8'hb0) ?
                              reg1548 : wire1534))));
                    end
                  if ($signed((reg1552[(3'h6):(1'h0)] ?
                      $unsigned((wire1534 && (8'ha5))) : ((forvar1557 ?
                              forvar1566 : reg1543) ?
                          $unsigned(reg1559) : (reg1554 ? reg1565 : reg1568)))))
                    begin
                      reg1570 <= ((|reg1558[(3'h4):(2'h3)]) ?
                          (-reg1545) : reg1554[(1'h0):(1'h0)]);
                      reg1571 <= reg1543;
                    end
                  else
                    begin
                      reg1570 <= $signed((-(+$signed(forvar1540))));
                    end
                end
            end
          for (forvar1572 = (1'h0); (forvar1572 < (1'h0)); forvar1572 = (forvar1572 + (1'h1)))
            begin
              if ((((&(wire1538 <= forvar1557)) ?
                  $unsigned((~|reg1556)) : (-reg1556[(2'h3):(1'h1)])) - (reg1543[(2'h3):(1'h0)] ?
                  $signed((8'ha1)) : ((reg1544 == reg1563) ?
                      (~&reg1564) : $signed((8'h9f))))))
                begin
                  reg1573 <= reg1565;
                  for (forvar1574 = (1'h0); (forvar1574 < (1'h1)); forvar1574 = (forvar1574 + (1'h1)))
                    begin
                      reg1575 <= {$unsigned(wire1539)};
                      reg1576 <= ((~|(reg1554[(3'h6):(1'h0)] <= $unsigned(reg1569))) ~^ ((~&$unsigned(reg1547)) != $signed((forvar1574 >> (8'had)))));
                      reg1577 <= (reg1552[(3'h4):(2'h3)] << (~&(reg1568 << (reg1568 <= wire1539))));
                      reg1578 <= {{$unsigned({(8'ha6)})}};
                    end
                  for (forvar1579 = (1'h0); (forvar1579 < (2'h2)); forvar1579 = (forvar1579 + (1'h1)))
                    begin
                      reg1580 <= (reg1578[(3'h6):(3'h4)] ?
                          reg1556[(2'h2):(1'h1)] : $signed({wire1537[(2'h2):(2'h2)]}));
                      reg1581 <= reg1556[(1'h0):(1'h0)];
                    end
                  for (forvar1582 = (1'h0); (forvar1582 < (2'h2)); forvar1582 = (forvar1582 + (1'h1)))
                    begin
                      reg1583 <= ((~|$unsigned($unsigned(forvar1541))) > ((^~forvar1541[(2'h3):(2'h3)]) ^ (~|$signed((8'h9c)))));
                      reg1584 <= $unsigned(($signed((wire1533 ^ (8'hb7))) ?
                          (!$signed((8'haa))) : {$signed(wire1536)}));
                      reg1585 <= (^~wire1535);
                      reg1586 <= (reg1577[(4'h9):(3'h4)] ?
                          $signed({{reg1571}}) : $unsigned(((-reg1575) >> (forvar1553 - reg1567))));
                    end
                end
              else
                begin
                  reg1573 <= ($unsigned(forvar1557[(3'h5):(1'h0)]) <<< ($unsigned(reg1564) ?
                      $signed(wire1538[(4'he):(2'h2)]) : (~^(reg1555 ?
                          forvar1579 : reg1576))));
                  for (forvar1574 = (1'h0); (forvar1574 < (2'h2)); forvar1574 = (forvar1574 + (1'h1)))
                    begin
                      reg1575 <= $signed(($unsigned($unsigned(forvar1566)) >>> (reg1567[(1'h0):(1'h0)] >>> (forvar1560 ?
                          (8'hae) : reg1573))));
                      reg1576 <= {($signed($unsigned(forvar1574)) ?
                              $signed((wire1539 ?
                                  forvar1542 : forvar1546)) : (8'h9c))};
                      reg1577 <= (~|reg1573[(3'h6):(1'h0)]);
                      reg1578 <= wire1538;
                    end
                  reg1579 <= $signed((^$signed(((8'hae) ? reg1549 : (8'h9c)))));
                end
              for (forvar1587 = (1'h0); (forvar1587 < (1'h1)); forvar1587 = (forvar1587 + (1'h1)))
                begin
                  for (forvar1588 = (1'h0); (forvar1588 < (1'h1)); forvar1588 = (forvar1588 + (1'h1)))
                    begin
                      reg1589 <= (8'hb1);
                      reg1590 <= ($unsigned(reg1575) != $signed((~^(wire1538 ?
                          (8'ha5) : reg1545))));
                      reg1591 <= reg1578;
                    end
                end
            end
          for (forvar1592 = (1'h0); (forvar1592 < (2'h3)); forvar1592 = (forvar1592 + (1'h1)))
            begin
              for (forvar1593 = (1'h0); (forvar1593 < (2'h3)); forvar1593 = (forvar1593 + (1'h1)))
                begin
                  reg1594 <= ($signed($signed(reg1565)) ?
                      ((reg1558[(1'h0):(1'h0)] ^ $unsigned((8'ha0))) <<< ($signed(reg1559) ?
                          (reg1542 ?
                              reg1573 : wire1533) : (8'hb5))) : $unsigned(reg1555));
                  reg1595 <= $signed({forvar1541});
                end
              reg1596 <= ($signed($unsigned($unsigned((8'hb0)))) != reg1563[(1'h1):(1'h0)]);
            end
          for (forvar1597 = (1'h0); (forvar1597 < (1'h0)); forvar1597 = (forvar1597 + (1'h1)))
            begin
              reg1598 <= $signed((+$signed((8'ha7))));
              if (reg1596)
                begin
                  for (forvar1599 = (1'h0); (forvar1599 < (1'h0)); forvar1599 = (forvar1599 + (1'h1)))
                    begin
                      reg1600 <= $unsigned(forvar1557);
                      reg1601 <= $signed((reg1595[(4'ha):(4'h9)] ^~ {((8'ha8) - reg1571)}));
                      reg1602 <= forvar1592;
                      reg1603 <= (|reg1555);
                    end
                  if ((((-reg1564) ?
                      $signed((~&wire1534)) : (~((8'ha1) ?
                          (8'had) : forvar1587))) >>> (reg1555[(3'h4):(1'h0)] >= (|forvar1588))))
                    begin
                      reg1604 <= (($unsigned(reg1559) ?
                          (^{(8'hb0)}) : ((reg1600 != forvar1592) ?
                              reg1601 : (^~forvar1592))) + $signed(reg1576));
                      reg1605 <= $unsigned({(forvar1557 && $signed(reg1571))});
                      reg1606 <= reg1552[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg1604 <= (~|{($unsigned(reg1595) != {reg1594})});
                      reg1605 <= wire1536;
                      reg1606 <= reg1558;
                      reg1607 <= ({$signed($unsigned(reg1590))} ?
                          {reg1584} : ((8'hab) ^ (~|(reg1603 & wire1539))));
                    end
                  for (forvar1608 = (1'h0); (forvar1608 < (1'h0)); forvar1608 = (forvar1608 + (1'h1)))
                    begin
                      reg1609 <= $signed($unsigned($unsigned((wire1537 & reg1570))));
                      reg1610 <= $signed($signed($unsigned((wire1535 ?
                          reg1591 : (8'hb5)))));
                      reg1611 <= reg1542[(3'h4):(2'h3)];
                    end
                  for (forvar1612 = (1'h0); (forvar1612 < (1'h1)); forvar1612 = (forvar1612 + (1'h1)))
                    begin
                      reg1613 <= reg1575[(4'ha):(3'h6)];
                      reg1614 <= $unsigned((reg1568[(2'h2):(1'h0)] ?
                          forvar1579[(4'h8):(4'h8)] : reg1595));
                      reg1615 <= reg1558[(3'h5):(2'h3)];
                      reg1616 <= ($signed((8'hba)) ?
                          forvar1566 : (~&reg1613[(3'h6):(3'h4)]));
                    end
                end
              else
                begin
                  if ((forvar1540 ^~ ((reg1602[(4'he):(3'h5)] & reg1613[(3'h4):(3'h4)]) ?
                      reg1542 : $unsigned(((8'ha7) ? (8'had) : reg1560)))))
                    begin
                      reg1599 <= {((~forvar1588) ?
                              ((~reg1575) ?
                                  ((8'ha5) < reg1544) : $unsigned(reg1550)) : (wire1533[(3'h4):(1'h0)] < (~&reg1585)))};
                      reg1600 <= $unsigned($signed({(reg1568 <= reg1570)}));
                      reg1601 <= ((|($signed(forvar1592) ?
                          $signed(reg1556) : reg1543[(1'h1):(1'h1)])) || ($signed($unsigned(forvar1574)) - {reg1569}));
                    end
                  else
                    begin
                      reg1599 <= (reg1602 >= (8'h9c));
                    end
                  if ((~&(!reg1549)))
                    begin
                      reg1602 <= reg1542;
                      reg1603 <= $unsigned((reg1556[(2'h2):(1'h1)] ?
                          $unsigned($signed(reg1605)) : (|$unsigned(wire1539))));
                      reg1604 <= ((($signed(wire1538) ?
                              reg1581[(4'h8):(1'h1)] : reg1579[(4'ha):(3'h6)]) <= reg1573) ?
                          $unsigned(($unsigned(reg1601) || $unsigned(forvar1572))) : $signed(reg1585));
                      reg1605 <= (reg1598 ?
                          $unsigned($unsigned($signed(reg1556))) : $unsigned($unsigned($unsigned(reg1601))));
                    end
                  else
                    begin
                      reg1602 <= (~^(~^forvar1574));
                      reg1603 <= $unsigned(forvar1560);
                      reg1604 <= $unsigned((forvar1566 ?
                          ((reg1614 != forvar1553) >= reg1575) : $signed($unsigned(reg1559))));
                    end
                end
              for (forvar1617 = (1'h0); (forvar1617 < (2'h3)); forvar1617 = (forvar1617 + (1'h1)))
                begin
                  for (forvar1618 = (1'h0); (forvar1618 < (1'h0)); forvar1618 = (forvar1618 + (1'h1)))
                    begin
                      reg1619 <= (((^(reg1550 ? forvar1541 : (8'hb0))) ?
                              $unsigned({forvar1597}) : {(wire1534 ?
                                      reg1589 : forvar1582)}) ?
                          $signed((~^reg1586[(2'h3):(2'h2)])) : {$signed($unsigned((8'h9c)))});
                      reg1620 <= ((reg1565[(3'h5):(1'h0)] < $unsigned($signed(forvar1557))) >> ((~(reg1581 >> (8'h9d))) >= reg1543));
                      reg1621 <= $signed($signed(reg1577));
                    end
                  for (forvar1622 = (1'h0); (forvar1622 < (1'h1)); forvar1622 = (forvar1622 + (1'h1)))
                    begin
                      reg1623 <= reg1594;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg1607[(4'hd):(3'h5)])
        begin
          if ((|$unsigned($signed((^~reg1619)))))
            begin
              for (forvar1624 = (1'h0); (forvar1624 < (1'h0)); forvar1624 = (forvar1624 + (1'h1)))
                begin
                  for (forvar1625 = (1'h0); (forvar1625 < (1'h1)); forvar1625 = (forvar1625 + (1'h1)))
                    begin
                      reg1626 <= forvar1624;
                      reg1627 <= reg1620;
                    end
                  for (forvar1628 = (1'h0); (forvar1628 < (2'h3)); forvar1628 = (forvar1628 + (1'h1)))
                    begin
                      reg1629 <= reg1548[(4'h8):(3'h5)];
                      reg1630 <= (8'h9f);
                      reg1631 <= $unsigned($signed(reg1565));
                      reg1632 <= $signed((~((reg1542 ^ reg1579) ^~ ((8'ha2) ~^ reg1585))));
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h3)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= (reg1576[(3'h6):(2'h2)] * ($signed((~&reg1549)) <= reg1581[(3'h7):(2'h2)]));
                      reg1635 <= (~({(+reg1616)} ?
                          ((^forvar1587) <<< (reg1571 <= reg1570)) : (-(|forvar1541))));
                      reg1636 <= (-forvar1553);
                      reg1637 <= (($unsigned(((8'hb9) ?
                          reg1564 : reg1555)) < $unsigned(forvar1617[(3'h6):(2'h3)])) >>> $unsigned(reg1631));
                    end
                  if (reg1570)
                    begin
                      reg1638 <= $signed((~&((reg1569 < forvar1579) | forvar1572[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg1638 <= (({$signed(reg1542)} | reg1589[(2'h2):(1'h0)]) ?
                          ((^{(8'hb7)}) != ((^reg1568) ^~ (^~reg1545))) : $signed({(forvar1599 ?
                                  reg1550 : reg1602)}));
                      reg1639 <= (8'hb6);
                      reg1640 <= wire1533[(4'h8):(2'h2)];
                    end
                end
              if (((^reg1584) ?
                  forvar1608[(3'h6):(2'h3)] : ((((8'ha3) ? reg1586 : reg1632) ?
                      reg1613 : $unsigned(reg1638)) == ((|reg1598) ?
                      $signed((8'hb5)) : $unsigned(reg1581)))))
                begin
                  if ((reg1590 + reg1575))
                    begin
                      reg1641 <= (!(&((~(8'haa)) ?
                          (reg1580 && reg1604) : forvar1579)));
                      reg1642 <= ({($unsigned(wire1535) ?
                                  (8'haf) : $unsigned(reg1567))} ?
                          (reg1621 & {$signed(forvar1618)}) : (+$unsigned((reg1554 > reg1640))));
                      reg1643 <= (forvar1572 - forvar1622);
                    end
                  else
                    begin
                      reg1641 <= {$unsigned(((|reg1606) ?
                              $unsigned(reg1590) : (^(8'hba))))};
                      reg1642 <= $signed($signed((reg1579[(3'h4):(1'h1)] ?
                          $unsigned(reg1643) : $signed(reg1594))));
                      reg1643 <= reg1632;
                    end
                  reg1644 <= reg1569;
                end
              else
                begin
                  for (forvar1641 = (1'h0); (forvar1641 < (2'h2)); forvar1641 = (forvar1641 + (1'h1)))
                    begin
                      reg1642 <= ((reg1611 ?
                              $signed(reg1559) : reg1571[(1'h1):(1'h0)]) ?
                          (forvar1592[(3'h6):(3'h5)] ?
                              reg1615 : forvar1579) : (~|(reg1555 ?
                              {reg1585} : {forvar1633})));
                      reg1643 <= (~&(~^reg1619[(1'h1):(1'h0)]));
                      reg1644 <= reg1583[(4'h8):(2'h3)];
                      reg1645 <= reg1555;
                    end
                  for (forvar1646 = (1'h0); (forvar1646 < (1'h1)); forvar1646 = (forvar1646 + (1'h1)))
                    begin
                      reg1647 <= $unsigned(($signed((~|wire1533)) > reg1638[(2'h3):(1'h0)]));
                      reg1648 <= $signed({(-forvar1612)});
                    end
                  for (forvar1649 = (1'h0); (forvar1649 < (2'h3)); forvar1649 = (forvar1649 + (1'h1)))
                    begin
                      reg1650 <= ($signed($unsigned(reg1548[(1'h1):(1'h0)])) ^ (($unsigned(reg1554) ?
                              (~|forvar1622) : $unsigned(forvar1625)) ?
                          ((reg1613 - forvar1542) | ((8'hb1) ?
                              reg1606 : reg1636)) : $unsigned($unsigned(forvar1624))));
                      reg1651 <= $unsigned(wire1538[(4'h9):(3'h5)]);
                      reg1652 <= $unsigned((~&reg1601[(3'h7):(3'h5)]));
                      reg1653 <= $unsigned($unsigned($signed(reg1558)));
                    end
                end
              reg1654 <= {reg1620[(4'hc):(4'hc)]};
            end
          else
            begin
              for (forvar1624 = (1'h0); (forvar1624 < (1'h1)); forvar1624 = (forvar1624 + (1'h1)))
                begin
                  if (((reg1644[(4'hb):(3'h7)] ?
                      $unsigned($unsigned(reg1632)) : ((reg1604 != reg1643) >= reg1555[(1'h1):(1'h1)])) >= wire1536[(3'h4):(1'h0)]))
                    begin
                      reg1625 <= $unsigned($unsigned(((~^forvar1588) ?
                          (forvar1612 >>> forvar1587) : reg1589)));
                      reg1626 <= $unsigned({(~^forvar1617[(4'h8):(3'h7)])});
                      reg1627 <= ((~&$signed($unsigned(forvar1588))) ?
                          (wire1537 ?
                              $signed(reg1568[(2'h3):(2'h2)]) : reg1552[(2'h2):(1'h1)]) : {$signed(reg1542[(2'h2):(1'h1)])});
                      reg1628 <= $signed(reg1640[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1625 <= forvar1628[(1'h0):(1'h0)];
                      reg1626 <= reg1579;
                    end
                  if (({{((8'ha4) ? reg1551 : reg1570)}} ?
                      $signed(reg1577[(3'h6):(3'h5)]) : forvar1579[(3'h4):(2'h3)]))
                    begin
                      reg1629 <= $signed((reg1571 ?
                          ((^~reg1545) ?
                              (wire1538 <<< (8'hb9)) : ((8'hb3) <<< (8'hb9))) : {(reg1570 ?
                                  forvar1553 : reg1626)}));
                    end
                  else
                    begin
                      reg1629 <= (($signed((reg1581 ~^ (8'haf))) && reg1628[(2'h3):(2'h3)]) ?
                          (&({reg1648} ?
                              (reg1577 <<< forvar1587) : reg1579[(4'he):(4'hc)])) : $unsigned(((wire1536 ?
                                  (8'h9c) : wire1537) ?
                              $unsigned(reg1558) : $signed(reg1580))));
                      reg1630 <= ((~&(-$signed(reg1600))) ?
                          reg1571 : (forvar1624[(2'h3):(1'h0)] ?
                              $unsigned((reg1603 <<< (8'h9d))) : $unsigned(wire1536)));
                      reg1631 <= reg1554[(3'h4):(3'h4)];
                      reg1632 <= (-$signed(($signed(reg1594) ?
                          {reg1564} : {reg1619})));
                    end
                end
              if ({(^~(reg1594[(3'h4):(2'h2)] ~^ $signed(reg1596)))})
                begin
                  reg1633 <= reg1638;
                end
              else
                begin
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h3)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= reg1543[(4'h8):(2'h3)];
                      reg1635 <= $signed($signed(reg1647[(4'he):(1'h0)]));
                      reg1636 <= $signed((|$signed(reg1643)));
                    end
                  for (forvar1637 = (1'h0); (forvar1637 < (1'h1)); forvar1637 = (forvar1637 + (1'h1)))
                    begin
                      reg1638 <= reg1558;
                      reg1639 <= (reg1607[(4'hc):(3'h5)] <= reg1629[(1'h0):(1'h0)]);
                      reg1640 <= $signed($unsigned(({(8'h9d)} - $signed(wire1535))));
                    end
                end
              for (forvar1641 = (1'h0); (forvar1641 < (2'h3)); forvar1641 = (forvar1641 + (1'h1)))
                begin
                  for (forvar1642 = (1'h0); (forvar1642 < (1'h0)); forvar1642 = (forvar1642 + (1'h1)))
                    begin
                      reg1643 <= (&$unsigned($unsigned($unsigned(forvar1574))));
                      reg1644 <= ($unsigned((!(forvar1541 ?
                          reg1584 : forvar1641))) <<< (($signed((8'hac)) >>> reg1610) >> reg1548[(1'h1):(1'h1)]));
                    end
                  reg1645 <= reg1586[(4'ha):(3'h7)];
                end
            end
          if ($unsigned(forvar1592))
            begin
              if (reg1623[(1'h0):(1'h0)])
                begin
                  if (reg1642)
                    begin
                      reg1655 <= $unsigned(reg1611[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1655 <= (+reg1550[(3'h5):(2'h2)]);
                      reg1656 <= {(~^(reg1560 ?
                              reg1569[(3'h5):(1'h0)] : forvar1622))};
                      reg1657 <= {(8'hb4)};
                    end
                  reg1658 <= (reg1638[(3'h4):(2'h2)] ?
                      {$signed((reg1556 | reg1571))} : reg1559);
                  for (forvar1659 = (1'h0); (forvar1659 < (2'h2)); forvar1659 = (forvar1659 + (1'h1)))
                    begin
                      reg1660 <= $unsigned($signed($signed($unsigned(reg1559))));
                      reg1661 <= ($unsigned(($unsigned(forvar1618) ?
                              reg1584 : $signed(wire1536))) ?
                          $unsigned(((reg1633 ?
                              reg1558 : forvar1553) >= $unsigned(wire1538))) : (~|{(&reg1605)}));
                      reg1662 <= (~^reg1579[(2'h2):(2'h2)]);
                    end
                end
              else
                begin
                  for (forvar1655 = (1'h0); (forvar1655 < (1'h0)); forvar1655 = (forvar1655 + (1'h1)))
                    begin
                      reg1656 <= {((~&{reg1583}) ?
                              reg1619 : ($unsigned(reg1644) == (^(8'ha4))))};
                    end
                  if (((&{(reg1543 <<< reg1610)}) ? reg1602 : $signed((8'ha0))))
                    begin
                      reg1657 <= {$signed(((reg1579 ^ forvar1593) ?
                              ((8'hb3) ?
                                  reg1567 : reg1621) : (reg1643 && reg1580)))};
                    end
                  else
                    begin
                      reg1657 <= ({reg1645[(3'h6):(1'h0)]} ?
                          (8'haf) : $signed($unsigned((8'hb1))));
                      reg1658 <= (~^(((forvar1642 >= reg1548) ~^ $signed(reg1549)) <<< reg1632));
                    end
                end
            end
          else
            begin
              if ((~(!(8'hb1))))
                begin
                  reg1655 <= (^$signed($signed(reg1642)));
                end
              else
                begin
                  for (forvar1655 = (1'h0); (forvar1655 < (1'h0)); forvar1655 = (forvar1655 + (1'h1)))
                    begin
                      reg1656 <= ((~^{(reg1554 < reg1619)}) ?
                          reg1640 : forvar1593[(1'h1):(1'h0)]);
                      reg1657 <= $signed(forvar1649[(4'hf):(4'h9)]);
                      reg1658 <= $signed({wire1534[(2'h3):(2'h2)]});
                    end
                  for (forvar1659 = (1'h0); (forvar1659 < (1'h1)); forvar1659 = (forvar1659 + (1'h1)))
                    begin
                      reg1660 <= (~|$signed(reg1595));
                      reg1661 <= (reg1565[(2'h2):(1'h1)] ?
                          (($signed(forvar1541) ?
                                  reg1644[(2'h2):(1'h1)] : reg1619[(4'hb):(2'h3)]) ?
                              $unsigned((forvar1622 * (8'hb0))) : (reg1598[(3'h4):(1'h0)] ?
                                  (reg1570 ?
                                      reg1550 : forvar1637) : $unsigned(reg1615))) : (reg1615[(3'h4):(1'h1)] ^~ $signed((~|reg1607))));
                      reg1662 <= (reg1632[(4'hf):(1'h0)] ?
                          $unsigned(((~^forvar1593) >= forvar1612)) : (!forvar1582));
                    end
                end
              for (forvar1663 = (1'h0); (forvar1663 < (2'h2)); forvar1663 = (forvar1663 + (1'h1)))
                begin
                  if ((!$signed(((|forvar1625) ^ $signed(reg1598)))))
                    begin
                      reg1664 <= ($unsigned(forvar1582) ?
                          forvar1655[(2'h2):(1'h1)] : reg1637[(4'hc):(1'h0)]);
                      reg1665 <= ((((reg1599 ? reg1585 : (8'haf)) ?
                              $unsigned(reg1567) : $signed(forvar1574)) <<< (reg1551 ?
                              (8'haf) : {forvar1612})) ?
                          reg1601[(2'h2):(2'h2)] : (!$signed((!(8'hae)))));
                      reg1666 <= forvar1593;
                    end
                  else
                    begin
                      reg1664 <= ($signed(reg1645[(1'h1):(1'h0)]) ~^ (8'hba));
                    end
                  reg1667 <= $unsigned(($unsigned($unsigned(reg1594)) ?
                      $unsigned(reg1604[(3'h4):(2'h3)]) : reg1661[(4'ha):(4'ha)]));
                end
            end
        end
      else
        begin
          for (forvar1624 = (1'h0); (forvar1624 < (2'h2)); forvar1624 = (forvar1624 + (1'h1)))
            begin
              reg1625 <= $unsigned((8'hb9));
              reg1626 <= (^~{(8'ha4)});
            end
          for (forvar1627 = (1'h0); (forvar1627 < (2'h3)); forvar1627 = (forvar1627 + (1'h1)))
            begin
              if (((~|(reg1564 >>> {reg1605})) ?
                  $signed(reg1635[(3'h4):(1'h1)]) : $unsigned(wire1538[(2'h2):(1'h1)])))
                begin
                  for (forvar1628 = (1'h0); (forvar1628 < (2'h3)); forvar1628 = (forvar1628 + (1'h1)))
                    begin
                      reg1629 <= $unsigned((^((~reg1626) ~^ (reg1554 == reg1542))));
                      reg1630 <= (8'hb4);
                    end
                  if ((+(($signed(forvar1633) ^ (reg1554 <= reg1641)) ~^ $signed((8'ha8)))))
                    begin
                      reg1631 <= reg1629;
                      reg1632 <= $signed($signed(forvar1625));
                    end
                  else
                    begin
                      reg1631 <= (8'h9f);
                      reg1632 <= reg1575[(4'h9):(3'h5)];
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h3)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= $unsigned((~|((reg1644 ? (8'ha5) : reg1654) ?
                          wire1538[(4'hc):(4'h8)] : (reg1637 ?
                              reg1630 : reg1560))));
                      reg1635 <= ($unsigned(forvar1641[(1'h1):(1'h0)]) ^~ reg1562);
                      reg1636 <= $signed((forvar1542[(1'h0):(1'h0)] != {(|reg1655)}));
                    end
                end
              else
                begin
                  reg1628 <= ($unsigned((~^((8'hac) ?
                      reg1636 : (8'hac)))) ^~ forvar1557);
                  for (forvar1629 = (1'h0); (forvar1629 < (1'h0)); forvar1629 = (forvar1629 + (1'h1)))
                    begin
                      reg1630 <= $signed(reg1586[(3'h5):(2'h2)]);
                      reg1631 <= reg1611;
                    end
                  for (forvar1632 = (1'h0); (forvar1632 < (2'h2)); forvar1632 = (forvar1632 + (1'h1)))
                    begin
                      reg1633 <= $signed({(~|$signed(reg1552))});
                      reg1634 <= forvar1608[(3'h7):(2'h2)];
                    end
                end
            end
          if ((8'haa))
            begin
              if ($unsigned($signed((~$unsigned(reg1658)))))
                begin
                  if (reg1603)
                    begin
                      reg1637 <= ($signed(reg1598) ?
                          reg1576[(3'h5):(2'h2)] : $unsigned(forvar1637));
                      reg1638 <= reg1660;
                      reg1639 <= (((~|reg1544[(2'h3):(2'h3)]) ?
                          ((forvar1557 <= (8'hb6)) >> $signed(reg1635)) : $unsigned(forvar1642)) ~^ (reg1559 ?
                          (!$signed(reg1630)) : (-$signed(reg1543))));
                    end
                  else
                    begin
                      reg1637 <= $signed((($unsigned(reg1554) != {reg1665}) >>> ({reg1560} ?
                          (reg1620 * forvar1637) : (reg1620 - reg1576))));
                      reg1638 <= forvar1637;
                    end
                end
              else
                begin
                  reg1637 <= reg1642;
                  reg1638 <= (reg1667[(4'hb):(2'h3)] <= (reg1633[(1'h0):(1'h0)] == ($signed(forvar1637) && $unsigned(reg1594))));
                  if ((^$signed($signed(reg1627))))
                    begin
                      reg1639 <= (reg1651[(3'h4):(2'h3)] > (($signed(forvar1612) >> (+forvar1612)) ?
                          reg1589 : ({wire1538} | $signed((8'h9f)))));
                      reg1640 <= ($unsigned(((reg1650 ?
                              reg1637 : forvar1593) <<< (reg1552 > reg1625))) ?
                          $unsigned(reg1658[(3'h5):(1'h0)]) : $signed($unsigned(wire1538)));
                    end
                  else
                    begin
                      reg1639 <= $signed(forvar1557[(3'h4):(1'h0)]);
                      reg1640 <= (^~$signed(reg1623));
                      reg1641 <= reg1661[(3'h5):(3'h5)];
                    end
                  reg1642 <= reg1571;
                end
              if ($unsigned(reg1598))
                begin
                  for (forvar1643 = (1'h0); (forvar1643 < (2'h3)); forvar1643 = (forvar1643 + (1'h1)))
                    begin
                      reg1644 <= ((reg1640[(1'h0):(1'h0)] ?
                          reg1555 : {(reg1571 > forvar1628)}) == ($signed(((8'ha9) ?
                              wire1536 : reg1581)) ?
                          (forvar1627[(2'h2):(2'h2)] ?
                              (!forvar1592) : $signed(reg1615)) : {(forvar1655 | reg1611)}));
                      reg1645 <= reg1543;
                      reg1646 <= {reg1654};
                    end
                  if ((8'hb7))
                    begin
                      reg1647 <= reg1548;
                      reg1648 <= ((^forvar1642[(1'h0):(1'h0)]) ?
                          (({(8'ha7)} - $signed(reg1602)) ^~ (reg1571[(2'h3):(1'h1)] != $signed(reg1648))) : $unsigned(forvar1643[(1'h0):(1'h0)]));
                      reg1649 <= reg1667;
                    end
                  else
                    begin
                      reg1647 <= reg1547[(2'h3):(1'h1)];
                      reg1648 <= (forvar1625[(2'h3):(2'h3)] ?
                          {(+$signed(reg1590))} : (^~reg1660[(2'h3):(2'h2)]));
                      reg1649 <= {(+reg1653[(3'h6):(1'h1)])};
                    end
                  if (($signed(forvar1617[(3'h6):(3'h6)]) ?
                      (-$signed((forvar1574 ?
                          (8'had) : reg1567))) : (~forvar1655)))
                    begin
                      reg1650 <= (8'hac);
                      reg1651 <= $unsigned(reg1621);
                    end
                  else
                    begin
                      reg1650 <= (&(|$unsigned(wire1536)));
                      reg1651 <= ({reg1569} & $unsigned(((reg1643 ?
                          reg1542 : reg1652) ~^ reg1610)));
                      reg1652 <= forvar1633;
                    end
                end
              else
                begin
                  reg1643 <= reg1600[(4'he):(4'hc)];
                  for (forvar1644 = (1'h0); (forvar1644 < (2'h2)); forvar1644 = (forvar1644 + (1'h1)))
                    begin
                      reg1645 <= reg1657;
                    end
                  reg1646 <= reg1627[(3'h7):(1'h1)];
                  for (forvar1647 = (1'h0); (forvar1647 < (2'h2)); forvar1647 = (forvar1647 + (1'h1)))
                    begin
                      reg1648 <= ($unsigned({$unsigned(forvar1587)}) ?
                          reg1644 : (8'hab));
                      reg1649 <= (|(reg1639[(4'h9):(4'h8)] ?
                          reg1636 : (+(forvar1629 ^ reg1555))));
                    end
                end
            end
          else
            begin
              reg1637 <= (($unsigned($signed(reg1584)) & (-(-forvar1540))) ?
                  reg1545[(2'h3):(2'h2)] : reg1595[(2'h3):(2'h2)]);
              for (forvar1638 = (1'h0); (forvar1638 < (1'h1)); forvar1638 = (forvar1638 + (1'h1)))
                begin
                  for (forvar1639 = (1'h0); (forvar1639 < (1'h0)); forvar1639 = (forvar1639 + (1'h1)))
                    begin
                      reg1640 <= wire1536[(2'h2):(1'h0)];
                      reg1641 <= reg1645[(1'h1):(1'h0)];
                      reg1642 <= ((^~(forvar1593[(3'h7):(3'h5)] << {reg1583})) ?
                          reg1647 : reg1641);
                      reg1643 <= forvar1632[(1'h0):(1'h0)];
                    end
                end
              if ($unsigned(wire1536))
                begin
                  for (forvar1644 = (1'h0); (forvar1644 < (1'h0)); forvar1644 = (forvar1644 + (1'h1)))
                    begin
                      reg1645 <= forvar1632;
                      reg1646 <= reg1640[(3'h6):(2'h3)];
                      reg1647 <= $signed(reg1555[(2'h3):(2'h2)]);
                      reg1648 <= ((+forvar1579[(4'h8):(2'h3)]) ?
                          $signed({forvar1632[(2'h2):(1'h1)]}) : wire1538);
                    end
                  if ($signed((8'hb4)))
                    begin
                      reg1649 <= ((^~$signed($signed(reg1646))) << (wire1533[(4'ha):(4'ha)] & ((+reg1667) ?
                          $signed(forvar1546) : (reg1581 >= reg1568))));
                      reg1650 <= (~&$signed((^~(reg1640 ?
                          reg1611 : forvar1592))));
                      reg1651 <= (($unsigned({(8'ha2)}) ~^ (&$signed((8'haa)))) ^~ $signed(forvar1638[(3'h6):(3'h5)]));
                      reg1652 <= {{reg1584[(4'ha):(2'h2)]}};
                    end
                  else
                    begin
                      reg1649 <= $unsigned(reg1619);
                    end
                  for (forvar1653 = (1'h0); (forvar1653 < (2'h2)); forvar1653 = (forvar1653 + (1'h1)))
                    begin
                      reg1654 <= $signed(({(forvar1642 ?
                              (8'hb9) : forvar1541)} >= reg1568[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  if ((((reg1568 ~^ (-(8'h9e))) ?
                      $unsigned((&forvar1541)) : reg1656[(1'h1):(1'h0)]) <= $signed($unsigned($signed(reg1667)))))
                    begin
                      reg1644 <= $signed(forvar1646);
                      reg1645 <= (reg1638 ?
                          wire1535 : ((~^(wire1537 >> reg1654)) ?
                              forvar1542 : reg1651));
                      reg1646 <= (^$unsigned(forvar1553));
                    end
                  else
                    begin
                      reg1644 <= {({forvar1541} ?
                              $signed((8'hae)) : ((reg1594 ?
                                      wire1536 : (8'hb3)) ?
                                  reg1603 : (reg1610 <<< reg1635)))};
                      reg1645 <= {(reg1644[(1'h1):(1'h1)] ?
                              (8'hb8) : reg1600[(4'hb):(4'h8)])};
                      reg1646 <= $unsigned($signed({(8'hb4)}));
                      reg1647 <= $unsigned(reg1584[(3'h7):(1'h1)]);
                    end
                  for (forvar1648 = (1'h0); (forvar1648 < (1'h1)); forvar1648 = (forvar1648 + (1'h1)))
                    begin
                      reg1649 <= reg1638;
                      reg1650 <= wire1533;
                      reg1651 <= $signed(reg1548[(3'h6):(3'h5)]);
                    end
                  if ($signed((~|forvar1648)))
                    begin
                      reg1652 <= {reg1547[(2'h3):(2'h3)]};
                      reg1653 <= {(^~((^(8'ha3)) != $signed(reg1552)))};
                      reg1654 <= {($unsigned((forvar1641 ?
                              wire1536 : (8'haf))) == (!forvar1597))};
                      reg1655 <= reg1590;
                    end
                  else
                    begin
                      reg1652 <= (forvar1542[(1'h1):(1'h0)] ?
                          $signed({{forvar1625}}) : $unsigned(((reg1594 == reg1600) >> {forvar1624})));
                      reg1653 <= ($signed((~&wire1534)) ?
                          {$signed($unsigned(forvar1541))} : reg1639);
                      reg1654 <= {$unsigned($signed({reg1639}))};
                    end
                  if ((8'ha3))
                    begin
                      reg1656 <= ($unsigned((!reg1569[(3'h6):(1'h1)])) ?
                          $unsigned(((forvar1592 ?
                              reg1583 : forvar1646) > (reg1643 ?
                              (8'ha7) : reg1590))) : forvar1637);
                      reg1657 <= (reg1667[(3'h6):(3'h4)] > (~&({forvar1653} < $signed(forvar1622))));
                      reg1658 <= reg1542;
                    end
                  else
                    begin
                      reg1656 <= $signed(reg1639[(4'ha):(3'h6)]);
                      reg1657 <= forvar1643[(2'h2):(1'h0)];
                    end
                end
              reg1659 <= (((|(~|(8'hb0))) * (|(reg1570 ?
                  reg1602 : reg1563))) & reg1662[(1'h1):(1'h0)]);
            end
        end
      for (forvar1668 = (1'h0); (forvar1668 < (2'h2)); forvar1668 = (forvar1668 + (1'h1)))
        begin
          reg1669 <= $signed(($unsigned((reg1652 | forvar1608)) ?
              forvar1622[(3'h6):(1'h1)] : forvar1643[(2'h3):(1'h1)]));
          if ($unsigned(reg1614[(1'h1):(1'h1)]))
            begin
              for (forvar1670 = (1'h0); (forvar1670 < (1'h0)); forvar1670 = (forvar1670 + (1'h1)))
                begin
                  for (forvar1671 = (1'h0); (forvar1671 < (2'h2)); forvar1671 = (forvar1671 + (1'h1)))
                    begin
                      reg1672 <= (^(forvar1587 || (~&$unsigned((8'hb0)))));
                      reg1673 <= $unsigned($unsigned(((reg1664 == forvar1655) ?
                          reg1548[(3'h5):(2'h3)] : $unsigned(reg1649))));
                    end
                  for (forvar1674 = (1'h0); (forvar1674 < (1'h0)); forvar1674 = (forvar1674 + (1'h1)))
                    begin
                      reg1675 <= $unsigned($unsigned(wire1533));
                      reg1676 <= (8'ha8);
                      reg1677 <= $signed(($unsigned(((8'hae) ?
                          reg1551 : reg1575)) * forvar1566[(4'h9):(4'h9)]));
                    end
                  if ($signed($signed($unsigned($unsigned(reg1675)))))
                    begin
                      reg1678 <= reg1640;
                      reg1679 <= {((reg1559 >>> ((8'ha7) ?
                              (8'hac) : (8'hb3))) <= reg1675)};
                      reg1680 <= reg1634[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg1678 <= forvar1628[(1'h1):(1'h0)];
                    end
                end
              if (forvar1671)
                begin
                  if ($signed(((~(reg1649 + reg1542)) - ({reg1643} ?
                      $unsigned(reg1586) : $unsigned(reg1620)))))
                    begin
                      reg1681 <= $signed(((|$signed(reg1666)) - ((-(8'hb4)) == forvar1642[(3'h4):(2'h3)])));
                      reg1682 <= $signed(({$unsigned(reg1604)} ?
                          ((forvar1593 && reg1558) ?
                              (reg1550 ?
                                  forvar1633 : reg1547) : forvar1648[(3'h7):(2'h3)]) : ((reg1638 * reg1645) << reg1675[(2'h2):(2'h2)])));
                      reg1683 <= reg1632[(2'h3):(2'h2)];
                      reg1684 <= (|$unsigned(reg1544));
                    end
                  else
                    begin
                      reg1681 <= reg1647[(4'hd):(1'h0)];
                      reg1682 <= (8'hb5);
                    end
                  for (forvar1685 = (1'h0); (forvar1685 < (1'h0)); forvar1685 = (forvar1685 + (1'h1)))
                    begin
                      reg1686 <= $unsigned(wire1538);
                      reg1687 <= ($unsigned(((+reg1675) ?
                          $unsigned(reg1606) : (~reg1558))) >> $signed({reg1556[(2'h2):(2'h2)]}));
                      reg1688 <= (reg1645[(2'h3):(1'h0)] ?
                          (reg1644[(2'h3):(1'h1)] ~^ reg1681) : reg1590[(3'h6):(1'h1)]);
                    end
                end
              else
                begin
                  if ($unsigned(reg1645))
                    begin
                      reg1681 <= {((!$unsigned((8'hae))) ?
                              ($unsigned(reg1542) ^~ {reg1619}) : (((8'hb1) != forvar1653) ^ $signed(forvar1648)))};
                      reg1682 <= forvar1622;
                      reg1683 <= (+$signed($unsigned(reg1563[(3'h6):(3'h6)])));
                    end
                  else
                    begin
                      reg1681 <= (8'ha2);
                    end
                  for (forvar1684 = (1'h0); (forvar1684 < (1'h1)); forvar1684 = (forvar1684 + (1'h1)))
                    begin
                      reg1685 <= $signed(({(~^forvar1588)} ^~ reg1602));
                    end
                  reg1686 <= forvar1618[(3'h4):(2'h2)];
                end
            end
          else
            begin
              if ((8'ha9))
                begin
                  reg1670 <= reg1688;
                end
              else
                begin
                  if ({$unsigned((&(forvar1633 >= reg1688)))})
                    begin
                      reg1670 <= $unsigned((8'ha3));
                      reg1671 <= (reg1644[(4'hd):(3'h4)] | reg1638[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg1670 <= $unsigned($unsigned(reg1664[(2'h2):(1'h1)]));
                      reg1671 <= (!$unsigned(((|reg1590) | reg1599)));
                      reg1672 <= reg1688[(3'h4):(2'h3)];
                      reg1673 <= $signed(((+reg1542) ?
                          $signed($unsigned(reg1585)) : forvar1663));
                    end
                  for (forvar1674 = (1'h0); (forvar1674 < (1'h0)); forvar1674 = (forvar1674 + (1'h1)))
                    begin
                      reg1675 <= $signed(((reg1636[(2'h2):(1'h1)] ?
                          (^~reg1602) : $signed((8'hba))) | $unsigned((reg1629 && reg1609))));
                      reg1676 <= reg1616;
                      reg1677 <= $signed($signed(reg1564[(4'he):(4'hd)]));
                    end
                end
            end
        end
      for (forvar1689 = (1'h0); (forvar1689 < (2'h2)); forvar1689 = (forvar1689 + (1'h1)))
        begin
          for (forvar1690 = (1'h0); (forvar1690 < (1'h0)); forvar1690 = (forvar1690 + (1'h1)))
            begin
              for (forvar1691 = (1'h0); (forvar1691 < (1'h0)); forvar1691 = (forvar1691 + (1'h1)))
                begin
                  for (forvar1692 = (1'h0); (forvar1692 < (1'h1)); forvar1692 = (forvar1692 + (1'h1)))
                    begin
                      reg1693 <= $unsigned({(+(reg1666 ? reg1639 : reg1653))});
                      reg1694 <= $signed(($unsigned((forvar1670 ?
                              forvar1624 : (8'hb4))) ?
                          forvar1637 : reg1594[(2'h3):(1'h0)]));
                    end
                end
              reg1695 <= $signed(({$signed(reg1611)} ?
                  (^~(forvar1542 - (8'hb3))) : $unsigned($unsigned(reg1640))));
              if (reg1552[(3'h5):(3'h4)])
                begin
                  for (forvar1696 = (1'h0); (forvar1696 < (1'h1)); forvar1696 = (forvar1696 + (1'h1)))
                    begin
                      reg1697 <= $unsigned($unsigned(reg1673));
                      reg1698 <= $signed(((reg1638[(3'h5):(2'h2)] <= wire1539) << $unsigned($unsigned(reg1631))));
                      reg1699 <= (8'hb7);
                      reg1700 <= $unsigned((^~reg1611[(2'h2):(1'h1)]));
                    end
                  if (reg1577[(1'h0):(1'h0)])
                    begin
                      reg1701 <= (forvar1622 ?
                          $signed(($signed(reg1688) ?
                              (reg1573 | (8'ha8)) : (reg1695 ?
                                  forvar1671 : reg1611))) : (|(reg1614 ?
                              reg1580[(4'ha):(3'h4)] : (~&reg1605))));
                      reg1702 <= ({({forvar1617} * (wire1533 << reg1609))} ?
                          reg1637[(4'h9):(1'h0)] : ((&reg1591[(1'h0):(1'h0)]) + reg1542[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg1701 <= {reg1631[(2'h3):(1'h0)]};
                    end
                end
              else
                begin
                  if ($signed(reg1642))
                    begin
                      reg1696 <= (~$unsigned(forvar1574[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1696 <= ($unsigned(forvar1633[(3'h7):(3'h6)]) - (((reg1687 ?
                              reg1570 : forvar1542) ?
                          reg1606[(3'h7):(3'h7)] : (reg1600 && wire1538)) >> reg1669[(4'hf):(4'hf)]));
                      reg1697 <= ($signed(reg1578) > forvar1633);
                      reg1698 <= reg1637;
                      reg1699 <= (~^reg1653);
                    end
                  if (forvar1639)
                    begin
                      reg1700 <= (reg1547 <<< ((~&reg1611) ?
                          forvar1627 : ((reg1598 ? forvar1582 : (8'hb3)) ?
                              $signed(forvar1624) : {forvar1670})));
                      reg1701 <= ({($signed(reg1680) >= $unsigned(reg1696))} - $signed($signed($unsigned(reg1552))));
                    end
                  else
                    begin
                      reg1700 <= {reg1636};
                      reg1701 <= (-(8'hb1));
                    end
                  for (forvar1702 = (1'h0); (forvar1702 < (1'h1)); forvar1702 = (forvar1702 + (1'h1)))
                    begin
                      reg1703 <= $unsigned($unsigned(((reg1654 ?
                              reg1683 : reg1577) ?
                          reg1658 : (reg1609 ? forvar1540 : wire1534))));
                      reg1704 <= (($signed($unsigned((8'ha5))) && reg1682[(4'h8):(3'h5)]) ?
                          reg1591 : forvar1659[(2'h3):(1'h0)]);
                      reg1705 <= $unsigned($unsigned(reg1563));
                    end
                end
              if ($unsigned($unsigned($signed($unsigned(wire1538)))))
                begin
                  if ((~|reg1544))
                    begin
                      reg1706 <= $signed($unsigned(reg1656[(1'h0):(1'h0)]));
                      reg1707 <= {reg1577};
                    end
                  else
                    begin
                      reg1706 <= $unsigned(($signed((+reg1601)) <= reg1672[(4'he):(4'h8)]));
                      reg1707 <= $signed(($signed({reg1573}) - (~reg1626)));
                      reg1708 <= $unsigned(forvar1668[(3'h5):(3'h5)]);
                    end
                  reg1709 <= ($signed({{(8'haa)}}) ^ ((&(~|reg1579)) ?
                      ((reg1682 ?
                          (8'had) : (8'ha8)) ^~ $unsigned(reg1596)) : $unsigned((reg1577 && reg1595))));
                  for (forvar1710 = (1'h0); (forvar1710 < (1'h1)); forvar1710 = (forvar1710 + (1'h1)))
                    begin
                      reg1711 <= (^~$signed(({reg1586} ?
                          (~reg1670) : $signed(forvar1668))));
                      reg1712 <= forvar1546[(3'h4):(1'h1)];
                    end
                end
              else
                begin
                  if (forvar1618[(3'h6):(2'h2)])
                    begin
                      reg1706 <= $signed(forvar1685[(4'hd):(3'h6)]);
                      reg1707 <= reg1658[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1706 <= (reg1637[(4'ha):(1'h0)] + reg1550[(4'hd):(4'h9)]);
                      reg1707 <= $unsigned($unsigned(reg1576[(1'h0):(1'h0)]));
                      reg1708 <= (reg1542 ?
                          {{reg1702}} : ($signed((|reg1602)) ?
                              {(8'ha7)} : ($unsigned((8'hab)) ?
                                  (+reg1565) : $unsigned(reg1547))));
                      reg1709 <= (+(reg1684 * $unsigned(reg1708[(1'h0):(1'h0)])));
                    end
                end
            end
          for (forvar1713 = (1'h0); (forvar1713 < (1'h0)); forvar1713 = (forvar1713 + (1'h1)))
            begin
              if (forvar1541[(3'h4):(1'h0)])
                begin
                  for (forvar1714 = (1'h0); (forvar1714 < (2'h2)); forvar1714 = (forvar1714 + (1'h1)))
                    begin
                      reg1715 <= (~$signed($signed($signed(reg1551))));
                      reg1716 <= (((forvar1612 + $unsigned(reg1627)) ?
                              (+reg1679) : (8'hb2)) ?
                          $unsigned(($unsigned(reg1616) | $signed(forvar1647))) : reg1568);
                      reg1717 <= $unsigned($signed({(forvar1557 ?
                              reg1626 : reg1620)}));
                    end
                  if ($unsigned((^$unsigned(((8'ha8) ? (8'hb7) : forvar1713)))))
                    begin
                      reg1718 <= $unsigned({(+{wire1536})});
                      reg1719 <= ({reg1671[(1'h1):(1'h1)]} ?
                          $unsigned((-(reg1709 ?
                              (8'ha6) : (8'ha8)))) : (8'h9e));
                      reg1720 <= reg1680;
                      reg1721 <= {{$unsigned(forvar1587)}};
                    end
                  else
                    begin
                      reg1718 <= $signed($unsigned(reg1549));
                      reg1719 <= (^~reg1696);
                      reg1720 <= $signed(($unsigned($unsigned(forvar1546)) >>> forvar1608));
                    end
                  for (forvar1722 = (1'h0); (forvar1722 < (2'h2)); forvar1722 = (forvar1722 + (1'h1)))
                    begin
                      reg1723 <= (({(-reg1704)} >= $unsigned($unsigned(reg1655))) <= (~(reg1639 ^~ (!(8'ha7)))));
                      reg1724 <= forvar1663;
                      reg1725 <= reg1665[(3'h4):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar1714 = (1'h0); (forvar1714 < (2'h2)); forvar1714 = (forvar1714 + (1'h1)))
                    begin
                      reg1715 <= ((((reg1632 ?
                              (8'hb2) : reg1699) || $unsigned(reg1580)) ~^ (!$unsigned((8'hb2)))) ?
                          reg1559 : $signed($unsigned((+reg1552))));
                      reg1716 <= ($signed(($signed((8'ha8)) & (!forvar1572))) ?
                          $signed({$unsigned(reg1647)}) : (^~$unsigned((forvar1557 ?
                              reg1687 : (8'ha6)))));
                      reg1717 <= $signed(forvar1655);
                    end
                  for (forvar1718 = (1'h0); (forvar1718 < (2'h3)); forvar1718 = (forvar1718 + (1'h1)))
                    begin
                      reg1719 <= $unsigned({({reg1649} ^~ {reg1698})});
                      reg1720 <= (~{((!reg1654) ?
                              (forvar1684 ?
                                  reg1596 : (8'h9e)) : reg1581[(3'h4):(1'h0)])});
                    end
                  reg1721 <= reg1629;
                  for (forvar1722 = (1'h0); (forvar1722 < (1'h0)); forvar1722 = (forvar1722 + (1'h1)))
                    begin
                      reg1723 <= reg1571;
                    end
                end
            end
          for (forvar1726 = (1'h0); (forvar1726 < (2'h2)); forvar1726 = (forvar1726 + (1'h1)))
            begin
              for (forvar1727 = (1'h0); (forvar1727 < (1'h1)); forvar1727 = (forvar1727 + (1'h1)))
                begin
                  if ((reg1589[(1'h0):(1'h0)] << {(reg1708[(1'h0):(1'h0)] ?
                          $signed(forvar1710) : ((8'ha6) ?
                              forvar1659 : reg1594))}))
                    begin
                      reg1728 <= reg1631[(3'h6):(3'h6)];
                      reg1729 <= $unsigned(({(~^reg1629)} <= reg1552));
                    end
                  else
                    begin
                      reg1728 <= $signed({{reg1680[(3'h4):(1'h0)]}});
                      reg1729 <= ($unsigned(forvar1702[(1'h1):(1'h1)]) | reg1570[(4'h9):(3'h6)]);
                    end
                end
              reg1730 <= (reg1652 ? reg1718 : {{reg1571[(1'h1):(1'h1)]}});
              reg1731 <= $unsigned(forvar1702[(2'h2):(1'h1)]);
              for (forvar1732 = (1'h0); (forvar1732 < (1'h1)); forvar1732 = (forvar1732 + (1'h1)))
                begin
                  reg1733 <= (reg1564[(4'h8):(1'h1)] < ((((8'haf) ~^ reg1577) ?
                          (reg1662 ? reg1590 : reg1602) : {wire1539}) ?
                      $unsigned((reg1603 | reg1643)) : reg1628[(4'h8):(4'h8)]));
                end
            end
        end
    end
  assign wire1734 = reg1662[(4'h9):(4'h8)];
  assign wire1735 = (8'hb3);
  assign wire1736 = ((8'hb8) ? (8'had) : reg1684[(3'h4):(1'h0)]);
  assign wire1737 = (~|reg1551[(5'h10):(3'h4)]);
  assign wire1738 = ($unsigned(((^~forvar1649) ?
                            $signed((8'ha2)) : {reg1616})) ?
                        $unsigned($signed((^~reg1733))) : reg1675);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3039  (y, clk, wire3040, wire3041, wire3042, wire3043, wire3044);
  output wire [(32'ha3b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire3040;
  input wire [(4'hf):(1'h0)] wire3041;
  input wire [(5'h10):(1'h0)] wire3042;
  input wire [(3'h7):(1'h0)] wire3043;
  input wire signed [(2'h3):(1'h0)] wire3044;
  reg [(4'hd):(1'h0)] reg3528 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3527 = (1'h0);
  reg [(4'he):(1'h0)] reg3526 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3525 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3524 = (1'h0);
  reg [(2'h2):(1'h0)] reg3523 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3522 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3521 = (1'h0);
  reg [(3'h4):(1'h0)] reg3520 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3519 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3518 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3517 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3516 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3515 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3514 = (1'h0);
  reg [(4'he):(1'h0)] reg3513 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3512 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3511 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3510 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3509 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3508 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3507 = (1'h0);
  reg [(4'ha):(1'h0)] reg3506 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3501 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3505 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3504 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3503 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3502 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3501 = (1'h0);
  reg [(3'h4):(1'h0)] reg3500 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3499 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3498 = (1'h0);
  reg [(3'h6):(1'h0)] reg3497 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3496 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3495 = (1'h0);
  reg [(4'hb):(1'h0)] reg3494 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3493 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3492 = (1'h0);
  reg [(4'he):(1'h0)] forvar3491 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3490 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3489 = (1'h0);
  reg [(4'h8):(1'h0)] reg3488 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3487 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3486 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3485 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3484 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3483 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3477 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3474 = (1'h0);
  reg [(4'hd):(1'h0)] reg3472 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3470 = (1'h0);
  reg [(2'h3):(1'h0)] reg3482 = (1'h0);
  reg [(3'h6):(1'h0)] reg3481 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3480 = (1'h0);
  reg [(4'hc):(1'h0)] reg3479 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3478 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3477 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3476 = (1'h0);
  reg [(4'h8):(1'h0)] reg3475 = (1'h0);
  reg [(4'hd):(1'h0)] reg3474 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3473 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3472 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3471 = (1'h0);
  reg [(4'hc):(1'h0)] reg3470 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3469 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3468 = (1'h0);
  reg [(3'h7):(1'h0)] reg3467 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3466 = (1'h0);
  reg [(2'h2):(1'h0)] reg3465 = (1'h0);
  reg [(4'he):(1'h0)] reg3464 = (1'h0);
  reg [(4'ha):(1'h0)] reg3463 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3462 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3461 = (1'h0);
  reg [(3'h7):(1'h0)] reg3460 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3457 = (1'h0);
  reg [(4'hf):(1'h0)] reg3459 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3458 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3457 = (1'h0);
  reg [(2'h3):(1'h0)] reg3456 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3455 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3454 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3453 = (1'h0);
  reg [(3'h5):(1'h0)] reg3452 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3451 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3450 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3449 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3448 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3447 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3446 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3445 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3444 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3443 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3435 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3429 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3428 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3425 = (1'h0);
  reg [(4'ha):(1'h0)] reg3423 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3420 = (1'h0);
  reg [(2'h3):(1'h0)] reg3419 = (1'h0);
  reg [(2'h2):(1'h0)] reg3416 = (1'h0);
  reg [(5'h10):(1'h0)] reg3436 = (1'h0);
  reg [(4'he):(1'h0)] reg3442 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3441 = (1'h0);
  reg [(4'hf):(1'h0)] reg3440 = (1'h0);
  reg [(5'h10):(1'h0)] reg3439 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3438 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3437 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3436 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3435 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3434 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3433 = (1'h0);
  reg [(4'he):(1'h0)] reg3432 = (1'h0);
  reg [(4'he):(1'h0)] reg3431 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3430 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3429 = (1'h0);
  reg [(4'ha):(1'h0)] reg3428 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3427 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3426 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3425 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3424 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3423 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3422 = (1'h0);
  reg [(2'h2):(1'h0)] reg3421 = (1'h0);
  reg [(4'hb):(1'h0)] reg3420 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3419 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3418 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3417 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3416 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3415 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3405 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3404 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3403 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3414 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3413 = (1'h0);
  reg [(4'hf):(1'h0)] reg3412 = (1'h0);
  reg [(4'hc):(1'h0)] reg3411 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3410 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3398 = (1'h0);
  reg [(4'hb):(1'h0)] reg3409 = (1'h0);
  reg [(4'hf):(1'h0)] reg3408 = (1'h0);
  reg [(3'h5):(1'h0)] reg3407 = (1'h0);
  reg [(4'ha):(1'h0)] reg3406 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3405 = (1'h0);
  reg [(3'h4):(1'h0)] reg3404 = (1'h0);
  reg [(4'hf):(1'h0)] reg3403 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3401 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3391 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3394 = (1'h0);
  reg [(2'h3):(1'h0)] reg3392 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3390 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3383 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3382 = (1'h0);
  reg [(4'h9):(1'h0)] reg3378 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3375 = (1'h0);
  reg [(3'h5):(1'h0)] reg3402 = (1'h0);
  reg [(4'h8):(1'h0)] reg3401 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3400 = (1'h0);
  reg [(2'h3):(1'h0)] reg3399 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3398 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3397 = (1'h0);
  reg [(3'h4):(1'h0)] reg3396 = (1'h0);
  reg [(3'h4):(1'h0)] reg3395 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3394 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3393 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3392 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3391 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3390 = (1'h0);
  reg [(2'h3):(1'h0)] reg3389 = (1'h0);
  reg [(4'hf):(1'h0)] reg3388 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3387 = (1'h0);
  reg [(4'ha):(1'h0)] reg3386 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3385 = (1'h0);
  reg [(3'h4):(1'h0)] reg3384 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3383 = (1'h0);
  reg [(3'h7):(1'h0)] reg3382 = (1'h0);
  reg [(4'hb):(1'h0)] reg3381 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3380 = (1'h0);
  reg [(5'h10):(1'h0)] reg3379 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3378 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3377 = (1'h0);
  reg [(3'h7):(1'h0)] reg3376 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3375 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3374 = (1'h0);
  reg [(4'hf):(1'h0)] reg3373 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3372 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire3371;
  wire signed [(2'h2):(1'h0)] wire3370;
  wire signed [(3'h4):(1'h0)] wire3369;
  wire signed [(3'h5):(1'h0)] wire3368;
  wire [(4'hc):(1'h0)] wire3045;
  wire signed [(4'he):(1'h0)] wire3046;
  wire [(4'he):(1'h0)] wire3047;
  wire [(4'h8):(1'h0)] wire3048;
  reg signed [(4'hc):(1'h0)] reg3049 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3050 = (1'h0);
  reg [(4'h8):(1'h0)] reg3051 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3050 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3052 = (1'h0);
  reg [(4'h8):(1'h0)] reg3053 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3054 = (1'h0);
  reg [(4'he):(1'h0)] reg3055 = (1'h0);
  reg [(4'h8):(1'h0)] reg3056 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3057 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3058 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3059 = (1'h0);
  reg [(4'h9):(1'h0)] reg3060 = (1'h0);
  reg [(3'h4):(1'h0)] reg3061 = (1'h0);
  reg [(4'h8):(1'h0)] reg3062 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3063 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3064 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3065 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3066 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3067 = (1'h0);
  reg [(4'hf):(1'h0)] reg3068 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3069 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3070 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3071 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3072 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3073 = (1'h0);
  reg [(3'h7):(1'h0)] reg3074 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3075 = (1'h0);
  reg [(3'h7):(1'h0)] reg3076 = (1'h0);
  reg [(2'h2):(1'h0)] reg3077 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3078 = (1'h0);
  reg [(3'h7):(1'h0)] reg3079 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3080 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3081 = (1'h0);
  reg [(2'h3):(1'h0)] reg3082 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3083 = (1'h0);
  reg [(4'h9):(1'h0)] reg3084 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3085 = (1'h0);
  reg [(4'he):(1'h0)] reg3086 = (1'h0);
  reg [(4'hf):(1'h0)] reg3087 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3088 = (1'h0);
  reg [(3'h5):(1'h0)] reg3089 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3090 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3091 = (1'h0);
  reg [(4'hb):(1'h0)] reg3092 = (1'h0);
  reg [(5'h10):(1'h0)] reg3093 = (1'h0);
  reg [(4'hf):(1'h0)] reg3094 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3095 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3081 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3082 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3085 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3087 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3088 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3091 = (1'h0);
  reg [(4'he):(1'h0)] reg3096 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3097 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3098 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3051 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3054 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3057 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3059 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3060 = (1'h0);
  reg [(3'h6):(1'h0)] reg3063 = (1'h0);
  reg [(4'h8):(1'h0)] reg3064 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3065 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3066 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3070 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3073 = (1'h0);
  reg [(4'he):(1'h0)] forvar3075 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3078 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3086 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3090 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3098 = (1'h0);
  reg [(3'h4):(1'h0)] reg3099 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3100 = (1'h0);
  reg [(3'h5):(1'h0)] reg3101 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3102 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3103 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3104 = (1'h0);
  reg [(4'ha):(1'h0)] reg3105 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3101 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3103 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3106 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3107 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3108 = (1'h0);
  reg [(3'h6):(1'h0)] reg3109 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3110 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3111 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3112 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3113 = (1'h0);
  reg [(3'h5):(1'h0)] reg3114 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3115 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3116 = (1'h0);
  wire [(4'hf):(1'h0)] wire3366;
  assign y = {reg3528,
                 reg3527,
                 reg3526,
                 reg3525,
                 forvar3524,
                 reg3523,
                 reg3522,
                 reg3521,
                 reg3520,
                 reg3519,
                 reg3518,
                 forvar3517,
                 forvar3516,
                 reg3515,
                 reg3514,
                 reg3513,
                 forvar3512,
                 reg3511,
                 forvar3510,
                 forvar3509,
                 forvar3508,
                 forvar3507,
                 reg3506,
                 reg3501,
                 reg3505,
                 forvar3504,
                 reg3503,
                 reg3502,
                 forvar3501,
                 reg3500,
                 reg3499,
                 reg3498,
                 reg3497,
                 reg3496,
                 forvar3495,
                 reg3494,
                 forvar3493,
                 reg3492,
                 forvar3491,
                 reg3490,
                 reg3489,
                 reg3488,
                 reg3487,
                 reg3486,
                 forvar3485,
                 forvar3484,
                 forvar3483,
                 reg3477,
                 forvar3474,
                 reg3472,
                 forvar3470,
                 reg3482,
                 reg3481,
                 reg3480,
                 reg3479,
                 reg3478,
                 forvar3477,
                 reg3476,
                 reg3475,
                 reg3474,
                 reg3473,
                 forvar3472,
                 forvar3471,
                 reg3470,
                 forvar3469,
                 reg3468,
                 reg3467,
                 forvar3466,
                 reg3465,
                 reg3464,
                 reg3463,
                 forvar3462,
                 reg3461,
                 reg3460,
                 forvar3457,
                 reg3459,
                 reg3458,
                 reg3457,
                 reg3456,
                 reg3455,
                 forvar3454,
                 forvar3453,
                 reg3452,
                 reg3451,
                 reg3450,
                 reg3449,
                 reg3448,
                 reg3447,
                 reg3446,
                 forvar3445,
                 forvar3444,
                 forvar3443,
                 forvar3435,
                 reg3429,
                 forvar3428,
                 forvar3425,
                 reg3423,
                 forvar3420,
                 reg3419,
                 reg3416,
                 reg3436,
                 reg3442,
                 reg3441,
                 reg3440,
                 reg3439,
                 reg3438,
                 reg3437,
                 forvar3436,
                 reg3435,
                 reg3434,
                 reg3433,
                 reg3432,
                 reg3431,
                 reg3430,
                 forvar3429,
                 reg3428,
                 reg3427,
                 reg3426,
                 reg3425,
                 reg3424,
                 forvar3423,
                 reg3422,
                 reg3421,
                 reg3420,
                 forvar3419,
                 reg3418,
                 reg3417,
                 forvar3416,
                 forvar3415,
                 reg3405,
                 forvar3404,
                 forvar3403,
                 reg3414,
                 reg3413,
                 reg3412,
                 reg3411,
                 forvar3410,
                 reg3398,
                 reg3409,
                 reg3408,
                 reg3407,
                 reg3406,
                 forvar3405,
                 reg3404,
                 reg3403,
                 forvar3401,
                 reg3391,
                 forvar3394,
                 reg3392,
                 reg3390,
                 reg3383,
                 forvar3382,
                 reg3378,
                 forvar3375,
                 reg3402,
                 reg3401,
                 reg3400,
                 reg3399,
                 forvar3398,
                 reg3397,
                 reg3396,
                 reg3395,
                 reg3394,
                 reg3393,
                 forvar3392,
                 forvar3391,
                 forvar3390,
                 reg3389,
                 reg3388,
                 reg3387,
                 reg3386,
                 reg3385,
                 reg3384,
                 forvar3383,
                 reg3382,
                 reg3381,
                 reg3380,
                 reg3379,
                 forvar3378,
                 reg3377,
                 reg3376,
                 reg3375,
                 forvar3374,
                 reg3373,
                 forvar3372,
                 wire3371,
                 wire3370,
                 wire3369,
                 wire3368,
                 wire3045,
                 wire3046,
                 wire3047,
                 wire3048,
                 reg3049,
                 reg3050,
                 reg3051,
                 forvar3050,
                 reg3052,
                 reg3053,
                 reg3054,
                 reg3055,
                 reg3056,
                 forvar3057,
                 reg3058,
                 reg3059,
                 reg3060,
                 reg3061,
                 reg3062,
                 forvar3063,
                 forvar3064,
                 reg3065,
                 reg3066,
                 reg3067,
                 reg3068,
                 reg3069,
                 forvar3070,
                 reg3071,
                 reg3072,
                 forvar3073,
                 reg3074,
                 reg3075,
                 reg3076,
                 reg3077,
                 reg3078,
                 reg3079,
                 reg3080,
                 forvar3081,
                 reg3082,
                 reg3083,
                 reg3084,
                 forvar3085,
                 reg3086,
                 reg3087,
                 forvar3088,
                 reg3089,
                 reg3090,
                 forvar3091,
                 reg3092,
                 reg3093,
                 reg3094,
                 reg3095,
                 reg3081,
                 forvar3082,
                 reg3085,
                 forvar3087,
                 reg3088,
                 reg3091,
                 reg3096,
                 reg3097,
                 reg3098,
                 forvar3051,
                 forvar3054,
                 reg3057,
                 forvar3059,
                 forvar3060,
                 reg3063,
                 reg3064,
                 forvar3065,
                 forvar3066,
                 reg3070,
                 reg3073,
                 forvar3075,
                 forvar3078,
                 forvar3086,
                 forvar3090,
                 forvar3098,
                 reg3099,
                 reg3100,
                 reg3101,
                 reg3102,
                 forvar3103,
                 reg3104,
                 reg3105,
                 forvar3101,
                 reg3103,
                 forvar3106,
                 forvar3107,
                 reg3108,
                 reg3109,
                 reg3110,
                 reg3111,
                 reg3112,
                 reg3113,
                 reg3114,
                 reg3115,
                 reg3116,
                 wire3366,
                 (1'h0)};
  assign wire3045 = (wire3041[(4'ha):(4'ha)] ?
                        wire3043 : $unsigned($unsigned(wire3042[(4'h9):(3'h6)])));
  assign wire3046 = (|{(-(wire3042 <<< wire3040))});
  assign wire3047 = ({(~(wire3046 ? wire3046 : wire3040))} ?
                        $signed(wire3043) : (({wire3046} >>> wire3045) ?
                            $unsigned((-wire3045)) : $unsigned(((8'haa) ?
                                (8'hba) : (8'had)))));
  assign wire3048 = $unsigned(wire3047[(4'hc):(4'hb)]);
  always
    @(posedge clk) begin
      reg3049 <= ($signed(wire3047[(3'h5):(2'h2)]) ?
          wire3047 : $unsigned({wire3040[(3'h6):(2'h3)]}));
      if ($unsigned({(8'h9f)}))
        begin
          if ($signed((~&$unsigned({wire3041}))))
            begin
              reg3050 <= $signed($signed(wire3047[(4'hb):(3'h6)]));
            end
          else
            begin
              if (($unsigned($signed($unsigned(reg3049))) ?
                  (8'ha0) : (|($unsigned(wire3046) ?
                      $unsigned((8'had)) : {reg3050}))))
                begin
                  reg3050 <= wire3046[(3'h4):(2'h3)];
                  reg3051 <= $signed(reg3049[(4'hb):(2'h2)]);
                end
              else
                begin
                  for (forvar3050 = (1'h0); (forvar3050 < (1'h0)); forvar3050 = (forvar3050 + (1'h1)))
                    begin
                      reg3051 <= $unsigned((8'hae));
                      reg3052 <= forvar3050[(4'h9):(3'h6)];
                    end
                  if ($signed(((reg3049[(3'h6):(3'h4)] ?
                      {reg3052} : wire3040) <= $unsigned((-(8'h9f))))))
                    begin
                      reg3053 <= wire3041;
                    end
                  else
                    begin
                      reg3053 <= ((^~$signed($unsigned(reg3052))) ?
                          forvar3050 : (~$signed(((8'h9d) >> wire3045))));
                      reg3054 <= wire3044[(2'h3):(1'h1)];
                      reg3055 <= wire3041;
                      reg3056 <= wire3042[(2'h3):(1'h0)];
                    end
                  for (forvar3057 = (1'h0); (forvar3057 < (1'h0)); forvar3057 = (forvar3057 + (1'h1)))
                    begin
                      reg3058 <= forvar3050;
                      reg3059 <= reg3055[(1'h1):(1'h1)];
                      reg3060 <= $unsigned(reg3052);
                      reg3061 <= ((&$signed(wire3044[(1'h0):(1'h0)])) ?
                          reg3050 : forvar3057);
                    end
                  reg3062 <= reg3051;
                end
              for (forvar3063 = (1'h0); (forvar3063 < (1'h0)); forvar3063 = (forvar3063 + (1'h1)))
                begin
                  for (forvar3064 = (1'h0); (forvar3064 < (1'h1)); forvar3064 = (forvar3064 + (1'h1)))
                    begin
                      reg3065 <= $unsigned($unsigned({(forvar3050 ?
                              wire3047 : forvar3050)}));
                    end
                  if ({wire3040})
                    begin
                      reg3066 <= $signed(reg3061);
                    end
                  else
                    begin
                      reg3066 <= (~&(~^($signed(wire3043) >> $unsigned(reg3066))));
                      reg3067 <= $signed($unsigned($signed((^reg3062))));
                      reg3068 <= (((8'hb7) ~^ $signed((^~reg3059))) ?
                          {$signed((wire3045 >> wire3044))} : (^~wire3043));
                      reg3069 <= $signed((~wire3046));
                    end
                  for (forvar3070 = (1'h0); (forvar3070 < (2'h2)); forvar3070 = (forvar3070 + (1'h1)))
                    begin
                      reg3071 <= (~^$unsigned($signed(wire3040[(1'h1):(1'h1)])));
                      reg3072 <= $signed(((^~(8'hab)) ~^ ({(8'hba)} ?
                          (-reg3054) : forvar3057)));
                    end
                end
              if ((reg3049 ?
                  wire3047 : ((reg3067 ?
                          reg3069[(3'h4):(2'h3)] : (wire3040 >= reg3062)) ?
                      ((reg3053 ?
                          wire3046 : forvar3050) >>> $unsigned(reg3067)) : {(wire3045 ?
                              wire3041 : forvar3070)})))
                begin
                  for (forvar3073 = (1'h0); (forvar3073 < (1'h0)); forvar3073 = (forvar3073 + (1'h1)))
                    begin
                      reg3074 <= {reg3059};
                      reg3075 <= $signed($signed($unsigned(reg3062[(2'h2):(2'h2)])));
                      reg3076 <= forvar3070[(3'h6):(2'h3)];
                    end
                  if ($signed(reg3067))
                    begin
                      reg3077 <= wire3048[(3'h5):(3'h4)];
                      reg3078 <= ($unsigned(forvar3070[(3'h6):(3'h5)]) & (&$unsigned({reg3074})));
                    end
                  else
                    begin
                      reg3077 <= wire3044[(1'h0):(1'h0)];
                      reg3078 <= {((^~((8'hb3) ?
                              reg3071 : reg3056)) | reg3053)};
                      reg3079 <= ((~(((8'ha2) ? forvar3063 : (8'hb7)) ?
                              (+reg3062) : (^reg3076))) ?
                          $unsigned({$unsigned(reg3062)}) : wire3040);
                      reg3080 <= $unsigned($unsigned((reg3060[(4'h9):(3'h7)] ?
                          $signed(reg3079) : (~|reg3060))));
                    end
                end
              else
                begin
                  for (forvar3073 = (1'h0); (forvar3073 < (2'h3)); forvar3073 = (forvar3073 + (1'h1)))
                    begin
                      reg3074 <= (~^wire3046);
                    end
                end
              if ((((~^$signed(reg3071)) ?
                  reg3062[(2'h2):(2'h2)] : (((8'ha7) * reg3074) ?
                      (reg3072 ?
                          wire3041 : reg3056) : $signed(wire3041))) ~^ {(wire3043 == wire3047[(3'h5):(2'h3)])}))
                begin
                  for (forvar3081 = (1'h0); (forvar3081 < (2'h2)); forvar3081 = (forvar3081 + (1'h1)))
                    begin
                      reg3082 <= (((+reg3074[(3'h5):(3'h4)]) ?
                          {reg3071} : reg3061) & (wire3048[(3'h4):(1'h1)] << reg3056[(2'h2):(2'h2)]));
                      reg3083 <= reg3061[(2'h3):(1'h0)];
                      reg3084 <= reg3062;
                    end
                  for (forvar3085 = (1'h0); (forvar3085 < (1'h1)); forvar3085 = (forvar3085 + (1'h1)))
                    begin
                      reg3086 <= (wire3043[(3'h4):(2'h2)] ?
                          (+wire3045[(4'hb):(4'h9)]) : $unsigned((^~$unsigned((8'hb9)))));
                      reg3087 <= (reg3065 << (^$unsigned(forvar3057)));
                    end
                  for (forvar3088 = (1'h0); (forvar3088 < (2'h2)); forvar3088 = (forvar3088 + (1'h1)))
                    begin
                      reg3089 <= (reg3056 << $unsigned($unsigned((wire3046 <= reg3052))));
                      reg3090 <= wire3040[(1'h0):(1'h0)];
                    end
                  for (forvar3091 = (1'h0); (forvar3091 < (1'h0)); forvar3091 = (forvar3091 + (1'h1)))
                    begin
                      reg3092 <= $unsigned(wire3044);
                      reg3093 <= {({{reg3089}} || wire3047)};
                      reg3094 <= (forvar3064 | forvar3063[(3'h6):(1'h0)]);
                      reg3095 <= (reg3068[(3'h4):(1'h1)] ^ (($signed((8'ha7)) > reg3058[(1'h0):(1'h0)]) << reg3068));
                    end
                end
              else
                begin
                  reg3081 <= ($unsigned(wire3042[(2'h3):(1'h1)]) < $signed(reg3054[(1'h1):(1'h0)]));
                  for (forvar3082 = (1'h0); (forvar3082 < (2'h3)); forvar3082 = (forvar3082 + (1'h1)))
                    begin
                      reg3083 <= (&$signed(((forvar3081 & forvar3070) ?
                          reg3093[(3'h5):(2'h3)] : (forvar3063 ^ wire3041))));
                      reg3084 <= (((reg3059[(3'h4):(1'h1)] ?
                              {forvar3063} : {forvar3050}) ?
                          reg3067[(4'hd):(3'h4)] : (8'ha6)) ^ reg3065[(4'he):(4'hb)]);
                      reg3085 <= (8'ha2);
                    end
                  reg3086 <= (forvar3064[(4'h9):(2'h2)] ?
                      reg3084 : $unsigned($unsigned(reg3090[(3'h7):(1'h0)])));
                  for (forvar3087 = (1'h0); (forvar3087 < (1'h0)); forvar3087 = (forvar3087 + (1'h1)))
                    begin
                      reg3088 <= $unsigned(({(~&(8'hac))} >> $signed($signed(reg3058))));
                      reg3089 <= ($unsigned($signed(reg3053)) ?
                          $unsigned((^~reg3088)) : (($unsigned(wire3046) ?
                              {(8'hb5)} : reg3081[(3'h7):(1'h0)]) | (-reg3051[(3'h4):(3'h4)])));
                      reg3090 <= {(-(|(|reg3060)))};
                      reg3091 <= reg3060;
                    end
                end
            end
          reg3096 <= {$signed((~^reg3054))};
          reg3097 <= (8'haf);
          reg3098 <= wire3047;
        end
      else
        begin
          if (wire3045[(4'ha):(1'h1)])
            begin
              reg3050 <= $signed(((8'hba) ?
                  $signed(wire3045) : ({reg3075} || $unsigned(reg3061))));
            end
          else
            begin
              for (forvar3050 = (1'h0); (forvar3050 < (2'h2)); forvar3050 = (forvar3050 + (1'h1)))
                begin
                  for (forvar3051 = (1'h0); (forvar3051 < (2'h3)); forvar3051 = (forvar3051 + (1'h1)))
                    begin
                      reg3052 <= wire3045[(2'h3):(1'h1)];
                      reg3053 <= ((((-reg3088) >= $unsigned(reg3080)) || ($unsigned(wire3042) ?
                          (|(8'hb6)) : (!wire3040))) - $signed((~&((8'ha3) ?
                          reg3082 : reg3059))));
                    end
                  for (forvar3054 = (1'h0); (forvar3054 < (2'h2)); forvar3054 = (forvar3054 + (1'h1)))
                    begin
                      reg3055 <= $signed((^wire3046));
                      reg3056 <= {reg3067};
                      reg3057 <= $unsigned($unsigned((reg3056 > {forvar3064})));
                      reg3058 <= $unsigned((~|$signed(reg3062)));
                    end
                end
              if ((8'hb9))
                begin
                  for (forvar3059 = (1'h0); (forvar3059 < (1'h0)); forvar3059 = (forvar3059 + (1'h1)))
                    begin
                      reg3060 <= {reg3080[(2'h2):(1'h0)]};
                    end
                end
              else
                begin
                  reg3059 <= (~&($signed($unsigned(wire3048)) < $unsigned($signed(reg3081))));
                  for (forvar3060 = (1'h0); (forvar3060 < (2'h2)); forvar3060 = (forvar3060 + (1'h1)))
                    begin
                      reg3061 <= reg3075[(1'h0):(1'h0)];
                      reg3062 <= ((reg3095[(3'h4):(2'h3)] ~^ ((reg3066 ?
                          forvar3082 : (8'ha2)) >>> {reg3076})) <<< ({$signed(reg3074)} ?
                          $unsigned((~(8'hb6))) : $signed((8'hb8))));
                      reg3063 <= {(reg3095 ? {(~&forvar3088)} : reg3076)};
                      reg3064 <= $unsigned(((~^forvar3054) == reg3067[(3'h7):(3'h5)]));
                    end
                end
              for (forvar3065 = (1'h0); (forvar3065 < (2'h2)); forvar3065 = (forvar3065 + (1'h1)))
                begin
                  for (forvar3066 = (1'h0); (forvar3066 < (2'h2)); forvar3066 = (forvar3066 + (1'h1)))
                    begin
                      reg3067 <= {$signed(({(8'had)} ?
                              forvar3060[(3'h5):(3'h4)] : $signed(reg3084)))};
                      reg3068 <= $signed((~&forvar3065));
                      reg3069 <= (8'hb2);
                      reg3070 <= reg3085[(2'h2):(1'h0)];
                    end
                  if (((~^$signed($unsigned(forvar3063))) ?
                      reg3085[(2'h2):(1'h1)] : $signed(forvar3087)))
                    begin
                      reg3071 <= reg3090[(4'ha):(1'h0)];
                      reg3072 <= reg3093;
                    end
                  else
                    begin
                      reg3071 <= (($signed((^~reg3092)) ?
                          $unsigned((reg3065 | forvar3059)) : wire3045[(2'h3):(1'h1)]) ^ (8'ha1));
                      reg3072 <= $unsigned($unsigned(reg3076));
                      reg3073 <= reg3072;
                      reg3074 <= (-$signed(($unsigned(forvar3073) ?
                          $unsigned(forvar3057) : {reg3064})));
                    end
                  for (forvar3075 = (1'h0); (forvar3075 < (1'h1)); forvar3075 = (forvar3075 + (1'h1)))
                    begin
                      reg3076 <= {forvar3051};
                      reg3077 <= ((forvar3063 ?
                          ((reg3068 ? (8'ha7) : (8'hb6)) ?
                              reg3084[(3'h7):(2'h2)] : ((8'h9d) - (8'hb9))) : ((~&reg3079) ?
                              $signed(forvar3054) : wire3040[(2'h2):(2'h2)])) ~^ $signed(reg3092));
                    end
                  for (forvar3078 = (1'h0); (forvar3078 < (1'h1)); forvar3078 = (forvar3078 + (1'h1)))
                    begin
                      reg3079 <= reg3088[(4'h8):(4'h8)];
                      reg3080 <= (forvar3078 ?
                          $signed((~|$unsigned((8'hb1)))) : (reg3055[(3'h7):(3'h7)] & $unsigned({wire3047})));
                      reg3081 <= ((-forvar3088) ?
                          reg3070[(4'hc):(4'h9)] : {(~&(~&(8'hae)))});
                    end
                end
              for (forvar3082 = (1'h0); (forvar3082 < (1'h1)); forvar3082 = (forvar3082 + (1'h1)))
                begin
                  if (forvar3057[(1'h1):(1'h0)])
                    begin
                      reg3083 <= $unsigned(reg3085[(1'h1):(1'h1)]);
                      reg3084 <= (8'hab);
                      reg3085 <= (!(8'hb0));
                    end
                  else
                    begin
                      reg3083 <= reg3058;
                      reg3084 <= (reg3071 ?
                          ($unsigned($unsigned(forvar3075)) >>> $unsigned(reg3069[(4'hb):(4'h9)])) : ((8'haa) ?
                              $signed(reg3095) : reg3049));
                      reg3085 <= reg3095[(2'h3):(2'h2)];
                    end
                end
            end
          if (reg3064[(2'h2):(1'h0)])
            begin
              for (forvar3086 = (1'h0); (forvar3086 < (2'h3)); forvar3086 = (forvar3086 + (1'h1)))
                begin
                  for (forvar3087 = (1'h0); (forvar3087 < (2'h2)); forvar3087 = (forvar3087 + (1'h1)))
                    begin
                      reg3088 <= {((^$signed(reg3092)) ?
                              wire3043[(3'h4):(3'h4)] : (^~{(8'hb3)}))};
                      reg3089 <= reg3081[(3'h5):(3'h4)];
                      reg3090 <= reg3049[(4'ha):(3'h5)];
                    end
                end
            end
          else
            begin
              if (reg3056[(1'h1):(1'h1)])
                begin
                  if (reg3056)
                    begin
                      reg3086 <= ($signed(wire3040) ?
                          $signed((+((8'hae) ?
                              reg3079 : forvar3063))) : $signed(reg3067[(4'ha):(3'h7)]));
                      reg3087 <= $signed((^$signed($unsigned((8'h9d)))));
                      reg3088 <= $signed(({$signed(reg3049)} ^ $unsigned($signed((8'hb8)))));
                      reg3089 <= $signed((~|((8'ha5) ?
                          reg3067[(2'h2):(1'h1)] : $unsigned((8'hb4)))));
                    end
                  else
                    begin
                      reg3086 <= (reg3072 ?
                          (reg3096 + $unsigned(reg3080)) : ((reg3065 ?
                                  {reg3094} : (forvar3065 ?
                                      (8'ha3) : reg3093)) ?
                              (reg3070[(4'h9):(3'h7)] ^~ $unsigned((8'hb4))) : {wire3048}));
                      reg3087 <= reg3089;
                      reg3088 <= (~$unsigned({$signed(wire3043)}));
                    end
                  for (forvar3090 = (1'h0); (forvar3090 < (1'h1)); forvar3090 = (forvar3090 + (1'h1)))
                    begin
                      reg3091 <= wire3048[(1'h1):(1'h0)];
                      reg3092 <= (8'ha8);
                      reg3093 <= (|$signed({reg3074[(2'h2):(2'h2)]}));
                      reg3094 <= forvar3070;
                    end
                  if ((~&($signed($unsigned(wire3045)) ?
                      wire3047[(1'h0):(1'h0)] : forvar3082[(2'h2):(1'h1)])))
                    begin
                      reg3095 <= ({$unsigned($signed((8'h9c)))} ~^ $signed(((~&reg3074) < {reg3096})));
                    end
                  else
                    begin
                      reg3095 <= (~&$signed(forvar3050[(4'h9):(1'h1)]));
                      reg3096 <= forvar3066;
                    end
                end
              else
                begin
                  for (forvar3086 = (1'h0); (forvar3086 < (1'h0)); forvar3086 = (forvar3086 + (1'h1)))
                    begin
                      reg3087 <= reg3056;
                      reg3088 <= ($unsigned(((forvar3078 << reg3091) >>> forvar3063[(3'h4):(1'h1)])) < reg3067);
                      reg3089 <= $unsigned({{{reg3098}}});
                    end
                  for (forvar3090 = (1'h0); (forvar3090 < (2'h2)); forvar3090 = (forvar3090 + (1'h1)))
                    begin
                      reg3091 <= $signed((~&(-(reg3050 ? (8'hb6) : wire3043))));
                      reg3092 <= {(+(-$unsigned(reg3093)))};
                      reg3093 <= $signed((({forvar3073} ?
                              (forvar3066 >= reg3097) : (reg3091 >> reg3096)) ?
                          ($unsigned(reg3049) ?
                              {forvar3073} : forvar3081[(3'h5):(2'h2)]) : (reg3088 ?
                              forvar3070[(3'h7):(3'h7)] : $signed(reg3053))));
                    end
                end
              reg3097 <= $unsigned(((8'ha7) ?
                  $signed(((8'ha1) ? reg3093 : reg3054)) : (^(reg3057 ?
                      reg3056 : reg3058))));
              if ($unsigned(($unsigned(forvar3064[(1'h1):(1'h1)]) ^~ ((~^wire3044) << $unsigned(reg3063)))))
                begin
                  for (forvar3098 = (1'h0); (forvar3098 < (1'h1)); forvar3098 = (forvar3098 + (1'h1)))
                    begin
                      reg3099 <= ((((8'ha7) | forvar3050) - forvar3086) ?
                          {$signed(forvar3060[(1'h1):(1'h1)])} : forvar3064[(1'h1):(1'h1)]);
                      reg3100 <= {reg3052};
                      reg3101 <= forvar3073[(2'h3):(2'h3)];
                      reg3102 <= reg3084;
                    end
                  for (forvar3103 = (1'h0); (forvar3103 < (1'h1)); forvar3103 = (forvar3103 + (1'h1)))
                    begin
                      reg3104 <= ({((wire3041 ~^ forvar3082) ?
                                  reg3084[(2'h3):(2'h2)] : (reg3099 ?
                                      reg3069 : (8'ha5)))} ?
                          $signed($unsigned(forvar3098)) : $signed(({forvar3066} ?
                              $signed(forvar3081) : forvar3082)));
                      reg3105 <= $unsigned(reg3071);
                    end
                end
              else
                begin
                  if ((~$unsigned(forvar3087[(4'hc):(4'h9)])))
                    begin
                      reg3098 <= forvar3078[(3'h4):(2'h3)];
                      reg3099 <= reg3089[(2'h3):(1'h0)];
                      reg3100 <= (((-$signed(forvar3082)) * (+(forvar3087 ?
                          forvar3087 : reg3059))) >>> reg3077);
                    end
                  else
                    begin
                      reg3098 <= (((&forvar3065[(1'h0):(1'h0)]) ^ (wire3047[(2'h2):(1'h1)] ?
                          $signed(reg3049) : (reg3084 >>> reg3049))) <<< (($unsigned(reg3053) >>> (reg3100 - (8'hba))) ?
                          (^(^~(8'hb6))) : $unsigned({reg3094})));
                    end
                  for (forvar3101 = (1'h0); (forvar3101 < (2'h3)); forvar3101 = (forvar3101 + (1'h1)))
                    begin
                      reg3102 <= forvar3098;
                      reg3103 <= $signed(((reg3084 >> $signed(forvar3054)) ?
                          {reg3076} : reg3057[(4'h8):(1'h1)]));
                      reg3104 <= reg3084[(2'h2):(1'h0)];
                      reg3105 <= (~|$unsigned((&((8'haf) == reg3097))));
                    end
                end
              for (forvar3106 = (1'h0); (forvar3106 < (1'h0)); forvar3106 = (forvar3106 + (1'h1)))
                begin
                  for (forvar3107 = (1'h0); (forvar3107 < (2'h2)); forvar3107 = (forvar3107 + (1'h1)))
                    begin
                      reg3108 <= ($signed({reg3102[(1'h0):(1'h0)]}) ?
                          forvar3086[(1'h0):(1'h0)] : (((!forvar3075) ^~ reg3090[(2'h3):(2'h2)]) < $signed((wire3046 ?
                              forvar3064 : wire3041))));
                      reg3109 <= reg3062;
                      reg3110 <= (((~^(~&reg3084)) >>> reg3059[(3'h6):(3'h6)]) ?
                          (8'hb0) : {((forvar3107 ? reg3055 : (8'h9d)) ?
                                  (reg3062 ?
                                      (8'ha2) : reg3073) : $unsigned((8'hb1)))});
                      reg3111 <= $signed($unsigned((8'hb3)));
                    end
                  if (reg3101[(2'h2):(1'h0)])
                    begin
                      reg3112 <= reg3086[(4'hc):(1'h0)];
                      reg3113 <= (!{($signed(wire3047) != $unsigned(forvar3090))});
                    end
                  else
                    begin
                      reg3112 <= ((^~((reg3080 ?
                          (8'ha5) : forvar3088) ~^ $signed(forvar3070))) << reg3105[(2'h3):(1'h1)]);
                      reg3113 <= (8'hb8);
                      reg3114 <= $unsigned(reg3063);
                      reg3115 <= (({forvar3064[(4'h9):(4'h9)]} ?
                              reg3052[(2'h3):(1'h0)] : reg3108) ?
                          reg3112[(4'h8):(3'h7)] : {{(+reg3081)}});
                    end
                end
            end
        end
      reg3116 <= (8'ha0);
    end
  module3117 modinst3367 (wire3366, clk, reg3050, forvar3078, forvar3073, reg3072, reg3070);
  assign wire3368 = forvar3075[(4'h9):(4'h9)];
  assign wire3369 = $unsigned(((wire3044[(1'h0):(1'h0)] ?
                            $signed((8'haf)) : (wire3366 ?
                                reg3101 : forvar3050)) ?
                        $unsigned(forvar3066[(3'h5):(3'h5)]) : $signed(reg3093)));
  assign wire3370 = $unsigned(reg3086[(3'h7):(2'h2)]);
  assign wire3371 = {$signed((^{reg3058}))};
  always
    @(posedge clk) begin
      for (forvar3372 = (1'h0); (forvar3372 < (2'h2)); forvar3372 = (forvar3372 + (1'h1)))
        begin
          reg3373 <= reg3078;
        end
      if ($signed((|((reg3087 > forvar3372) >>> {(8'haf)}))))
        begin
          for (forvar3374 = (1'h0); (forvar3374 < (1'h0)); forvar3374 = (forvar3374 + (1'h1)))
            begin
              if (((((wire3044 ?
                      reg3088 : forvar3073) >> $signed((8'ha1))) != forvar3050) ?
                  $unsigned(reg3094) : wire3044[(1'h0):(1'h0)]))
                begin
                  if (reg3064[(2'h3):(2'h3)])
                    begin
                      reg3375 <= (reg3105[(4'h9):(2'h3)] ?
                          (8'h9f) : $signed({{reg3063}}));
                      reg3376 <= $unsigned((&$unsigned((wire3368 ?
                          (8'had) : forvar3078))));
                      reg3377 <= {(-$signed($unsigned(reg3109)))};
                    end
                  else
                    begin
                      reg3375 <= (!$unsigned(((reg3058 ? reg3115 : (8'hb9)) ?
                          wire3045[(2'h2):(2'h2)] : $signed(reg3070))));
                      reg3376 <= $unsigned((((!reg3109) ?
                              $unsigned(reg3054) : (+wire3371)) ?
                          (+forvar3090) : forvar3091[(2'h2):(2'h2)]));
                    end
                  for (forvar3378 = (1'h0); (forvar3378 < (2'h2)); forvar3378 = (forvar3378 + (1'h1)))
                    begin
                      reg3379 <= (~|(+reg3057));
                      reg3380 <= $signed((forvar3070[(3'h7):(1'h0)] ^ forvar3057));
                      reg3381 <= (wire3045[(3'h4):(2'h2)] ?
                          forvar3078[(4'hb):(4'h9)] : $signed((!(reg3069 >= forvar3051))));
                    end
                  reg3382 <= forvar3063;
                end
              else
                begin
                  if (reg3064)
                    begin
                      reg3375 <= forvar3065[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3375 <= reg3074;
                      reg3376 <= reg3376[(3'h7):(2'h3)];
                      reg3377 <= (~|$unsigned(($unsigned(forvar3106) & $signed(reg3064))));
                    end
                  for (forvar3378 = (1'h0); (forvar3378 < (2'h3)); forvar3378 = (forvar3378 + (1'h1)))
                    begin
                      reg3379 <= reg3072;
                      reg3380 <= forvar3065[(4'hc):(4'hb)];
                      reg3381 <= forvar3066;
                      reg3382 <= (|{$signed((^reg3110))});
                    end
                  for (forvar3383 = (1'h0); (forvar3383 < (1'h1)); forvar3383 = (forvar3383 + (1'h1)))
                    begin
                      reg3384 <= reg3062[(3'h6):(1'h1)];
                      reg3385 <= {$signed(((+reg3114) ?
                              $unsigned(reg3081) : forvar3073[(4'h8):(3'h6)]))};
                    end
                  if ((forvar3107 >> $signed(reg3070)))
                    begin
                      reg3386 <= ((($signed(wire3041) ?
                              wire3048[(3'h5):(3'h5)] : (&reg3089)) ?
                          ({forvar3066} ?
                              (+reg3073) : $signed(reg3084)) : (^~forvar3060)) > forvar3088);
                      reg3387 <= ((reg3060[(3'h6):(3'h5)] ?
                              (wire3042[(3'h5):(2'h2)] ?
                                  reg3072 : $signed(wire3043)) : forvar3051[(3'h5):(1'h0)]) ?
                          ((~$unsigned((8'h9f))) & $unsigned(reg3376)) : (reg3067[(4'hc):(4'hb)] && ($unsigned(reg3375) ?
                              ((8'hac) ? reg3104 : reg3099) : wire3042)));
                      reg3388 <= $signed(wire3045);
                    end
                  else
                    begin
                      reg3386 <= forvar3057[(1'h1):(1'h0)];
                      reg3387 <= (|(8'hb9));
                    end
                end
            end
          reg3389 <= reg3062[(4'h8):(3'h7)];
          for (forvar3390 = (1'h0); (forvar3390 < (2'h3)); forvar3390 = (forvar3390 + (1'h1)))
            begin
              for (forvar3391 = (1'h0); (forvar3391 < (2'h3)); forvar3391 = (forvar3391 + (1'h1)))
                begin
                  for (forvar3392 = (1'h0); (forvar3392 < (1'h1)); forvar3392 = (forvar3392 + (1'h1)))
                    begin
                      reg3393 <= $unsigned(((reg3385[(1'h1):(1'h1)] >>> (reg3113 + forvar3087)) > (((8'ha9) ?
                          (8'hae) : reg3057) ^ $unsigned(forvar3103))));
                      reg3394 <= reg3388;
                    end
                  if (forvar3374[(2'h3):(2'h3)])
                    begin
                      reg3395 <= ($signed(wire3043[(2'h2):(2'h2)]) <= (~^(+$unsigned(reg3073))));
                      reg3396 <= forvar3390[(3'h6):(3'h6)];
                      reg3397 <= (forvar3060[(2'h2):(1'h0)] + {$unsigned((wire3371 ?
                              (8'ha0) : forvar3090))});
                    end
                  else
                    begin
                      reg3395 <= forvar3075[(1'h1):(1'h1)];
                    end
                  for (forvar3398 = (1'h0); (forvar3398 < (1'h0)); forvar3398 = (forvar3398 + (1'h1)))
                    begin
                      reg3399 <= (~|$unsigned((8'hb9)));
                      reg3400 <= $unsigned((reg3377[(3'h5):(2'h2)] ?
                          (reg3077 < wire3370) : ((reg3049 + (8'ha4)) ?
                              $unsigned(wire3370) : (~^(8'hb4)))));
                    end
                  reg3401 <= (~&reg3111[(2'h3):(1'h1)]);
                end
              reg3402 <= $signed((8'ha2));
            end
        end
      else
        begin
          for (forvar3374 = (1'h0); (forvar3374 < (1'h1)); forvar3374 = (forvar3374 + (1'h1)))
            begin
              for (forvar3375 = (1'h0); (forvar3375 < (1'h0)); forvar3375 = (forvar3375 + (1'h1)))
                begin
                  if ($signed(reg3055[(4'h8):(3'h5)]))
                    begin
                      reg3376 <= {((reg3397[(2'h2):(2'h2)] <= ((8'hba) ?
                              (8'hb9) : (8'ha7))) | $unsigned(reg3379))};
                      reg3377 <= $signed(forvar3070);
                      reg3378 <= $signed(((-(reg3393 ?
                          forvar3078 : forvar3085)) < (+reg3057[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg3376 <= wire3048;
                      reg3377 <= $unsigned((wire3041[(4'h8):(3'h7)] == ($unsigned(reg3069) < (~reg3105))));
                      reg3378 <= ((8'hae) ?
                          ($unsigned($signed(reg3075)) ?
                              wire3369 : {forvar3392}) : ((~|$signed(reg3099)) << $unsigned(((8'hb8) << wire3368))));
                      reg3379 <= reg3384[(2'h2):(1'h1)];
                    end
                  if ((($unsigned($signed((8'hba))) ?
                      ({(8'hab)} ?
                          $signed(reg3379) : (reg3051 ?
                              reg3102 : reg3400)) : (((8'hb3) <= reg3074) ?
                          (reg3376 ?
                              forvar3082 : reg3073) : $signed(reg3384))) <<< (~|$signed((~^reg3073)))))
                    begin
                      reg3380 <= {$signed(reg3088)};
                      reg3381 <= {$signed(((^~forvar3060) ?
                              {reg3080} : (reg3395 || reg3088)))};
                    end
                  else
                    begin
                      reg3380 <= ((reg3077[(1'h0):(1'h0)] << ((~^reg3104) << $unsigned(reg3380))) && (reg3103[(2'h2):(1'h1)] ?
                          $unsigned((8'ha2)) : (^~forvar3091[(3'h5):(2'h3)])));
                      reg3381 <= (($signed(reg3098) ?
                          (+(|forvar3078)) : $signed(reg3050)) - $unsigned(((reg3073 ?
                              reg3384 : (8'ha9)) ?
                          {wire3045} : forvar3060)));
                    end
                end
              for (forvar3382 = (1'h0); (forvar3382 < (2'h2)); forvar3382 = (forvar3382 + (1'h1)))
                begin
                  if ((&($unsigned((8'hb8)) ?
                      $unsigned(((8'had) >= reg3396)) : (forvar3392 ?
                          (8'hb0) : $signed(reg3094)))))
                    begin
                      reg3383 <= $unsigned(($unsigned(reg3109[(2'h3):(2'h3)]) <= (reg3399 ?
                          (reg3081 == reg3395) : (8'ha5))));
                      reg3384 <= (reg3096 + $unsigned(($unsigned(wire3042) == {reg3060})));
                      reg3385 <= (&(wire3048[(3'h7):(3'h4)] >> reg3056));
                      reg3386 <= $unsigned(((forvar3391 < (reg3375 && (8'h9d))) ?
                          {$unsigned(reg3375)} : reg3381));
                    end
                  else
                    begin
                      reg3383 <= reg3088;
                    end
                  if ($signed(reg3099))
                    begin
                      reg3387 <= ($signed(($signed(forvar3059) ?
                              $signed(reg3052) : $unsigned(reg3073))) ?
                          $signed(reg3093[(4'hc):(4'h9)]) : forvar3060[(3'h5):(3'h5)]);
                      reg3388 <= $signed((-$signed($signed(reg3396))));
                      reg3389 <= ($unsigned(reg3099) & (((reg3074 == reg3387) ^~ (reg3076 <<< reg3060)) ?
                          ((forvar3088 ? reg3060 : forvar3070) ?
                              (wire3370 ^~ (8'ha8)) : reg3094) : ($signed(reg3102) ~^ (forvar3091 ?
                              reg3378 : reg3388))));
                    end
                  else
                    begin
                      reg3387 <= (forvar3082 << ((^((8'h9d) ?
                              reg3067 : reg3079)) ?
                          reg3395 : ((forvar3057 ? forvar3390 : wire3041) ?
                              (~^forvar3070) : (reg3383 <<< reg3056))));
                    end
                end
              reg3390 <= $unsigned(forvar3050[(1'h1):(1'h1)]);
              if (forvar3375[(3'h6):(1'h0)])
                begin
                  for (forvar3391 = (1'h0); (forvar3391 < (1'h1)); forvar3391 = (forvar3391 + (1'h1)))
                    begin
                      reg3392 <= $unsigned({{((8'ha3) ? wire3370 : reg3098)}});
                      reg3393 <= $signed($unsigned((reg3115 ~^ (reg3072 & reg3082))));
                    end
                  for (forvar3394 = (1'h0); (forvar3394 < (1'h1)); forvar3394 = (forvar3394 + (1'h1)))
                    begin
                      reg3395 <= {forvar3059};
                      reg3396 <= {$signed(reg3386[(3'h6):(1'h1)])};
                    end
                  reg3397 <= (8'hae);
                end
              else
                begin
                  if (reg3082[(1'h1):(1'h1)])
                    begin
                      reg3391 <= (8'hb6);
                      reg3392 <= forvar3070[(4'h8):(2'h3)];
                      reg3393 <= reg3378;
                    end
                  else
                    begin
                      reg3391 <= reg3072;
                      reg3392 <= (~&reg3053[(1'h0):(1'h0)]);
                      reg3393 <= ($signed((~|(forvar3398 ?
                              wire3042 : reg3072))) ?
                          $signed(reg3110) : (((forvar3050 ^ reg3089) ?
                                  reg3083[(2'h3):(1'h1)] : $unsigned(reg3062)) ?
                              {((8'ha2) ?
                                      reg3394 : reg3402)} : $unsigned((~|reg3090))));
                      reg3394 <= (((!(reg3060 ?
                          forvar3063 : (8'had))) >= reg3073) & (+$unsigned({(8'ha7)})));
                    end
                end
            end
          if (((!$unsigned($unsigned((8'ha4)))) ?
              forvar3054[(4'h8):(3'h6)] : $signed((^~reg3379[(4'ha):(4'ha)]))))
            begin
              if (forvar3098[(4'h8):(4'h8)])
                begin
                  for (forvar3398 = (1'h0); (forvar3398 < (1'h0)); forvar3398 = (forvar3398 + (1'h1)))
                    begin
                      reg3399 <= (^~{(forvar3106 ?
                              forvar3078[(4'h9):(1'h0)] : $unsigned(reg3377))});
                      reg3400 <= reg3063;
                    end
                  for (forvar3401 = (1'h0); (forvar3401 < (1'h1)); forvar3401 = (forvar3401 + (1'h1)))
                    begin
                      reg3402 <= $unsigned({forvar3073[(1'h0):(1'h0)]});
                      reg3403 <= $unsigned({reg3055[(4'h8):(2'h2)]});
                      reg3404 <= (^~{(reg3071[(4'h9):(3'h7)] <= reg3376[(3'h7):(2'h3)])});
                    end
                  for (forvar3405 = (1'h0); (forvar3405 < (2'h3)); forvar3405 = (forvar3405 + (1'h1)))
                    begin
                      reg3406 <= (reg3111[(3'h4):(3'h4)] ?
                          forvar3390[(1'h1):(1'h1)] : ($signed((~^(8'hab))) ?
                              {reg3078[(2'h3):(1'h1)]} : $unsigned((reg3090 ?
                                  (8'ha5) : reg3092))));
                      reg3407 <= $unsigned($signed($unsigned(wire3366[(2'h3):(2'h2)])));
                      reg3408 <= $unsigned((-({reg3062} != (~^wire3040))));
                    end
                  reg3409 <= (|$signed(forvar3075));
                end
              else
                begin
                  reg3398 <= (reg3050 ?
                      (reg3083[(2'h3):(2'h3)] ~^ $unsigned(forvar3372[(4'he):(4'h8)])) : reg3080[(1'h0):(1'h0)]);
                  reg3399 <= $unsigned($unsigned((reg3062[(1'h0):(1'h0)] && (reg3377 - forvar3392))));
                end
              for (forvar3410 = (1'h0); (forvar3410 < (1'h1)); forvar3410 = (forvar3410 + (1'h1)))
                begin
                  if (((reg3086 ? {{wire3046}} : (^~reg3089)) - forvar3378))
                    begin
                      reg3411 <= ((~|(reg3068[(2'h3):(2'h3)] ?
                              ((8'ha6) | reg3108) : forvar3075)) ?
                          (((forvar3086 >> reg3101) ?
                              ((8'hb9) != reg3049) : (reg3074 ?
                                  reg3061 : forvar3065)) <= {reg3085}) : $unsigned(((~&forvar3090) ?
                              $unsigned((8'h9d)) : $signed(forvar3066))));
                      reg3412 <= $unsigned((forvar3410[(3'h4):(2'h2)] ?
                          ((reg3378 < reg3408) == $signed(reg3076)) : wire3369));
                      reg3413 <= (|(~^(reg3402[(2'h2):(1'h1)] || $signed(reg3388))));
                    end
                  else
                    begin
                      reg3411 <= (!(8'ha0));
                      reg3412 <= forvar3390;
                    end
                end
              reg3414 <= $unsigned(forvar3073);
            end
          else
            begin
              if ($signed($signed(($signed(reg3382) ?
                  forvar3088 : $signed(reg3112)))))
                begin
                  if (forvar3064[(4'h8):(3'h6)])
                    begin
                      reg3398 <= $signed((+((8'hac) == reg3060)));
                      reg3399 <= (8'h9f);
                      reg3400 <= (reg3392[(2'h3):(2'h3)] ?
                          reg3386[(1'h0):(1'h0)] : (reg3402 ?
                              (~wire3368[(1'h1):(1'h1)]) : $unsigned($unsigned(forvar3098))));
                      reg3401 <= forvar3088;
                    end
                  else
                    begin
                      reg3398 <= forvar3107[(4'hb):(3'h4)];
                      reg3399 <= ((8'hae) > {({forvar3081} << (wire3369 ~^ wire3040))});
                      reg3400 <= reg3058[(2'h3):(2'h3)];
                      reg3401 <= $signed($signed((~|(+reg3068))));
                    end
                end
              else
                begin
                  for (forvar3398 = (1'h0); (forvar3398 < (1'h0)); forvar3398 = (forvar3398 + (1'h1)))
                    begin
                      reg3399 <= ($signed($signed((~|reg3408))) ?
                          {{(reg3074 >= wire3370)}} : forvar3398[(3'h6):(1'h0)]);
                      reg3400 <= ((-forvar3405) ?
                          ((((8'ha3) && (8'hac)) ? (8'hb3) : (~^forvar3051)) ?
                              reg3373 : forvar3378) : $unsigned(wire3042[(4'h8):(3'h6)]));
                      reg3401 <= $unsigned($unsigned(forvar3391));
                      reg3402 <= (reg3088[(3'h7):(1'h0)] <<< $signed(({reg3110} ?
                          (8'hb9) : reg3377[(1'h0):(1'h0)])));
                    end
                end
              for (forvar3403 = (1'h0); (forvar3403 < (2'h3)); forvar3403 = (forvar3403 + (1'h1)))
                begin
                  for (forvar3404 = (1'h0); (forvar3404 < (1'h1)); forvar3404 = (forvar3404 + (1'h1)))
                    begin
                      reg3405 <= $unsigned((reg3067 ?
                          (((8'ha8) ?
                              reg3402 : reg3059) ~^ (reg3381 ^ reg3113)) : $unsigned((~^forvar3374))));
                      reg3406 <= (+reg3398);
                    end
                  if (((&(^~$unsigned(reg3064))) >>> (~^(~|(reg3407 ?
                      reg3375 : reg3052)))))
                    begin
                      reg3407 <= (~{{$unsigned(forvar3405)}});
                      reg3408 <= reg3083[(3'h6):(3'h6)];
                    end
                  else
                    begin
                      reg3407 <= (!$unsigned($unsigned((~&reg3373))));
                      reg3408 <= reg3088[(4'he):(3'h7)];
                      reg3409 <= $unsigned((+$signed((forvar3065 ?
                          wire3046 : forvar3081))));
                    end
                  for (forvar3410 = (1'h0); (forvar3410 < (2'h2)); forvar3410 = (forvar3410 + (1'h1)))
                    begin
                      reg3411 <= reg3079;
                      reg3412 <= {{forvar3391[(3'h7):(3'h5)]}};
                      reg3413 <= wire3043[(1'h0):(1'h0)];
                    end
                end
            end
          if ({reg3400})
            begin
              for (forvar3415 = (1'h0); (forvar3415 < (1'h1)); forvar3415 = (forvar3415 + (1'h1)))
                begin
                  for (forvar3416 = (1'h0); (forvar3416 < (1'h1)); forvar3416 = (forvar3416 + (1'h1)))
                    begin
                      reg3417 <= ($unsigned(reg3054) ?
                          ((-((8'ha2) < forvar3065)) ?
                              $unsigned(reg3111[(2'h2):(2'h2)]) : (((8'h9e) ?
                                      forvar3404 : (8'hb4)) ?
                                  reg3076 : (~&reg3091))) : $unsigned((^(forvar3398 ?
                              (8'hba) : (8'hb8)))));
                      reg3418 <= ($unsigned(reg3071) ?
                          ($signed($signed(reg3386)) & (~&$unsigned((8'hae)))) : $unsigned({reg3379[(4'h9):(3'h7)]}));
                    end
                  for (forvar3419 = (1'h0); (forvar3419 < (1'h1)); forvar3419 = (forvar3419 + (1'h1)))
                    begin
                      reg3420 <= $unsigned($signed(forvar3103));
                      reg3421 <= reg3087;
                      reg3422 <= $unsigned(reg3078);
                    end
                  for (forvar3423 = (1'h0); (forvar3423 < (2'h3)); forvar3423 = (forvar3423 + (1'h1)))
                    begin
                      reg3424 <= $signed(((-$signed(reg3413)) >>> $unsigned($unsigned((8'ha7)))));
                      reg3425 <= (reg3393 >> ((~&(|reg3108)) ?
                          reg3091 : ((forvar3401 > reg3080) && (reg3065 ?
                              wire3366 : wire3042))));
                      reg3426 <= (({wire3366} ?
                          $signed({(8'ha7)}) : $signed(forvar3405[(2'h3):(1'h0)])) & forvar3403[(2'h3):(1'h0)]);
                      reg3427 <= (~forvar3060[(4'h9):(2'h3)]);
                    end
                end
              if (((($signed(reg3385) ?
                  {forvar3057} : {reg3077}) >= ((forvar3057 | reg3063) && $unsigned((8'hb2)))) <= reg3050))
                begin
                  reg3428 <= $unsigned(((forvar3107 == (|(8'hab))) ?
                      $signed((&(8'h9f))) : (|reg3424[(1'h0):(1'h0)])));
                end
              else
                begin
                  reg3428 <= (~|$unsigned((^{(8'hae)})));
                  for (forvar3429 = (1'h0); (forvar3429 < (1'h0)); forvar3429 = (forvar3429 + (1'h1)))
                    begin
                      reg3430 <= (~^(8'ha6));
                      reg3431 <= (-reg3079);
                      reg3432 <= ((~$signed($unsigned(reg3095))) - $unsigned($signed((~|forvar3054))));
                      reg3433 <= reg3112;
                    end
                end
              if (($signed(($unsigned(reg3376) == forvar3075[(4'h9):(3'h6)])) * forvar3378[(4'hb):(1'h1)]))
                begin
                  if ((^($unsigned({reg3095}) ?
                      reg3078 : (|(reg3412 <= reg3059)))))
                    begin
                      reg3434 <= reg3389;
                      reg3435 <= ($signed($unsigned($unsigned((8'h9d)))) ?
                          ($unsigned(forvar3087[(3'h4):(1'h0)]) ?
                              ((!reg3391) >= (wire3048 && forvar3410)) : ((reg3081 ?
                                      reg3113 : forvar3082) ?
                                  (forvar3103 > reg3074) : (wire3368 ?
                                      forvar3081 : reg3091))) : forvar3090);
                    end
                  else
                    begin
                      reg3434 <= ((!((+reg3113) <= {reg3383})) <= ($unsigned((reg3395 ?
                              reg3430 : (8'hb6))) ?
                          reg3116[(3'h6):(1'h0)] : ($signed(forvar3382) ?
                              (reg3431 ?
                                  reg3049 : forvar3382) : $signed(reg3073))));
                      reg3435 <= ($unsigned(reg3432) <= (-reg3108));
                    end
                  for (forvar3436 = (1'h0); (forvar3436 < (1'h1)); forvar3436 = (forvar3436 + (1'h1)))
                    begin
                      reg3437 <= $unsigned(reg3109[(2'h3):(2'h2)]);
                      reg3438 <= reg3082[(2'h3):(1'h1)];
                    end
                  if (reg3076)
                    begin
                      reg3439 <= (!reg3068);
                    end
                  else
                    begin
                      reg3439 <= wire3048[(3'h5):(2'h3)];
                      reg3440 <= {$unsigned(reg3071)};
                      reg3441 <= forvar3091[(2'h2):(2'h2)];
                      reg3442 <= ({reg3086} ?
                          $unsigned(($unsigned(reg3387) + (reg3062 ?
                              (8'h9e) : wire3041))) : {reg3109});
                    end
                end
              else
                begin
                  if (forvar3394)
                    begin
                      reg3434 <= ({(~|(^reg3082))} ?
                          wire3044 : reg3384[(1'h0):(1'h0)]);
                      reg3435 <= (~$signed(forvar3064));
                      reg3436 <= $signed((reg3426[(1'h0):(1'h0)] ?
                          $signed((~^reg3385)) : wire3041));
                      reg3437 <= reg3428;
                    end
                  else
                    begin
                      reg3434 <= forvar3064[(2'h3):(2'h3)];
                      reg3435 <= (($unsigned(reg3096) ?
                          (reg3111[(1'h0):(1'h0)] ^ forvar3088[(3'h4):(1'h0)]) : (~^reg3112[(1'h1):(1'h1)])) != ((reg3088[(4'ha):(4'h8)] <<< (reg3375 ?
                              reg3432 : reg3090)) ?
                          ((forvar3392 ? forvar3085 : reg3396) ?
                              reg3072 : $unsigned(reg3074)) : $unsigned((+reg3050))));
                      reg3436 <= $unsigned(reg3408);
                    end
                  if ($unsigned($signed($unsigned($signed(forvar3419)))))
                    begin
                      reg3438 <= ((^($unsigned(forvar3106) >= (~|reg3402))) | reg3057[(4'h8):(3'h7)]);
                    end
                  else
                    begin
                      reg3438 <= ($signed({((8'hb1) ?
                              wire3044 : reg3104)}) || {(reg3414[(2'h3):(2'h3)] <= (~^reg3383))});
                      reg3439 <= $unsigned(($signed(reg3088[(4'hb):(2'h3)]) ?
                          reg3440 : (~|(-reg3109))));
                    end
                end
            end
          else
            begin
              for (forvar3415 = (1'h0); (forvar3415 < (2'h3)); forvar3415 = (forvar3415 + (1'h1)))
                begin
                  if ((+(reg3085 >>> ({reg3401} - reg3100))))
                    begin
                      reg3416 <= reg3111;
                      reg3417 <= forvar3436;
                      reg3418 <= {$unsigned(forvar3429[(2'h3):(2'h3)])};
                      reg3419 <= reg3092[(4'h9):(2'h3)];
                    end
                  else
                    begin
                      reg3416 <= ((forvar3054[(2'h2):(1'h1)] ?
                              $unsigned(forvar3398[(3'h7):(3'h7)]) : $signed((reg3416 > reg3100))) ?
                          ((reg3072[(3'h4):(2'h3)] ?
                                  (reg3408 ~^ forvar3410) : {reg3437}) ?
                              reg3055 : ($signed(forvar3054) >= $signed(reg3092))) : (reg3109[(2'h2):(1'h0)] ?
                              $unsigned((~|reg3406)) : ($unsigned(forvar3060) ?
                                  (wire3046 ?
                                      (8'h9d) : reg3101) : $unsigned(wire3041))));
                    end
                  for (forvar3420 = (1'h0); (forvar3420 < (1'h1)); forvar3420 = (forvar3420 + (1'h1)))
                    begin
                      reg3421 <= ((reg3112 >>> reg3067[(3'h6):(2'h2)]) ?
                          (~|reg3401[(3'h5):(3'h4)]) : reg3383);
                      reg3422 <= $unsigned($signed(reg3405[(1'h1):(1'h1)]));
                      reg3423 <= {({(reg3396 ? reg3082 : wire3369)} ?
                              $unsigned((reg3397 < reg3400)) : $unsigned((-reg3433)))};
                      reg3424 <= {reg3442};
                    end
                  for (forvar3425 = (1'h0); (forvar3425 < (1'h1)); forvar3425 = (forvar3425 + (1'h1)))
                    begin
                      reg3426 <= $signed($unsigned(forvar3050[(3'h4):(1'h0)]));
                    end
                  reg3427 <= $signed($unsigned($signed((8'haf))));
                end
              for (forvar3428 = (1'h0); (forvar3428 < (2'h3)); forvar3428 = (forvar3428 + (1'h1)))
                begin
                  if (((&reg3072[(2'h2):(1'h0)]) != $signed($signed($unsigned(wire3046)))))
                    begin
                      reg3429 <= ($signed({(reg3087 ? reg3435 : (8'ha3))}) ?
                          $signed(reg3400[(3'h5):(2'h3)]) : {$signed((reg3052 ?
                                  forvar3087 : reg3068))});
                      reg3430 <= (8'ha7);
                      reg3431 <= {reg3096};
                    end
                  else
                    begin
                      reg3429 <= wire3047[(4'h9):(3'h6)];
                      reg3430 <= $signed((reg3105 ?
                          (reg3076[(3'h6):(2'h2)] ?
                              (forvar3066 ^~ (8'hb3)) : (forvar3098 >= reg3392)) : ((-reg3075) ?
                              (~^(8'hb1)) : $unsigned(forvar3059))));
                      reg3431 <= ((8'hb4) ?
                          ((|$unsigned(reg3423)) >>> reg3409[(4'ha):(4'ha)]) : (^reg3416));
                    end
                  if (((~^{(reg3387 << reg3428)}) ?
                      reg3438 : $signed($unsigned(reg3071[(2'h3):(1'h1)]))))
                    begin
                      reg3432 <= reg3092;
                      reg3433 <= (8'hb1);
                      reg3434 <= ($signed((^reg3060[(3'h4):(1'h1)])) ?
                          ((~^(~reg3097)) + reg3082) : {reg3387[(4'hf):(3'h5)]});
                    end
                  else
                    begin
                      reg3432 <= ($signed($unsigned(reg3049)) ^~ (8'h9c));
                    end
                  for (forvar3435 = (1'h0); (forvar3435 < (1'h0)); forvar3435 = (forvar3435 + (1'h1)))
                    begin
                      reg3436 <= forvar3404[(2'h3):(1'h1)];
                      reg3437 <= forvar3082[(3'h7):(1'h0)];
                    end
                  if ((({reg3430[(4'h9):(3'h6)]} && ((~^(8'hba)) ?
                          reg3382 : (wire3041 <<< reg3399))) ?
                      $unsigned((-(forvar3107 << forvar3378))) : (($signed(reg3432) & (reg3430 + forvar3404)) ?
                          ($unsigned(reg3403) ?
                              forvar3051[(4'hb):(4'h8)] : $signed(forvar3404)) : $unsigned((reg3393 ?
                              reg3392 : forvar3410)))))
                    begin
                      reg3438 <= (+{(!$unsigned(reg3396))});
                      reg3439 <= (~^($unsigned($signed(forvar3391)) <= (~^reg3405)));
                      reg3440 <= $unsigned(((|$signed(reg3435)) ?
                          ((-reg3402) >= reg3411[(4'hc):(3'h6)]) : ((reg3436 ?
                              forvar3085 : (8'ha6)) + (+(8'hb1)))));
                      reg3441 <= (forvar3404[(3'h5):(1'h0)] <<< reg3109);
                    end
                  else
                    begin
                      reg3438 <= reg3116[(4'ha):(1'h0)];
                      reg3439 <= (-forvar3098[(3'h4):(2'h3)]);
                      reg3440 <= (forvar3090 & $unsigned((^~{reg3087})));
                    end
                end
              reg3442 <= (reg3386[(4'ha):(1'h1)] || reg3099[(2'h3):(1'h0)]);
            end
          for (forvar3443 = (1'h0); (forvar3443 < (1'h0)); forvar3443 = (forvar3443 + (1'h1)))
            begin
              for (forvar3444 = (1'h0); (forvar3444 < (1'h1)); forvar3444 = (forvar3444 + (1'h1)))
                begin
                  for (forvar3445 = (1'h0); (forvar3445 < (1'h0)); forvar3445 = (forvar3445 + (1'h1)))
                    begin
                      reg3446 <= {{(reg3389[(2'h2):(2'h2)] ?
                                  reg3111[(1'h1):(1'h1)] : (forvar3075 <<< reg3426))}};
                      reg3447 <= reg3054[(3'h5):(3'h5)];
                    end
                  if (forvar3419)
                    begin
                      reg3448 <= (8'ha0);
                      reg3449 <= $signed({(^(reg3088 ? (8'hb8) : reg3062))});
                    end
                  else
                    begin
                      reg3448 <= ({((~|(8'hb9)) ?
                              (reg3405 != reg3393) : ((8'ha2) ?
                                  (8'ha7) : reg3416))} + reg3382[(2'h2):(1'h1)]);
                      reg3449 <= (+(((reg3093 ?
                              reg3091 : forvar3403) <<< (~^reg3063)) ?
                          reg3427[(2'h2):(2'h2)] : $unsigned(reg3071)));
                    end
                end
              reg3450 <= (($unsigned(forvar3444) * (^$unsigned(reg3414))) ?
                  $unsigned((8'hae)) : (8'ha4));
              reg3451 <= (-(+forvar3416[(2'h3):(2'h3)]));
            end
        end
      reg3452 <= $signed((((reg3089 <<< reg3115) ?
          $signed(reg3069) : (reg3400 != (8'hb6))) != ((+reg3373) ?
          (reg3412 >= reg3093) : (~&(8'ha8)))));
    end
  always
    @(posedge clk) begin
      for (forvar3453 = (1'h0); (forvar3453 < (1'h1)); forvar3453 = (forvar3453 + (1'h1)))
        begin
          if ((($unsigned($signed(reg3395)) == reg3397) ?
              {(|(!reg3434))} : reg3437))
            begin
              for (forvar3454 = (1'h0); (forvar3454 < (2'h2)); forvar3454 = (forvar3454 + (1'h1)))
                begin
                  if ($signed(reg3377))
                    begin
                      reg3455 <= {{$unsigned((forvar3392 << reg3391))}};
                    end
                  else
                    begin
                      reg3455 <= forvar3060[(3'h4):(2'h3)];
                    end
                  if ($signed(($signed(reg3376) ~^ (reg3087 ?
                      (reg3400 << (8'hba)) : reg3375))))
                    begin
                      reg3456 <= $unsigned($unsigned(($signed(forvar3085) ?
                          {reg3452} : (8'hb5))));
                      reg3457 <= $unsigned($unsigned(({reg3086} ^~ forvar3445)));
                      reg3458 <= ((((~reg3115) ?
                              (~|(8'ha8)) : (reg3381 && forvar3078)) ?
                          (!(wire3041 << reg3055)) : $signed(((8'hb7) ?
                              reg3062 : forvar3428))) - (reg3084[(3'h7):(1'h0)] ?
                          (-$unsigned(reg3091)) : $unsigned(reg3057[(4'h8):(3'h7)])));
                      reg3459 <= (reg3431[(3'h6):(1'h0)] * reg3457);
                    end
                  else
                    begin
                      reg3456 <= reg3096[(4'h9):(2'h3)];
                    end
                end
            end
          else
            begin
              if (reg3066)
                begin
                  for (forvar3454 = (1'h0); (forvar3454 < (1'h1)); forvar3454 = (forvar3454 + (1'h1)))
                    begin
                      reg3455 <= reg3380[(1'h0):(1'h0)];
                      reg3456 <= $unsigned($signed(((reg3433 ?
                          reg3111 : (8'hb2)) ^~ (+reg3419))));
                      reg3457 <= $unsigned((8'ha4));
                    end
                  reg3458 <= $unsigned((^~($signed(reg3069) != $signed(reg3375))));
                end
              else
                begin
                  for (forvar3454 = (1'h0); (forvar3454 < (2'h3)); forvar3454 = (forvar3454 + (1'h1)))
                    begin
                      reg3455 <= $signed((~&((reg3064 >= reg3071) <= (reg3113 ?
                          forvar3415 : reg3062))));
                      reg3456 <= $signed($unsigned({(8'hb0)}));
                    end
                  for (forvar3457 = (1'h0); (forvar3457 < (1'h0)); forvar3457 = (forvar3457 + (1'h1)))
                    begin
                      reg3458 <= $unsigned(($signed($unsigned(wire3371)) ?
                          ($unsigned(forvar3403) != (forvar3443 ?
                              forvar3075 : wire3044)) : (~(forvar3457 ?
                              reg3393 : (8'haf)))));
                      reg3459 <= {reg3430[(3'h4):(3'h4)]};
                      reg3460 <= (($unsigned($signed(reg3114)) ?
                              $signed((reg3116 ?
                                  forvar3425 : reg3406)) : {$unsigned(reg3060)}) ?
                          (forvar3087[(3'h4):(1'h1)] ?
                              reg3059[(2'h3):(1'h0)] : $signed($unsigned((8'ha0)))) : reg3052);
                    end
                  reg3461 <= forvar3086[(1'h1):(1'h1)];
                end
              for (forvar3462 = (1'h0); (forvar3462 < (1'h1)); forvar3462 = (forvar3462 + (1'h1)))
                begin
                  if ((~|($signed((&reg3105)) ? reg3435 : (!reg3451))))
                    begin
                      reg3463 <= $unsigned({$unsigned(forvar3392[(4'he):(2'h2)])});
                      reg3464 <= (reg3446[(4'hd):(2'h3)] || (8'hb5));
                      reg3465 <= ((reg3108 | ($unsigned(reg3083) << $unsigned((8'ha2)))) > (8'ha6));
                    end
                  else
                    begin
                      reg3463 <= $unsigned($signed(reg3391[(2'h3):(1'h0)]));
                    end
                  for (forvar3466 = (1'h0); (forvar3466 < (2'h3)); forvar3466 = (forvar3466 + (1'h1)))
                    begin
                      reg3467 <= reg3389[(2'h2):(2'h2)];
                      reg3468 <= (reg3100[(4'hf):(3'h7)] != (({reg3386} << (~forvar3403)) >= (~(!reg3452))));
                    end
                end
            end
        end
      for (forvar3469 = (1'h0); (forvar3469 < (1'h0)); forvar3469 = (forvar3469 + (1'h1)))
        begin
          if (reg3094)
            begin
              reg3470 <= (reg3401[(3'h4):(1'h1)] ?
                  reg3450[(2'h2):(1'h1)] : forvar3419[(2'h3):(1'h1)]);
              for (forvar3471 = (1'h0); (forvar3471 < (1'h0)); forvar3471 = (forvar3471 + (1'h1)))
                begin
                  for (forvar3472 = (1'h0); (forvar3472 < (2'h3)); forvar3472 = (forvar3472 + (1'h1)))
                    begin
                      reg3473 <= forvar3073[(1'h0):(1'h0)];
                      reg3474 <= (reg3079[(3'h6):(3'h5)] ?
                          $unsigned((8'hb0)) : (8'hb0));
                      reg3475 <= (!forvar3066[(4'hb):(4'hb)]);
                      reg3476 <= reg3470[(1'h0):(1'h0)];
                    end
                end
              for (forvar3477 = (1'h0); (forvar3477 < (1'h0)); forvar3477 = (forvar3477 + (1'h1)))
                begin
                  if ((^~(^$signed(forvar3090))))
                    begin
                      reg3478 <= $signed(reg3098[(1'h0):(1'h0)]);
                      reg3479 <= $signed(($unsigned(reg3433) || ((^forvar3466) ?
                          reg3459 : (forvar3457 ? (8'ha9) : reg3459))));
                      reg3480 <= ((~^(~|(reg3050 ? forvar3064 : forvar3428))) ?
                          (((8'hab) ?
                              (~|reg3385) : forvar3086) <= $signed((reg3432 ?
                              reg3419 : forvar3462))) : forvar3070);
                    end
                  else
                    begin
                      reg3478 <= (forvar3372 ?
                          (~&((8'h9f) >> (~|(8'hb9)))) : $unsigned((reg3070 ^~ reg3412[(2'h2):(1'h0)])));
                      reg3479 <= $signed(($unsigned(reg3064) ?
                          (|reg3100[(3'h7):(3'h6)]) : (-(8'ha5))));
                      reg3480 <= ({$signed(reg3417[(1'h1):(1'h1)])} ?
                          (-(8'ha9)) : ($signed($unsigned((8'ha8))) ?
                              reg3060[(3'h7):(3'h7)] : forvar3471[(4'h8):(1'h0)]));
                      reg3481 <= wire3371;
                    end
                end
              reg3482 <= {reg3417};
            end
          else
            begin
              for (forvar3470 = (1'h0); (forvar3470 < (1'h0)); forvar3470 = (forvar3470 + (1'h1)))
                begin
                  for (forvar3471 = (1'h0); (forvar3471 < (1'h0)); forvar3471 = (forvar3471 + (1'h1)))
                    begin
                      reg3472 <= reg3080[(1'h1):(1'h0)];
                    end
                  reg3473 <= (8'hb3);
                  for (forvar3474 = (1'h0); (forvar3474 < (2'h2)); forvar3474 = (forvar3474 + (1'h1)))
                    begin
                      reg3475 <= {(8'h9d)};
                      reg3476 <= ((reg3077[(1'h1):(1'h0)] ?
                              $signed((reg3419 || (8'hba))) : $signed((-forvar3394))) ?
                          (~&$unsigned((forvar3419 ?
                              reg3480 : reg3105))) : (forvar3436[(4'hd):(4'h9)] ?
                              forvar3405[(2'h2):(1'h0)] : ((reg3460 ?
                                  reg3412 : forvar3390) >>> (reg3061 ?
                                  forvar3065 : forvar3435))));
                    end
                  if (reg3104[(3'h7):(3'h6)])
                    begin
                      reg3477 <= $unsigned((forvar3435[(1'h1):(1'h1)] ?
                          {((8'ha0) ?
                                  reg3049 : reg3435)} : $unsigned($signed(forvar3462))));
                      reg3478 <= (8'hab);
                      reg3479 <= reg3081;
                    end
                  else
                    begin
                      reg3477 <= (reg3398 ?
                          $unsigned(wire3368) : ($signed((8'h9f)) <= $signed((reg3402 * reg3404))));
                      reg3478 <= reg3474;
                      reg3479 <= (8'hae);
                    end
                end
            end
          for (forvar3483 = (1'h0); (forvar3483 < (1'h1)); forvar3483 = (forvar3483 + (1'h1)))
            begin
              for (forvar3484 = (1'h0); (forvar3484 < (1'h0)); forvar3484 = (forvar3484 + (1'h1)))
                begin
                  for (forvar3485 = (1'h0); (forvar3485 < (1'h1)); forvar3485 = (forvar3485 + (1'h1)))
                    begin
                      reg3486 <= ($unsigned($unsigned(((8'hb9) ?
                              reg3104 : reg3460))) ?
                          reg3092[(2'h3):(2'h2)] : {(^$signed(reg3384))});
                      reg3487 <= ({$unsigned((reg3377 - wire3044))} ?
                          ($unsigned(reg3382) << reg3067) : (8'ha4));
                      reg3488 <= ((&((-(8'hb2)) <= forvar3405)) & reg3074[(3'h6):(3'h5)]);
                      reg3489 <= $signed(reg3399[(1'h1):(1'h0)]);
                    end
                  reg3490 <= $unsigned($unsigned(reg3489));
                  for (forvar3491 = (1'h0); (forvar3491 < (2'h2)); forvar3491 = (forvar3491 + (1'h1)))
                    begin
                      reg3492 <= $signed($unsigned(($unsigned(forvar3060) >= (reg3377 < forvar3477))));
                    end
                end
              for (forvar3493 = (1'h0); (forvar3493 < (1'h1)); forvar3493 = (forvar3493 + (1'h1)))
                begin
                  reg3494 <= (((+{reg3061}) == ((reg3442 ?
                      reg3437 : (8'haf)) > $unsigned((8'ha6)))) ^~ (&reg3446));
                  for (forvar3495 = (1'h0); (forvar3495 < (1'h1)); forvar3495 = (forvar3495 + (1'h1)))
                    begin
                      reg3496 <= (-(^(forvar3436 ?
                          (!forvar3091) : (~reg3092))));
                      reg3497 <= ((^$signed((reg3407 <<< forvar3394))) == (($unsigned(forvar3420) ?
                              (^(8'hb5)) : (reg3422 ? reg3416 : reg3109)) ?
                          reg3460 : (forvar3444 ?
                              (8'hb9) : $unsigned(reg3100))));
                      reg3498 <= ($unsigned(($signed((8'ha3)) ?
                          (forvar3087 <<< forvar3428) : reg3070)) & forvar3078);
                    end
                  reg3499 <= (((forvar3403[(1'h1):(1'h0)] ^ (reg3380 ?
                      (8'hb2) : reg3425)) <<< (|{reg3449})) > (^forvar3435[(2'h2):(1'h0)]));
                end
              reg3500 <= (&forvar3383);
              if ((-reg3473))
                begin
                  for (forvar3501 = (1'h0); (forvar3501 < (1'h0)); forvar3501 = (forvar3501 + (1'h1)))
                    begin
                      reg3502 <= (-((~&$signed(reg3391)) > {forvar3484[(1'h1):(1'h0)]}));
                      reg3503 <= $unsigned(reg3465);
                    end
                  for (forvar3504 = (1'h0); (forvar3504 < (1'h1)); forvar3504 = (forvar3504 + (1'h1)))
                    begin
                      reg3505 <= reg3387;
                    end
                end
              else
                begin
                  reg3501 <= (!reg3482);
                end
            end
          reg3506 <= $signed(forvar3404[(4'h8):(1'h0)]);
        end
      for (forvar3507 = (1'h0); (forvar3507 < (2'h3)); forvar3507 = (forvar3507 + (1'h1)))
        begin
          for (forvar3508 = (1'h0); (forvar3508 < (2'h3)); forvar3508 = (forvar3508 + (1'h1)))
            begin
              for (forvar3509 = (1'h0); (forvar3509 < (1'h0)); forvar3509 = (forvar3509 + (1'h1)))
                begin
                  for (forvar3510 = (1'h0); (forvar3510 < (2'h3)); forvar3510 = (forvar3510 + (1'h1)))
                    begin
                      reg3511 <= {(-forvar3470[(1'h1):(1'h0)])};
                    end
                  for (forvar3512 = (1'h0); (forvar3512 < (1'h0)); forvar3512 = (forvar3512 + (1'h1)))
                    begin
                      reg3513 <= ({(8'ha1)} <<< $signed((reg3412 ?
                          $unsigned((8'ha8)) : $signed(reg3084))));
                    end
                end
              if (reg3430[(1'h0):(1'h0)])
                begin
                  reg3514 <= ({(reg3422[(3'h4):(1'h1)] ?
                          (forvar3091 > forvar3070) : (~forvar3065))} << $signed($signed(forvar3392[(4'hf):(1'h0)])));
                end
              else
                begin
                  reg3514 <= ({((8'ha4) ?
                          (reg3056 >> forvar3493) : (forvar3054 > reg3436))} * {{reg3435}});
                  reg3515 <= ((~|forvar3073) ~^ $unsigned((-{forvar3075})));
                end
              for (forvar3516 = (1'h0); (forvar3516 < (2'h3)); forvar3516 = (forvar3516 + (1'h1)))
                begin
                  for (forvar3517 = (1'h0); (forvar3517 < (2'h3)); forvar3517 = (forvar3517 + (1'h1)))
                    begin
                      reg3518 <= $signed({(^$signed((8'haf)))});
                      reg3519 <= $signed({$signed($signed(reg3378))});
                    end
                  if ($signed($signed((forvar3470 ?
                      $signed(reg3093) : reg3070[(3'h6):(1'h0)]))))
                    begin
                      reg3520 <= (wire3371 <<< $signed((~|{reg3113})));
                      reg3521 <= (+({(reg3520 ~^ reg3447)} ?
                          reg3473[(1'h1):(1'h1)] : reg3055));
                      reg3522 <= {$unsigned({(reg3096 ? reg3069 : (8'ha3))})};
                      reg3523 <= $unsigned(forvar3085);
                    end
                  else
                    begin
                      reg3520 <= (($signed((reg3067 ?
                          reg3395 : reg3390)) << ((^reg3114) ?
                          $signed((8'hb1)) : $signed(reg3458))) ^ reg3063);
                      reg3521 <= (forvar3088[(1'h0):(1'h0)] | (!(((8'h9c) ?
                          forvar3382 : reg3473) <= {(8'ha1)})));
                    end
                  for (forvar3524 = (1'h0); (forvar3524 < (1'h0)); forvar3524 = (forvar3524 + (1'h1)))
                    begin
                      reg3525 <= $unsigned(reg3097);
                    end
                end
            end
          reg3526 <= {$unsigned(reg3073)};
          reg3527 <= (((^(forvar3484 && reg3100)) ?
                  reg3503[(1'h1):(1'h0)] : {(wire3366 ?
                          reg3064 : forvar3425)}) ?
              $signed($signed(reg3473[(1'h0):(1'h0)])) : (({reg3449} >= (reg3063 ?
                      reg3464 : forvar3509)) ?
                  (reg3086[(3'h4):(1'h1)] << forvar3517[(2'h2):(2'h2)]) : forvar3445[(2'h3):(1'h1)]));
          reg3528 <= (|({(&reg3063)} && ({reg3070} && (^~forvar3398))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2361
#( parameter param3034 = ((-(((8'ha7) ? (8'ha9) : (8'ha5)) << ((8'hb8) ? (8'haa) : (8'h9e)))) ? ((-(|(8'hb2))) ? ({(8'ha5)} >> {(8'hb6)}) : (((8'hac) ^ (8'ha2)) - ((8'had) + (8'hb7)))) : {(((8'hae) + (8'h9d)) ~^ (~(8'ha0)))}) )
(y, clk, wire2366, wire2365, wire2364, wire2363, wire2362);
  output wire [(32'h4ee):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire2366;
  input wire signed [(3'h7):(1'h0)] wire2365;
  input wire [(4'h8):(1'h0)] wire2364;
  input wire [(4'hb):(1'h0)] wire2363;
  input wire signed [(4'hf):(1'h0)] wire2362;
  wire signed [(4'hc):(1'h0)] wire3033;
  wire signed [(4'he):(1'h0)] wire3032;
  reg signed [(4'he):(1'h0)] reg3031 = (1'h0);
  reg [(3'h7):(1'h0)] reg3030 = (1'h0);
  reg [(2'h3):(1'h0)] reg3029 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3028 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3027 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3026 = (1'h0);
  reg [(3'h5):(1'h0)] reg3025 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3024 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3023 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3022 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3021 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3020 = (1'h0);
  reg [(3'h6):(1'h0)] reg3019 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3018 = (1'h0);
  reg [(4'he):(1'h0)] reg3017 = (1'h0);
  reg [(4'hb):(1'h0)] reg3016 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3015 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3010 = (1'h0);
  reg [(4'hc):(1'h0)] reg3008 = (1'h0);
  reg [(3'h4):(1'h0)] reg3015 = (1'h0);
  reg [(4'ha):(1'h0)] reg3014 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3013 = (1'h0);
  reg [(2'h3):(1'h0)] reg3012 = (1'h0);
  reg [(5'h10):(1'h0)] reg3011 = (1'h0);
  reg [(3'h7):(1'h0)] reg3010 = (1'h0);
  reg [(4'hf):(1'h0)] reg3009 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3008 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3007 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3006 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2998 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3005 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3004 = (1'h0);
  reg [(4'hd):(1'h0)] reg3003 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3002 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3001 = (1'h0);
  reg [(4'hd):(1'h0)] reg3000 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2999 = (1'h0);
  reg [(4'ha):(1'h0)] reg2998 = (1'h0);
  reg [(4'he):(1'h0)] reg2997 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2996 = (1'h0);
  reg [(2'h3):(1'h0)] reg2995 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2994 = (1'h0);
  reg [(5'h10):(1'h0)] reg2993 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2992 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2991 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2986 = (1'h0);
  reg [(4'he):(1'h0)] reg2983 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2982 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2979 = (1'h0);
  reg [(4'h8):(1'h0)] reg2978 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2977 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2974 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2964 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2963 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2959 = (1'h0);
  reg [(2'h3):(1'h0)] reg2992 = (1'h0);
  reg [(3'h6):(1'h0)] reg2991 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2990 = (1'h0);
  reg [(4'he):(1'h0)] reg2989 = (1'h0);
  reg [(3'h5):(1'h0)] reg2988 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2987 = (1'h0);
  reg [(2'h2):(1'h0)] reg2986 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2985 = (1'h0);
  reg [(5'h10):(1'h0)] reg2984 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2983 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2982 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2981 = (1'h0);
  reg [(2'h2):(1'h0)] reg2980 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2979 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2978 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2965 = (1'h0);
  reg [(4'ha):(1'h0)] reg2977 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2976 = (1'h0);
  reg [(4'hd):(1'h0)] reg2975 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2974 = (1'h0);
  reg [(4'he):(1'h0)] reg2973 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2972 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2971 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2970 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2969 = (1'h0);
  reg [(5'h10):(1'h0)] reg2968 = (1'h0);
  reg [(3'h4):(1'h0)] reg2967 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2966 = (1'h0);
  reg [(4'h9):(1'h0)] reg2965 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2960 = (1'h0);
  reg [(3'h5):(1'h0)] reg2958 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2964 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2963 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2962 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2961 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2960 = (1'h0);
  reg [(4'ha):(1'h0)] reg2959 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2958 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2957 = (1'h0);
  reg [(4'h9):(1'h0)] reg2956 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2955 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2954 = (1'h0);
  reg [(4'h9):(1'h0)] reg2953 = (1'h0);
  reg [(2'h3):(1'h0)] reg2952 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2951 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2950 = (1'h0);
  reg [(4'hf):(1'h0)] reg2949 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2948 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2947 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2946 = (1'h0);
  reg [(4'h8):(1'h0)] reg2945 = (1'h0);
  reg [(4'hd):(1'h0)] reg2944 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2943 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2942 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2941 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2940 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2939 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2938 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2937 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2936 = (1'h0);
  reg [(3'h4):(1'h0)] reg2935 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2934 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2933 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2932 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2931 = (1'h0);
  reg [(4'hc):(1'h0)] reg2930 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2929 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2928 = (1'h0);
  reg [(4'he):(1'h0)] reg2927 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2926 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2925 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2924 = (1'h0);
  reg [(4'he):(1'h0)] forvar2923 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2922 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2921 = (1'h0);
  reg [(4'hb):(1'h0)] reg2920 = (1'h0);
  wire [(3'h5):(1'h0)] wire2918;
  wire signed [(4'hd):(1'h0)] wire2369;
  wire [(4'ha):(1'h0)] wire2368;
  wire signed [(3'h5):(1'h0)] wire2367;
  assign y = {wire3033,
                 wire3032,
                 reg3031,
                 reg3030,
                 reg3029,
                 reg3028,
                 forvar3027,
                 forvar3026,
                 reg3025,
                 reg3024,
                 reg3023,
                 forvar3022,
                 reg3021,
                 forvar3020,
                 reg3019,
                 reg3018,
                 reg3017,
                 reg3016,
                 forvar3015,
                 forvar3010,
                 reg3008,
                 reg3015,
                 reg3014,
                 forvar3013,
                 reg3012,
                 reg3011,
                 reg3010,
                 reg3009,
                 forvar3008,
                 forvar3007,
                 forvar3006,
                 forvar2998,
                 reg3005,
                 reg3004,
                 reg3003,
                 reg3002,
                 forvar3001,
                 reg3000,
                 reg2999,
                 reg2998,
                 reg2997,
                 reg2996,
                 reg2995,
                 reg2994,
                 reg2993,
                 forvar2992,
                 forvar2991,
                 forvar2986,
                 reg2983,
                 reg2982,
                 reg2979,
                 reg2978,
                 forvar2977,
                 reg2974,
                 forvar2964,
                 forvar2963,
                 forvar2959,
                 reg2992,
                 reg2991,
                 reg2990,
                 reg2989,
                 reg2988,
                 reg2987,
                 reg2986,
                 reg2985,
                 reg2984,
                 forvar2983,
                 forvar2982,
                 reg2981,
                 reg2980,
                 forvar2979,
                 forvar2978,
                 forvar2965,
                 reg2977,
                 reg2976,
                 reg2975,
                 forvar2974,
                 reg2973,
                 reg2972,
                 reg2971,
                 forvar2970,
                 reg2969,
                 reg2968,
                 reg2967,
                 reg2966,
                 reg2965,
                 forvar2960,
                 reg2958,
                 reg2964,
                 reg2963,
                 reg2962,
                 reg2961,
                 reg2960,
                 reg2959,
                 forvar2958,
                 forvar2957,
                 reg2956,
                 reg2955,
                 reg2954,
                 reg2953,
                 reg2952,
                 forvar2951,
                 reg2950,
                 reg2949,
                 forvar2948,
                 reg2947,
                 reg2946,
                 reg2945,
                 reg2944,
                 forvar2943,
                 reg2942,
                 reg2941,
                 reg2940,
                 reg2939,
                 forvar2938,
                 forvar2937,
                 forvar2936,
                 reg2935,
                 reg2934,
                 reg2933,
                 forvar2932,
                 forvar2931,
                 reg2930,
                 forvar2929,
                 reg2928,
                 reg2927,
                 reg2926,
                 reg2925,
                 forvar2924,
                 forvar2923,
                 reg2922,
                 forvar2921,
                 reg2920,
                 wire2918,
                 wire2369,
                 wire2368,
                 wire2367,
                 (1'h0)};
  assign wire2367 = {$signed(((wire2362 ? (8'hb2) : wire2365) ?
                            wire2363[(4'h8):(1'h0)] : $unsigned(wire2366)))};
  assign wire2368 = wire2362[(4'h8):(3'h7)];
  assign wire2369 = wire2364[(1'h0):(1'h0)];
  module2370 modinst2919 (wire2918, clk, wire2364, wire2362, wire2363, wire2369);
  always
    @(posedge clk) begin
      reg2920 <= wire2365;
      for (forvar2921 = (1'h0); (forvar2921 < (1'h0)); forvar2921 = (forvar2921 + (1'h1)))
        begin
          reg2922 <= (8'ha6);
          for (forvar2923 = (1'h0); (forvar2923 < (2'h2)); forvar2923 = (forvar2923 + (1'h1)))
            begin
              for (forvar2924 = (1'h0); (forvar2924 < (2'h3)); forvar2924 = (forvar2924 + (1'h1)))
                begin
                  if ($unsigned($unsigned($signed((wire2364 == wire2367)))))
                    begin
                      reg2925 <= (!reg2922);
                      reg2926 <= ($signed($signed((8'haf))) <<< (-(+$unsigned(wire2369))));
                      reg2927 <= (wire2364 >>> $unsigned($unsigned(wire2365)));
                      reg2928 <= ($signed((((8'ha4) <= forvar2921) ?
                              (&(8'hab)) : $signed(wire2369))) ?
                          wire2362 : $unsigned((((8'hae) && reg2922) ?
                              $unsigned((8'h9d)) : forvar2921)));
                    end
                  else
                    begin
                      reg2925 <= reg2922[(3'h4):(3'h4)];
                      reg2926 <= $unsigned(((+(wire2364 ?
                          (8'hab) : (8'ha7))) << ((reg2927 ?
                              wire2369 : (8'ha6)) ?
                          (!reg2920) : wire2362[(4'hc):(4'h9)])));
                      reg2927 <= (^(($signed(forvar2921) ~^ $signed(wire2369)) ?
                          $unsigned($unsigned(reg2928)) : $unsigned($unsigned(forvar2924))));
                    end
                  for (forvar2929 = (1'h0); (forvar2929 < (2'h2)); forvar2929 = (forvar2929 + (1'h1)))
                    begin
                      reg2930 <= $signed($signed((wire2918[(3'h4):(2'h2)] < (wire2367 ?
                          forvar2929 : wire2365))));
                    end
                end
              for (forvar2931 = (1'h0); (forvar2931 < (1'h0)); forvar2931 = (forvar2931 + (1'h1)))
                begin
                  for (forvar2932 = (1'h0); (forvar2932 < (1'h1)); forvar2932 = (forvar2932 + (1'h1)))
                    begin
                      reg2933 <= wire2364[(3'h4):(2'h2)];
                    end
                  if (wire2918[(2'h3):(2'h3)])
                    begin
                      reg2934 <= ((($unsigned(forvar2921) ?
                              wire2363 : wire2366) != ($unsigned((8'ha3)) ?
                              wire2366[(1'h0):(1'h0)] : ((8'hb4) ?
                                  wire2363 : wire2918))) ?
                          (~^$unsigned((+(8'hb3)))) : {((wire2366 ?
                                      reg2922 : forvar2932) ?
                                  forvar2924 : (wire2365 ?
                                      wire2366 : wire2364))});
                    end
                  else
                    begin
                      reg2934 <= {{($unsigned(wire2362) - (!reg2934))}};
                      reg2935 <= (+wire2368);
                    end
                end
            end
        end
      for (forvar2936 = (1'h0); (forvar2936 < (1'h1)); forvar2936 = (forvar2936 + (1'h1)))
        begin
          for (forvar2937 = (1'h0); (forvar2937 < (2'h2)); forvar2937 = (forvar2937 + (1'h1)))
            begin
              for (forvar2938 = (1'h0); (forvar2938 < (1'h0)); forvar2938 = (forvar2938 + (1'h1)))
                begin
                  reg2939 <= $unsigned({$unsigned((8'hb1))});
                end
              if (wire2369[(3'h6):(1'h1)])
                begin
                  if (wire2363)
                    begin
                      reg2940 <= $unsigned(forvar2936);
                      reg2941 <= (8'haf);
                    end
                  else
                    begin
                      reg2940 <= reg2940;
                      reg2941 <= $signed(($signed((reg2928 ?
                              reg2935 : wire2369)) ?
                          (|(wire2368 ?
                              reg2934 : wire2364)) : reg2934[(2'h3):(2'h3)]));
                      reg2942 <= reg2930;
                    end
                  for (forvar2943 = (1'h0); (forvar2943 < (2'h2)); forvar2943 = (forvar2943 + (1'h1)))
                    begin
                      reg2944 <= forvar2932[(1'h1):(1'h0)];
                      reg2945 <= reg2942;
                      reg2946 <= (~|$signed(reg2934));
                      reg2947 <= (~|$unsigned(((forvar2931 - reg2935) << (reg2928 < (8'hb8)))));
                    end
                  for (forvar2948 = (1'h0); (forvar2948 < (2'h3)); forvar2948 = (forvar2948 + (1'h1)))
                    begin
                      reg2949 <= $unsigned((((wire2369 * reg2920) && $signed(wire2367)) > {$unsigned(wire2365)}));
                      reg2950 <= {{forvar2936[(2'h3):(1'h0)]}};
                    end
                  for (forvar2951 = (1'h0); (forvar2951 < (1'h1)); forvar2951 = (forvar2951 + (1'h1)))
                    begin
                      reg2952 <= $unsigned(((~^(wire2366 >>> reg2940)) ?
                          (~^(wire2362 > reg2949)) : ((!reg2930) >= (8'had))));
                      reg2953 <= ((8'hb0) ?
                          (~&$signed((wire2365 >> (8'ha7)))) : reg2934[(2'h2):(1'h1)]);
                      reg2954 <= $signed((reg2953[(4'h8):(3'h4)] ?
                          reg2928[(1'h0):(1'h0)] : $unsigned((forvar2932 ?
                              wire2368 : forvar2948))));
                      reg2955 <= (reg2940 >> ($signed(reg2925) ?
                          (&(forvar2948 ?
                              (8'haf) : forvar2931)) : $unsigned((reg2927 ?
                              reg2922 : reg2953))));
                    end
                end
              else
                begin
                  if ($signed((&forvar2951[(4'h8):(3'h6)])))
                    begin
                      reg2940 <= {forvar2931[(3'h7):(1'h0)]};
                      reg2941 <= ((+($unsigned(reg2920) ?
                          (8'h9d) : (!forvar2951))) >>> $unsigned(wire2368[(3'h6):(2'h2)]));
                    end
                  else
                    begin
                      reg2940 <= (|$unsigned($unsigned((reg2922 ?
                          wire2369 : forvar2932))));
                      reg2941 <= reg2935;
                      reg2942 <= $signed((reg2955 && (+(reg2950 >> forvar2936))));
                    end
                end
            end
          reg2956 <= (8'hb2);
        end
      if ((&wire2362[(2'h2):(1'h1)]))
        begin
          for (forvar2957 = (1'h0); (forvar2957 < (2'h2)); forvar2957 = (forvar2957 + (1'h1)))
            begin
              if ($unsigned($signed(reg2952[(1'h0):(1'h0)])))
                begin
                  for (forvar2958 = (1'h0); (forvar2958 < (1'h0)); forvar2958 = (forvar2958 + (1'h1)))
                    begin
                      reg2959 <= $unsigned({{(wire2369 ?
                                  forvar2931 : wire2363)}});
                      reg2960 <= $unsigned((forvar2924 ?
                          ($unsigned(forvar2958) <= {reg2946}) : reg2930));
                    end
                  if ($signed(($signed((wire2363 ^~ reg2949)) & wire2366)))
                    begin
                      reg2961 <= (!((&$signed((8'hb7))) < {(|(8'hba))}));
                    end
                  else
                    begin
                      reg2961 <= $signed({(+$signed(forvar2931))});
                      reg2962 <= $unsigned(reg2935);
                      reg2963 <= (8'ha2);
                      reg2964 <= {reg2955};
                    end
                end
              else
                begin
                  reg2958 <= ($unsigned({forvar2958}) && reg2963);
                  reg2959 <= $signed($unsigned($signed(forvar2943[(3'h7):(3'h5)])));
                  for (forvar2960 = (1'h0); (forvar2960 < (1'h1)); forvar2960 = (forvar2960 + (1'h1)))
                    begin
                      reg2961 <= reg2927[(1'h0):(1'h0)];
                      reg2962 <= reg2955[(3'h5):(1'h1)];
                      reg2963 <= reg2950[(3'h6):(2'h3)];
                      reg2964 <= forvar2938;
                    end
                end
              if ((8'h9f))
                begin
                  reg2965 <= reg2942;
                  if (forvar2936[(2'h3):(1'h1)])
                    begin
                      reg2966 <= (wire2918[(1'h0):(1'h0)] ?
                          reg2947 : $signed((reg2961[(1'h1):(1'h1)] ?
                              reg2934[(2'h3):(2'h3)] : $unsigned(reg2963))));
                      reg2967 <= (^reg2961[(3'h5):(1'h1)]);
                      reg2968 <= {($signed($signed(forvar2943)) ?
                              (-{forvar2943}) : (+reg2965[(2'h2):(1'h0)]))};
                      reg2969 <= reg2935;
                    end
                  else
                    begin
                      reg2966 <= $unsigned((~|((!reg2965) * (reg2963 ?
                          forvar2921 : reg2958))));
                      reg2967 <= forvar2957[(1'h0):(1'h0)];
                      reg2968 <= $unsigned((reg2922[(2'h2):(1'h1)] >>> {(reg2926 ?
                              reg2941 : reg2953)}));
                      reg2969 <= {{((wire2362 >= reg2966) ?
                                  {forvar2957} : wire2367[(2'h2):(1'h1)])}};
                    end
                  for (forvar2970 = (1'h0); (forvar2970 < (1'h0)); forvar2970 = (forvar2970 + (1'h1)))
                    begin
                      reg2971 <= $unsigned($signed(((wire2366 == (8'hb9)) ?
                          $signed(reg2962) : reg2928[(1'h0):(1'h0)])));
                      reg2972 <= $signed((forvar2921[(1'h1):(1'h1)] ?
                          (reg2969[(3'h5):(2'h2)] ?
                              (reg2939 ?
                                  reg2928 : reg2956) : {reg2946}) : ((~^(8'hb7)) ?
                              $signed(forvar2936) : forvar2931[(1'h1):(1'h0)])));
                      reg2973 <= (($signed((reg2944 == (8'hb9))) ?
                          reg2935[(1'h0):(1'h0)] : (~&(wire2918 ?
                              (8'hba) : reg2958))) <= forvar2957);
                    end
                  for (forvar2974 = (1'h0); (forvar2974 < (2'h3)); forvar2974 = (forvar2974 + (1'h1)))
                    begin
                      reg2975 <= reg2939;
                      reg2976 <= reg2946;
                      reg2977 <= (8'hb0);
                    end
                end
              else
                begin
                  for (forvar2965 = (1'h0); (forvar2965 < (2'h2)); forvar2965 = (forvar2965 + (1'h1)))
                    begin
                      reg2966 <= forvar2943[(1'h1):(1'h0)];
                      reg2967 <= (($unsigned({reg2941}) ?
                          ($unsigned(wire2362) ?
                              (~reg2935) : (reg2955 ?
                                  forvar2948 : reg2962)) : reg2975[(4'h8):(3'h5)]) < {$unsigned((reg2954 || reg2972))});
                    end
                end
              for (forvar2978 = (1'h0); (forvar2978 < (2'h3)); forvar2978 = (forvar2978 + (1'h1)))
                begin
                  for (forvar2979 = (1'h0); (forvar2979 < (1'h0)); forvar2979 = (forvar2979 + (1'h1)))
                    begin
                      reg2980 <= reg2961;
                      reg2981 <= forvar2936;
                    end
                end
              for (forvar2982 = (1'h0); (forvar2982 < (1'h0)); forvar2982 = (forvar2982 + (1'h1)))
                begin
                  for (forvar2983 = (1'h0); (forvar2983 < (1'h0)); forvar2983 = (forvar2983 + (1'h1)))
                    begin
                      reg2984 <= $unsigned(((+(+forvar2957)) ?
                          $signed($signed(reg2942)) : wire2369));
                      reg2985 <= {$unsigned($unsigned((reg2928 ?
                              wire2368 : (8'hba))))};
                      reg2986 <= ((forvar2970[(3'h5):(3'h5)] ?
                          reg2946 : ((^reg2939) == forvar2932[(1'h0):(1'h0)])) || (&$unsigned($signed(reg2920))));
                      reg2987 <= ((($signed(reg2966) <= (reg2940 ?
                                  reg2940 : reg2964)) ?
                              (reg2961 ?
                                  (~&reg2954) : $unsigned(reg2954)) : ($signed(forvar2979) ?
                                  (8'hba) : (~|(8'hb2)))) ?
                          ((forvar2948[(1'h1):(1'h0)] << wire2365) ?
                              ($signed(forvar2924) < reg2966) : $signed(forvar2948)) : reg2960);
                    end
                  if (reg2977)
                    begin
                      reg2988 <= reg2930[(4'h9):(3'h4)];
                      reg2989 <= reg2972;
                      reg2990 <= ((^$signed(reg2920[(2'h2):(2'h2)])) ?
                          (|forvar2958) : $signed(wire2363[(4'h8):(4'h8)]));
                    end
                  else
                    begin
                      reg2988 <= ((~|$unsigned((reg2956 ? reg2939 : reg2925))) ?
                          reg2989 : $signed(reg2975[(4'hc):(3'h5)]));
                      reg2989 <= $unsigned(reg2964[(4'h9):(2'h2)]);
                      reg2990 <= $signed((8'hb3));
                      reg2991 <= reg2961[(3'h5):(2'h2)];
                    end
                  reg2992 <= reg2987[(2'h2):(1'h0)];
                end
            end
        end
      else
        begin
          for (forvar2957 = (1'h0); (forvar2957 < (1'h1)); forvar2957 = (forvar2957 + (1'h1)))
            begin
              for (forvar2958 = (1'h0); (forvar2958 < (2'h3)); forvar2958 = (forvar2958 + (1'h1)))
                begin
                  for (forvar2959 = (1'h0); (forvar2959 < (2'h3)); forvar2959 = (forvar2959 + (1'h1)))
                    begin
                      reg2960 <= $signed(reg2954[(4'he):(4'ha)]);
                      reg2961 <= $unsigned(($unsigned(reg2990) ?
                          {(reg2945 ?
                                  reg2966 : reg2966)} : reg2925[(2'h3):(2'h3)]));
                      reg2962 <= {(~|$unsigned(reg2992[(2'h3):(1'h0)]))};
                    end
                end
            end
          for (forvar2963 = (1'h0); (forvar2963 < (2'h3)); forvar2963 = (forvar2963 + (1'h1)))
            begin
              for (forvar2964 = (1'h0); (forvar2964 < (1'h0)); forvar2964 = (forvar2964 + (1'h1)))
                begin
                  for (forvar2965 = (1'h0); (forvar2965 < (2'h3)); forvar2965 = (forvar2965 + (1'h1)))
                    begin
                      reg2966 <= $unsigned({$signed((~(8'ha0)))});
                      reg2967 <= ((~&(reg2977[(4'h9):(4'h9)] ?
                          (wire2368 <<< reg2952) : (-(8'hb5)))) >= $signed({forvar2924}));
                      reg2968 <= (~(|($unsigned(forvar2963) ?
                          $unsigned(reg2985) : reg2988[(3'h4):(2'h2)])));
                      reg2969 <= (($unsigned($unsigned(forvar2948)) ?
                              $signed({reg2920}) : $signed($unsigned(reg2968))) ?
                          reg2986[(1'h1):(1'h0)] : $unsigned(($signed(reg2940) < reg2926)));
                    end
                  for (forvar2970 = (1'h0); (forvar2970 < (2'h3)); forvar2970 = (forvar2970 + (1'h1)))
                    begin
                      reg2971 <= ($signed({$unsigned(reg2950)}) << $signed((reg2920[(3'h4):(2'h3)] ?
                          $unsigned(reg2968) : ((8'ha2) != (8'hb0)))));
                      reg2972 <= $unsigned({(8'hb6)});
                    end
                  if (forvar2938)
                    begin
                      reg2973 <= $unsigned((forvar2957[(1'h0):(1'h0)] ?
                          {$signed((8'ha2))} : reg2969));
                      reg2974 <= (+(&($signed(reg2965) ^~ (8'hb8))));
                      reg2975 <= forvar2932[(2'h2):(1'h0)];
                      reg2976 <= $unsigned(forvar2924[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg2973 <= (8'hb0);
                      reg2974 <= (~&(~^($unsigned(forvar2974) != (8'ha4))));
                      reg2975 <= reg2920;
                      reg2976 <= $unsigned($signed($signed((reg2989 ^~ reg2981))));
                    end
                  for (forvar2977 = (1'h0); (forvar2977 < (2'h2)); forvar2977 = (forvar2977 + (1'h1)))
                    begin
                      reg2978 <= $signed($unsigned(($unsigned(reg2950) ^~ (forvar2936 ?
                          (8'had) : reg2988))));
                      reg2979 <= wire2364;
                      reg2980 <= (~{($signed(reg2965) || (forvar2924 ?
                              reg2981 : forvar2948))});
                    end
                end
              reg2981 <= reg2930[(4'h8):(1'h0)];
              reg2982 <= $unsigned((forvar2979[(1'h1):(1'h1)] ?
                  (8'had) : $signed($signed(reg2928))));
              if ((forvar2938[(1'h0):(1'h0)] ?
                  $unsigned((~&$signed(forvar2970))) : $unsigned({(&(8'hb1))})))
                begin
                  if (wire2368)
                    begin
                      reg2983 <= {$signed((^$signed(forvar2964)))};
                    end
                  else
                    begin
                      reg2983 <= {(+$signed($unsigned(forvar2931)))};
                      reg2984 <= ({(&forvar2965[(3'h7):(3'h4)])} >= {reg2942});
                    end
                  if ($signed($signed($unsigned($signed(reg2955)))))
                    begin
                      reg2985 <= ($unsigned($signed((reg2980 >>> reg2940))) ?
                          reg2962 : reg2925);
                      reg2986 <= $unsigned(forvar2936);
                    end
                  else
                    begin
                      reg2985 <= ((^reg2986) ? {(8'ha6)} : (8'h9c));
                    end
                  if (reg2960)
                    begin
                      reg2987 <= (((reg2949 > $signed(forvar2943)) ?
                          $unsigned((~&reg2958)) : reg2964[(4'hb):(3'h7)]) <= $unsigned((reg2955[(2'h2):(2'h2)] == reg2989)));
                      reg2988 <= forvar2923;
                      reg2989 <= (+((reg2941 ?
                          {reg2950} : (8'hba)) || (|reg2974)));
                      reg2990 <= ((+reg2992[(1'h0):(1'h0)]) || reg2933[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2987 <= $signed($unsigned({forvar2921[(2'h3):(2'h2)]}));
                    end
                end
              else
                begin
                  if (((8'ha2) && $signed(reg2962[(4'he):(4'h9)])))
                    begin
                      reg2983 <= $unsigned(((-wire2368) ?
                          $unsigned(reg2976[(4'hf):(3'h5)]) : $signed($unsigned(reg2989))));
                      reg2984 <= forvar2923[(1'h0):(1'h0)];
                      reg2985 <= (~|(reg2986 * ((!reg2960) == $signed(reg2973))));
                    end
                  else
                    begin
                      reg2983 <= forvar2938;
                    end
                  for (forvar2986 = (1'h0); (forvar2986 < (1'h0)); forvar2986 = (forvar2986 + (1'h1)))
                    begin
                      reg2987 <= (+wire2368);
                      reg2988 <= $unsigned((^~$signed($signed((8'h9d)))));
                    end
                  reg2989 <= (($unsigned(forvar2970[(3'h7):(3'h6)]) << (&(reg2925 ?
                          reg2922 : reg2926))) ?
                      $unsigned($unsigned(wire2366[(1'h1):(1'h0)])) : $unsigned($signed((reg2933 && reg2971))));
                end
            end
          for (forvar2991 = (1'h0); (forvar2991 < (1'h0)); forvar2991 = (forvar2991 + (1'h1)))
            begin
              if (reg2952[(1'h0):(1'h0)])
                begin
                  for (forvar2992 = (1'h0); (forvar2992 < (1'h0)); forvar2992 = (forvar2992 + (1'h1)))
                    begin
                      reg2993 <= (^reg2978[(1'h0):(1'h0)]);
                      reg2994 <= $unsigned($unsigned(reg2940[(2'h3):(1'h0)]));
                      reg2995 <= $signed((reg2976 ^ wire2365));
                    end
                  reg2996 <= (((reg2933[(1'h1):(1'h1)] >> $signed((8'hb9))) ?
                          reg2960[(2'h2):(2'h2)] : $unsigned((forvar2938 != reg2976))) ?
                      reg2958[(1'h0):(1'h0)] : forvar2951);
                  if ($unsigned(reg2928[(1'h1):(1'h1)]))
                    begin
                      reg2997 <= ($unsigned((8'hac)) ?
                          (+{(8'hae)}) : (reg2985 ?
                              $signed(((8'ha5) ?
                                  forvar2936 : reg2961)) : $unsigned((reg2920 ?
                                  reg2956 : forvar2982))));
                      reg2998 <= forvar2991;
                      reg2999 <= $unsigned(reg2986[(1'h0):(1'h0)]);
                      reg3000 <= reg2956[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2997 <= reg2992[(1'h0):(1'h0)];
                      reg2998 <= (reg2920 ?
                          reg2972[(4'h8):(4'h8)] : (~|{reg2953}));
                      reg2999 <= ($signed({(reg2982 ~^ forvar2970)}) < $unsigned((-(!reg2946))));
                    end
                  for (forvar3001 = (1'h0); (forvar3001 < (1'h1)); forvar3001 = (forvar3001 + (1'h1)))
                    begin
                      reg3002 <= forvar2977[(3'h6):(3'h4)];
                      reg3003 <= ({$signed((forvar2931 ?
                                  forvar2983 : reg2947))} ?
                          (&((reg2946 || reg2941) ?
                              ((8'ha6) ?
                                  forvar2958 : wire2918) : $signed(reg2940))) : wire2367);
                      reg3004 <= ((((reg2986 < reg2928) >= $signed(forvar2982)) - ((|wire2369) ?
                          ((8'hb0) ?
                              forvar2957 : reg2990) : $unsigned(reg2968))) > (forvar2932[(2'h2):(1'h0)] || ((reg2993 >= reg2978) ?
                          $signed(forvar2921) : reg2935[(3'h4):(1'h0)])));
                      reg3005 <= $signed(($signed($signed(reg2965)) ?
                          (-$signed(forvar2932)) : $signed(forvar2964)));
                    end
                end
              else
                begin
                  for (forvar2992 = (1'h0); (forvar2992 < (2'h3)); forvar2992 = (forvar2992 + (1'h1)))
                    begin
                      reg2993 <= ($signed((!$signed(forvar3001))) ^~ $signed($signed($signed(forvar2974))));
                      reg2994 <= forvar3001[(1'h0):(1'h0)];
                    end
                  if ({((8'hb2) & (!forvar2970))})
                    begin
                      reg2995 <= (~^{((reg2995 ? wire2363 : (8'ha6)) ?
                              (|forvar2974) : reg2984)});
                    end
                  else
                    begin
                      reg2995 <= reg2947[(3'h7):(3'h5)];
                      reg2996 <= ((~&$unsigned(forvar2964[(3'h6):(1'h0)])) ?
                          ((^~(reg2941 ?
                              (8'hb1) : reg2958)) >>> $signed((reg2997 ?
                              forvar2958 : reg2967))) : (wire2918 * forvar2958[(3'h6):(3'h4)]));
                      reg2997 <= ((reg3005[(1'h1):(1'h1)] ?
                          $unsigned((reg2926 >>> (8'ha8))) : $unsigned($signed((8'ha6)))) + $unsigned(((8'hac) ?
                          (8'had) : forvar2977[(3'h5):(3'h4)])));
                    end
                  for (forvar2998 = (1'h0); (forvar2998 < (1'h1)); forvar2998 = (forvar2998 + (1'h1)))
                    begin
                      reg2999 <= $signed($unsigned((reg2941 ?
                          (8'h9f) : ((8'ha6) ? (8'hb7) : (8'ha6)))));
                      reg3000 <= reg2983;
                    end
                  for (forvar3001 = (1'h0); (forvar3001 < (1'h1)); forvar3001 = (forvar3001 + (1'h1)))
                    begin
                      reg3002 <= ($unsigned((~^{reg2933})) << $signed(reg2992));
                      reg3003 <= forvar2964[(3'h6):(2'h2)];
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar3006 = (1'h0); (forvar3006 < (1'h1)); forvar3006 = (forvar3006 + (1'h1)))
        begin
          for (forvar3007 = (1'h0); (forvar3007 < (2'h3)); forvar3007 = (forvar3007 + (1'h1)))
            begin
              if (forvar2932[(2'h3):(2'h2)])
                begin
                  for (forvar3008 = (1'h0); (forvar3008 < (2'h2)); forvar3008 = (forvar3008 + (1'h1)))
                    begin
                      reg3009 <= (forvar2957[(2'h2):(1'h0)] ~^ reg2963);
                      reg3010 <= forvar2991[(3'h4):(2'h3)];
                      reg3011 <= $unsigned(forvar2957);
                    end
                  reg3012 <= $unsigned(reg2956[(4'h9):(1'h1)]);
                  for (forvar3013 = (1'h0); (forvar3013 < (1'h1)); forvar3013 = (forvar3013 + (1'h1)))
                    begin
                      reg3014 <= (+($unsigned($signed(forvar2936)) >> (8'had)));
                      reg3015 <= $signed($unsigned(wire2363));
                    end
                end
              else
                begin
                  if ((reg2935 ? reg2954 : $unsigned(reg2952)))
                    begin
                      reg3008 <= $unsigned((($signed(reg2986) ?
                              (8'hab) : (-wire2365)) ?
                          {(~^reg2947)} : {(wire2366 ^ reg3010)}));
                      reg3009 <= $unsigned(($unsigned(forvar2921[(1'h0):(1'h0)]) ?
                          $unsigned(reg2949) : {(reg2979 * reg3015)}));
                    end
                  else
                    begin
                      reg3008 <= $unsigned(($signed($unsigned((8'ha0))) >> $unsigned($unsigned(forvar2982))));
                    end
                  for (forvar3010 = (1'h0); (forvar3010 < (1'h0)); forvar3010 = (forvar3010 + (1'h1)))
                    begin
                      reg3011 <= (^$unsigned($signed(reg2959)));
                      reg3012 <= $signed((forvar2978 ?
                          (forvar2977[(2'h3):(1'h1)] == reg2933) : reg2976));
                    end
                  for (forvar3013 = (1'h0); (forvar3013 < (2'h2)); forvar3013 = (forvar3013 + (1'h1)))
                    begin
                      reg3014 <= forvar2921[(3'h4):(3'h4)];
                    end
                  for (forvar3015 = (1'h0); (forvar3015 < (2'h2)); forvar3015 = (forvar3015 + (1'h1)))
                    begin
                      reg3016 <= ((^~(reg2991 ?
                          (^reg2927) : (reg2983 ?
                              (8'hb2) : reg2964))) < (^((forvar2963 <<< reg2998) ?
                          {forvar2965} : reg2928[(2'h3):(1'h1)])));
                      reg3017 <= $unsigned($unsigned((~(reg2985 ?
                          reg2980 : reg2994))));
                      reg3018 <= $unsigned(reg2964);
                      reg3019 <= forvar2977;
                    end
                end
              for (forvar3020 = (1'h0); (forvar3020 < (1'h0)); forvar3020 = (forvar3020 + (1'h1)))
                begin
                  reg3021 <= reg2986[(1'h1):(1'h0)];
                  for (forvar3022 = (1'h0); (forvar3022 < (2'h3)); forvar3022 = (forvar3022 + (1'h1)))
                    begin
                      reg3023 <= $unsigned(reg2989[(4'h9):(3'h4)]);
                      reg3024 <= forvar2923;
                    end
                end
              reg3025 <= ($signed({(^~forvar2963)}) ?
                  $signed($signed(reg3012)) : forvar2948);
              for (forvar3026 = (1'h0); (forvar3026 < (2'h3)); forvar3026 = (forvar3026 + (1'h1)))
                begin
                  for (forvar3027 = (1'h0); (forvar3027 < (2'h3)); forvar3027 = (forvar3027 + (1'h1)))
                    begin
                      reg3028 <= forvar2938[(1'h1):(1'h1)];
                      reg3029 <= $signed((~|$signed((reg2920 ?
                          reg2998 : reg3016))));
                      reg3030 <= (forvar3027[(3'h6):(3'h5)] << {($signed(reg2944) >= (8'hb9))});
                      reg3031 <= (~reg2922[(3'h4):(2'h2)]);
                    end
                end
            end
        end
    end
  assign wire3032 = reg3024;
  assign wire3033 = (~&reg2961);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2370
#( parameter param2917 = ((&(~^(8'ha1))) ? ((((8'hb1) + (8'ha9)) ^ (|(8'hae))) ? (!(~|(8'hac))) : (|(^(8'hac)))) : (({(8'hba)} ~^ ((8'ha4) != (8'ha0))) <= {(~(8'ha2))})) )
(y, clk, wire2374, wire2373, wire2372, wire2371);
  output wire [(32'h174e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire2374;
  input wire signed [(4'hd):(1'h0)] wire2373;
  input wire signed [(3'h6):(1'h0)] wire2372;
  input wire [(3'h5):(1'h0)] wire2371;
  reg signed [(5'h10):(1'h0)] reg2916 = (1'h0);
  reg [(4'he):(1'h0)] reg2915 = (1'h0);
  reg [(4'hf):(1'h0)] reg2914 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2913 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2912 = (1'h0);
  reg [(4'hc):(1'h0)] reg2909 = (1'h0);
  reg [(4'hb):(1'h0)] reg2907 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2906 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2903 = (1'h0);
  reg [(4'he):(1'h0)] reg2900 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2898 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2895 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2886 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2892 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2890 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2888 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2887 = (1'h0);
  reg [(3'h4):(1'h0)] reg2912 = (1'h0);
  reg [(4'ha):(1'h0)] reg2911 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2910 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2909 = (1'h0);
  reg [(4'he):(1'h0)] reg2908 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2907 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2906 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2905 = (1'h0);
  reg [(4'ha):(1'h0)] reg2904 = (1'h0);
  reg [(4'hb):(1'h0)] reg2903 = (1'h0);
  reg [(2'h2):(1'h0)] reg2902 = (1'h0);
  reg [(3'h5):(1'h0)] reg2901 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2900 = (1'h0);
  reg [(4'hf):(1'h0)] reg2899 = (1'h0);
  reg [(4'he):(1'h0)] reg2898 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2897 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2896 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2895 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2894 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2893 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2892 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2891 = (1'h0);
  reg [(4'hc):(1'h0)] reg2890 = (1'h0);
  reg [(3'h5):(1'h0)] reg2889 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2888 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2887 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2886 = (1'h0);
  reg [(5'h10):(1'h0)] reg2872 = (1'h0);
  reg [(4'he):(1'h0)] reg2885 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2884 = (1'h0);
  reg [(3'h5):(1'h0)] reg2883 = (1'h0);
  reg [(3'h7):(1'h0)] reg2882 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2881 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2880 = (1'h0);
  reg [(4'hc):(1'h0)] reg2879 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2878 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2877 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2876 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2875 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2874 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2873 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2872 = (1'h0);
  reg [(2'h3):(1'h0)] reg2871 = (1'h0);
  reg [(3'h6):(1'h0)] reg2870 = (1'h0);
  reg [(3'h6):(1'h0)] reg2869 = (1'h0);
  reg [(3'h5):(1'h0)] reg2868 = (1'h0);
  reg [(4'hd):(1'h0)] reg2867 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2866 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2865 = (1'h0);
  reg [(2'h2):(1'h0)] reg2864 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2863 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2862 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2861 = (1'h0);
  reg [(4'ha):(1'h0)] reg2860 = (1'h0);
  reg [(3'h6):(1'h0)] reg2859 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2858 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2853 = (1'h0);
  reg [(3'h5):(1'h0)] reg2852 = (1'h0);
  reg [(3'h5):(1'h0)] reg2857 = (1'h0);
  reg [(5'h10):(1'h0)] reg2856 = (1'h0);
  reg [(4'hf):(1'h0)] reg2855 = (1'h0);
  reg [(4'h9):(1'h0)] reg2854 = (1'h0);
  reg [(3'h6):(1'h0)] reg2853 = (1'h0);
  reg [(4'he):(1'h0)] forvar2852 = (1'h0);
  reg [(3'h7):(1'h0)] reg2851 = (1'h0);
  reg [(4'hd):(1'h0)] reg2850 = (1'h0);
  reg [(4'hf):(1'h0)] reg2849 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2848 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2847 = (1'h0);
  reg [(4'he):(1'h0)] reg2846 = (1'h0);
  reg [(4'hf):(1'h0)] reg2845 = (1'h0);
  reg [(3'h7):(1'h0)] reg2844 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2843 = (1'h0);
  reg [(4'h9):(1'h0)] reg2842 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2841 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2840 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2839 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2824 = (1'h0);
  reg [(4'hb):(1'h0)] reg2823 = (1'h0);
  reg [(4'hd):(1'h0)] reg2821 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2816 = (1'h0);
  reg [(4'he):(1'h0)] reg2838 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2837 = (1'h0);
  reg [(4'hf):(1'h0)] reg2836 = (1'h0);
  reg [(3'h6):(1'h0)] reg2835 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2834 = (1'h0);
  reg [(5'h10):(1'h0)] reg2833 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2832 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2831 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2830 = (1'h0);
  reg [(4'hb):(1'h0)] reg2829 = (1'h0);
  reg [(2'h3):(1'h0)] reg2828 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2827 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2826 = (1'h0);
  reg [(3'h7):(1'h0)] reg2825 = (1'h0);
  reg [(2'h2):(1'h0)] reg2824 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2823 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2822 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2821 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2820 = (1'h0);
  reg [(3'h6):(1'h0)] reg2819 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2818 = (1'h0);
  reg [(2'h2):(1'h0)] reg2817 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2816 = (1'h0);
  reg [(2'h3):(1'h0)] reg2815 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2814 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2813 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2812 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2811 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2810 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2809 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2808 = (1'h0);
  reg [(4'he):(1'h0)] reg2807 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2806 = (1'h0);
  reg [(3'h4):(1'h0)] reg2805 = (1'h0);
  reg [(2'h2):(1'h0)] reg2804 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2803 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2802 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2801 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2800 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2799 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2798 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2797 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2796 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2795 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2794 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2792 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2785 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2783 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2793 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2792 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2791 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2790 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2787 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2784 = (1'h0);
  reg [(5'h10):(1'h0)] reg2773 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2767 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2760 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2759 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2763 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2761 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2756 = (1'h0);
  reg [(4'hc):(1'h0)] reg2777 = (1'h0);
  reg [(4'hc):(1'h0)] reg2790 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2789 = (1'h0);
  reg [(3'h6):(1'h0)] reg2788 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2787 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2786 = (1'h0);
  reg [(3'h5):(1'h0)] reg2785 = (1'h0);
  reg [(4'hf):(1'h0)] reg2784 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2783 = (1'h0);
  reg [(2'h2):(1'h0)] reg2782 = (1'h0);
  reg [(5'h10):(1'h0)] reg2781 = (1'h0);
  reg [(3'h4):(1'h0)] reg2780 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2779 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2778 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2777 = (1'h0);
  reg [(4'hf):(1'h0)] reg2776 = (1'h0);
  reg [(4'h8):(1'h0)] reg2775 = (1'h0);
  reg [(4'hf):(1'h0)] reg2774 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2773 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2772 = (1'h0);
  reg [(2'h2):(1'h0)] reg2771 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2770 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2769 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2768 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2767 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2766 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2765 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2764 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2763 = (1'h0);
  reg [(3'h5):(1'h0)] reg2762 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2761 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2760 = (1'h0);
  reg [(4'he):(1'h0)] reg2759 = (1'h0);
  reg [(4'hd):(1'h0)] reg2758 = (1'h0);
  reg [(4'hf):(1'h0)] reg2757 = (1'h0);
  reg [(4'hf):(1'h0)] reg2756 = (1'h0);
  reg [(4'he):(1'h0)] reg2755 = (1'h0);
  reg [(4'h8):(1'h0)] reg2754 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2753 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2752 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2751 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2750 = (1'h0);
  reg [(4'hf):(1'h0)] reg2749 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2748 = (1'h0);
  reg [(2'h2):(1'h0)] reg2747 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2746 = (1'h0);
  reg [(4'he):(1'h0)] forvar2744 = (1'h0);
  reg [(4'h9):(1'h0)] reg2742 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2739 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2746 = (1'h0);
  reg [(4'ha):(1'h0)] reg2745 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2744 = (1'h0);
  reg [(4'h9):(1'h0)] reg2743 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2742 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2741 = (1'h0);
  reg [(4'h9):(1'h0)] reg2740 = (1'h0);
  reg [(5'h10):(1'h0)] reg2739 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2738 = (1'h0);
  reg [(2'h2):(1'h0)] reg2737 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2736 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2734 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2735 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2734 = (1'h0);
  reg [(5'h10):(1'h0)] reg2733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2732 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2731 = (1'h0);
  reg [(2'h2):(1'h0)] reg2730 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2729 = (1'h0);
  reg [(5'h10):(1'h0)] reg2729 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2728 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2720 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2727 = (1'h0);
  reg [(4'hf):(1'h0)] reg2726 = (1'h0);
  reg [(4'ha):(1'h0)] reg2725 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2721 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2717 = (1'h0);
  reg [(3'h4):(1'h0)] reg2716 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2703 = (1'h0);
  reg [(4'hf):(1'h0)] reg2697 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2694 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2687 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2683 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2682 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2680 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2676 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2673 = (1'h0);
  reg [(2'h2):(1'h0)] reg2672 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2724 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2723 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2722 = (1'h0);
  reg [(3'h7):(1'h0)] reg2721 = (1'h0);
  reg [(4'hf):(1'h0)] reg2720 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2719 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2718 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2711 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2706 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2702 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2698 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2693 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2689 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2688 = (1'h0);
  reg [(3'h4):(1'h0)] reg2717 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2716 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2715 = (1'h0);
  reg [(4'hb):(1'h0)] reg2714 = (1'h0);
  reg [(4'hf):(1'h0)] reg2713 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2712 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2711 = (1'h0);
  reg [(3'h4):(1'h0)] reg2710 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2708 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2704 = (1'h0);
  reg [(4'hd):(1'h0)] reg2709 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2708 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2707 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2706 = (1'h0);
  reg [(4'ha):(1'h0)] reg2705 = (1'h0);
  reg [(4'ha):(1'h0)] reg2704 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2703 = (1'h0);
  reg [(4'he):(1'h0)] forvar2702 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2701 = (1'h0);
  reg [(3'h7):(1'h0)] reg2700 = (1'h0);
  reg [(4'he):(1'h0)] reg2699 = (1'h0);
  reg [(3'h4):(1'h0)] reg2698 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2697 = (1'h0);
  reg [(3'h4):(1'h0)] reg2696 = (1'h0);
  reg [(3'h6):(1'h0)] reg2695 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2694 = (1'h0);
  reg [(4'he):(1'h0)] forvar2693 = (1'h0);
  reg [(3'h5):(1'h0)] reg2692 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2691 = (1'h0);
  reg [(4'h8):(1'h0)] reg2690 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2689 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2688 = (1'h0);
  reg [(3'h5):(1'h0)] reg2687 = (1'h0);
  reg [(4'hf):(1'h0)] reg2686 = (1'h0);
  reg [(5'h10):(1'h0)] reg2685 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2684 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2683 = (1'h0);
  reg [(2'h3):(1'h0)] reg2682 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2678 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2677 = (1'h0);
  reg [(4'he):(1'h0)] reg2674 = (1'h0);
  reg [(4'he):(1'h0)] reg2681 = (1'h0);
  reg [(4'ha):(1'h0)] reg2680 = (1'h0);
  reg [(4'hd):(1'h0)] reg2679 = (1'h0);
  reg [(2'h2):(1'h0)] reg2678 = (1'h0);
  reg [(4'he):(1'h0)] forvar2677 = (1'h0);
  reg [(3'h4):(1'h0)] reg2676 = (1'h0);
  reg [(4'ha):(1'h0)] reg2675 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2674 = (1'h0);
  reg [(4'hd):(1'h0)] reg2673 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2672 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2671 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2671 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2670 = (1'h0);
  reg [(4'h9):(1'h0)] reg2669 = (1'h0);
  reg [(3'h5):(1'h0)] reg2668 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2667 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2666 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2665 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2664 = (1'h0);
  reg [(3'h5):(1'h0)] reg2663 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2662 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2661 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2660 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2659 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2658 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2657 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2656 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2655 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2654 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2653 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2651 = (1'h0);
  reg [(3'h4):(1'h0)] reg2652 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2651 = (1'h0);
  reg [(2'h3):(1'h0)] reg2650 = (1'h0);
  reg [(3'h6):(1'h0)] reg2649 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2648 = (1'h0);
  reg [(4'h8):(1'h0)] reg2647 = (1'h0);
  reg [(4'hb):(1'h0)] reg2646 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2645 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2644 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2643 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2642 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2641 = (1'h0);
  reg [(3'h6):(1'h0)] reg2640 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2639 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2639 = (1'h0);
  reg [(4'hd):(1'h0)] reg2638 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2637 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2636 = (1'h0);
  reg [(4'hc):(1'h0)] reg2635 = (1'h0);
  reg [(5'h10):(1'h0)] reg2634 = (1'h0);
  reg [(4'hf):(1'h0)] reg2633 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2632 = (1'h0);
  reg [(5'h10):(1'h0)] reg2631 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2630 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2629 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2628 = (1'h0);
  reg [(4'he):(1'h0)] forvar2627 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2559 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2556 = (1'h0);
  reg [(4'hb):(1'h0)] reg2553 = (1'h0);
  reg [(4'he):(1'h0)] forvar2552 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2546 = (1'h0);
  reg [(4'hf):(1'h0)] reg2544 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2618 = (1'h0);
  reg [(4'ha):(1'h0)] reg2616 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2611 = (1'h0);
  reg [(4'hf):(1'h0)] reg2606 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2608 = (1'h0);
  reg [(4'hd):(1'h0)] reg2601 = (1'h0);
  reg [(3'h4):(1'h0)] reg2600 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2626 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2625 = (1'h0);
  reg [(3'h4):(1'h0)] reg2624 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2623 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2622 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2621 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2612 = (1'h0);
  reg [(3'h5):(1'h0)] reg2620 = (1'h0);
  reg [(4'hf):(1'h0)] reg2619 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2618 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2617 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2616 = (1'h0);
  reg [(3'h5):(1'h0)] reg2615 = (1'h0);
  reg [(4'h8):(1'h0)] reg2614 = (1'h0);
  reg [(4'h8):(1'h0)] reg2613 = (1'h0);
  reg [(4'hf):(1'h0)] reg2612 = (1'h0);
  reg [(4'ha):(1'h0)] reg2611 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2610 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2609 = (1'h0);
  reg [(3'h6):(1'h0)] reg2608 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2607 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2606 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2605 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2604 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2603 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2602 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2601 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2600 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2598 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2597 = (1'h0);
  reg [(2'h3):(1'h0)] reg2593 = (1'h0);
  reg [(2'h2):(1'h0)] reg2599 = (1'h0);
  reg [(3'h6):(1'h0)] reg2598 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2597 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2596 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2595 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2594 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2593 = (1'h0);
  reg [(4'hd):(1'h0)] reg2592 = (1'h0);
  reg [(5'h10):(1'h0)] reg2591 = (1'h0);
  reg [(4'hb):(1'h0)] reg2590 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2589 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2588 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2587 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2586 = (1'h0);
  reg [(3'h5):(1'h0)] reg2585 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2584 = (1'h0);
  reg [(3'h7):(1'h0)] reg2584 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2583 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2582 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2581 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2580 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2579 = (1'h0);
  reg [(2'h3):(1'h0)] reg2578 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2577 = (1'h0);
  reg [(4'hf):(1'h0)] reg2576 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2575 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2574 = (1'h0);
  reg [(4'hc):(1'h0)] reg2573 = (1'h0);
  reg [(3'h7):(1'h0)] reg2572 = (1'h0);
  reg [(4'h8):(1'h0)] reg2571 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2570 = (1'h0);
  reg [(3'h4):(1'h0)] reg2569 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2567 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2564 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2561 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2558 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2557 = (1'h0);
  reg [(3'h4):(1'h0)] reg2566 = (1'h0);
  reg [(5'h10):(1'h0)] reg2565 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2564 = (1'h0);
  reg [(4'he):(1'h0)] reg2563 = (1'h0);
  reg [(2'h3):(1'h0)] reg2562 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2561 = (1'h0);
  reg [(4'hb):(1'h0)] reg2560 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2559 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2558 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2557 = (1'h0);
  reg [(3'h4):(1'h0)] reg2556 = (1'h0);
  reg [(4'hf):(1'h0)] reg2555 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2554 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2553 = (1'h0);
  reg [(2'h2):(1'h0)] reg2552 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2551 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2550 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2549 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2548 = (1'h0);
  reg [(3'h4):(1'h0)] reg2547 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2546 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2545 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2544 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2521 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2518 = (1'h0);
  reg [(3'h6):(1'h0)] reg2529 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2527 = (1'h0);
  reg [(4'ha):(1'h0)] reg2525 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2524 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2516 = (1'h0);
  reg [(4'hb):(1'h0)] reg2543 = (1'h0);
  reg [(3'h4):(1'h0)] reg2542 = (1'h0);
  reg [(4'ha):(1'h0)] reg2541 = (1'h0);
  reg [(4'hb):(1'h0)] reg2540 = (1'h0);
  reg [(4'hc):(1'h0)] reg2539 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2537 = (1'h0);
  reg [(4'h9):(1'h0)] reg2536 = (1'h0);
  reg [(2'h3):(1'h0)] reg2538 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2537 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2536 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2535 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2534 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2533 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2532 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2531 = (1'h0);
  reg [(3'h5):(1'h0)] reg2530 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2529 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2528 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2527 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2526 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2525 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2524 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2523 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2522 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2521 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2520 = (1'h0);
  reg [(4'hf):(1'h0)] reg2519 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2518 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2517 = (1'h0);
  reg [(3'h5):(1'h0)] reg2516 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2515 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire2514;
  wire signed [(2'h2):(1'h0)] wire2513;
  wire [(4'ha):(1'h0)] wire2512;
  wire [(4'he):(1'h0)] wire2511;
  reg [(4'hf):(1'h0)] reg2510 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2509 = (1'h0);
  reg [(3'h7):(1'h0)] reg2508 = (1'h0);
  reg [(3'h6):(1'h0)] reg2507 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2506 = (1'h0);
  reg [(4'hf):(1'h0)] reg2505 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2504 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2503 = (1'h0);
  reg [(3'h4):(1'h0)] reg2502 = (1'h0);
  reg [(4'h8):(1'h0)] reg2501 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2500 = (1'h0);
  reg [(4'hc):(1'h0)] reg2499 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2498 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2497 = (1'h0);
  reg [(4'h8):(1'h0)] reg2496 = (1'h0);
  reg [(4'hf):(1'h0)] reg2495 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2493 = (1'h0);
  reg [(3'h6):(1'h0)] reg2494 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2493 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2489 = (1'h0);
  reg [(4'hd):(1'h0)] reg2492 = (1'h0);
  reg [(4'hf):(1'h0)] reg2491 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2490 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2489 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2488 = (1'h0);
  reg [(4'h8):(1'h0)] reg2487 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2486 = (1'h0);
  reg [(4'hd):(1'h0)] reg2478 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2476 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2475 = (1'h0);
  reg [(2'h2):(1'h0)] reg2473 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2469 = (1'h0);
  reg [(4'h9):(1'h0)] reg2468 = (1'h0);
  reg [(4'hf):(1'h0)] reg2465 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2458 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2485 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2484 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2483 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2482 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2481 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2480 = (1'h0);
  reg [(3'h7):(1'h0)] reg2479 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2478 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2477 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2476 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2475 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2474 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2473 = (1'h0);
  reg [(4'ha):(1'h0)] reg2472 = (1'h0);
  reg [(4'h9):(1'h0)] reg2471 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2470 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2469 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2468 = (1'h0);
  reg [(4'hb):(1'h0)] reg2467 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2466 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2465 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2464 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2463 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2462 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2461 = (1'h0);
  reg [(4'he):(1'h0)] reg2460 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2459 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2458 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2457 = (1'h0);
  reg [(4'he):(1'h0)] reg2456 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2455 = (1'h0);
  reg [(4'hf):(1'h0)] reg2454 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2453 = (1'h0);
  reg [(3'h7):(1'h0)] reg2452 = (1'h0);
  reg [(4'hb):(1'h0)] reg2451 = (1'h0);
  reg [(4'he):(1'h0)] reg2450 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2449 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2448 = (1'h0);
  reg [(2'h2):(1'h0)] reg2447 = (1'h0);
  reg [(4'hc):(1'h0)] reg2446 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2445 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2444 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2443 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2442 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2441 = (1'h0);
  reg [(4'hf):(1'h0)] reg2440 = (1'h0);
  reg [(2'h2):(1'h0)] reg2439 = (1'h0);
  reg [(4'he):(1'h0)] reg2438 = (1'h0);
  reg [(4'h9):(1'h0)] reg2437 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2436 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2435 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2434 = (1'h0);
  reg [(4'hb):(1'h0)] reg2433 = (1'h0);
  reg [(4'hc):(1'h0)] reg2432 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2431 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2427 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2426 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2430 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2429 = (1'h0);
  reg [(4'hb):(1'h0)] reg2428 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2427 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2426 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2425 = (1'h0);
  reg [(4'h8):(1'h0)] reg2424 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2423 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2422 = (1'h0);
  reg [(2'h2):(1'h0)] reg2421 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2420 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2419 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2418 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2417 = (1'h0);
  reg [(4'he):(1'h0)] reg2409 = (1'h0);
  reg [(4'hd):(1'h0)] reg2407 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2406 = (1'h0);
  reg [(4'hd):(1'h0)] reg2416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2415 = (1'h0);
  reg [(4'hb):(1'h0)] reg2414 = (1'h0);
  reg [(4'hf):(1'h0)] reg2413 = (1'h0);
  reg [(5'h10):(1'h0)] reg2412 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2411 = (1'h0);
  reg [(4'h8):(1'h0)] reg2410 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2409 = (1'h0);
  reg [(4'h8):(1'h0)] reg2408 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2407 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2406 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2405 = (1'h0);
  reg [(4'hc):(1'h0)] reg2404 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2403 = (1'h0);
  reg [(2'h3):(1'h0)] reg2402 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2401 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2400 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2399 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2398 = (1'h0);
  reg [(3'h7):(1'h0)] reg2397 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2396 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2395 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2394 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2393 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2392 = (1'h0);
  reg [(4'hc):(1'h0)] reg2391 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2390 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2389 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2388 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2383 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2381 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2387 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2386 = (1'h0);
  reg [(3'h6):(1'h0)] reg2385 = (1'h0);
  reg [(4'hb):(1'h0)] reg2384 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2383 = (1'h0);
  reg [(4'he):(1'h0)] reg2382 = (1'h0);
  reg [(3'h5):(1'h0)] reg2381 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2380 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2379 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire2378;
  wire signed [(4'h8):(1'h0)] wire2377;
  wire [(4'hf):(1'h0)] wire2376;
  wire [(4'hb):(1'h0)] wire2375;
  assign y = {reg2916,
                 reg2915,
                 reg2914,
                 forvar2913,
                 forvar2912,
                 reg2909,
                 reg2907,
                 forvar2906,
                 forvar2903,
                 reg2900,
                 forvar2898,
                 reg2895,
                 forvar2886,
                 reg2892,
                 forvar2890,
                 reg2888,
                 reg2887,
                 reg2912,
                 reg2911,
                 reg2910,
                 forvar2909,
                 reg2908,
                 forvar2907,
                 reg2906,
                 forvar2905,
                 reg2904,
                 reg2903,
                 reg2902,
                 reg2901,
                 forvar2900,
                 reg2899,
                 reg2898,
                 reg2897,
                 reg2896,
                 forvar2895,
                 forvar2894,
                 reg2893,
                 forvar2892,
                 reg2891,
                 reg2890,
                 reg2889,
                 forvar2888,
                 forvar2887,
                 reg2886,
                 reg2872,
                 reg2885,
                 reg2884,
                 reg2883,
                 reg2882,
                 forvar2881,
                 reg2880,
                 reg2879,
                 reg2878,
                 reg2877,
                 reg2876,
                 reg2875,
                 reg2874,
                 forvar2873,
                 forvar2872,
                 reg2871,
                 reg2870,
                 reg2869,
                 reg2868,
                 reg2867,
                 forvar2866,
                 reg2865,
                 reg2864,
                 forvar2863,
                 reg2862,
                 reg2861,
                 reg2860,
                 reg2859,
                 forvar2858,
                 forvar2853,
                 reg2852,
                 reg2857,
                 reg2856,
                 reg2855,
                 reg2854,
                 reg2853,
                 forvar2852,
                 reg2851,
                 reg2850,
                 reg2849,
                 forvar2848,
                 forvar2847,
                 reg2846,
                 reg2845,
                 reg2844,
                 reg2843,
                 reg2842,
                 forvar2841,
                 forvar2840,
                 forvar2839,
                 forvar2824,
                 reg2823,
                 reg2821,
                 reg2816,
                 reg2838,
                 forvar2837,
                 reg2836,
                 reg2835,
                 reg2834,
                 reg2833,
                 reg2832,
                 forvar2831,
                 forvar2830,
                 reg2829,
                 reg2828,
                 reg2827,
                 reg2826,
                 reg2825,
                 reg2824,
                 forvar2823,
                 reg2822,
                 forvar2821,
                 forvar2820,
                 reg2819,
                 reg2818,
                 reg2817,
                 forvar2816,
                 reg2815,
                 reg2814,
                 reg2813,
                 reg2812,
                 forvar2811,
                 forvar2810,
                 reg2809,
                 reg2808,
                 reg2807,
                 reg2806,
                 reg2805,
                 reg2804,
                 reg2803,
                 forvar2802,
                 reg2801,
                 forvar2800,
                 forvar2799,
                 reg2798,
                 reg2797,
                 reg2796,
                 reg2795,
                 forvar2794,
                 forvar2792,
                 forvar2785,
                 reg2783,
                 reg2793,
                 reg2792,
                 reg2791,
                 forvar2790,
                 reg2787,
                 forvar2784,
                 reg2773,
                 forvar2767,
                 reg2760,
                 forvar2759,
                 forvar2763,
                 reg2761,
                 forvar2756,
                 reg2777,
                 reg2790,
                 reg2789,
                 reg2788,
                 forvar2787,
                 reg2786,
                 reg2785,
                 reg2784,
                 forvar2783,
                 reg2782,
                 reg2781,
                 reg2780,
                 reg2779,
                 forvar2778,
                 forvar2777,
                 reg2776,
                 reg2775,
                 reg2774,
                 forvar2773,
                 reg2772,
                 reg2771,
                 reg2770,
                 reg2769,
                 forvar2768,
                 reg2767,
                 reg2766,
                 reg2765,
                 reg2764,
                 reg2763,
                 reg2762,
                 forvar2761,
                 forvar2760,
                 reg2759,
                 reg2758,
                 reg2757,
                 reg2756,
                 reg2755,
                 reg2754,
                 forvar2753,
                 forvar2752,
                 forvar2751,
                 reg2750,
                 reg2749,
                 reg2748,
                 reg2747,
                 forvar2746,
                 forvar2744,
                 reg2742,
                 forvar2739,
                 reg2746,
                 reg2745,
                 reg2744,
                 reg2743,
                 forvar2742,
                 reg2741,
                 reg2740,
                 reg2739,
                 forvar2738,
                 reg2737,
                 reg2736,
                 forvar2734,
                 reg2735,
                 reg2734,
                 reg2733,
                 reg2732,
                 reg2731,
                 reg2730,
                 forvar2729,
                 reg2729,
                 forvar2728,
                 forvar2720,
                 reg2727,
                 reg2726,
                 reg2725,
                 forvar2721,
                 forvar2717,
                 reg2716,
                 forvar2703,
                 reg2697,
                 forvar2694,
                 forvar2687,
                 reg2683,
                 forvar2682,
                 forvar2680,
                 forvar2676,
                 forvar2673,
                 reg2672,
                 reg2724,
                 reg2723,
                 reg2722,
                 reg2721,
                 reg2720,
                 reg2719,
                 reg2718,
                 forvar2711,
                 forvar2706,
                 reg2702,
                 forvar2698,
                 reg2693,
                 forvar2689,
                 forvar2688,
                 reg2717,
                 forvar2716,
                 reg2715,
                 reg2714,
                 reg2713,
                 reg2712,
                 reg2711,
                 reg2710,
                 reg2708,
                 forvar2704,
                 reg2709,
                 forvar2708,
                 reg2707,
                 reg2706,
                 reg2705,
                 reg2704,
                 reg2703,
                 forvar2702,
                 reg2701,
                 reg2700,
                 reg2699,
                 reg2698,
                 forvar2697,
                 reg2696,
                 reg2695,
                 reg2694,
                 forvar2693,
                 reg2692,
                 reg2691,
                 reg2690,
                 reg2689,
                 reg2688,
                 reg2687,
                 reg2686,
                 reg2685,
                 reg2684,
                 forvar2683,
                 reg2682,
                 forvar2678,
                 reg2677,
                 reg2674,
                 reg2681,
                 reg2680,
                 reg2679,
                 reg2678,
                 forvar2677,
                 reg2676,
                 reg2675,
                 forvar2674,
                 reg2673,
                 forvar2672,
                 forvar2671,
                 reg2671,
                 reg2670,
                 reg2669,
                 reg2668,
                 reg2667,
                 forvar2666,
                 reg2665,
                 reg2664,
                 reg2663,
                 reg2662,
                 forvar2661,
                 reg2660,
                 reg2659,
                 reg2658,
                 reg2657,
                 forvar2656,
                 forvar2655,
                 reg2654,
                 reg2653,
                 reg2651,
                 reg2652,
                 forvar2651,
                 reg2650,
                 reg2649,
                 reg2648,
                 reg2647,
                 reg2646,
                 reg2645,
                 reg2644,
                 forvar2643,
                 reg2642,
                 reg2641,
                 reg2640,
                 forvar2639,
                 reg2639,
                 reg2638,
                 reg2637,
                 reg2636,
                 reg2635,
                 reg2634,
                 reg2633,
                 reg2632,
                 reg2631,
                 reg2630,
                 forvar2629,
                 forvar2628,
                 forvar2627,
                 forvar2559,
                 forvar2556,
                 reg2553,
                 forvar2552,
                 forvar2546,
                 reg2544,
                 forvar2618,
                 reg2616,
                 forvar2611,
                 reg2606,
                 forvar2608,
                 reg2601,
                 reg2600,
                 reg2626,
                 reg2625,
                 reg2624,
                 reg2623,
                 forvar2622,
                 forvar2621,
                 forvar2612,
                 reg2620,
                 reg2619,
                 reg2618,
                 reg2617,
                 forvar2616,
                 reg2615,
                 reg2614,
                 reg2613,
                 reg2612,
                 reg2611,
                 reg2610,
                 reg2609,
                 reg2608,
                 reg2607,
                 forvar2606,
                 reg2605,
                 reg2604,
                 reg2603,
                 reg2602,
                 forvar2601,
                 forvar2600,
                 forvar2598,
                 reg2597,
                 reg2593,
                 reg2599,
                 reg2598,
                 forvar2597,
                 reg2596,
                 reg2595,
                 reg2594,
                 forvar2593,
                 reg2592,
                 reg2591,
                 reg2590,
                 forvar2589,
                 reg2588,
                 reg2587,
                 forvar2586,
                 reg2585,
                 forvar2584,
                 reg2584,
                 forvar2583,
                 reg2582,
                 reg2581,
                 reg2580,
                 reg2579,
                 reg2578,
                 forvar2577,
                 reg2576,
                 reg2575,
                 reg2574,
                 reg2573,
                 reg2572,
                 reg2571,
                 reg2570,
                 reg2569,
                 reg2568,
                 reg2567,
                 reg2564,
                 forvar2561,
                 reg2558,
                 forvar2557,
                 reg2566,
                 reg2565,
                 forvar2564,
                 reg2563,
                 reg2562,
                 reg2561,
                 reg2560,
                 reg2559,
                 forvar2558,
                 reg2557,
                 reg2556,
                 reg2555,
                 reg2554,
                 forvar2553,
                 reg2552,
                 reg2551,
                 reg2550,
                 reg2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 forvar2545,
                 forvar2544,
                 forvar2521,
                 forvar2518,
                 reg2529,
                 reg2527,
                 reg2525,
                 reg2524,
                 forvar2516,
                 reg2543,
                 reg2542,
                 reg2541,
                 reg2540,
                 reg2539,
                 forvar2537,
                 reg2536,
                 reg2538,
                 reg2537,
                 forvar2536,
                 reg2535,
                 forvar2534,
                 reg2533,
                 reg2532,
                 reg2531,
                 reg2530,
                 forvar2529,
                 reg2528,
                 forvar2527,
                 reg2526,
                 forvar2525,
                 forvar2524,
                 reg2523,
                 reg2522,
                 reg2521,
                 reg2520,
                 reg2519,
                 reg2518,
                 reg2517,
                 reg2516,
                 forvar2515,
                 wire2514,
                 wire2513,
                 wire2512,
                 wire2511,
                 reg2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 forvar2506,
                 reg2505,
                 forvar2504,
                 reg2503,
                 reg2502,
                 reg2501,
                 reg2500,
                 reg2499,
                 reg2498,
                 forvar2497,
                 reg2496,
                 reg2495,
                 reg2493,
                 reg2494,
                 forvar2493,
                 forvar2489,
                 reg2492,
                 reg2491,
                 reg2490,
                 reg2489,
                 forvar2488,
                 reg2487,
                 forvar2486,
                 reg2478,
                 forvar2476,
                 forvar2475,
                 reg2473,
                 forvar2469,
                 reg2468,
                 reg2465,
                 reg2458,
                 reg2485,
                 reg2484,
                 reg2483,
                 reg2482,
                 reg2481,
                 reg2480,
                 reg2479,
                 forvar2478,
                 reg2477,
                 reg2476,
                 reg2475,
                 reg2474,
                 forvar2473,
                 reg2472,
                 reg2471,
                 reg2470,
                 reg2469,
                 forvar2468,
                 reg2467,
                 reg2466,
                 forvar2465,
                 reg2464,
                 reg2463,
                 reg2462,
                 forvar2461,
                 reg2460,
                 reg2459,
                 forvar2458,
                 reg2457,
                 reg2456,
                 reg2455,
                 reg2454,
                 forvar2453,
                 reg2452,
                 reg2451,
                 reg2450,
                 forvar2449,
                 forvar2448,
                 reg2447,
                 reg2446,
                 reg2445,
                 reg2444,
                 reg2443,
                 forvar2442,
                 reg2441,
                 reg2440,
                 reg2439,
                 reg2438,
                 reg2437,
                 forvar2436,
                 forvar2435,
                 reg2434,
                 reg2433,
                 reg2432,
                 reg2431,
                 reg2427,
                 forvar2426,
                 reg2430,
                 reg2429,
                 reg2428,
                 forvar2427,
                 reg2426,
                 reg2425,
                 reg2424,
                 reg2423,
                 reg2422,
                 reg2421,
                 forvar2420,
                 forvar2419,
                 forvar2418,
                 reg2417,
                 reg2409,
                 reg2407,
                 forvar2406,
                 reg2416,
                 reg2415,
                 reg2414,
                 reg2413,
                 reg2412,
                 reg2411,
                 reg2410,
                 forvar2409,
                 reg2408,
                 forvar2407,
                 reg2406,
                 reg2405,
                 reg2404,
                 reg2403,
                 reg2402,
                 forvar2401,
                 reg2400,
                 forvar2399,
                 reg2398,
                 reg2397,
                 forvar2396,
                 forvar2395,
                 forvar2394,
                 reg2393,
                 reg2392,
                 reg2391,
                 reg2390,
                 forvar2389,
                 reg2388,
                 reg2383,
                 forvar2381,
                 reg2387,
                 reg2386,
                 reg2385,
                 reg2384,
                 forvar2383,
                 reg2382,
                 reg2381,
                 forvar2380,
                 forvar2379,
                 wire2378,
                 wire2377,
                 wire2376,
                 wire2375,
                 (1'h0)};
  assign wire2375 = ((^$unsigned((^wire2373))) | ($unsigned((wire2373 <<< (8'hb3))) >= $signed({wire2372})));
  assign wire2376 = ((-($signed(wire2371) | wire2373[(3'h5):(1'h0)])) * (~&wire2373[(2'h2):(1'h1)]));
  assign wire2377 = $signed(wire2376[(2'h3):(1'h1)]);
  assign wire2378 = wire2376;
  always
    @(posedge clk) begin
      for (forvar2379 = (1'h0); (forvar2379 < (2'h3)); forvar2379 = (forvar2379 + (1'h1)))
        begin
          for (forvar2380 = (1'h0); (forvar2380 < (2'h2)); forvar2380 = (forvar2380 + (1'h1)))
            begin
              if ((forvar2380 | wire2378))
                begin
                  if (((wire2374 ? wire2374[(2'h2):(1'h0)] : wire2378) ?
                      wire2372[(3'h6):(2'h2)] : (($unsigned(wire2372) ?
                              $signed((8'ha4)) : (+wire2377)) ?
                          {(wire2372 < wire2378)} : ((!wire2375) | wire2374[(2'h2):(1'h0)]))))
                    begin
                      reg2381 <= wire2378[(2'h2):(1'h0)];
                      reg2382 <= ($unsigned((^~((8'ha7) ?
                          wire2372 : forvar2379))) + wire2371[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg2381 <= wire2375[(4'h8):(3'h5)];
                    end
                  for (forvar2383 = (1'h0); (forvar2383 < (2'h3)); forvar2383 = (forvar2383 + (1'h1)))
                    begin
                      reg2384 <= wire2372[(2'h3):(1'h1)];
                      reg2385 <= wire2375[(3'h4):(3'h4)];
                      reg2386 <= wire2374;
                      reg2387 <= {{reg2384}};
                    end
                end
              else
                begin
                  for (forvar2381 = (1'h0); (forvar2381 < (2'h2)); forvar2381 = (forvar2381 + (1'h1)))
                    begin
                      reg2382 <= (reg2385 << {wire2376});
                      reg2383 <= wire2378[(2'h2):(1'h1)];
                      reg2384 <= ((&$signed(wire2377[(1'h1):(1'h1)])) ?
                          $signed(wire2371[(2'h3):(2'h3)]) : forvar2381[(4'h9):(4'h8)]);
                      reg2385 <= $signed({$unsigned(wire2373)});
                    end
                  if ((((~&(~&reg2387)) ?
                      ($signed(wire2371) ~^ reg2385) : reg2387) || ((+{wire2374}) ?
                      $unsigned(forvar2381[(1'h0):(1'h0)]) : $signed(reg2385))))
                    begin
                      reg2386 <= $signed(forvar2379[(3'h4):(1'h0)]);
                      reg2387 <= {((^~(+forvar2381)) ?
                              {forvar2379} : (wire2371 ?
                                  forvar2380[(1'h0):(1'h0)] : (|(8'ha2))))};
                    end
                  else
                    begin
                      reg2386 <= reg2387;
                      reg2387 <= $unsigned(wire2376[(4'ha):(2'h2)]);
                      reg2388 <= $unsigned((~$signed($unsigned((8'hb0)))));
                    end
                  for (forvar2389 = (1'h0); (forvar2389 < (2'h3)); forvar2389 = (forvar2389 + (1'h1)))
                    begin
                      reg2390 <= forvar2389;
                      reg2391 <= $signed(reg2384[(1'h0):(1'h0)]);
                      reg2392 <= forvar2383[(3'h6):(3'h6)];
                      reg2393 <= $unsigned({({reg2392} ?
                              (forvar2389 || reg2392) : reg2392[(1'h1):(1'h1)])});
                    end
                end
            end
          for (forvar2394 = (1'h0); (forvar2394 < (1'h0)); forvar2394 = (forvar2394 + (1'h1)))
            begin
              for (forvar2395 = (1'h0); (forvar2395 < (2'h3)); forvar2395 = (forvar2395 + (1'h1)))
                begin
                  for (forvar2396 = (1'h0); (forvar2396 < (2'h2)); forvar2396 = (forvar2396 + (1'h1)))
                    begin
                      reg2397 <= ((8'h9e) >= $signed(forvar2381[(3'h7):(1'h0)]));
                      reg2398 <= (~^(~|reg2388[(2'h3):(1'h1)]));
                    end
                end
              for (forvar2399 = (1'h0); (forvar2399 < (1'h1)); forvar2399 = (forvar2399 + (1'h1)))
                begin
                  reg2400 <= $unsigned((^~{(reg2392 ? forvar2389 : wire2378)}));
                  for (forvar2401 = (1'h0); (forvar2401 < (1'h1)); forvar2401 = (forvar2401 + (1'h1)))
                    begin
                      reg2402 <= forvar2381[(2'h3):(1'h0)];
                      reg2403 <= $unsigned($signed($unsigned((^reg2388))));
                      reg2404 <= reg2387[(3'h5):(2'h2)];
                    end
                end
              if (reg2397)
                begin
                  if ((^~({reg2382} < (reg2388 >= (reg2387 ?
                      wire2373 : wire2378)))))
                    begin
                      reg2405 <= (forvar2379[(3'h4):(2'h3)] - (((8'ha2) * (forvar2381 ?
                          (8'ha8) : forvar2389)) ^ forvar2396));
                    end
                  else
                    begin
                      reg2405 <= $unsigned((reg2397[(2'h2):(2'h2)] ^~ forvar2394[(1'h0):(1'h0)]));
                      reg2406 <= (|(^{reg2404}));
                    end
                  for (forvar2407 = (1'h0); (forvar2407 < (2'h2)); forvar2407 = (forvar2407 + (1'h1)))
                    begin
                      reg2408 <= forvar2401[(3'h7):(3'h5)];
                    end
                  for (forvar2409 = (1'h0); (forvar2409 < (1'h1)); forvar2409 = (forvar2409 + (1'h1)))
                    begin
                      reg2410 <= (&(~&(^reg2385[(3'h5):(3'h4)])));
                      reg2411 <= (wire2373[(2'h3):(2'h2)] ?
                          $signed($signed((|reg2397))) : $signed({(wire2377 ?
                                  (8'hb9) : (8'ha8))}));
                      reg2412 <= reg2387;
                    end
                  if (wire2377[(2'h2):(1'h0)])
                    begin
                      reg2413 <= (~$unsigned(($unsigned(reg2405) - forvar2407)));
                      reg2414 <= ($unsigned(reg2388) ?
                          forvar2381[(2'h3):(2'h2)] : $unsigned($signed((reg2391 || reg2398))));
                      reg2415 <= reg2393;
                      reg2416 <= (($signed(reg2415) > {(-forvar2383)}) + ($unsigned($unsigned((8'ha1))) >= $signed($unsigned(forvar2389))));
                    end
                  else
                    begin
                      reg2413 <= (|reg2398);
                    end
                end
              else
                begin
                  reg2405 <= reg2402[(2'h2):(2'h2)];
                  for (forvar2406 = (1'h0); (forvar2406 < (2'h3)); forvar2406 = (forvar2406 + (1'h1)))
                    begin
                      reg2407 <= $unsigned({({(8'ha5)} - reg2405[(4'h9):(1'h0)])});
                      reg2408 <= ((~|$signed(reg2385[(3'h5):(1'h0)])) ?
                          (-(~&(~forvar2380))) : (~(((8'hb8) ?
                              reg2387 : wire2375) == (forvar2407 == reg2398))));
                      reg2409 <= wire2378[(3'h5):(3'h4)];
                      reg2410 <= {($unsigned((~&forvar2399)) ?
                              {(+forvar2380)} : $signed((-reg2398)))};
                    end
                  if ((reg2404[(4'hb):(4'h9)] > forvar2389))
                    begin
                      reg2411 <= {(^(~^(reg2408 ? reg2390 : reg2411)))};
                      reg2412 <= {$signed(($signed((8'hac)) > reg2416))};
                    end
                  else
                    begin
                      reg2411 <= {$signed({$unsigned(reg2405)})};
                      reg2412 <= $unsigned({(|reg2416)});
                      reg2413 <= (~&({(wire2378 ^~ reg2404)} >>> $signed(wire2376[(2'h2):(2'h2)])));
                      reg2414 <= reg2403;
                    end
                end
            end
        end
      reg2417 <= $signed(wire2375[(4'h8):(3'h7)]);
      for (forvar2418 = (1'h0); (forvar2418 < (2'h3)); forvar2418 = (forvar2418 + (1'h1)))
        begin
          for (forvar2419 = (1'h0); (forvar2419 < (2'h3)); forvar2419 = (forvar2419 + (1'h1)))
            begin
              for (forvar2420 = (1'h0); (forvar2420 < (2'h3)); forvar2420 = (forvar2420 + (1'h1)))
                begin
                  if (({((~&forvar2395) >>> forvar2407[(3'h6):(2'h3)])} ?
                      wire2374 : reg2409))
                    begin
                      reg2421 <= ($signed((8'h9f)) ?
                          reg2417 : $unsigned((forvar2395 ?
                              (8'hb7) : (reg2382 ? reg2404 : reg2388))));
                      reg2422 <= forvar2379;
                    end
                  else
                    begin
                      reg2421 <= reg2417[(1'h1):(1'h1)];
                      reg2422 <= (+wire2376[(2'h2):(1'h0)]);
                    end
                  if (((^reg2400) >>> reg2409))
                    begin
                      reg2423 <= $unsigned(reg2398);
                      reg2424 <= reg2414;
                      reg2425 <= forvar2381[(3'h7):(2'h2)];
                    end
                  else
                    begin
                      reg2423 <= ((~&$unsigned(forvar2409[(4'ha):(3'h6)])) ?
                          $unsigned({reg2410}) : reg2410);
                    end
                end
              if (($unsigned(({(8'haf)} || forvar2409)) <<< ($signed($signed(reg2416)) ^ $signed($signed(reg2388)))))
                begin
                  reg2426 <= ($signed(($signed(reg2403) ?
                          forvar2396[(4'h8):(3'h4)] : {reg2383})) ?
                      {$unsigned((~^reg2425))} : $signed(wire2374[(1'h0):(1'h0)]));
                  for (forvar2427 = (1'h0); (forvar2427 < (1'h1)); forvar2427 = (forvar2427 + (1'h1)))
                    begin
                      reg2428 <= $signed($signed($signed({forvar2395})));
                      reg2429 <= $unsigned($unsigned(((+reg2381) ?
                          (wire2374 ? forvar2407 : reg2416) : reg2388)));
                      reg2430 <= forvar2401[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar2426 = (1'h0); (forvar2426 < (1'h1)); forvar2426 = (forvar2426 + (1'h1)))
                    begin
                      reg2427 <= $signed($unsigned((8'h9f)));
                      reg2428 <= $unsigned((-{(reg2398 >>> forvar2419)}));
                      reg2429 <= (($unsigned($signed(forvar2383)) - reg2416[(4'ha):(4'h8)]) >> $unsigned($signed((8'ha3))));
                      reg2430 <= ($unsigned((|reg2381[(1'h1):(1'h0)])) ?
                          (^~(8'ha7)) : $signed(((reg2400 || reg2387) ?
                              reg2400 : (forvar2401 ? reg2408 : reg2421))));
                    end
                  reg2431 <= (+(reg2393 <<< (~|(^~reg2421))));
                  reg2432 <= reg2413[(4'hb):(3'h4)];
                  if ((|(~(+reg2382[(3'h5):(1'h0)]))))
                    begin
                      reg2433 <= $unsigned(($unsigned($signed(reg2429)) ?
                          $unsigned($unsigned((8'h9d))) : (&{reg2390})));
                    end
                  else
                    begin
                      reg2433 <= ((+wire2378[(4'h8):(3'h7)]) ?
                          forvar2407 : (($unsigned(reg2423) > (reg2405 >> reg2400)) ?
                              reg2381 : forvar2379));
                      reg2434 <= reg2406;
                    end
                end
              for (forvar2435 = (1'h0); (forvar2435 < (1'h1)); forvar2435 = (forvar2435 + (1'h1)))
                begin
                  for (forvar2436 = (1'h0); (forvar2436 < (2'h3)); forvar2436 = (forvar2436 + (1'h1)))
                    begin
                      reg2437 <= ($unsigned({{forvar2406}}) - $signed(reg2423));
                    end
                  if ($signed(reg2388[(1'h0):(1'h0)]))
                    begin
                      reg2438 <= $signed((-$unsigned($signed((8'hba)))));
                      reg2439 <= ($unsigned(reg2385) << $unsigned(reg2400[(3'h6):(3'h4)]));
                      reg2440 <= reg2417[(4'h9):(3'h7)];
                      reg2441 <= forvar2396[(4'h9):(3'h7)];
                    end
                  else
                    begin
                      reg2438 <= (wire2376[(3'h6):(3'h4)] || $signed($signed(((8'ha7) ?
                          reg2438 : forvar2395))));
                      reg2439 <= (&$unsigned($signed(reg2417[(3'h6):(1'h1)])));
                    end
                  for (forvar2442 = (1'h0); (forvar2442 < (2'h2)); forvar2442 = (forvar2442 + (1'h1)))
                    begin
                      reg2443 <= ((forvar2379 ?
                              ($unsigned(wire2375) ~^ $unsigned(forvar2379)) : $signed((-reg2416))) ?
                          ($signed($unsigned(reg2384)) && ({reg2433} ?
                              (~forvar2379) : (~&reg2400))) : (+((forvar2381 < reg2417) ?
                              $unsigned((8'hb8)) : $signed(reg2439))));
                      reg2444 <= (-(&$signed($unsigned((8'ha4)))));
                      reg2445 <= (wire2373 | {(&reg2443[(1'h0):(1'h0)])});
                      reg2446 <= reg2403;
                    end
                end
              reg2447 <= (|(-{(forvar2401 >>> reg2408)}));
            end
          for (forvar2448 = (1'h0); (forvar2448 < (1'h1)); forvar2448 = (forvar2448 + (1'h1)))
            begin
              for (forvar2449 = (1'h0); (forvar2449 < (2'h3)); forvar2449 = (forvar2449 + (1'h1)))
                begin
                  if ((8'hb4))
                    begin
                      reg2450 <= {forvar2407};
                    end
                  else
                    begin
                      reg2450 <= $unsigned((((reg2411 ^ reg2386) || {(8'ha2)}) + ((^~reg2447) * (reg2447 * forvar2448))));
                      reg2451 <= $unsigned(($unsigned({forvar2418}) ?
                          ((8'hb5) * reg2403) : $unsigned(((8'haa) ?
                              (8'ha1) : forvar2380))));
                      reg2452 <= $signed({(|$signed(forvar2380))});
                    end
                end
            end
          if (reg2383)
            begin
              if ($signed({$signed((wire2372 & (8'ha0)))}))
                begin
                  for (forvar2453 = (1'h0); (forvar2453 < (2'h3)); forvar2453 = (forvar2453 + (1'h1)))
                    begin
                      reg2454 <= $unsigned($signed(forvar2419));
                      reg2455 <= ((^~((reg2430 ? forvar2406 : reg2425) ?
                              (reg2416 ?
                                  forvar2448 : forvar2427) : (|reg2454))) ?
                          (wire2375[(3'h5):(2'h2)] == (~reg2417)) : $unsigned($unsigned(reg2422)));
                      reg2456 <= $signed(reg2455);
                      reg2457 <= (!reg2451[(2'h3):(2'h2)]);
                    end
                end
              else
                begin
                  for (forvar2453 = (1'h0); (forvar2453 < (1'h0)); forvar2453 = (forvar2453 + (1'h1)))
                    begin
                      reg2454 <= forvar2436[(1'h0):(1'h0)];
                      reg2455 <= $signed(reg2457);
                      reg2456 <= $signed(($unsigned($signed(forvar2442)) ?
                          reg2434[(4'hb):(3'h5)] : $unsigned($unsigned(reg2456))));
                      reg2457 <= {(reg2457[(4'h8):(1'h0)] ?
                              forvar2399[(4'he):(2'h2)] : $unsigned((reg2440 ?
                                  forvar2419 : reg2386)))};
                    end
                  for (forvar2458 = (1'h0); (forvar2458 < (2'h2)); forvar2458 = (forvar2458 + (1'h1)))
                    begin
                      reg2459 <= (($unsigned(((8'ha5) <= reg2398)) >>> $unsigned($unsigned((8'ha3)))) ?
                          $unsigned({reg2457[(4'h8):(3'h6)]}) : $unsigned(((~(8'ha2)) ?
                              forvar2453 : (reg2426 ? forvar2396 : (8'had)))));
                      reg2460 <= (|((^wire2375[(4'h8):(2'h3)]) ?
                          ((8'ha2) << (forvar2436 ?
                              reg2447 : reg2424)) : (forvar2419 < ((8'ha9) ?
                              reg2409 : (8'ha9)))));
                    end
                end
              for (forvar2461 = (1'h0); (forvar2461 < (2'h3)); forvar2461 = (forvar2461 + (1'h1)))
                begin
                  if ($signed((reg2414 + {{reg2417}})))
                    begin
                      reg2462 <= ($signed(reg2427[(3'h6):(3'h4)]) ?
                          $unsigned((forvar2458[(1'h1):(1'h0)] | (reg2404 ?
                              (8'hb1) : forvar2426))) : $unsigned((&{forvar2436})));
                      reg2463 <= wire2373[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg2462 <= forvar2395[(1'h0):(1'h0)];
                      reg2463 <= (+reg2452);
                      reg2464 <= (+reg2423);
                    end
                  for (forvar2465 = (1'h0); (forvar2465 < (2'h2)); forvar2465 = (forvar2465 + (1'h1)))
                    begin
                      reg2466 <= (~|(reg2384 <= (!((8'hab) >= reg2410))));
                      reg2467 <= $signed($signed($unsigned($unsigned(reg2400))));
                    end
                end
              if ((({{(8'hb9)}} > ($signed(reg2416) ?
                      reg2467 : forvar2419[(4'h9):(1'h1)])) ?
                  $unsigned(forvar2449) : ({reg2392[(4'h9):(1'h0)]} | $unsigned($signed(reg2402)))))
                begin
                  for (forvar2468 = (1'h0); (forvar2468 < (2'h3)); forvar2468 = (forvar2468 + (1'h1)))
                    begin
                      reg2469 <= (+(8'ha3));
                      reg2470 <= (^$signed(((forvar2409 ~^ reg2450) && (~reg2431))));
                    end
                end
              else
                begin
                  for (forvar2468 = (1'h0); (forvar2468 < (2'h3)); forvar2468 = (forvar2468 + (1'h1)))
                    begin
                      reg2469 <= $signed((((reg2445 ~^ reg2410) ?
                          {reg2462} : forvar2426[(1'h0):(1'h0)]) || forvar2380));
                      reg2470 <= reg2414;
                      reg2471 <= reg2459;
                      reg2472 <= (+((forvar2442[(1'h1):(1'h1)] | (reg2454 || reg2383)) ?
                          (forvar2442 > {(8'hb7)}) : wire2372[(2'h3):(1'h1)]));
                    end
                  for (forvar2473 = (1'h0); (forvar2473 < (1'h1)); forvar2473 = (forvar2473 + (1'h1)))
                    begin
                      reg2474 <= reg2416;
                      reg2475 <= (&(+forvar2465[(2'h2):(1'h1)]));
                      reg2476 <= ((8'hb3) ? reg2404 : reg2425);
                      reg2477 <= (~|$signed((~(8'hb9))));
                    end
                end
              if (((8'ha6) ? reg2386 : ((~&reg2411) && reg2470[(1'h0):(1'h0)])))
                begin
                  for (forvar2478 = (1'h0); (forvar2478 < (2'h3)); forvar2478 = (forvar2478 + (1'h1)))
                    begin
                      reg2479 <= $signed($signed((reg2466 > reg2405)));
                      reg2480 <= ({$unsigned($unsigned(reg2426))} <<< forvar2383);
                    end
                  if (reg2467[(4'h9):(2'h3)])
                    begin
                      reg2481 <= ($unsigned($unsigned((-reg2427))) - (($unsigned(reg2455) ?
                              $unsigned(forvar2394) : (-reg2390)) ?
                          ((~^reg2392) ?
                              (reg2439 ?
                                  reg2445 : reg2409) : (8'h9d)) : ($signed(forvar2409) << $signed(reg2407))));
                      reg2482 <= reg2439[(2'h2):(1'h0)];
                      reg2483 <= (((reg2422 < {(8'ha8)}) ?
                              $signed({reg2402}) : reg2477[(3'h4):(3'h4)]) ?
                          (forvar2426[(2'h2):(2'h2)] ?
                              $signed((reg2428 < forvar2449)) : ($signed((8'hb5)) ?
                                  $signed(reg2451) : reg2430[(1'h1):(1'h0)])) : $signed((~^(^~reg2382))));
                    end
                  else
                    begin
                      reg2481 <= (((-$unsigned(reg2417)) != (~wire2372[(3'h6):(3'h6)])) && ($unsigned($signed(forvar2420)) ?
                          reg2480[(1'h0):(1'h0)] : ($signed(reg2426) && (reg2425 != (8'hae)))));
                      reg2482 <= reg2482[(2'h3):(1'h1)];
                      reg2483 <= ($unsigned((reg2457[(4'h9):(2'h3)] | $signed(forvar2468))) <<< ((~(reg2474 ?
                          forvar2418 : reg2402)) || (reg2383[(4'hc):(4'h8)] && $unsigned(reg2398))));
                      reg2484 <= $signed($signed(((^~reg2443) ?
                          reg2471 : (8'hab))));
                    end
                  reg2485 <= (reg2484[(3'h5):(3'h5)] ~^ (reg2426 ?
                      $signed((-forvar2399)) : $signed(reg2463)));
                end
              else
                begin
                  for (forvar2478 = (1'h0); (forvar2478 < (1'h0)); forvar2478 = (forvar2478 + (1'h1)))
                    begin
                      reg2479 <= $unsigned(reg2471);
                    end
                  if ((^~$signed((reg2469[(1'h1):(1'h0)] ^ (reg2451 * reg2392)))))
                    begin
                      reg2480 <= $signed(reg2445[(2'h2):(1'h0)]);
                      reg2481 <= (~{(!$unsigned(reg2407))});
                      reg2482 <= $unsigned(reg2424);
                      reg2483 <= (reg2427[(3'h5):(2'h2)] ?
                          (!forvar2394[(2'h3):(1'h1)]) : $signed($unsigned(forvar2380)));
                    end
                  else
                    begin
                      reg2480 <= (((reg2417 ?
                              {reg2463} : reg2485[(3'h4):(1'h0)]) + $signed($unsigned(reg2417))) ?
                          (~reg2476[(1'h0):(1'h0)]) : {(forvar2478[(4'h8):(3'h6)] ?
                                  ((8'hb5) - reg2406) : ((8'hb4) & reg2460))});
                      reg2481 <= (({$unsigned(forvar2458)} ?
                              forvar2399[(2'h2):(2'h2)] : $signed(wire2375)) ?
                          (+$signed((reg2441 >> reg2440))) : ($signed((!reg2415)) ?
                              ($signed(reg2444) < wire2372) : ($signed(reg2416) != (reg2443 ?
                                  reg2412 : (8'ha2)))));
                    end
                end
            end
          else
            begin
              for (forvar2453 = (1'h0); (forvar2453 < (1'h1)); forvar2453 = (forvar2453 + (1'h1)))
                begin
                  if ($signed($signed(wire2374[(2'h2):(1'h1)])))
                    begin
                      reg2454 <= reg2439;
                    end
                  else
                    begin
                      reg2454 <= (^reg2407[(4'hd):(3'h4)]);
                      reg2455 <= $signed(({{forvar2465}} + (!$signed(reg2433))));
                      reg2456 <= $unsigned(reg2410);
                      reg2457 <= ((reg2424[(4'h8):(4'h8)] ?
                              $signed(forvar2461[(4'hb):(1'h1)]) : $signed(reg2472)) ?
                          (!reg2400) : (!reg2441[(3'h4):(2'h3)]));
                    end
                  if ((reg2437 ?
                      $unsigned(($unsigned((8'h9d)) && reg2437)) : (((8'hab) << $unsigned(reg2431)) ?
                          reg2480 : $unsigned(reg2481[(2'h3):(1'h1)]))))
                    begin
                      reg2458 <= $unsigned(reg2384);
                      reg2459 <= (&((^forvar2461[(4'h9):(3'h6)]) << ((reg2456 * reg2392) ?
                          reg2384[(1'h1):(1'h1)] : $signed(reg2432))));
                    end
                  else
                    begin
                      reg2458 <= $signed(reg2450[(4'hc):(2'h3)]);
                    end
                  if (forvar2379)
                    begin
                      reg2460 <= forvar2458;
                    end
                  else
                    begin
                      reg2460 <= reg2398[(3'h5):(1'h0)];
                    end
                end
              for (forvar2461 = (1'h0); (forvar2461 < (1'h0)); forvar2461 = (forvar2461 + (1'h1)))
                begin
                  if (reg2427)
                    begin
                      reg2462 <= (&reg2406[(1'h1):(1'h1)]);
                      reg2463 <= $unsigned($unsigned((~(reg2440 & reg2382))));
                    end
                  else
                    begin
                      reg2462 <= reg2471;
                    end
                  if ((~^forvar2427[(4'h8):(3'h6)]))
                    begin
                      reg2464 <= reg2403[(4'hb):(3'h4)];
                      reg2465 <= ($signed(($signed(reg2426) | $unsigned(reg2429))) ?
                          $unsigned(($signed(wire2378) ?
                              forvar2478[(4'hf):(4'hf)] : forvar2419[(3'h5):(3'h5)])) : reg2391[(1'h0):(1'h0)]);
                      reg2466 <= wire2376[(4'hf):(4'hf)];
                      reg2467 <= (~|((reg2479 == wire2375) ?
                          reg2425[(2'h2):(1'h1)] : ($unsigned((8'ha0)) ?
                              $signed(reg2407) : (reg2447 >>> reg2440))));
                    end
                  else
                    begin
                      reg2464 <= (($signed(reg2438[(3'h6):(2'h2)]) >> $unsigned((reg2444 >= (8'haa)))) <<< (~&(((8'ha1) & reg2469) ?
                          (reg2417 ?
                              reg2383 : reg2407) : (forvar2409 ^~ forvar2395))));
                      reg2465 <= (((~&forvar2383[(2'h3):(2'h2)]) == ($unsigned(reg2413) ?
                          reg2405 : {(8'hab)})) << (~^({(8'h9c)} == (forvar2473 != forvar2381))));
                      reg2466 <= $signed(reg2414);
                    end
                  reg2468 <= forvar2418[(1'h1):(1'h1)];
                  for (forvar2469 = (1'h0); (forvar2469 < (2'h3)); forvar2469 = (forvar2469 + (1'h1)))
                    begin
                      reg2470 <= (~&($unsigned({reg2390}) >>> ((~^reg2433) ?
                          $signed(reg2467) : $signed(reg2468))));
                      reg2471 <= $unsigned(($signed((-reg2444)) < {(reg2438 >>> reg2417)}));
                      reg2472 <= $signed(({reg2437[(2'h2):(1'h1)]} || $signed({reg2415})));
                      reg2473 <= $unsigned($unsigned(((&reg2445) ~^ reg2427)));
                    end
                end
              reg2474 <= reg2462[(2'h2):(1'h0)];
              for (forvar2475 = (1'h0); (forvar2475 < (1'h0)); forvar2475 = (forvar2475 + (1'h1)))
                begin
                  for (forvar2476 = (1'h0); (forvar2476 < (2'h2)); forvar2476 = (forvar2476 + (1'h1)))
                    begin
                      reg2477 <= (~|$signed((&forvar2406)));
                      reg2478 <= (((+reg2450) ^~ (reg2477 ?
                              $signed(reg2408) : $signed(forvar2394))) ?
                          ($signed(reg2444[(4'hb):(4'hb)]) ?
                              (+(reg2482 - reg2425)) : (wire2375[(3'h6):(3'h4)] ?
                                  $signed(reg2467) : $unsigned(reg2476))) : $signed(forvar2476));
                      reg2479 <= reg2446;
                    end
                  if ((wire2377[(2'h3):(1'h0)] << ((~|forvar2380) ?
                      (!(^reg2480)) : {((8'ha2) ? reg2428 : forvar2401)})))
                    begin
                      reg2480 <= $unsigned($unsigned((wire2372[(2'h3):(1'h0)] ?
                          (^~reg2423) : (~^reg2483))));
                      reg2481 <= ((|({reg2464} >>> reg2410[(3'h7):(3'h4)])) ?
                          $unsigned((((8'haa) ^ reg2454) ^ $signed(reg2426))) : $unsigned((~|$signed(reg2465))));
                    end
                  else
                    begin
                      reg2480 <= $signed((~|(reg2451 ?
                          (reg2440 ? reg2387 : reg2434) : $unsigned(reg2479))));
                    end
                  if (({(reg2455 << {forvar2442})} ?
                      reg2432 : $unsigned($unsigned((reg2400 | (8'hb9))))))
                    begin
                      reg2482 <= ({$signed($signed(reg2481))} ?
                          ($signed((&reg2403)) != (reg2407 ?
                              $signed(reg2468) : (8'ha9))) : (^~$unsigned(reg2383[(1'h0):(1'h0)])));
                      reg2483 <= (|{(|reg2450[(3'h7):(3'h7)])});
                      reg2484 <= ($unsigned(((^forvar2420) ?
                              reg2404[(4'ha):(4'h9)] : $signed(wire2373))) ?
                          $unsigned($signed((reg2484 | (8'haa)))) : $signed(($unsigned(reg2478) ?
                              (reg2423 ?
                                  forvar2478 : reg2427) : $signed(reg2441))));
                      reg2485 <= $signed($unsigned((-$signed(reg2421))));
                    end
                  else
                    begin
                      reg2482 <= (^~reg2444[(4'ha):(1'h1)]);
                    end
                  for (forvar2486 = (1'h0); (forvar2486 < (2'h3)); forvar2486 = (forvar2486 + (1'h1)))
                    begin
                      reg2487 <= reg2422;
                    end
                end
            end
          for (forvar2488 = (1'h0); (forvar2488 < (2'h3)); forvar2488 = (forvar2488 + (1'h1)))
            begin
              if ($unsigned((8'h9f)))
                begin
                  if (((~&(reg2480[(2'h3):(1'h1)] > $unsigned(reg2469))) < $unsigned($unsigned((reg2424 ?
                      reg2383 : reg2383)))))
                    begin
                      reg2489 <= (&$unsigned($signed($signed((8'hb2)))));
                      reg2490 <= ((8'hb0) >> (forvar2469 ?
                          reg2447 : {reg2409[(4'h8):(3'h4)]}));
                      reg2491 <= $signed({(-(forvar2406 == (8'hb4)))});
                      reg2492 <= (forvar2427 & (((~|forvar2469) ?
                          wire2373[(2'h3):(1'h1)] : $signed(forvar2469)) >> (8'ha8)));
                    end
                  else
                    begin
                      reg2489 <= $unsigned((forvar2435[(3'h6):(1'h1)] >>> $signed(reg2386[(2'h3):(1'h0)])));
                      reg2490 <= $unsigned(forvar2406);
                      reg2491 <= (-reg2454[(4'hb):(2'h2)]);
                    end
                end
              else
                begin
                  for (forvar2489 = (1'h0); (forvar2489 < (1'h0)); forvar2489 = (forvar2489 + (1'h1)))
                    begin
                      reg2490 <= $unsigned(($unsigned(forvar2436) ?
                          ((~^reg2447) ?
                              $signed(forvar2449) : $unsigned(reg2402)) : (forvar2399 | (8'ha5))));
                    end
                end
              if ((|forvar2380))
                begin
                  for (forvar2493 = (1'h0); (forvar2493 < (2'h3)); forvar2493 = (forvar2493 + (1'h1)))
                    begin
                      reg2494 <= (^reg2390);
                    end
                end
              else
                begin
                  if (($unsigned(({reg2412} <= $signed(forvar2419))) ?
                      {$unsigned($signed(reg2422))} : $unsigned(reg2414)))
                    begin
                      reg2493 <= (~&reg2472[(3'h5):(3'h5)]);
                      reg2494 <= {{(-(reg2457 ^~ forvar2468))}};
                      reg2495 <= $unsigned((~|{(~&(8'hb1))}));
                    end
                  else
                    begin
                      reg2493 <= ((^~$signed($signed(reg2468))) <<< ((reg2443 ?
                          (8'hb0) : $unsigned(reg2429)) < ($signed(forvar2396) ?
                          forvar2420[(3'h4):(2'h2)] : (reg2455 ?
                              wire2373 : forvar2473))));
                      reg2494 <= (&reg2397);
                      reg2495 <= $signed((^forvar2458));
                      reg2496 <= $signed((~&$unsigned((~|forvar2394))));
                    end
                  for (forvar2497 = (1'h0); (forvar2497 < (2'h3)); forvar2497 = (forvar2497 + (1'h1)))
                    begin
                      reg2498 <= reg2456;
                      reg2499 <= (({(forvar2380 ?
                                  reg2425 : reg2424)} && {(reg2438 <= reg2416)}) ?
                          ((&reg2416) <= (^forvar2468[(3'h7):(2'h2)])) : $signed(reg2473[(1'h0):(1'h0)]));
                      reg2500 <= reg2495;
                    end
                  if ((($signed((forvar2453 ? forvar2426 : reg2388)) ?
                          forvar2488 : $signed((reg2384 <= (8'hac)))) ?
                      $unsigned($signed($unsigned(reg2450))) : (|$unsigned(reg2455[(4'hc):(4'h9)]))))
                    begin
                      reg2501 <= (($signed($signed(reg2450)) ?
                          forvar2427 : reg2432[(4'hb):(2'h2)]) < (-$unsigned((~|reg2416))));
                      reg2502 <= reg2384[(3'h7):(3'h6)];
                      reg2503 <= (~$signed($signed(reg2494[(3'h6):(1'h0)])));
                    end
                  else
                    begin
                      reg2501 <= reg2457[(4'h9):(4'h9)];
                      reg2502 <= $unsigned(reg2474[(1'h1):(1'h0)]);
                      reg2503 <= forvar2465;
                    end
                  for (forvar2504 = (1'h0); (forvar2504 < (1'h0)); forvar2504 = (forvar2504 + (1'h1)))
                    begin
                      reg2505 <= reg2426[(2'h2):(2'h2)];
                    end
                end
              for (forvar2506 = (1'h0); (forvar2506 < (1'h1)); forvar2506 = (forvar2506 + (1'h1)))
                begin
                  if ((!((8'ha1) < (^~$unsigned(reg2432)))))
                    begin
                      reg2507 <= forvar2488;
                      reg2508 <= {reg2455};
                      reg2509 <= reg2400;
                      reg2510 <= forvar2448;
                    end
                  else
                    begin
                      reg2507 <= $unsigned($unsigned(reg2414));
                      reg2508 <= ((~$signed($signed(reg2452))) ~^ (((&forvar2420) ?
                              $signed(reg2487) : (forvar2465 ?
                                  reg2447 : forvar2448)) ?
                          $signed((reg2464 ?
                              (8'ha3) : reg2388)) : $signed(reg2421)));
                      reg2509 <= reg2407;
                    end
                end
            end
        end
    end
  assign wire2511 = reg2385[(3'h4):(2'h2)];
  assign wire2512 = $unsigned(reg2479[(3'h6):(2'h2)]);
  assign wire2513 = reg2489[(1'h1):(1'h1)];
  assign wire2514 = $signed(reg2428[(3'h7):(1'h0)]);
  always
    @(posedge clk) begin
      if ((~^(|wire2511)))
        begin
          if ($unsigned((reg2471 ?
              ($unsigned((8'ha6)) - (reg2485 - (8'hab))) : ((forvar2396 ?
                  reg2414 : reg2439) - $unsigned(forvar2395)))))
            begin
              for (forvar2515 = (1'h0); (forvar2515 < (2'h2)); forvar2515 = (forvar2515 + (1'h1)))
                begin
                  if ($signed($signed(reg2393)))
                    begin
                      reg2516 <= $signed(((8'h9d) ?
                          (^~(reg2503 ?
                              reg2428 : wire2373)) : {$signed((8'hba))}));
                      reg2517 <= forvar2395[(2'h3):(1'h1)];
                      reg2518 <= ({(^reg2422)} | ($unsigned((~^reg2482)) > reg2481));
                      reg2519 <= $signed(reg2405);
                    end
                  else
                    begin
                      reg2516 <= {($signed($signed(reg2446)) ?
                              ($signed(reg2444) >>> (8'h9d)) : reg2468)};
                      reg2517 <= $unsigned((&{reg2495}));
                    end
                  if (($signed($signed(reg2479[(3'h5):(1'h0)])) ?
                      forvar2383[(2'h3):(1'h0)] : $unsigned(reg2407)))
                    begin
                      reg2520 <= ({reg2510} != {$signed((reg2400 ?
                              reg2510 : reg2423))});
                      reg2521 <= $unsigned((reg2481 ?
                          (forvar2488[(3'h6):(3'h5)] * forvar2396[(4'hb):(3'h6)]) : (reg2439 ^ (~^reg2516))));
                      reg2522 <= reg2478;
                      reg2523 <= $signed({((forvar2406 ?
                              reg2425 : (8'hb0)) >= $unsigned((8'ha7)))});
                    end
                  else
                    begin
                      reg2520 <= ({{reg2471[(2'h3):(2'h3)]}} == $signed($unsigned(((8'ha4) <<< reg2390))));
                    end
                end
              for (forvar2524 = (1'h0); (forvar2524 < (1'h0)); forvar2524 = (forvar2524 + (1'h1)))
                begin
                  for (forvar2525 = (1'h0); (forvar2525 < (2'h2)); forvar2525 = (forvar2525 + (1'h1)))
                    begin
                      reg2526 <= (($unsigned(reg2479) ?
                              reg2517 : $signed((reg2516 ?
                                  reg2492 : (8'hac)))) ?
                          reg2479 : $signed((~|{wire2511})));
                    end
                  for (forvar2527 = (1'h0); (forvar2527 < (1'h1)); forvar2527 = (forvar2527 + (1'h1)))
                    begin
                      reg2528 <= {$unsigned(forvar2493)};
                    end
                end
              for (forvar2529 = (1'h0); (forvar2529 < (2'h2)); forvar2529 = (forvar2529 + (1'h1)))
                begin
                  if ((8'hab))
                    begin
                      reg2530 <= ((({reg2455} ?
                              (reg2431 ?
                                  forvar2461 : reg2422) : $signed(reg2482)) ?
                          reg2480 : reg2390) | $signed(forvar2486));
                      reg2531 <= (reg2430[(3'h5):(2'h2)] ^~ reg2443);
                      reg2532 <= (~&reg2522);
                      reg2533 <= reg2384;
                    end
                  else
                    begin
                      reg2530 <= (({$signed(forvar2506)} ?
                              $signed($unsigned(forvar2458)) : $signed($signed(forvar2381))) ?
                          {$signed($signed(reg2528))} : forvar2396);
                      reg2531 <= forvar2383[(2'h2):(2'h2)];
                      reg2532 <= reg2528[(2'h3):(1'h0)];
                      reg2533 <= $unsigned($unsigned(forvar2469[(2'h3):(2'h3)]));
                    end
                end
              if ({forvar2475[(2'h3):(2'h3)]})
                begin
                  for (forvar2534 = (1'h0); (forvar2534 < (1'h0)); forvar2534 = (forvar2534 + (1'h1)))
                    begin
                      reg2535 <= (~|(!reg2489[(2'h2):(1'h1)]));
                    end
                  for (forvar2536 = (1'h0); (forvar2536 < (1'h0)); forvar2536 = (forvar2536 + (1'h1)))
                    begin
                      reg2537 <= ((~&reg2487) ?
                          (|((reg2402 ?
                              (8'hb2) : reg2408) || $signed(reg2455))) : $signed(reg2460[(4'hd):(2'h3)]));
                      reg2538 <= $signed(($unsigned(reg2516[(1'h1):(1'h1)]) <<< $unsigned(forvar2383)));
                    end
                end
              else
                begin
                  for (forvar2534 = (1'h0); (forvar2534 < (2'h3)); forvar2534 = (forvar2534 + (1'h1)))
                    begin
                      reg2535 <= ((reg2535 ?
                          $signed(forvar2395) : $signed($unsigned(reg2430))) < {wire2375});
                      reg2536 <= ((-(8'ha6)) ?
                          (~&forvar2453[(2'h3):(2'h2)]) : ((+$unsigned(forvar2389)) ?
                              forvar2399[(2'h3):(1'h0)] : reg2440[(1'h0):(1'h0)]));
                    end
                  for (forvar2537 = (1'h0); (forvar2537 < (2'h2)); forvar2537 = (forvar2537 + (1'h1)))
                    begin
                      reg2538 <= $unsigned(reg2505);
                      reg2539 <= $unsigned((wire2511 ?
                          (^(^reg2470)) : {$signed(reg2537)}));
                      reg2540 <= $unsigned((((reg2465 & reg2400) > forvar2476) ?
                          $unsigned((reg2400 < reg2406)) : ($unsigned(wire2376) * reg2508)));
                      reg2541 <= (((reg2441 != ((8'haf) ? wire2375 : reg2463)) ?
                              $signed((+reg2473)) : reg2410[(1'h0):(1'h0)]) ?
                          (reg2536[(1'h0):(1'h0)] ^~ $unsigned($signed((8'hae)))) : reg2423);
                    end
                  if ($unsigned($unsigned($signed((reg2467 | reg2434)))))
                    begin
                      reg2542 <= $unsigned((-(8'hab)));
                      reg2543 <= $unsigned(reg2495[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg2542 <= $signed(($unsigned($signed(reg2493)) ?
                          (-$signed(reg2456)) : $signed(forvar2465[(3'h6):(2'h3)])));
                    end
                end
            end
          else
            begin
              for (forvar2515 = (1'h0); (forvar2515 < (1'h0)); forvar2515 = (forvar2515 + (1'h1)))
                begin
                  for (forvar2516 = (1'h0); (forvar2516 < (2'h2)); forvar2516 = (forvar2516 + (1'h1)))
                    begin
                      reg2517 <= (((reg2466 ? (-reg2481) : (~^reg2501)) ?
                              $unsigned($signed(reg2406)) : reg2430) ?
                          forvar2504[(4'h9):(3'h6)] : $signed($unsigned((reg2478 ?
                              reg2412 : (8'had)))));
                    end
                  reg2518 <= {$signed({$signed(reg2387)})};
                  reg2519 <= reg2473;
                  reg2520 <= $signed({wire2376});
                end
            end
        end
      else
        begin
          for (forvar2515 = (1'h0); (forvar2515 < (2'h3)); forvar2515 = (forvar2515 + (1'h1)))
            begin
              for (forvar2516 = (1'h0); (forvar2516 < (2'h2)); forvar2516 = (forvar2516 + (1'h1)))
                begin
                  reg2517 <= (((reg2414 ?
                          reg2505 : $unsigned(wire2511)) ^~ reg2464[(3'h4):(2'h2)]) ?
                      ($signed(reg2432[(1'h1):(1'h1)]) ?
                          reg2501[(2'h3):(2'h3)] : $unsigned((&forvar2448))) : (&(~((8'ha4) == reg2490))));
                end
              if ((~&$signed((^~$signed(reg2441)))))
                begin
                  if ($unsigned(reg2450[(1'h0):(1'h0)]))
                    begin
                      reg2518 <= (!$signed(((forvar2515 ?
                              forvar2469 : reg2477) ?
                          (wire2514 ? forvar2486 : reg2475) : forvar2420)));
                      reg2519 <= (+$signed(reg2454));
                      reg2520 <= $unsigned((reg2538[(1'h1):(1'h0)] > ($unsigned((8'h9e)) < $signed(reg2411))));
                    end
                  else
                    begin
                      reg2518 <= ($signed((reg2498 * $signed(reg2402))) ?
                          $signed(({(8'h9c)} ?
                              (wire2511 <= reg2535) : $signed(reg2404))) : (&{{forvar2418}}));
                      reg2519 <= reg2520[(2'h2):(1'h1)];
                      reg2520 <= reg2500[(2'h3):(2'h2)];
                    end
                  if ($unsigned($signed((~|$unsigned(reg2501)))))
                    begin
                      reg2521 <= reg2428;
                      reg2522 <= reg2479[(2'h2):(1'h1)];
                      reg2523 <= (forvar2506 ?
                          ((-reg2472[(4'ha):(3'h5)]) ?
                              (~&(reg2421 ?
                                  (8'hae) : reg2423)) : ($signed(forvar2536) ^~ (forvar2516 ^ (8'ha2)))) : (((|(8'hb2)) ?
                              forvar2448[(1'h1):(1'h1)] : (~&reg2475)) & ({wire2376} == reg2479)));
                      reg2524 <= (((8'hb7) ?
                          $unsigned($unsigned(reg2463)) : $unsigned(reg2444)) >> ({(-wire2511)} | ((forvar2516 + reg2517) & (reg2516 ?
                          (8'hb8) : forvar2442))));
                    end
                  else
                    begin
                      reg2521 <= forvar2435;
                      reg2522 <= (reg2533 ?
                          ((reg2412[(3'h6):(3'h4)] * reg2383) ?
                              (reg2483 ?
                                  (reg2443 ?
                                      reg2428 : reg2441) : $unsigned(reg2520)) : reg2493[(4'h8):(1'h0)]) : $signed(forvar2536[(2'h2):(2'h2)]));
                    end
                  reg2525 <= {((reg2431[(4'he):(4'h9)] ?
                              (^reg2500) : (reg2492 ^ reg2492)) ?
                          {(reg2487 ~^ reg2417)} : reg2458[(1'h0):(1'h0)])};
                  if (reg2427)
                    begin
                      reg2526 <= $signed({$unsigned(reg2482)});
                      reg2527 <= $unsigned($unsigned((+$unsigned((8'hb3)))));
                      reg2528 <= ({{reg2501[(1'h0):(1'h0)]}} ?
                          $signed(($signed(reg2479) ?
                              (reg2423 ~^ reg2405) : reg2444)) : $signed($unsigned(wire2375[(4'ha):(1'h1)])));
                      reg2529 <= (^~forvar2383);
                    end
                  else
                    begin
                      reg2526 <= forvar2401;
                      reg2527 <= ($unsigned(reg2491[(4'h9):(3'h4)]) ?
                          (^~($signed(reg2477) ?
                              reg2490[(3'h5):(3'h4)] : $signed(reg2457))) : $unsigned(reg2482[(2'h2):(1'h1)]));
                    end
                end
              else
                begin
                  for (forvar2518 = (1'h0); (forvar2518 < (1'h0)); forvar2518 = (forvar2518 + (1'h1)))
                    begin
                      reg2519 <= ((|forvar2409[(1'h1):(1'h1)]) - (((reg2412 ?
                          forvar2458 : forvar2489) && reg2439[(2'h2):(2'h2)]) + wire2372[(3'h4):(3'h4)]));
                      reg2520 <= (reg2464 ?
                          $unsigned((-$unsigned(forvar2486))) : $unsigned({(-reg2530)}));
                    end
                  for (forvar2521 = (1'h0); (forvar2521 < (2'h2)); forvar2521 = (forvar2521 + (1'h1)))
                    begin
                      reg2522 <= forvar2458[(2'h3):(2'h2)];
                      reg2523 <= (^~(8'ha9));
                    end
                end
            end
        end
      if ($signed($unsigned($signed((8'ha2)))))
        begin
          for (forvar2544 = (1'h0); (forvar2544 < (2'h3)); forvar2544 = (forvar2544 + (1'h1)))
            begin
              for (forvar2545 = (1'h0); (forvar2545 < (2'h3)); forvar2545 = (forvar2545 + (1'h1)))
                begin
                  if ($signed({($signed(reg2434) >= $unsigned(reg2465))}))
                    begin
                      reg2546 <= ({forvar2475} > ((&forvar2401) ?
                          {reg2510} : (reg2509 ? (!reg2430) : {forvar2435})));
                      reg2547 <= $signed(forvar2389);
                      reg2548 <= $unsigned($signed(wire2514));
                    end
                  else
                    begin
                      reg2546 <= $signed(reg2498[(2'h2):(1'h0)]);
                      reg2547 <= $unsigned((~(((8'hb2) ?
                          reg2387 : reg2502) ^ {reg2384})));
                      reg2548 <= ((reg2384[(4'ha):(2'h2)] >>> {(^reg2425)}) >= ($unsigned(forvar2476[(3'h4):(1'h1)]) ?
                          (8'hb2) : (((8'ha8) ?
                              (8'hb2) : reg2411) || $unsigned(wire2376))));
                    end
                  if ($signed(forvar2401[(1'h1):(1'h1)]))
                    begin
                      reg2549 <= $signed($signed({((8'haa) << forvar2518)}));
                      reg2550 <= (reg2445 ?
                          ($unsigned((8'ha7)) ?
                              ((~&reg2546) ?
                                  $signed(forvar2383) : $signed((8'ha0))) : $unsigned({reg2492})) : $signed($unsigned(((8'ha7) ^~ (8'h9f)))));
                    end
                  else
                    begin
                      reg2549 <= $signed((&(&$unsigned(reg2450))));
                      reg2550 <= forvar2381[(3'h6):(3'h6)];
                      reg2551 <= (forvar2537 ?
                          $signed((~|(forvar2527 ?
                              reg2466 : forvar2524))) : (reg2547[(1'h1):(1'h0)] ?
                              $unsigned((reg2539 ?
                                  forvar2419 : (8'hb6))) : ({reg2447} >= reg2429[(1'h0):(1'h0)])));
                    end
                  reg2552 <= (({{reg2451}} ~^ {(~&reg2537)}) ?
                      forvar2545 : forvar2468);
                  for (forvar2553 = (1'h0); (forvar2553 < (2'h3)); forvar2553 = (forvar2553 + (1'h1)))
                    begin
                      reg2554 <= $signed((reg2456 > ($unsigned(forvar2469) ?
                          (reg2425 || reg2477) : {(8'hb7)})));
                      reg2555 <= $signed((~|(reg2421[(2'h2):(2'h2)] ?
                          forvar2399[(3'h4):(2'h2)] : (forvar2448 ?
                              reg2551 : forvar2399))));
                    end
                end
              reg2556 <= reg2493;
              if (($unsigned($signed((|reg2400))) ?
                  (!(reg2516[(3'h4):(2'h2)] | $unsigned(reg2454))) : reg2393[(3'h5):(1'h1)]))
                begin
                  reg2557 <= (~reg2454[(2'h3):(2'h3)]);
                  for (forvar2558 = (1'h0); (forvar2558 < (2'h3)); forvar2558 = (forvar2558 + (1'h1)))
                    begin
                      reg2559 <= forvar2426[(2'h2):(2'h2)];
                      reg2560 <= $signed((-reg2424));
                      reg2561 <= ((^~(forvar2529[(4'ha):(2'h3)] ?
                          (~reg2460) : reg2403)) >= $signed((|(forvar2465 >>> reg2402))));
                      reg2562 <= $unsigned((8'ha5));
                    end
                  reg2563 <= $signed(((~&reg2526) ?
                      reg2423 : reg2466[(3'h5):(1'h0)]));
                  for (forvar2564 = (1'h0); (forvar2564 < (2'h2)); forvar2564 = (forvar2564 + (1'h1)))
                    begin
                      reg2565 <= (^((^~$signed(forvar2553)) > {forvar2506[(4'hb):(4'hb)]}));
                      reg2566 <= reg2483;
                    end
                end
              else
                begin
                  for (forvar2557 = (1'h0); (forvar2557 < (2'h2)); forvar2557 = (forvar2557 + (1'h1)))
                    begin
                      reg2558 <= (+forvar2515);
                      reg2559 <= (^((8'hb4) ?
                          reg2404[(4'hc):(1'h1)] : $signed($signed((8'ha7)))));
                      reg2560 <= reg2563[(2'h2):(2'h2)];
                    end
                  for (forvar2561 = (1'h0); (forvar2561 < (1'h0)); forvar2561 = (forvar2561 + (1'h1)))
                    begin
                      reg2562 <= ({((reg2387 ? (8'ha7) : reg2500) ?
                              reg2537[(1'h0):(1'h0)] : {(8'ha7)})} <= (&reg2492[(3'h6):(2'h3)]));
                      reg2563 <= ({$unsigned($signed(wire2376))} - reg2549);
                      reg2564 <= reg2542;
                      reg2565 <= ((8'hac) ?
                          (~&((forvar2453 > reg2566) * reg2547[(1'h1):(1'h1)])) : forvar2383[(2'h2):(1'h1)]);
                    end
                  if ((reg2423 * $unsigned($signed({forvar2478}))))
                    begin
                      reg2566 <= forvar2518;
                      reg2567 <= $signed({$unsigned((~&(8'hac)))});
                      reg2568 <= ({$unsigned($signed(reg2527))} > ($signed($unsigned(reg2452)) <= (|(reg2528 - reg2391))));
                      reg2569 <= (~^{$unsigned(forvar2406[(2'h3):(1'h1)])});
                    end
                  else
                    begin
                      reg2566 <= {wire2375[(4'h8):(3'h6)]};
                      reg2567 <= $unsigned(($signed($signed(forvar2381)) == ($signed(reg2421) ^ wire2375)));
                    end
                  if (reg2429[(2'h3):(2'h2)])
                    begin
                      reg2570 <= (8'h9c);
                      reg2571 <= $signed(reg2471);
                    end
                  else
                    begin
                      reg2570 <= (8'hb3);
                      reg2571 <= reg2558[(2'h3):(1'h1)];
                      reg2572 <= (~&reg2546);
                    end
                end
              if ({$signed({reg2480})})
                begin
                  if ((8'hb1))
                    begin
                      reg2573 <= (&((^~$signed(reg2450)) ?
                          $unsigned($signed(forvar2515)) : (^~(forvar2545 ?
                              reg2547 : reg2391))));
                      reg2574 <= reg2471;
                      reg2575 <= (($unsigned((8'ha8)) ~^ ((reg2400 ?
                              reg2574 : forvar2515) ?
                          (reg2384 == forvar2557) : (forvar2504 <= forvar2537))) > $unsigned({(reg2552 ?
                              reg2405 : (8'haa))}));
                    end
                  else
                    begin
                      reg2573 <= ($unsigned($unsigned($signed(forvar2518))) ?
                          $signed($unsigned(reg2446)) : forvar2524);
                      reg2574 <= $unsigned($signed((reg2429 ?
                          $unsigned(reg2571) : reg2484[(3'h6):(2'h2)])));
                      reg2575 <= {$unsigned((~(reg2558 ? reg2526 : reg2567)))};
                      reg2576 <= (-(reg2403 ?
                          reg2494[(1'h1):(1'h0)] : $signed($unsigned(forvar2465))));
                    end
                  for (forvar2577 = (1'h0); (forvar2577 < (1'h1)); forvar2577 = (forvar2577 + (1'h1)))
                    begin
                      reg2578 <= ($signed($unsigned((~&reg2441))) ?
                          reg2498[(1'h0):(1'h0)] : {{(~&wire2511)}});
                      reg2579 <= ({(reg2384[(4'h8):(2'h3)] <= $signed(reg2519))} ?
                          {{{reg2438}}} : ($signed(((8'hb5) ^ (8'hab))) ~^ ($unsigned(reg2484) || (reg2500 ?
                              reg2439 : reg2402))));
                      reg2580 <= {(^(~^(|wire2375)))};
                      reg2581 <= $signed(reg2496[(3'h6):(3'h5)]);
                    end
                end
              else
                begin
                  reg2573 <= {(|forvar2476[(3'h5):(2'h2)])};
                end
            end
          reg2582 <= {(^(forvar2418[(3'h4):(1'h0)] ^ reg2546))};
          for (forvar2583 = (1'h0); (forvar2583 < (1'h0)); forvar2583 = (forvar2583 + (1'h1)))
            begin
              if (({(forvar2488[(2'h3):(2'h3)] + $unsigned(reg2525))} ?
                  forvar2461 : $unsigned((forvar2486[(3'h6):(1'h1)] * (reg2452 != (8'hb3))))))
                begin
                  reg2584 <= $unsigned(reg2566[(1'h1):(1'h0)]);
                end
              else
                begin
                  for (forvar2584 = (1'h0); (forvar2584 < (1'h0)); forvar2584 = (forvar2584 + (1'h1)))
                    begin
                      reg2585 <= $unsigned($signed(reg2387[(3'h7):(1'h0)]));
                    end
                  for (forvar2586 = (1'h0); (forvar2586 < (1'h1)); forvar2586 = (forvar2586 + (1'h1)))
                    begin
                      reg2587 <= $signed(reg2499);
                      reg2588 <= ($unsigned($unsigned((reg2521 ?
                          reg2552 : (8'ha8)))) << $unsigned(reg2582));
                    end
                  for (forvar2589 = (1'h0); (forvar2589 < (2'h2)); forvar2589 = (forvar2589 + (1'h1)))
                    begin
                      reg2590 <= reg2518[(1'h0):(1'h0)];
                      reg2591 <= $unsigned(forvar2583[(4'h9):(2'h3)]);
                    end
                  reg2592 <= reg2398;
                end
              if ($signed($signed(forvar2489[(3'h4):(1'h1)])))
                begin
                  for (forvar2593 = (1'h0); (forvar2593 < (2'h3)); forvar2593 = (forvar2593 + (1'h1)))
                    begin
                      reg2594 <= (($signed(((8'hba) || reg2474)) ?
                              forvar2473 : reg2384[(1'h0):(1'h0)]) ?
                          ($signed(reg2410) >= {(reg2415 ?
                                  reg2590 : reg2381)}) : reg2540[(2'h2):(1'h1)]);
                      reg2595 <= (^~$signed(((+reg2525) ?
                          (!forvar2593) : $signed((8'haf)))));
                      reg2596 <= reg2524;
                    end
                  for (forvar2597 = (1'h0); (forvar2597 < (1'h1)); forvar2597 = (forvar2597 + (1'h1)))
                    begin
                      reg2598 <= ($signed(reg2446) ?
                          $unsigned((^reg2464)) : reg2381);
                      reg2599 <= (reg2425 ? $unsigned(reg2433) : reg2433);
                    end
                end
              else
                begin
                  if ($signed($signed($unsigned((reg2548 >= reg2558)))))
                    begin
                      reg2593 <= $signed(($unsigned((reg2575 - reg2574)) ?
                          $unsigned((^(8'hb5))) : $unsigned((reg2569 ?
                              (8'ha7) : forvar2448))));
                      reg2594 <= reg2423[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2593 <= $signed((((forvar2478 ? reg2538 : reg2492) ?
                          $unsigned(reg2578) : (reg2584 ?
                              forvar2534 : (8'ha4))) != ((!forvar2506) ?
                          (~(8'ha8)) : (reg2414 && forvar2435))));
                    end
                  if ({($signed(reg2524) ?
                          ((+reg2405) >= {reg2443}) : {(^~reg2382)})})
                    begin
                      reg2595 <= ((8'h9d) ?
                          reg2520[(4'hc):(3'h5)] : $unsigned($unsigned(reg2571)));
                      reg2596 <= (8'haf);
                      reg2597 <= (($unsigned({reg2539}) ?
                              forvar2521[(1'h0):(1'h0)] : $unsigned($signed(reg2525))) ?
                          $unsigned($unsigned((reg2384 - (8'hb7)))) : $signed(({forvar2518} != (forvar2536 * reg2531))));
                    end
                  else
                    begin
                      reg2595 <= {((|reg2591) * $unsigned(reg2388))};
                    end
                  for (forvar2598 = (1'h0); (forvar2598 < (1'h1)); forvar2598 = (forvar2598 + (1'h1)))
                    begin
                      reg2599 <= (&reg2585);
                    end
                end
            end
          if (((~&((&wire2512) ? reg2454[(4'ha):(3'h5)] : $signed(reg2422))) ?
              (8'hb3) : reg2518[(2'h3):(1'h0)]))
            begin
              for (forvar2600 = (1'h0); (forvar2600 < (2'h3)); forvar2600 = (forvar2600 + (1'h1)))
                begin
                  for (forvar2601 = (1'h0); (forvar2601 < (1'h0)); forvar2601 = (forvar2601 + (1'h1)))
                    begin
                      reg2602 <= forvar2564;
                      reg2603 <= $unsigned(($signed((^reg2414)) < ((^~(8'hb1)) ?
                          (reg2587 <<< forvar2600) : (reg2538 ?
                              reg2590 : reg2566))));
                      reg2604 <= reg2550;
                      reg2605 <= ((8'hac) <<< ($signed($unsigned(reg2404)) || reg2466[(4'h9):(3'h6)]));
                    end
                  for (forvar2606 = (1'h0); (forvar2606 < (1'h1)); forvar2606 = (forvar2606 + (1'h1)))
                    begin
                      reg2607 <= reg2587;
                      reg2608 <= $unsigned(reg2471);
                      reg2609 <= {((forvar2395[(3'h5):(3'h4)] ?
                                  {reg2602} : reg2475[(1'h0):(1'h0)]) ?
                              forvar2407 : (!(&reg2527)))};
                    end
                end
              reg2610 <= {$signed(reg2402)};
              if (reg2410[(3'h6):(2'h2)])
                begin
                  reg2611 <= (~|$signed($signed(forvar2449)));
                  if ($unsigned((((&reg2548) && $signed((8'ha3))) & forvar2420[(1'h0):(1'h0)])))
                    begin
                      reg2612 <= ($unsigned($unsigned((reg2481 ?
                          reg2549 : (8'ha1)))) >= reg2489[(1'h0):(1'h0)]);
                      reg2613 <= ((~|$signed((^~forvar2395))) ^ {{reg2445[(3'h5):(1'h1)]}});
                      reg2614 <= ((~&(|$unsigned(reg2467))) ?
                          $signed(forvar2564) : (reg2430[(1'h1):(1'h1)] ?
                              $signed((reg2492 ?
                                  forvar2396 : reg2575)) : ($signed(reg2446) ?
                                  (reg2499 ?
                                      forvar2586 : (8'ha5)) : $unsigned(reg2520))));
                    end
                  else
                    begin
                      reg2612 <= reg2492[(2'h2):(1'h0)];
                      reg2613 <= reg2447[(1'h0):(1'h0)];
                      reg2614 <= $signed($unsigned(reg2499[(4'hc):(3'h7)]));
                    end
                  reg2615 <= forvar2577;
                  for (forvar2616 = (1'h0); (forvar2616 < (2'h3)); forvar2616 = (forvar2616 + (1'h1)))
                    begin
                      reg2617 <= ($signed($unsigned($unsigned(reg2403))) || wire2377[(3'h7):(3'h6)]);
                      reg2618 <= (forvar2593[(3'h6):(2'h3)] ?
                          $signed({(|(8'ha0))}) : reg2500);
                      reg2619 <= $unsigned($signed($signed(reg2560[(2'h2):(2'h2)])));
                      reg2620 <= $unsigned($unsigned($signed((~&reg2416))));
                    end
                end
              else
                begin
                  reg2611 <= $signed(reg2593);
                  for (forvar2612 = (1'h0); (forvar2612 < (1'h0)); forvar2612 = (forvar2612 + (1'h1)))
                    begin
                      reg2613 <= $unsigned(reg2525[(4'ha):(3'h4)]);
                    end
                end
              for (forvar2621 = (1'h0); (forvar2621 < (2'h3)); forvar2621 = (forvar2621 + (1'h1)))
                begin
                  for (forvar2622 = (1'h0); (forvar2622 < (1'h1)); forvar2622 = (forvar2622 + (1'h1)))
                    begin
                      reg2623 <= reg2459[(3'h5):(2'h3)];
                    end
                  if ({(~|(8'ha2))})
                    begin
                      reg2624 <= $unsigned((&wire2372));
                      reg2625 <= reg2565[(4'hf):(4'hc)];
                      reg2626 <= forvar2468;
                    end
                  else
                    begin
                      reg2624 <= ((|forvar2497[(1'h1):(1'h1)]) ?
                          $unsigned(($unsigned(reg2452) < {(8'had)})) : (~^$unsigned(reg2456)));
                    end
                end
            end
          else
            begin
              reg2600 <= reg2575[(3'h5):(1'h0)];
              if ({reg2415[(3'h5):(3'h5)]})
                begin
                  reg2601 <= (|$unsigned({forvar2394}));
                  if ((!((^{forvar2527}) ? {(~reg2457)} : {reg2441})))
                    begin
                      reg2602 <= reg2522;
                      reg2603 <= forvar2379[(2'h3):(1'h0)];
                      reg2604 <= (&(~|($unsigned(forvar2506) >> $signed(reg2498))));
                      reg2605 <= $unsigned($signed((^~$unsigned(forvar2468))));
                    end
                  else
                    begin
                      reg2602 <= reg2392[(1'h1):(1'h1)];
                      reg2603 <= $unsigned((&$signed($signed(forvar2515))));
                    end
                end
              else
                begin
                  for (forvar2601 = (1'h0); (forvar2601 < (2'h2)); forvar2601 = (forvar2601 + (1'h1)))
                    begin
                      reg2602 <= ($unsigned((~&(reg2626 & reg2463))) >= $unsigned(($unsigned(reg2580) >= $signed(reg2421))));
                      reg2603 <= (~&($unsigned($signed(reg2403)) > reg2561[(3'h5):(3'h5)]));
                      reg2604 <= wire2371[(1'h0):(1'h0)];
                    end
                end
              if ((reg2476 ?
                  forvar2475[(2'h3):(1'h0)] : (((8'h9f) <= (^~reg2455)) ?
                      $signed((~^reg2592)) : $unsigned(reg2542))))
                begin
                  for (forvar2606 = (1'h0); (forvar2606 < (1'h1)); forvar2606 = (forvar2606 + (1'h1)))
                    begin
                      reg2607 <= $unsigned($signed(reg2391));
                    end
                  for (forvar2608 = (1'h0); (forvar2608 < (2'h2)); forvar2608 = (forvar2608 + (1'h1)))
                    begin
                      reg2609 <= $signed((reg2556 | reg2452[(2'h3):(2'h3)]));
                      reg2610 <= reg2423[(4'ha):(3'h7)];
                    end
                end
              else
                begin
                  if ((8'ha0))
                    begin
                      reg2606 <= {((reg2425 <<< (-reg2584)) ?
                              ((~^(8'hb6)) != forvar2409[(3'h7):(1'h0)]) : reg2387[(4'h9):(1'h0)])};
                      reg2607 <= (8'ha4);
                      reg2608 <= (^~(((forvar2489 >>> reg2610) ?
                          (!reg2525) : reg2609) >> forvar2427[(3'h4):(3'h4)]));
                      reg2609 <= {{$signed((~&reg2452))}};
                    end
                  else
                    begin
                      reg2606 <= $signed(((reg2517[(2'h2):(1'h1)] & $unsigned(reg2510)) + {(reg2525 <<< reg2584)}));
                      reg2607 <= $signed(reg2430[(1'h1):(1'h1)]);
                      reg2608 <= (reg2564 ?
                          reg2537[(3'h5):(1'h0)] : ((8'haa) ^ reg2444[(4'hd):(1'h1)]));
                      reg2609 <= (8'hb5);
                    end
                end
              if ((~^reg2517[(2'h3):(1'h1)]))
                begin
                  for (forvar2611 = (1'h0); (forvar2611 < (2'h3)); forvar2611 = (forvar2611 + (1'h1)))
                    begin
                      reg2612 <= reg2468[(2'h3):(2'h2)];
                      reg2613 <= reg2462;
                    end
                  if ((8'hb8))
                    begin
                      reg2614 <= ({((forvar2436 ? (8'ha2) : forvar2557) ?
                                  reg2530[(3'h4):(2'h2)] : (reg2552 ?
                                      reg2428 : reg2507))} ?
                          $signed(reg2494[(3'h5):(1'h1)]) : $unsigned($signed($signed(reg2540))));
                      reg2615 <= $signed(({$signed(forvar2598)} == reg2572));
                      reg2616 <= {$unsigned(reg2563[(1'h1):(1'h0)])};
                    end
                  else
                    begin
                      reg2614 <= (8'ha4);
                      reg2615 <= reg2559[(2'h3):(1'h0)];
                      reg2616 <= ((~$unsigned({wire2375})) ?
                          forvar2442[(1'h1):(1'h1)] : $unsigned(((forvar2458 << forvar2486) - {wire2373})));
                      reg2617 <= forvar2593;
                    end
                  for (forvar2618 = (1'h0); (forvar2618 < (2'h2)); forvar2618 = (forvar2618 + (1'h1)))
                    begin
                      reg2619 <= ({(-$signed(reg2557))} ~^ {{reg2527}});
                    end
                end
              else
                begin
                  reg2611 <= (reg2605[(3'h5):(2'h2)] | $signed((8'haf)));
                  for (forvar2612 = (1'h0); (forvar2612 < (1'h1)); forvar2612 = (forvar2612 + (1'h1)))
                    begin
                      reg2613 <= (8'hb5);
                    end
                end
            end
        end
      else
        begin
          if (forvar2524[(3'h4):(2'h3)])
            begin
              reg2544 <= $signed((~^(reg2536[(1'h1):(1'h0)] == (forvar2406 ?
                  (8'haa) : (8'hb8)))));
              for (forvar2545 = (1'h0); (forvar2545 < (1'h1)); forvar2545 = (forvar2545 + (1'h1)))
                begin
                  for (forvar2546 = (1'h0); (forvar2546 < (2'h2)); forvar2546 = (forvar2546 + (1'h1)))
                    begin
                      reg2547 <= $signed((~|(reg2596[(3'h6):(3'h6)] <<< (reg2408 >>> forvar2488))));
                      reg2548 <= ((((reg2426 >>> forvar2420) ~^ (-reg2615)) ?
                          (^$unsigned(forvar2583)) : $unsigned(reg2530[(1'h1):(1'h1)])) >= ($unsigned($unsigned(forvar2561)) == (|(reg2403 ?
                          reg2540 : reg2503))));
                      reg2549 <= ($unsigned($unsigned($signed((8'ha3)))) ?
                          forvar2396[(3'h5):(3'h4)] : $unsigned((~|(&(8'hac)))));
                      reg2550 <= (&reg2406[(2'h3):(1'h1)]);
                    end
                  reg2551 <= $unsigned({forvar2478[(4'hc):(3'h6)]});
                  for (forvar2552 = (1'h0); (forvar2552 < (2'h2)); forvar2552 = (forvar2552 + (1'h1)))
                    begin
                      reg2553 <= (({reg2617} >> reg2528[(4'he):(4'h8)]) ?
                          reg2479[(3'h6):(2'h2)] : $unsigned({(reg2385 ?
                                  forvar2544 : forvar2621)}));
                      reg2554 <= {(~&reg2598[(2'h3):(2'h3)])};
                      reg2555 <= (+(~$unsigned((reg2519 ? reg2539 : reg2438))));
                    end
                end
              for (forvar2556 = (1'h0); (forvar2556 < (2'h2)); forvar2556 = (forvar2556 + (1'h1)))
                begin
                  for (forvar2557 = (1'h0); (forvar2557 < (1'h0)); forvar2557 = (forvar2557 + (1'h1)))
                    begin
                      reg2558 <= $unsigned(($unsigned(((8'h9d) ?
                              (8'ha7) : reg2539)) ?
                          wire2375 : (8'ha3)));
                    end
                  for (forvar2559 = (1'h0); (forvar2559 < (1'h1)); forvar2559 = (forvar2559 + (1'h1)))
                    begin
                      reg2560 <= ((8'h9e) * forvar2598);
                      reg2561 <= $unsigned((($unsigned((8'h9e)) << {reg2596}) ?
                          $signed((reg2447 | forvar2606)) : ($unsigned(forvar2486) >>> (~|(8'haa)))));
                    end
                end
            end
          else
            begin
              for (forvar2544 = (1'h0); (forvar2544 < (1'h0)); forvar2544 = (forvar2544 + (1'h1)))
                begin
                  for (forvar2545 = (1'h0); (forvar2545 < (2'h3)); forvar2545 = (forvar2545 + (1'h1)))
                    begin
                      reg2546 <= $unsigned((8'ha8));
                      reg2547 <= reg2533[(2'h2):(1'h1)];
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2627 = (1'h0); (forvar2627 < (1'h1)); forvar2627 = (forvar2627 + (1'h1)))
        begin
          for (forvar2628 = (1'h0); (forvar2628 < (1'h1)); forvar2628 = (forvar2628 + (1'h1)))
            begin
              for (forvar2629 = (1'h0); (forvar2629 < (2'h2)); forvar2629 = (forvar2629 + (1'h1)))
                begin
                  reg2630 <= (+(($unsigned(reg2470) > (&reg2614)) - $unsigned((reg2593 >>> reg2468))));
                  if ($unsigned(reg2548))
                    begin
                      reg2631 <= $signed({$signed((reg2585 ?
                              reg2604 : (8'ha6)))});
                      reg2632 <= ((({reg2421} ?
                              reg2524[(1'h1):(1'h1)] : (~^reg2592)) ?
                          ((forvar2383 ? forvar2593 : reg2539) ~^ (reg2446 ?
                              reg2487 : forvar2553)) : (^(reg2605 ?
                              forvar2468 : reg2530))) >>> (!$unsigned($signed(reg2432))));
                    end
                  else
                    begin
                      reg2631 <= $unsigned((((~reg2608) & (forvar2559 <<< (8'ha5))) ~^ (~|$signed(reg2556))));
                      reg2632 <= ($unsigned(((reg2482 ^~ reg2434) ?
                              $unsigned((8'haf)) : {forvar2418})) ?
                          ($unsigned((reg2409 | wire2374)) ~^ (reg2602 ~^ $signed(reg2456))) : reg2624);
                      reg2633 <= ($signed((8'had)) ^ $unsigned((!((8'ha4) ?
                          reg2456 : forvar2601))));
                      reg2634 <= reg2611;
                    end
                  if ($signed(($unsigned($signed(reg2519)) && $unsigned(reg2383))))
                    begin
                      reg2635 <= reg2501[(3'h7):(2'h2)];
                      reg2636 <= $signed((~^(-(reg2470 ? reg2541 : reg2501))));
                      reg2637 <= reg2571[(4'h8):(3'h6)];
                      reg2638 <= $signed((({forvar2493} ?
                              reg2547[(3'h4):(3'h4)] : forvar2380) ?
                          reg2406[(1'h1):(1'h1)] : forvar2409));
                    end
                  else
                    begin
                      reg2635 <= $unsigned(reg2634);
                      reg2636 <= (reg2430[(1'h1):(1'h1)] ^~ $unsigned($signed((reg2631 ?
                          reg2444 : (8'ha9)))));
                      reg2637 <= $signed((~^forvar2486));
                    end
                end
              if ($unsigned({$unsigned((forvar2516 ? (8'ha4) : reg2439))}))
                begin
                  reg2639 <= forvar2622;
                end
              else
                begin
                  for (forvar2639 = (1'h0); (forvar2639 < (1'h0)); forvar2639 = (forvar2639 + (1'h1)))
                    begin
                      reg2640 <= (((^(reg2600 + reg2433)) ?
                              (-{reg2575}) : (~$signed(reg2434))) ?
                          (~((reg2585 <= reg2434) - (reg2412 ?
                              reg2639 : reg2566))) : (reg2536 >> {((8'hb5) ?
                                  (8'hab) : (8'ha1))}));
                      reg2641 <= reg2559[(1'h1):(1'h1)];
                      reg2642 <= $unsigned(($unsigned((reg2492 ?
                              reg2479 : reg2600)) ?
                          $unsigned((reg2398 ?
                              reg2444 : (8'hb4))) : forvar2584[(1'h1):(1'h1)]));
                    end
                  for (forvar2643 = (1'h0); (forvar2643 < (2'h3)); forvar2643 = (forvar2643 + (1'h1)))
                    begin
                      reg2644 <= {($signed((^(8'h9e))) ?
                              $signed((~&reg2482)) : ((forvar2473 << forvar2583) > reg2625[(4'hf):(4'he)]))};
                      reg2645 <= ($unsigned($unsigned((reg2587 ?
                              reg2625 : reg2570))) ?
                          ((reg2413[(3'h7):(2'h2)] && $unsigned(forvar2527)) ?
                              ((|reg2562) >= {reg2571}) : (forvar2622 <<< $unsigned(forvar2552))) : {$signed($signed(reg2603))});
                      reg2646 <= (!reg2519[(4'h8):(1'h0)]);
                    end
                  if (reg2386)
                    begin
                      reg2647 <= $signed((~^($signed((8'hb0)) > (forvar2468 ^ forvar2556))));
                      reg2648 <= reg2510[(4'ha):(1'h0)];
                    end
                  else
                    begin
                      reg2647 <= (+(~(reg2519 << $unsigned(forvar2586))));
                      reg2648 <= (~&reg2417);
                      reg2649 <= ((reg2445[(2'h3):(1'h1)] ?
                          (forvar2559 ?
                              (forvar2524 | reg2439) : (forvar2488 - reg2572)) : ($signed(forvar2616) ?
                              (8'hb5) : {reg2426})) <= {$signed((~&reg2537))});
                      reg2650 <= ((((~^reg2522) ? reg2468 : forvar2401) ?
                              {$signed(reg2427)} : ((reg2458 | reg2561) >= $unsigned(reg2466))) ?
                          forvar2561 : $signed($unsigned((reg2597 <<< reg2463))));
                    end
                end
              if ((+({(reg2602 ? reg2447 : reg2633)} ?
                  reg2476 : (~|$unsigned(reg2531)))))
                begin
                  for (forvar2651 = (1'h0); (forvar2651 < (1'h0)); forvar2651 = (forvar2651 + (1'h1)))
                    begin
                      reg2652 <= $unsigned({$signed($unsigned(forvar2409))});
                    end
                end
              else
                begin
                  if ($unsigned($signed(({reg2650} >>> (reg2617 ?
                      reg2444 : reg2631)))))
                    begin
                      reg2651 <= forvar2497[(2'h3):(2'h2)];
                      reg2652 <= (~|(((&reg2592) ?
                              (~reg2385) : ((8'ha2) > reg2400)) ?
                          $signed((&reg2496)) : {forvar2589[(2'h3):(2'h3)]}));
                    end
                  else
                    begin
                      reg2651 <= $unsigned(($signed({(8'hab)}) <= $signed((forvar2559 >>> wire2376))));
                      reg2652 <= reg2459[(1'h0):(1'h0)];
                      reg2653 <= {(|($unsigned((8'ha0)) <<< reg2590))};
                      reg2654 <= $signed((~|$unsigned({(8'ha4)})));
                    end
                end
            end
          for (forvar2655 = (1'h0); (forvar2655 < (2'h2)); forvar2655 = (forvar2655 + (1'h1)))
            begin
              for (forvar2656 = (1'h0); (forvar2656 < (1'h1)); forvar2656 = (forvar2656 + (1'h1)))
                begin
                  if ((~|$unsigned(reg2516)))
                    begin
                      reg2657 <= forvar2651[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2657 <= reg2470;
                      reg2658 <= $unsigned($signed({((8'hb5) ?
                              reg2484 : (8'hb5))}));
                      reg2659 <= (reg2631[(5'h10):(4'hd)] != reg2519);
                    end
                  if ({(8'hba)})
                    begin
                      reg2660 <= ((^~$unsigned(reg2619)) >>> $signed((reg2550[(1'h0):(1'h0)] && (reg2547 | reg2456))));
                    end
                  else
                    begin
                      reg2660 <= $signed(reg2426);
                    end
                end
              for (forvar2661 = (1'h0); (forvar2661 < (2'h3)); forvar2661 = (forvar2661 + (1'h1)))
                begin
                  reg2662 <= (forvar2473[(2'h2):(1'h1)] ?
                      $unsigned(reg2554) : ($unsigned((reg2529 ?
                          reg2565 : (8'ha7))) > ((8'hb7) >>> $signed(reg2552))));
                  if ($signed((reg2565 >>> $signed(reg2406[(1'h1):(1'h0)]))))
                    begin
                      reg2663 <= (reg2433[(2'h2):(1'h0)] + forvar2468);
                      reg2664 <= reg2604;
                      reg2665 <= ({(reg2381[(1'h0):(1'h0)] && (^~forvar2486))} ?
                          (((forvar2598 || forvar2584) ~^ $unsigned(reg2508)) ?
                              $signed((reg2590 ?
                                  forvar2606 : reg2647)) : $signed(reg2523)) : forvar2612);
                    end
                  else
                    begin
                      reg2663 <= wire2378;
                    end
                  for (forvar2666 = (1'h0); (forvar2666 < (1'h0)); forvar2666 = (forvar2666 + (1'h1)))
                    begin
                      reg2667 <= $signed((!($unsigned(forvar2401) ?
                          {forvar2442} : (reg2427 != reg2647))));
                      reg2668 <= (8'ha4);
                      reg2669 <= forvar2583[(3'h5):(3'h4)];
                      reg2670 <= ({(reg2480 ?
                              (forvar2493 ?
                                  reg2409 : reg2503) : $unsigned(reg2543))} && ($signed(forvar2427) ?
                          (-reg2570[(2'h2):(1'h0)]) : $unsigned((forvar2558 ?
                              reg2477 : forvar2449))));
                    end
                end
            end
        end
      if ((8'ha1))
        begin
          if (reg2576)
            begin
              reg2671 <= reg2630;
            end
          else
            begin
              for (forvar2671 = (1'h0); (forvar2671 < (1'h1)); forvar2671 = (forvar2671 + (1'h1)))
                begin
                  for (forvar2672 = (1'h0); (forvar2672 < (1'h1)); forvar2672 = (forvar2672 + (1'h1)))
                    begin
                      reg2673 <= (^reg2402);
                    end
                end
              if (forvar2448)
                begin
                  for (forvar2674 = (1'h0); (forvar2674 < (2'h2)); forvar2674 = (forvar2674 + (1'h1)))
                    begin
                      reg2675 <= ($unsigned(wire2513[(2'h2):(2'h2)]) ^~ reg2402);
                      reg2676 <= $unsigned($signed((reg2528[(2'h2):(2'h2)] ^~ reg2555)));
                    end
                  for (forvar2677 = (1'h0); (forvar2677 < (2'h3)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= $unsigned({reg2503});
                      reg2679 <= forvar2593;
                      reg2680 <= (^($signed(wire2374[(2'h2):(1'h1)]) ?
                          reg2562 : $unsigned(reg2595)));
                      reg2681 <= ((!$unsigned(((8'h9f) ? reg2503 : (8'hb5)))) ?
                          {((reg2633 != (8'hb8)) ?
                                  (&reg2547) : (8'hb8))} : ($signed((reg2590 ?
                              reg2463 : reg2521)) > $unsigned($unsigned(reg2619))));
                    end
                end
              else
                begin
                  reg2674 <= (forvar2606 ~^ $signed($signed(reg2493)));
                  if ($unsigned(($unsigned((forvar2407 ?
                      reg2642 : reg2495)) && $signed(((8'ha8) ?
                      reg2555 : reg2579)))))
                    begin
                      reg2675 <= ($signed((-forvar2627[(3'h7):(1'h1)])) ?
                          (|((reg2445 ?
                              reg2678 : reg2598) - (reg2422 >>> reg2566))) : reg2505);
                      reg2676 <= ((($signed(reg2669) ?
                              (reg2605 ? reg2572 : reg2598) : ((8'h9f) ?
                                  forvar2409 : reg2437)) < (8'ha0)) ?
                          {reg2558} : (reg2484 ?
                              {forvar2473} : $signed(reg2569[(1'h1):(1'h1)])));
                      reg2677 <= reg2423[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2675 <= (!(8'hae));
                      reg2676 <= $unsigned(reg2480[(2'h2):(1'h1)]);
                    end
                  for (forvar2678 = (1'h0); (forvar2678 < (2'h2)); forvar2678 = (forvar2678 + (1'h1)))
                    begin
                      reg2679 <= $unsigned($unsigned(reg2554));
                      reg2680 <= {(forvar2465[(1'h1):(1'h0)] - $signed({reg2408}))};
                      reg2681 <= $signed($unsigned(reg2398));
                      reg2682 <= $unsigned($signed($unsigned((8'hb6))));
                    end
                  for (forvar2683 = (1'h0); (forvar2683 < (1'h0)); forvar2683 = (forvar2683 + (1'h1)))
                    begin
                      reg2684 <= {reg2439[(1'h1):(1'h1)]};
                      reg2685 <= forvar2383[(1'h0):(1'h0)];
                      reg2686 <= {$signed($unsigned(forvar2473))};
                      reg2687 <= (((^(reg2468 ? (8'hab) : (8'ha2))) ?
                          (~|$unsigned(forvar2672)) : $unsigned($unsigned(reg2625))) == {$signed($unsigned(reg2560))});
                    end
                end
            end
          if (((reg2483 ?
                  (8'ha7) : $unsigned((reg2564 ? reg2613 : forvar2427))) ?
              reg2477 : {forvar2478}))
            begin
              if (forvar2537)
                begin
                  if ($unsigned(reg2633))
                    begin
                      reg2688 <= (8'ha6);
                      reg2689 <= {reg2597};
                      reg2690 <= {{((reg2579 || (8'hab)) > $unsigned(reg2574))}};
                      reg2691 <= ((($unsigned(reg2425) ?
                              reg2498 : reg2599[(1'h0):(1'h0)]) >> {(8'hba)}) ?
                          $unsigned(forvar2629) : reg2531);
                    end
                  else
                    begin
                      reg2688 <= ($signed((-reg2434)) ?
                          $unsigned($signed({(8'h9d)})) : reg2558[(1'h0):(1'h0)]);
                      reg2689 <= $signed({reg2610[(4'hc):(4'h8)]});
                    end
                  if ((^~$signed(reg2604[(2'h3):(2'h2)])))
                    begin
                      reg2692 <= $signed(forvar2527);
                    end
                  else
                    begin
                      reg2692 <= ({(!(-reg2662))} || $unsigned($signed((reg2400 != forvar2674))));
                    end
                end
              else
                begin
                  if ((((reg2638[(1'h1):(1'h1)] && wire2374[(1'h1):(1'h0)]) - $signed(reg2474[(1'h1):(1'h0)])) ?
                      (^~reg2573) : (((^forvar2534) ?
                              (|reg2587) : $unsigned(wire2373)) ?
                          (&(reg2691 * reg2484)) : ((~&(8'h9d)) ?
                              reg2392[(2'h2):(2'h2)] : (|forvar2628)))))
                    begin
                      reg2688 <= reg2458;
                      reg2689 <= {$unsigned($signed({reg2414}))};
                      reg2690 <= (&$unsigned((~^{reg2681})));
                    end
                  else
                    begin
                      reg2688 <= ($unsigned($unsigned(forvar2583)) + $unsigned(((~^reg2570) ?
                          $unsigned(reg2493) : reg2646)));
                      reg2689 <= forvar2597[(1'h1):(1'h1)];
                    end
                end
              for (forvar2693 = (1'h0); (forvar2693 < (2'h2)); forvar2693 = (forvar2693 + (1'h1)))
                begin
                  if ($unsigned(reg2689[(4'hc):(4'hb)]))
                    begin
                      reg2694 <= $signed((reg2469[(1'h0):(1'h0)] && (+(~^reg2623))));
                      reg2695 <= (|$signed({(reg2386 <<< reg2567)}));
                      reg2696 <= (reg2483[(1'h1):(1'h1)] ?
                          reg2602 : ($signed($signed(reg2591)) ?
                              $unsigned((+reg2452)) : forvar2401));
                    end
                  else
                    begin
                      reg2694 <= forvar2478;
                      reg2695 <= ({((~^reg2571) ?
                                  (forvar2515 ?
                                      reg2561 : forvar2583) : $unsigned(reg2560))} ?
                          $unsigned($signed($signed(forvar2381))) : {$unsigned($unsigned(reg2571))});
                    end
                  for (forvar2697 = (1'h0); (forvar2697 < (2'h2)); forvar2697 = (forvar2697 + (1'h1)))
                    begin
                      reg2698 <= $signed((forvar2394 <= reg2503[(3'h5):(2'h3)]));
                      reg2699 <= ($unsigned((~$unsigned(reg2505))) ?
                          $signed({(~reg2609)}) : $signed(((reg2604 >> reg2413) ^ (reg2499 ?
                              reg2398 : reg2525))));
                      reg2700 <= {$unsigned((~$signed(reg2688)))};
                    end
                  if ($unsigned({{$unsigned(reg2459)}}))
                    begin
                      reg2701 <= $unsigned(($signed($signed((8'ha5))) ?
                          ($unsigned((8'h9d)) ?
                              $unsigned(forvar2529) : $unsigned((8'ha8))) : reg2455[(4'hb):(3'h4)]));
                    end
                  else
                    begin
                      reg2701 <= (~&((+(wire2374 ? reg2381 : (8'ha9))) ?
                          forvar2395[(1'h0):(1'h0)] : reg2393));
                    end
                  for (forvar2702 = (1'h0); (forvar2702 < (1'h0)); forvar2702 = (forvar2702 + (1'h1)))
                    begin
                      reg2703 <= ($unsigned(reg2483) ?
                          $signed($unsigned(forvar2552[(4'h8):(2'h2)])) : reg2470[(1'h0):(1'h0)]);
                    end
                end
              if ((reg2644 ? reg2649[(2'h3):(1'h0)] : (8'ha1)))
                begin
                  if (($unsigned($signed($unsigned(forvar2506))) ~^ $unsigned(reg2457[(4'h8):(1'h1)])))
                    begin
                      reg2704 <= (8'had);
                      reg2705 <= {(!((reg2533 >> reg2585) ?
                              (reg2463 ~^ reg2390) : (forvar2702 ?
                                  (8'hb1) : (8'ha7))))};
                      reg2706 <= reg2467[(4'hb):(4'h8)];
                      reg2707 <= $unsigned(forvar2504[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg2704 <= (8'hb4);
                    end
                  for (forvar2708 = (1'h0); (forvar2708 < (2'h3)); forvar2708 = (forvar2708 + (1'h1)))
                    begin
                      reg2709 <= $unsigned(($signed((!reg2468)) > $unsigned((forvar2506 > forvar2708))));
                    end
                end
              else
                begin
                  for (forvar2704 = (1'h0); (forvar2704 < (1'h1)); forvar2704 = (forvar2704 + (1'h1)))
                    begin
                      reg2705 <= $unsigned(((forvar2476 ?
                          (reg2654 ^ (8'hb6)) : ((8'hba) ?
                              reg2564 : (8'ha3))) ~^ forvar2546[(4'hd):(3'h7)]));
                      reg2706 <= reg2701[(3'h6):(2'h2)];
                      reg2707 <= $unsigned((-{(|(8'hb4))}));
                      reg2708 <= $signed(forvar2396[(4'hb):(3'h5)]);
                    end
                  if (($signed((~|$unsigned(reg2535))) ?
                      $unsigned(forvar2584[(2'h3):(2'h3)]) : $signed(reg2452[(3'h4):(1'h1)])))
                    begin
                      reg2709 <= (($signed(reg2383) ?
                              $signed(reg2565[(2'h2):(1'h1)]) : ((forvar2553 + reg2525) ?
                                  (reg2524 ^~ forvar2606) : {reg2650})) ?
                          {(~^forvar2435)} : ($signed(reg2500) ?
                              {reg2631} : forvar2678[(4'ha):(2'h2)]));
                      reg2710 <= reg2525;
                      reg2711 <= ((8'hb6) ?
                          forvar2476 : forvar2697[(3'h7):(1'h1)]);
                    end
                  else
                    begin
                      reg2709 <= ($signed((&reg2647[(2'h2):(2'h2)])) ?
                          reg2590[(3'h6):(3'h4)] : (reg2424[(2'h2):(1'h0)] - $signed($unsigned(reg2659))));
                      reg2710 <= $signed(($unsigned({reg2490}) ?
                          (reg2473[(2'h2):(1'h0)] ^ (forvar2558 > forvar2586)) : ($unsigned(reg2652) ?
                              $unsigned(reg2524) : (forvar2597 || reg2620))));
                      reg2711 <= (forvar2426 ?
                          reg2599[(1'h0):(1'h0)] : (($signed((8'hae)) ?
                              (8'ha0) : (reg2499 > reg2613)) - ((reg2691 ?
                              (8'hb0) : reg2591) >>> $unsigned(reg2565))));
                    end
                  if ({$signed(($unsigned(forvar2536) << $unsigned((8'hab))))})
                    begin
                      reg2712 <= $signed(forvar2616[(1'h1):(1'h0)]);
                      reg2713 <= (reg2585[(2'h3):(1'h1)] ~^ $unsigned(($unsigned((8'h9d)) >= $unsigned(forvar2420))));
                      reg2714 <= $unsigned($unsigned(reg2464));
                      reg2715 <= ({(^~{reg2477})} != {$unsigned((~&reg2548))});
                    end
                  else
                    begin
                      reg2712 <= (({$signed(reg2568)} ?
                              $signed(forvar2557) : $unsigned((!reg2706))) ?
                          ({(reg2615 >> forvar2465)} ?
                              ((reg2454 || reg2597) >>> (reg2673 ?
                                  forvar2389 : reg2569)) : reg2550) : ($signed(reg2607[(4'hc):(4'hc)]) ?
                              {(reg2457 <= (8'ha0))} : reg2664[(2'h3):(2'h3)]));
                    end
                  for (forvar2716 = (1'h0); (forvar2716 < (2'h3)); forvar2716 = (forvar2716 + (1'h1)))
                    begin
                      reg2717 <= reg2647;
                    end
                end
            end
          else
            begin
              for (forvar2688 = (1'h0); (forvar2688 < (2'h2)); forvar2688 = (forvar2688 + (1'h1)))
                begin
                  for (forvar2689 = (1'h0); (forvar2689 < (1'h1)); forvar2689 = (forvar2689 + (1'h1)))
                    begin
                      reg2690 <= $unsigned($signed(reg2500));
                      reg2691 <= reg2424;
                      reg2692 <= ((|forvar2583[(4'ha):(3'h5)]) ?
                          (~&$unsigned(reg2441[(2'h2):(1'h0)])) : ((reg2632[(2'h2):(1'h1)] ^ (~|reg2701)) ?
                              (~|reg2517[(2'h3):(1'h1)]) : $unsigned((forvar2546 ?
                                  reg2703 : reg2626))));
                    end
                  if ($signed($unsigned($signed($signed(reg2491)))))
                    begin
                      reg2693 <= (8'hb3);
                      reg2694 <= $unsigned((!(&$unsigned(reg2654))));
                    end
                  else
                    begin
                      reg2693 <= ((!$unsigned($unsigned(reg2692))) ?
                          {$signed(reg2684)} : {($unsigned(reg2404) ?
                                  reg2602[(4'ha):(3'h6)] : $unsigned(reg2636))});
                      reg2694 <= (~^($unsigned(reg2509[(2'h3):(1'h0)]) || reg2478));
                    end
                  reg2695 <= forvar2672;
                end
              reg2696 <= ($unsigned(reg2601[(4'h9):(4'h8)]) <= ({$unsigned(forvar2611)} ?
                  (~^{reg2387}) : $signed(reg2413)));
              for (forvar2697 = (1'h0); (forvar2697 < (2'h3)); forvar2697 = (forvar2697 + (1'h1)))
                begin
                  for (forvar2698 = (1'h0); (forvar2698 < (1'h0)); forvar2698 = (forvar2698 + (1'h1)))
                    begin
                      reg2699 <= $unsigned($signed(reg2555));
                    end
                  if (((reg2386[(1'h1):(1'h1)] ^ $signed((reg2477 ~^ reg2535))) ?
                      $signed(reg2559[(1'h0):(1'h0)]) : forvar2545[(3'h4):(2'h2)]))
                    begin
                      reg2700 <= $signed(((forvar2583 ?
                              {reg2416} : reg2386[(1'h0):(1'h0)]) ?
                          $signed({(8'h9e)}) : (^(reg2428 <= forvar2465))));
                      reg2701 <= $unsigned(reg2507);
                    end
                  else
                    begin
                      reg2700 <= (^(reg2570[(1'h1):(1'h1)] + (|(reg2590 ?
                          reg2520 : reg2429))));
                      reg2701 <= $signed((~^(~reg2474[(4'hd):(4'hb)])));
                      reg2702 <= ((8'haa) ?
                          ($unsigned({reg2531}) ?
                              ({(8'ha9)} ?
                                  (^~forvar2407) : {forvar2465}) : reg2582[(2'h3):(2'h2)]) : forvar2418);
                      reg2703 <= $unsigned(((-{forvar2627}) <<< $unsigned($unsigned(reg2500))));
                    end
                  for (forvar2704 = (1'h0); (forvar2704 < (2'h3)); forvar2704 = (forvar2704 + (1'h1)))
                    begin
                      reg2705 <= ((8'h9d) || {$unsigned($signed(forvar2693))});
                    end
                  for (forvar2706 = (1'h0); (forvar2706 < (2'h3)); forvar2706 = (forvar2706 + (1'h1)))
                    begin
                      reg2707 <= $signed((8'hb9));
                      reg2708 <= reg2440;
                      reg2709 <= $unsigned($signed({(forvar2458 ?
                              forvar2677 : reg2437)}));
                      reg2710 <= reg2567[(1'h1):(1'h1)];
                    end
                end
              if (({(|(reg2630 ? forvar2683 : (8'h9d)))} ?
                  reg2427 : forvar2683[(4'hd):(4'h8)]))
                begin
                  for (forvar2711 = (1'h0); (forvar2711 < (2'h3)); forvar2711 = (forvar2711 + (1'h1)))
                    begin
                      reg2712 <= (forvar2545[(3'h6):(2'h3)] ?
                          ((forvar2655[(1'h1):(1'h1)] == ((8'hb2) ?
                                  forvar2608 : reg2630)) ?
                              reg2673 : ($signed(forvar2401) * reg2646[(3'h7):(2'h3)])) : reg2630);
                    end
                  reg2713 <= $unsigned(({{reg2557}} >> {(reg2437 && forvar2486)}));
                end
              else
                begin
                  for (forvar2711 = (1'h0); (forvar2711 < (1'h1)); forvar2711 = (forvar2711 + (1'h1)))
                    begin
                      reg2712 <= reg2479[(1'h1):(1'h0)];
                      reg2713 <= $signed(reg2409[(3'h6):(3'h6)]);
                      reg2714 <= ({$unsigned($unsigned(reg2521))} >> (~^(8'ha2)));
                      reg2715 <= ((!forvar2515[(2'h2):(1'h0)]) - ({(reg2556 ?
                              reg2434 : reg2479)} | (&forvar2601[(2'h2):(2'h2)])));
                    end
                  for (forvar2716 = (1'h0); (forvar2716 < (1'h0)); forvar2716 = (forvar2716 + (1'h1)))
                    begin
                      reg2717 <= wire2375;
                      reg2718 <= $signed(({(|reg2650)} ?
                          (+(reg2495 ? forvar2616 : reg2427)) : reg2421));
                      reg2719 <= {reg2421};
                      reg2720 <= ($unsigned((forvar2488[(3'h7):(3'h4)] ?
                          $unsigned(reg2658) : ((8'hb6) & reg2631))) | reg2548[(3'h7):(3'h6)]);
                    end
                  if (reg2425[(1'h0):(1'h0)])
                    begin
                      reg2721 <= {forvar2678};
                      reg2722 <= reg2499;
                      reg2723 <= reg2507[(3'h5):(1'h0)];
                      reg2724 <= {(~|reg2669)};
                    end
                  else
                    begin
                      reg2721 <= $signed($signed($signed($unsigned(forvar2589))));
                      reg2722 <= $unsigned($unsigned({$signed(reg2685)}));
                    end
                end
            end
        end
      else
        begin
          if (reg2510[(1'h0):(1'h0)])
            begin
              for (forvar2671 = (1'h0); (forvar2671 < (1'h0)); forvar2671 = (forvar2671 + (1'h1)))
                begin
                  reg2672 <= (-$signed($signed(reg2651)));
                  for (forvar2673 = (1'h0); (forvar2673 < (1'h1)); forvar2673 = (forvar2673 + (1'h1)))
                    begin
                      reg2674 <= ((reg2653 || (!(reg2676 ?
                              reg2714 : reg2563))) ?
                          ($signed($unsigned(reg2636)) | reg2580) : reg2705[(3'h7):(3'h5)]);
                      reg2675 <= $signed($signed((reg2393 ?
                          {reg2714} : (reg2539 ? reg2402 : forvar2427))));
                    end
                  for (forvar2676 = (1'h0); (forvar2676 < (2'h3)); forvar2676 = (forvar2676 + (1'h1)))
                    begin
                      reg2677 <= ($unsigned($unsigned({forvar2407})) ?
                          $signed(reg2445[(3'h5):(1'h1)]) : {((-reg2664) ?
                                  {reg2522} : ((8'hb2) ? (8'h9d) : reg2722))});
                      reg2678 <= ((~forvar2676[(2'h3):(1'h1)]) ?
                          $unsigned((+(reg2411 & forvar2497))) : $signed($unsigned($signed(reg2525))));
                      reg2679 <= $signed($signed($signed(reg2570[(1'h0):(1'h0)])));
                    end
                end
              for (forvar2680 = (1'h0); (forvar2680 < (1'h0)); forvar2680 = (forvar2680 + (1'h1)))
                begin
                  reg2681 <= (!$signed(reg2483));
                  for (forvar2682 = (1'h0); (forvar2682 < (1'h0)); forvar2682 = (forvar2682 + (1'h1)))
                    begin
                      reg2683 <= reg2658;
                    end
                  if ((+$signed(reg2679)))
                    begin
                      reg2684 <= (8'hab);
                      reg2685 <= reg2457;
                    end
                  else
                    begin
                      reg2684 <= $signed((reg2409 ?
                          ((^~forvar2577) ?
                              forvar2577[(3'h6):(3'h4)] : $unsigned((8'ha1))) : (~&(~&reg2642))));
                    end
                  reg2686 <= forvar2420[(3'h4):(1'h0)];
                end
              for (forvar2687 = (1'h0); (forvar2687 < (1'h1)); forvar2687 = (forvar2687 + (1'h1)))
                begin
                  for (forvar2688 = (1'h0); (forvar2688 < (2'h2)); forvar2688 = (forvar2688 + (1'h1)))
                    begin
                      reg2689 <= (reg2381 ?
                          (reg2527[(3'h6):(3'h6)] <= forvar2597) : reg2426[(3'h4):(2'h2)]);
                      reg2690 <= ((($signed((8'hb0)) ?
                          (forvar2468 ?
                              (8'h9d) : reg2646) : $unsigned(forvar2673)) + (reg2484[(3'h4):(2'h3)] ~^ (^reg2529))) << (&($signed(wire2511) ?
                          (~&reg2593) : reg2468[(1'h0):(1'h0)])));
                    end
                  if (((8'hb9) ?
                      ((~reg2718[(1'h0):(1'h0)]) ?
                          (~^forvar2379[(1'h1):(1'h0)]) : reg2541) : $signed((reg2703[(4'h8):(1'h0)] ?
                          (^forvar2401) : (reg2610 >>> reg2475)))))
                    begin
                      reg2691 <= $unsigned({{$signed(reg2690)}});
                      reg2692 <= forvar2469;
                    end
                  else
                    begin
                      reg2691 <= (8'hb8);
                    end
                  reg2693 <= (~^$signed(((~reg2596) == $signed(forvar2426))));
                end
              for (forvar2694 = (1'h0); (forvar2694 < (2'h2)); forvar2694 = (forvar2694 + (1'h1)))
                begin
                  reg2695 <= {(8'hab)};
                  if ({$signed((~|wire2372))})
                    begin
                      reg2696 <= (^reg2439[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2696 <= ((^forvar2655) ?
                          $unsigned((~(^reg2541))) : (|reg2423[(5'h10):(4'hf)]));
                      reg2697 <= reg2466;
                    end
                  for (forvar2698 = (1'h0); (forvar2698 < (1'h1)); forvar2698 = (forvar2698 + (1'h1)))
                    begin
                      reg2699 <= ((^({(8'hb9)} ?
                              reg2509 : reg2464[(4'hf):(4'he)])) ?
                          reg2560[(1'h1):(1'h1)] : (~forvar2688[(1'h0):(1'h0)]));
                      reg2700 <= $signed($signed($unsigned($unsigned(forvar2711))));
                      reg2701 <= {(((forvar2612 ?
                                  reg2410 : (8'ha8)) < reg2455) ?
                              $unsigned((~|forvar2680)) : $unsigned($unsigned((8'hb9))))};
                    end
                  reg2702 <= reg2561[(3'h7):(2'h3)];
                end
            end
          else
            begin
              if ($signed((((~^forvar2486) <<< $signed(forvar2553)) >>> ((~^reg2404) || (&reg2501)))))
                begin
                  reg2671 <= {({$unsigned(reg2509)} ?
                          reg2505 : {((8'h9f) || reg2719)})};
                end
              else
                begin
                  reg2671 <= ({((-reg2568) < $unsigned(wire2373))} ?
                      $signed((~&$signed(reg2553))) : reg2528[(3'h7):(3'h4)]);
                  if (reg2466[(4'h8):(2'h2)])
                    begin
                      reg2672 <= (reg2570[(1'h0):(1'h0)] ^~ reg2417);
                      reg2673 <= $unsigned($signed(($signed(reg2719) ?
                          $unsigned(reg2574) : ((8'hb4) ?
                              forvar2493 : reg2642))));
                    end
                  else
                    begin
                      reg2672 <= $unsigned(forvar2584);
                      reg2673 <= (~|$unsigned({(reg2551 ? reg2527 : (8'haf))}));
                      reg2674 <= (^~$signed({$signed(reg2718)}));
                      reg2675 <= (~|reg2662[(3'h4):(2'h2)]);
                    end
                  reg2676 <= reg2387[(1'h1):(1'h1)];
                end
            end
          for (forvar2703 = (1'h0); (forvar2703 < (1'h0)); forvar2703 = (forvar2703 + (1'h1)))
            begin
              for (forvar2704 = (1'h0); (forvar2704 < (2'h3)); forvar2704 = (forvar2704 + (1'h1)))
                begin
                  reg2705 <= (~|$unsigned(((reg2597 < reg2548) ?
                      $signed(reg2482) : $signed(reg2703))));
                  if ((~&$signed(((~^reg2524) || (reg2604 ~^ (8'ha5))))))
                    begin
                      reg2706 <= reg2665[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg2706 <= (forvar2593[(4'h9):(3'h4)] | {$unsigned((^(8'hb8)))});
                      reg2707 <= {(~$signed($signed(reg2686)))};
                      reg2708 <= reg2539[(3'h7):(2'h2)];
                      reg2709 <= ((forvar2689 ?
                          ({reg2532} <= ((8'hab) ?
                              reg2601 : reg2617)) : ((reg2460 ?
                              forvar2706 : (8'ha6)) ^~ (reg2481 != wire2376))) <<< forvar2688[(1'h0):(1'h0)]);
                    end
                  if (reg2450)
                    begin
                      reg2710 <= (!$signed($signed(((8'h9f) ?
                          (8'haf) : forvar2584))));
                      reg2711 <= {forvar2672[(3'h6):(3'h4)]};
                      reg2712 <= $unsigned(forvar2559[(3'h6):(3'h6)]);
                    end
                  else
                    begin
                      reg2710 <= reg2546;
                      reg2711 <= reg2495;
                      reg2712 <= reg2599[(1'h0):(1'h0)];
                    end
                  if ($signed((+($signed(forvar2608) ?
                      (reg2521 >>> reg2407) : (forvar2689 ?
                          reg2710 : (8'hb1))))))
                    begin
                      reg2713 <= $unsigned(reg2489[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2713 <= ((~reg2434[(2'h2):(1'h0)]) << $signed($unsigned($unsigned(reg2689))));
                      reg2714 <= reg2554[(1'h0):(1'h0)];
                      reg2715 <= ($signed(reg2588[(3'h4):(2'h3)]) >> ((^(reg2569 + reg2462)) == forvar2564));
                      reg2716 <= $unsigned(forvar2426);
                    end
                end
              if ({reg2392[(3'h5):(3'h5)]})
                begin
                  for (forvar2717 = (1'h0); (forvar2717 < (2'h2)); forvar2717 = (forvar2717 + (1'h1)))
                    begin
                      reg2718 <= (($signed(reg2473) || (|(!reg2567))) <<< $signed(forvar2666));
                      reg2719 <= ((reg2463[(1'h0):(1'h0)] + {{reg2705}}) << ($signed(((8'hb4) ?
                              reg2493 : forvar2504)) ?
                          wire2375 : (8'hb9)));
                      reg2720 <= (($unsigned(forvar2504) >>> {(^~forvar2643)}) ?
                          (8'h9d) : (-$unsigned(reg2465[(4'hc):(2'h2)])));
                    end
                  for (forvar2721 = (1'h0); (forvar2721 < (1'h1)); forvar2721 = (forvar2721 + (1'h1)))
                    begin
                      reg2722 <= (($signed($unsigned(reg2676)) ?
                          forvar2683[(4'h9):(3'h5)] : (reg2476[(2'h2):(1'h0)] ?
                              (&reg2584) : (~|reg2650))) | (-$signed($signed(reg2527))));
                      reg2723 <= (+$unsigned((reg2456[(3'h4):(1'h0)] != $signed(reg2594))));
                      reg2724 <= reg2671;
                      reg2725 <= ((8'ha9) == {{(reg2386 ?
                                  wire2372 : reg2502)}});
                    end
                  reg2726 <= (~(((reg2670 != reg2677) ?
                      (reg2590 ? reg2706 : reg2480) : reg2473) + reg2490));
                  reg2727 <= reg2438[(1'h1):(1'h1)];
                end
              else
                begin
                  for (forvar2717 = (1'h0); (forvar2717 < (1'h1)); forvar2717 = (forvar2717 + (1'h1)))
                    begin
                      reg2718 <= $signed($unsigned((8'ha8)));
                      reg2719 <= reg2560[(3'h4):(2'h2)];
                    end
                  for (forvar2720 = (1'h0); (forvar2720 < (2'h2)); forvar2720 = (forvar2720 + (1'h1)))
                    begin
                      reg2721 <= (~|$signed($signed((forvar2475 ?
                          reg2669 : forvar2656))));
                      reg2722 <= reg2498;
                      reg2723 <= {forvar2488};
                      reg2724 <= reg2491[(1'h1):(1'h1)];
                    end
                end
            end
        end
      for (forvar2728 = (1'h0); (forvar2728 < (1'h1)); forvar2728 = (forvar2728 + (1'h1)))
        begin
          if (reg2431)
            begin
              reg2729 <= (8'hb6);
            end
          else
            begin
              if (forvar2564)
                begin
                  for (forvar2729 = (1'h0); (forvar2729 < (1'h0)); forvar2729 = (forvar2729 + (1'h1)))
                    begin
                      reg2730 <= (~&$unsigned(forvar2527));
                      reg2731 <= (({(reg2507 | reg2489)} == ((8'h9f) >= reg2687)) ?
                          forvar2478 : ((reg2671[(3'h7):(3'h7)] << (forvar2639 ?
                              forvar2698 : reg2496)) < (reg2523[(2'h2):(1'h0)] ?
                              ((8'hb5) ?
                                  forvar2436 : reg2667) : reg2667[(3'h5):(2'h3)])));
                    end
                  if ((~&(((~|reg2498) & reg2631[(3'h5):(3'h4)]) - ($signed(reg2727) && (reg2465 + reg2437)))))
                    begin
                      reg2732 <= ((^forvar2584[(1'h1):(1'h1)]) ~^ reg2498[(3'h4):(2'h2)]);
                      reg2733 <= ($unsigned((+forvar2552[(2'h3):(1'h1)])) ?
                          reg2606 : {(+reg2701[(1'h1):(1'h0)])});
                    end
                  else
                    begin
                      reg2732 <= ({({(8'ha4)} < $unsigned((8'h9f)))} < forvar2473);
                      reg2733 <= (~|reg2411[(1'h0):(1'h0)]);
                      reg2734 <= ($unsigned((8'ha4)) ?
                          {(~(reg2408 * (8'hba)))} : reg2682[(2'h3):(2'h2)]);
                      reg2735 <= ((($signed((8'h9d)) ?
                              $unsigned(forvar2674) : $unsigned(reg2469)) <<< reg2574[(3'h5):(2'h3)]) ?
                          reg2575[(4'ha):(4'h9)] : (reg2553 ^ reg2697));
                    end
                end
              else
                begin
                  if (reg2528[(1'h0):(1'h0)])
                    begin
                      reg2729 <= ({{$signed(reg2703)}} ?
                          (^~(~^((8'hba) ?
                              reg2591 : reg2552))) : (((forvar2702 ^~ (8'h9e)) ?
                                  $signed(reg2458) : $signed(reg2479)) ?
                              ((reg2387 >= reg2602) ?
                                  $unsigned(reg2678) : $signed(forvar2418)) : ($unsigned(reg2505) ?
                                  reg2549 : (reg2390 ? reg2476 : forvar2655))));
                      reg2730 <= (({$unsigned(forvar2506)} || $signed(reg2452)) ?
                          ($unsigned($unsigned((8'had))) < (forvar2525[(3'h4):(2'h3)] ?
                              (&reg2718) : $unsigned(reg2703))) : $unsigned({$unsigned(reg2432)}));
                      reg2731 <= (+$signed((~&reg2578[(2'h2):(1'h1)])));
                      reg2732 <= $unsigned($unsigned($signed((forvar2545 || reg2650))));
                    end
                  else
                    begin
                      reg2729 <= (~(8'hb7));
                    end
                  reg2733 <= reg2597[(4'hc):(3'h6)];
                  for (forvar2734 = (1'h0); (forvar2734 < (2'h3)); forvar2734 = (forvar2734 + (1'h1)))
                    begin
                      reg2735 <= ($unsigned(reg2684) > $signed($signed($signed(reg2551))));
                      reg2736 <= forvar2516[(2'h2):(1'h0)];
                      reg2737 <= $signed(forvar2708);
                    end
                end
            end
          if (((reg2636[(2'h2):(2'h2)] * (^(~^reg2430))) & reg2618[(4'h8):(2'h2)]))
            begin
              for (forvar2738 = (1'h0); (forvar2738 < (1'h0)); forvar2738 = (forvar2738 + (1'h1)))
                begin
                  if (forvar2703[(2'h3):(1'h0)])
                    begin
                      reg2739 <= (~|(~&((forvar2534 * forvar2476) ~^ (reg2445 || forvar2720))));
                      reg2740 <= ((~&(~^forvar2616[(1'h1):(1'h1)])) >= {forvar2427});
                      reg2741 <= ((~^((reg2568 | reg2697) ?
                              (reg2558 & reg2649) : reg2686[(1'h1):(1'h1)])) ?
                          ((reg2425[(4'ha):(4'h9)] ?
                              (reg2611 ^ reg2557) : reg2423[(3'h5):(2'h3)]) <= (~^reg2574[(2'h3):(2'h2)])) : (~|(-$unsigned(reg2735))));
                    end
                  else
                    begin
                      reg2739 <= reg2386[(1'h0):(1'h0)];
                    end
                  for (forvar2742 = (1'h0); (forvar2742 < (2'h2)); forvar2742 = (forvar2742 + (1'h1)))
                    begin
                      reg2743 <= ($signed({reg2426}) ?
                          $unsigned($unsigned({reg2732})) : (reg2430 << ($unsigned(reg2523) ?
                              ((8'ha1) << reg2633) : forvar2583)));
                      reg2744 <= (($signed($unsigned(forvar2577)) ?
                          $signed((reg2569 ?
                              forvar2546 : reg2388)) : reg2450[(3'h5):(3'h5)]) || $unsigned((reg2475 ?
                          {(8'had)} : $signed(reg2658))));
                      reg2745 <= (!$unsigned({(|reg2541)}));
                      reg2746 <= ($unsigned($signed($signed(reg2674))) ?
                          $signed((~((8'hb0) << forvar2651))) : $signed((8'hb3)));
                    end
                end
            end
          else
            begin
              for (forvar2738 = (1'h0); (forvar2738 < (2'h3)); forvar2738 = (forvar2738 + (1'h1)))
                begin
                  for (forvar2739 = (1'h0); (forvar2739 < (1'h1)); forvar2739 = (forvar2739 + (1'h1)))
                    begin
                      reg2740 <= $signed((-(forvar2420[(2'h2):(1'h1)] == (reg2625 < (8'haf)))));
                      reg2741 <= (((+$signed(forvar2717)) >>> {$signed(forvar2639)}) ?
                          $unsigned(reg2639) : ((!$unsigned(reg2638)) ?
                              ({forvar2618} ?
                                  forvar2721[(1'h1):(1'h1)] : $signed(reg2704)) : (reg2642 * $signed(reg2564))));
                    end
                end
              if ($unsigned(reg2432[(1'h1):(1'h1)]))
                begin
                  reg2742 <= (!(reg2550[(1'h1):(1'h0)] * ({forvar2655} < (!(8'hb7)))));
                  reg2743 <= $signed($signed($signed($signed(reg2703))));
                  for (forvar2744 = (1'h0); (forvar2744 < (2'h2)); forvar2744 = (forvar2744 + (1'h1)))
                    begin
                      reg2745 <= reg2579[(3'h4):(2'h2)];
                    end
                  for (forvar2746 = (1'h0); (forvar2746 < (2'h3)); forvar2746 = (forvar2746 + (1'h1)))
                    begin
                      reg2747 <= $unsigned(reg2533[(3'h6):(1'h0)]);
                      reg2748 <= $unsigned((&($signed(forvar2552) ?
                          $unsigned(reg2382) : $signed(reg2708))));
                      reg2749 <= ((|reg2605) ?
                          (reg2416 - ($signed(forvar2674) ?
                              ((8'ha3) >= wire2375) : $signed((8'hab)))) : {(-(8'hba))});
                      reg2750 <= reg2466[(4'hf):(4'ha)];
                    end
                end
              else
                begin
                  reg2742 <= (($unsigned(((8'hb9) > forvar2680)) ?
                          $unsigned({wire2375}) : ($unsigned(forvar2521) ?
                              $signed((8'hb4)) : {reg2505})) ?
                      {(!reg2388[(1'h1):(1'h1)])} : (-(8'haa)));
                  reg2743 <= reg2475;
                end
            end
        end
      if (((~((~^reg2619) ?
          (+reg2526) : ((8'hb4) ?
              reg2750 : reg2598))) != $signed(($signed(reg2530) && (reg2397 == forvar2468)))))
        begin
          for (forvar2751 = (1'h0); (forvar2751 < (1'h1)); forvar2751 = (forvar2751 + (1'h1)))
            begin
              for (forvar2752 = (1'h0); (forvar2752 < (2'h3)); forvar2752 = (forvar2752 + (1'h1)))
                begin
                  for (forvar2753 = (1'h0); (forvar2753 < (1'h1)); forvar2753 = (forvar2753 + (1'h1)))
                    begin
                      reg2754 <= forvar2742[(3'h5):(2'h2)];
                    end
                  if (($unsigned(reg2683[(3'h6):(3'h4)]) & forvar2544[(3'h5):(2'h2)]))
                    begin
                      reg2755 <= ($unsigned($unsigned($unsigned(reg2729))) ?
                          $signed(((~^reg2562) - $unsigned(reg2609))) : ({(8'hab)} ?
                              reg2604[(1'h1):(1'h1)] : (~forvar2583[(3'h6):(3'h6)])));
                      reg2756 <= reg2732[(4'h9):(4'h9)];
                      reg2757 <= reg2544[(4'hb):(3'h5)];
                      reg2758 <= forvar2611[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg2755 <= forvar2475[(1'h1):(1'h1)];
                    end
                end
            end
          reg2759 <= $unsigned(($signed(forvar2728[(2'h2):(2'h2)]) >= reg2411[(1'h0):(1'h0)]));
          for (forvar2760 = (1'h0); (forvar2760 < (1'h1)); forvar2760 = (forvar2760 + (1'h1)))
            begin
              for (forvar2761 = (1'h0); (forvar2761 < (2'h2)); forvar2761 = (forvar2761 + (1'h1)))
                begin
                  reg2762 <= {((reg2386[(3'h4):(3'h4)] ?
                          (!forvar2389) : {reg2440}) <<< {reg2680})};
                  reg2763 <= reg2704;
                  if (({({(8'had)} > (8'haf))} ?
                      forvar2639 : wire2375[(3'h4):(1'h1)]))
                    begin
                      reg2764 <= reg2649[(1'h0):(1'h0)];
                      reg2765 <= reg2756;
                      reg2766 <= (!(forvar2561[(2'h2):(1'h0)] * (8'hb7)));
                    end
                  else
                    begin
                      reg2764 <= (~&((+{(8'ha5)}) > $signed((reg2668 >>> reg2764))));
                      reg2765 <= (&(~(~&{forvar2453})));
                      reg2766 <= reg2571;
                    end
                end
              reg2767 <= (8'hba);
              for (forvar2768 = (1'h0); (forvar2768 < (1'h0)); forvar2768 = (forvar2768 + (1'h1)))
                begin
                  reg2769 <= $unsigned(reg2662);
                  if ($signed({(^~(~|(8'ha5)))}))
                    begin
                      reg2770 <= ($unsigned({(8'ha9)}) ?
                          ($signed(reg2386) ?
                              (wire2377[(3'h6):(3'h4)] << {reg2484}) : $signed(reg2533)) : ((~^{reg2685}) ?
                              ($signed(wire2512) ?
                                  $signed(reg2411) : (^~reg2692)) : $signed($signed(reg2736))));
                    end
                  else
                    begin
                      reg2770 <= (((~|(~^reg2494)) ?
                          forvar2556[(1'h0):(1'h0)] : (-reg2675)) != $signed(reg2535));
                      reg2771 <= $signed((&($signed(reg2529) - forvar2674[(1'h0):(1'h0)])));
                      reg2772 <= ((&(8'hb6)) >= forvar2488);
                    end
                  for (forvar2773 = (1'h0); (forvar2773 < (2'h2)); forvar2773 = (forvar2773 + (1'h1)))
                    begin
                      reg2774 <= reg2688[(4'hc):(4'ha)];
                      reg2775 <= reg2406;
                      reg2776 <= {$signed({(^~forvar2753)})};
                    end
                end
            end
          if ((~|(-forvar2518)))
            begin
              for (forvar2777 = (1'h0); (forvar2777 < (1'h1)); forvar2777 = (forvar2777 + (1'h1)))
                begin
                  for (forvar2778 = (1'h0); (forvar2778 < (1'h1)); forvar2778 = (forvar2778 + (1'h1)))
                    begin
                      reg2779 <= $signed(reg2493);
                      reg2780 <= (reg2705[(3'h7):(1'h0)] ?
                          (((wire2513 ? forvar2721 : reg2509) * {reg2384}) ?
                              ($signed(reg2479) ?
                                  (forvar2689 << reg2509) : (wire2511 ?
                                      reg2765 : reg2549)) : reg2588) : (~|forvar2427));
                      reg2781 <= $signed((reg2392[(1'h1):(1'h0)] ?
                          reg2406[(1'h1):(1'h1)] : reg2407));
                      reg2782 <= ($signed($signed((+reg2564))) ?
                          (^~reg2702[(3'h6):(3'h6)]) : (8'haa));
                    end
                  for (forvar2783 = (1'h0); (forvar2783 < (2'h2)); forvar2783 = (forvar2783 + (1'h1)))
                    begin
                      reg2784 <= ({$signed((!forvar2465))} ?
                          (-(forvar2612[(2'h2):(1'h0)] ?
                              reg2403 : $signed((8'had)))) : reg2417[(3'h4):(2'h2)]);
                      reg2785 <= $unsigned(forvar2612[(1'h0):(1'h0)]);
                      reg2786 <= ((reg2691 ?
                          ({forvar2702} ?
                              $unsigned((8'h9d)) : (reg2779 > forvar2783)) : {$unsigned(reg2680)}) ^~ $signed((+$signed(reg2452))));
                    end
                  for (forvar2787 = (1'h0); (forvar2787 < (1'h0)); forvar2787 = (forvar2787 + (1'h1)))
                    begin
                      reg2788 <= $signed((($signed(reg2725) ?
                              {reg2526} : reg2647[(1'h0):(1'h0)]) ?
                          ($signed(forvar2401) < (|(8'hb8))) : $signed(forvar2729)));
                      reg2789 <= ((!(reg2775 * $unsigned(forvar2536))) ?
                          ({(reg2723 ^ reg2404)} * ((8'ha6) >> forvar2577[(2'h3):(2'h3)])) : (wire2375 ?
                              {(reg2730 ?
                                      forvar2687 : reg2502)} : reg2573[(1'h0):(1'h0)]));
                    end
                end
              reg2790 <= ({$unsigned($signed((8'hb8)))} ?
                  $unsigned(forvar2427) : $unsigned((forvar2627 != $signed(reg2710))));
            end
          else
            begin
              reg2777 <= forvar2673[(2'h3):(2'h3)];
            end
        end
      else
        begin
          for (forvar2751 = (1'h0); (forvar2751 < (2'h3)); forvar2751 = (forvar2751 + (1'h1)))
            begin
              for (forvar2752 = (1'h0); (forvar2752 < (1'h0)); forvar2752 = (forvar2752 + (1'h1)))
                begin
                  for (forvar2753 = (1'h0); (forvar2753 < (1'h0)); forvar2753 = (forvar2753 + (1'h1)))
                    begin
                      reg2754 <= reg2785[(2'h3):(1'h0)];
                      reg2755 <= $unsigned(reg2777[(4'hb):(1'h1)]);
                    end
                  for (forvar2756 = (1'h0); (forvar2756 < (2'h3)); forvar2756 = (forvar2756 + (1'h1)))
                    begin
                      reg2757 <= reg2677;
                    end
                  reg2758 <= $signed(($signed(reg2756) == ($signed((8'hb9)) > reg2565[(2'h2):(1'h0)])));
                end
              if (($unsigned((reg2591[(3'h6):(2'h3)] ?
                      (^~(8'hb3)) : $unsigned(forvar2618))) ?
                  $signed($signed((forvar2678 >>> forvar2651))) : (+((reg2564 | forvar2678) << $unsigned(forvar2597)))))
                begin
                  reg2759 <= forvar2552;
                  for (forvar2760 = (1'h0); (forvar2760 < (1'h1)); forvar2760 = (forvar2760 + (1'h1)))
                    begin
                      reg2761 <= reg2434[(3'h7):(2'h3)];
                      reg2762 <= forvar2518[(4'ha):(4'ha)];
                    end
                  for (forvar2763 = (1'h0); (forvar2763 < (1'h1)); forvar2763 = (forvar2763 + (1'h1)))
                    begin
                      reg2764 <= $signed(((+reg2426) ?
                          (^forvar2716[(1'h1):(1'h0)]) : ((!forvar2553) > reg2675)));
                      reg2765 <= {$signed($signed($unsigned(reg2758)))};
                      reg2766 <= reg2705[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar2759 = (1'h0); (forvar2759 < (1'h0)); forvar2759 = (forvar2759 + (1'h1)))
                    begin
                      reg2760 <= $signed(reg2391[(3'h6):(2'h3)]);
                      reg2761 <= reg2743;
                      reg2762 <= $unsigned((~^{(~|forvar2537)}));
                    end
                  for (forvar2763 = (1'h0); (forvar2763 < (2'h3)); forvar2763 = (forvar2763 + (1'h1)))
                    begin
                      reg2764 <= (forvar2379 ?
                          ((reg2532[(1'h1):(1'h1)] ?
                                  forvar2729[(1'h1):(1'h0)] : $unsigned(forvar2763)) ?
                              $signed((8'ha0)) : reg2615) : (($unsigned(forvar2516) ?
                                  (reg2659 && reg2602) : (forvar2473 ?
                                      reg2747 : (8'h9e))) ?
                              $unsigned({reg2491}) : forvar2564));
                      reg2765 <= $unsigned(reg2536);
                      reg2766 <= forvar2666[(3'h7):(3'h4)];
                    end
                end
              for (forvar2767 = (1'h0); (forvar2767 < (2'h2)); forvar2767 = (forvar2767 + (1'h1)))
                begin
                  for (forvar2768 = (1'h0); (forvar2768 < (1'h0)); forvar2768 = (forvar2768 + (1'h1)))
                    begin
                      reg2769 <= (reg2676[(1'h1):(1'h1)] ?
                          reg2516 : forvar2473[(1'h0):(1'h0)]);
                      reg2770 <= (reg2749 ?
                          {(reg2689[(4'h9):(3'h7)] >> $unsigned(reg2466))} : {(8'ha7)});
                      reg2771 <= $signed((~|reg2750));
                      reg2772 <= reg2624[(1'h1):(1'h0)];
                    end
                  if (($unsigned($signed((~^reg2406))) ?
                      reg2541 : $signed(((!(8'ha2)) + $signed((8'ha2))))))
                    begin
                      reg2773 <= ((forvar2536 <<< $unsigned((forvar2556 + forvar2379))) ?
                          wire2372[(2'h3):(1'h0)] : (~&{(forvar2760 ?
                                  reg2416 : forvar2761)}));
                      reg2774 <= (!(-(reg2636[(1'h1):(1'h0)] | {forvar2407})));
                      reg2775 <= $unsigned({forvar2761});
                    end
                  else
                    begin
                      reg2773 <= ($unsigned((-forvar2597)) ?
                          $signed(reg2426[(1'h1):(1'h1)]) : forvar2621);
                      reg2774 <= (-(reg2580 >> {reg2587[(3'h6):(3'h6)]}));
                      reg2775 <= $unsigned(reg2757[(4'hc):(4'hc)]);
                      reg2776 <= reg2784[(4'hf):(2'h2)];
                    end
                  reg2777 <= ($signed((^~$signed((8'ha0)))) ?
                      ({(reg2651 >> (8'h9c))} > reg2487[(3'h7):(3'h4)]) : {((forvar2558 && reg2779) ?
                              reg2755[(4'h9):(3'h7)] : (+reg2675))});
                  for (forvar2778 = (1'h0); (forvar2778 < (2'h2)); forvar2778 = (forvar2778 + (1'h1)))
                    begin
                      reg2779 <= {{(8'had)}};
                      reg2780 <= wire2374[(1'h0):(1'h0)];
                      reg2781 <= $signed((&$unsigned((~reg2560))));
                      reg2782 <= ($unsigned(($unsigned(reg2714) ?
                              (forvar2628 && reg2523) : (reg2585 < forvar2389))) ?
                          ((-(!reg2510)) >> ((-reg2601) <= reg2491)) : $signed(reg2683));
                    end
                end
            end
          if (forvar2525[(3'h5):(3'h5)])
            begin
              for (forvar2783 = (1'h0); (forvar2783 < (1'h0)); forvar2783 = (forvar2783 + (1'h1)))
                begin
                  for (forvar2784 = (1'h0); (forvar2784 < (2'h3)); forvar2784 = (forvar2784 + (1'h1)))
                    begin
                      reg2785 <= $unsigned(forvar2544);
                      reg2786 <= reg2733[(3'h5):(3'h5)];
                      reg2787 <= (~reg2618);
                      reg2788 <= forvar2756[(1'h0):(1'h0)];
                    end
                  reg2789 <= $unsigned($signed($unsigned(reg2731[(2'h2):(1'h1)])));
                  for (forvar2790 = (1'h0); (forvar2790 < (2'h2)); forvar2790 = (forvar2790 + (1'h1)))
                    begin
                      reg2791 <= reg2760[(1'h1):(1'h0)];
                      reg2792 <= $signed(reg2747[(2'h2):(1'h0)]);
                    end
                  reg2793 <= {($unsigned($unsigned((8'h9f))) ?
                          $signed($signed(reg2711)) : ($signed((8'ha2)) ^~ reg2451))};
                end
            end
          else
            begin
              reg2783 <= (((reg2715 ^ (reg2646 ?
                  reg2637 : forvar2639)) || {reg2503}) < $unsigned((^~$signed(reg2464))));
              for (forvar2784 = (1'h0); (forvar2784 < (2'h2)); forvar2784 = (forvar2784 + (1'h1)))
                begin
                  for (forvar2785 = (1'h0); (forvar2785 < (2'h2)); forvar2785 = (forvar2785 + (1'h1)))
                    begin
                      reg2786 <= (($unsigned(forvar2516[(2'h2):(2'h2)]) * (reg2421[(2'h2):(1'h0)] ?
                              forvar2656[(3'h5):(3'h5)] : {wire2511})) ?
                          {{{reg2771}}} : ((8'h9c) ?
                              forvar2778 : forvar2516[(3'h6):(2'h3)]));
                      reg2787 <= {(~^$signed($unsigned((8'had))))};
                      reg2788 <= $signed((($unsigned(reg2675) ?
                              $signed(reg2465) : $signed((8'ha4))) ?
                          reg2495 : (~forvar2558)));
                    end
                  if (forvar2738)
                    begin
                      reg2789 <= forvar2790[(2'h2):(1'h0)];
                      reg2790 <= forvar2458;
                      reg2791 <= (((reg2718 ?
                          (forvar2739 >>> forvar2651) : ((8'hac) & reg2557)) | reg2542) * reg2684);
                    end
                  else
                    begin
                      reg2789 <= (forvar2616[(1'h1):(1'h0)] > (forvar2476[(3'h4):(3'h4)] - reg2662[(3'h6):(3'h6)]));
                    end
                  for (forvar2792 = (1'h0); (forvar2792 < (1'h1)); forvar2792 = (forvar2792 + (1'h1)))
                    begin
                      reg2793 <= $unsigned(forvar2728[(3'h4):(3'h4)]);
                    end
                end
              for (forvar2794 = (1'h0); (forvar2794 < (2'h3)); forvar2794 = (forvar2794 + (1'h1)))
                begin
                  if (reg2445)
                    begin
                      reg2795 <= ($signed(reg2650[(1'h0):(1'h0)]) || $unsigned({(reg2492 ?
                              (8'hac) : reg2657)}));
                      reg2796 <= reg2654;
                    end
                  else
                    begin
                      reg2795 <= ({$unsigned(((8'ha8) ^~ (8'h9f)))} ?
                          $signed($signed(reg2455[(1'h1):(1'h0)])) : wire2511[(4'hd):(2'h3)]);
                    end
                  if ($unsigned((((forvar2486 ^ reg2645) ?
                          $unsigned(reg2540) : (~&reg2498)) ?
                      $signed((|reg2489)) : ((forvar2767 ?
                              forvar2794 : reg2671) ?
                          $unsigned((8'hb9)) : $signed(forvar2475)))))
                    begin
                      reg2797 <= (~^forvar2524);
                    end
                  else
                    begin
                      reg2797 <= (($unsigned((^~reg2482)) && (|forvar2426[(2'h2):(1'h1)])) ?
                          ((8'ha9) + (((8'ha3) || reg2527) && $signed(reg2454))) : reg2428[(3'h5):(2'h3)]);
                      reg2798 <= ({((&reg2767) <<< reg2660)} ?
                          $signed(reg2459[(3'h5):(3'h4)]) : (reg2714[(4'h8):(2'h2)] != (^forvar2751)));
                    end
                end
              for (forvar2799 = (1'h0); (forvar2799 < (1'h0)); forvar2799 = (forvar2799 + (1'h1)))
                begin
                  for (forvar2800 = (1'h0); (forvar2800 < (2'h2)); forvar2800 = (forvar2800 + (1'h1)))
                    begin
                      reg2801 <= $signed(reg2713[(2'h2):(2'h2)]);
                    end
                  for (forvar2802 = (1'h0); (forvar2802 < (2'h3)); forvar2802 = (forvar2802 + (1'h1)))
                    begin
                      reg2803 <= reg2385[(2'h3):(1'h1)];
                      reg2804 <= reg2789;
                    end
                  if ((8'ha6))
                    begin
                      reg2805 <= ((8'haf) ?
                          $signed(forvar2516) : (~^$signed((~reg2527))));
                      reg2806 <= ({reg2645[(1'h1):(1'h1)]} * $unsigned($unsigned($unsigned(reg2605))));
                      reg2807 <= reg2567[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2805 <= reg2425;
                      reg2806 <= $signed(({(^~wire2377)} > (reg2480 >> (reg2721 && forvar2716))));
                      reg2807 <= ($unsigned((reg2410[(3'h7):(1'h1)] ?
                              $unsigned(reg2531) : (reg2641 * (8'ha0)))) ?
                          (8'ha2) : ((reg2541[(1'h1):(1'h0)] ?
                              $unsigned(reg2433) : $unsigned(forvar2720)) & $unsigned({reg2386})));
                      reg2808 <= reg2715[(3'h5):(2'h3)];
                    end
                  reg2809 <= {reg2648[(1'h1):(1'h0)]};
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2810 = (1'h0); (forvar2810 < (1'h0)); forvar2810 = (forvar2810 + (1'h1)))
        begin
          if ($unsigned($unsigned(($unsigned((8'ha9)) & {reg2574}))))
            begin
              for (forvar2811 = (1'h0); (forvar2811 < (1'h0)); forvar2811 = (forvar2811 + (1'h1)))
                begin
                  if (reg2465[(4'ha):(2'h2)])
                    begin
                      reg2812 <= $signed($unsigned($unsigned({forvar2761})));
                      reg2813 <= $unsigned((!$unsigned($unsigned(forvar2627))));
                      reg2814 <= ((~^reg2467) ?
                          reg2659 : (~^(^$signed(forvar2734))));
                      reg2815 <= (^~($signed((reg2721 << reg2443)) ?
                          ((^forvar2380) & reg2548[(4'he):(3'h7)]) : (reg2471 < forvar2783[(3'h7):(3'h4)])));
                    end
                  else
                    begin
                      reg2812 <= $unsigned(forvar2676);
                      reg2813 <= $signed((+(reg2671 ?
                          {forvar2601} : $unsigned(reg2807))));
                    end
                  for (forvar2816 = (1'h0); (forvar2816 < (2'h3)); forvar2816 = (forvar2816 + (1'h1)))
                    begin
                      reg2817 <= reg2542;
                      reg2818 <= $signed(forvar2703);
                      reg2819 <= (($signed(reg2469) ?
                          $signed((~&reg2388)) : wire2375[(3'h7):(3'h5)]) << {$signed($signed((8'hb5)))});
                    end
                end
              for (forvar2820 = (1'h0); (forvar2820 < (1'h0)); forvar2820 = (forvar2820 + (1'h1)))
                begin
                  for (forvar2821 = (1'h0); (forvar2821 < (2'h2)); forvar2821 = (forvar2821 + (1'h1)))
                    begin
                      reg2822 <= forvar2557[(1'h1):(1'h0)];
                    end
                  for (forvar2823 = (1'h0); (forvar2823 < (2'h3)); forvar2823 = (forvar2823 + (1'h1)))
                    begin
                      reg2824 <= {reg2772[(1'h0):(1'h0)]};
                    end
                  if ($signed(reg2762[(3'h4):(2'h3)]))
                    begin
                      reg2825 <= {(^~reg2578)};
                      reg2826 <= $signed($signed(reg2465));
                      reg2827 <= reg2554[(2'h2):(1'h1)];
                      reg2828 <= $unsigned(reg2518);
                    end
                  else
                    begin
                      reg2825 <= {((^~(forvar2564 * forvar2744)) <= reg2654)};
                      reg2826 <= $unsigned($signed(reg2441[(3'h7):(2'h2)]));
                      reg2827 <= $signed($signed(((reg2498 ?
                              reg2430 : (8'haa)) ?
                          $unsigned(reg2434) : (reg2707 ?
                              forvar2688 : (8'hab)))));
                      reg2828 <= reg2387[(1'h1):(1'h0)];
                    end
                  reg2829 <= (~|reg2793);
                end
              for (forvar2830 = (1'h0); (forvar2830 < (2'h2)); forvar2830 = (forvar2830 + (1'h1)))
                begin
                  for (forvar2831 = (1'h0); (forvar2831 < (1'h0)); forvar2831 = (forvar2831 + (1'h1)))
                    begin
                      reg2832 <= $signed(((&reg2700) ?
                          $unsigned($signed(forvar2426)) : reg2392));
                    end
                  if ({(^~(~|reg2598[(2'h3):(2'h2)]))})
                    begin
                      reg2833 <= (|(($signed(reg2698) || {reg2539}) ?
                          $signed($unsigned(forvar2598)) : $signed({reg2391})));
                      reg2834 <= reg2474;
                      reg2835 <= ($unsigned(($unsigned(reg2727) <<< {reg2654})) ~^ reg2813);
                    end
                  else
                    begin
                      reg2833 <= $signed(reg2817[(1'h1):(1'h1)]);
                    end
                  reg2836 <= forvar2628;
                end
              for (forvar2837 = (1'h0); (forvar2837 < (2'h2)); forvar2837 = (forvar2837 + (1'h1)))
                begin
                  reg2838 <= {forvar2465[(1'h0):(1'h0)]};
                end
            end
          else
            begin
              if ((^~reg2793[(2'h2):(1'h1)]))
                begin
                  for (forvar2811 = (1'h0); (forvar2811 < (1'h0)); forvar2811 = (forvar2811 + (1'h1)))
                    begin
                      reg2812 <= reg2616;
                      reg2813 <= $signed($signed((~|$signed((8'hb7)))));
                      reg2814 <= {$signed($unsigned(reg2537))};
                      reg2815 <= $signed((($unsigned(wire2372) && $unsigned(reg2439)) ?
                          ((+(8'h9d)) >= (reg2509 ?
                              reg2546 : forvar2527)) : forvar2785));
                    end
                  if (forvar2577[(2'h3):(1'h1)])
                    begin
                      reg2816 <= $signed(reg2510);
                      reg2817 <= ((|reg2630[(4'he):(2'h3)]) != ($unsigned((8'haf)) ?
                          ((reg2710 ? reg2538 : reg2782) ?
                              $signed((8'hba)) : (reg2438 > reg2819)) : $unsigned(reg2569)));
                      reg2818 <= reg2392;
                      reg2819 <= $signed((($signed(reg2604) >= (~reg2456)) == forvar2752));
                    end
                  else
                    begin
                      reg2816 <= forvar2489[(1'h0):(1'h0)];
                    end
                  for (forvar2820 = (1'h0); (forvar2820 < (1'h1)); forvar2820 = (forvar2820 + (1'h1)))
                    begin
                      reg2821 <= ((($signed((8'hb0)) ?
                              $unsigned(reg2520) : reg2721[(2'h2):(2'h2)]) && (|$unsigned(reg2430))) ?
                          reg2462 : ((~^$unsigned(reg2724)) ?
                              $signed(reg2687) : forvar2678));
                      reg2822 <= ($signed($unsigned($unsigned(reg2527))) ?
                          $signed(wire2372) : (((reg2663 == forvar2683) <= (reg2408 & reg2718)) == $signed(reg2662[(3'h6):(3'h6)])));
                      reg2823 <= $unsigned(forvar2394);
                    end
                end
              else
                begin
                  for (forvar2811 = (1'h0); (forvar2811 < (2'h3)); forvar2811 = (forvar2811 + (1'h1)))
                    begin
                      reg2812 <= (~^$signed(((~reg2771) ?
                          forvar2830 : (forvar2656 ? reg2567 : (8'hb2)))));
                    end
                end
              for (forvar2824 = (1'h0); (forvar2824 < (1'h1)); forvar2824 = (forvar2824 + (1'h1)))
                begin
                  reg2825 <= reg2633[(4'hb):(4'h8)];
                  if ($signed($unsigned($signed((|forvar2486)))))
                    begin
                      reg2826 <= {($signed({forvar2536}) ?
                              ((8'h9e) && reg2630) : forvar2734)};
                      reg2827 <= reg2822;
                    end
                  else
                    begin
                      reg2826 <= {{(reg2756[(1'h0):(1'h0)] - {reg2425})}};
                      reg2827 <= $unsigned($unsigned(({reg2731} ^~ {reg2660})));
                      reg2828 <= (~^$unsigned(($signed(reg2428) ?
                          reg2693 : reg2757[(2'h2):(2'h2)])));
                    end
                end
            end
          for (forvar2839 = (1'h0); (forvar2839 < (1'h1)); forvar2839 = (forvar2839 + (1'h1)))
            begin
              for (forvar2840 = (1'h0); (forvar2840 < (2'h2)); forvar2840 = (forvar2840 + (1'h1)))
                begin
                  for (forvar2841 = (1'h0); (forvar2841 < (1'h0)); forvar2841 = (forvar2841 + (1'h1)))
                    begin
                      reg2842 <= $signed(($signed($signed(forvar2697)) ?
                          (~^((8'ha0) ?
                              reg2544 : reg2460)) : ($signed((8'hb1)) ?
                              reg2561[(4'h8):(1'h0)] : (8'hab))));
                      reg2843 <= (&(~^(forvar2380 ?
                          $signed((8'hab)) : $unsigned((8'hab)))));
                      reg2844 <= reg2832;
                      reg2845 <= reg2476[(3'h5):(1'h0)];
                    end
                  reg2846 <= reg2457[(2'h3):(1'h1)];
                end
              for (forvar2847 = (1'h0); (forvar2847 < (1'h0)); forvar2847 = (forvar2847 + (1'h1)))
                begin
                  for (forvar2848 = (1'h0); (forvar2848 < (2'h3)); forvar2848 = (forvar2848 + (1'h1)))
                    begin
                      reg2849 <= $signed({((reg2774 ?
                              reg2502 : (8'ha3)) >>> (forvar2785 < forvar2486))});
                      reg2850 <= forvar2611;
                      reg2851 <= forvar2760;
                    end
                end
              if ((!(^$unsigned(reg2460[(4'ha):(3'h6)]))))
                begin
                  for (forvar2852 = (1'h0); (forvar2852 < (2'h3)); forvar2852 = (forvar2852 + (1'h1)))
                    begin
                      reg2853 <= (8'hb0);
                    end
                  if (reg2771[(2'h2):(1'h0)])
                    begin
                      reg2854 <= ((reg2717[(2'h2):(1'h0)] ?
                          reg2677 : (~&(reg2843 ^ forvar2600))) >= ((8'h9f) ?
                          $signed((8'hb4)) : reg2452));
                      reg2855 <= reg2430;
                      reg2856 <= (reg2659 != ((8'hb3) > $unsigned({reg2829})));
                    end
                  else
                    begin
                      reg2854 <= $unsigned($signed($signed($unsigned((8'hb0)))));
                    end
                  reg2857 <= $unsigned((~^$unsigned((reg2612 ?
                      reg2615 : forvar2406))));
                end
              else
                begin
                  reg2852 <= reg2682[(1'h1):(1'h0)];
                  for (forvar2853 = (1'h0); (forvar2853 < (2'h3)); forvar2853 = (forvar2853 + (1'h1)))
                    begin
                      reg2854 <= ($unsigned($signed(reg2785)) & (($signed(forvar2751) & (forvar2677 >>> reg2521)) ?
                          $unsigned((~&reg2651)) : (~|$signed(reg2790))));
                      reg2855 <= (~^($unsigned((~&forvar2544)) * ($signed((8'hb4)) < $signed(forvar2820))));
                      reg2856 <= reg2599;
                      reg2857 <= (^(($unsigned(reg2784) ?
                              reg2763[(2'h2):(1'h1)] : (forvar2394 ?
                                  forvar2639 : reg2508)) ?
                          $signed($signed(reg2507)) : ((reg2480 && forvar2521) ?
                              forvar2787[(1'h1):(1'h1)] : ((8'ha8) ?
                                  reg2443 : forvar2739))));
                    end
                end
              for (forvar2858 = (1'h0); (forvar2858 < (1'h1)); forvar2858 = (forvar2858 + (1'h1)))
                begin
                  if ((^forvar2687))
                    begin
                      reg2859 <= ($unsigned({(forvar2800 - reg2570)}) ?
                          reg2481 : (8'ha0));
                    end
                  else
                    begin
                      reg2859 <= $signed($signed(((|reg2835) << {forvar2703})));
                      reg2860 <= (^~(($unsigned((8'hb8)) <<< (forvar2671 || reg2485)) ?
                          forvar2746[(2'h2):(2'h2)] : reg2795[(1'h1):(1'h0)]));
                      reg2861 <= forvar2381;
                      reg2862 <= $unsigned((&forvar2702));
                    end
                  for (forvar2863 = (1'h0); (forvar2863 < (1'h1)); forvar2863 = (forvar2863 + (1'h1)))
                    begin
                      reg2864 <= reg2679[(2'h2):(1'h1)];
                      reg2865 <= reg2720;
                    end
                  for (forvar2866 = (1'h0); (forvar2866 < (1'h1)); forvar2866 = (forvar2866 + (1'h1)))
                    begin
                      reg2867 <= ($unsigned((8'hac)) ?
                          {reg2472} : $unsigned(reg2518[(3'h4):(1'h0)]));
                      reg2868 <= $signed(reg2383);
                      reg2869 <= $unsigned(reg2592[(2'h2):(2'h2)]);
                      reg2870 <= reg2438[(4'hb):(4'h8)];
                    end
                end
            end
          reg2871 <= reg2836;
          if ($unsigned(forvar2802[(2'h2):(1'h1)]))
            begin
              for (forvar2872 = (1'h0); (forvar2872 < (1'h0)); forvar2872 = (forvar2872 + (1'h1)))
                begin
                  for (forvar2873 = (1'h0); (forvar2873 < (1'h0)); forvar2873 = (forvar2873 + (1'h1)))
                    begin
                      reg2874 <= $unsigned({({(8'ha1)} + forvar2694)});
                      reg2875 <= (+$signed({$signed(reg2714)}));
                      reg2876 <= (8'h9e);
                      reg2877 <= (8'hb7);
                    end
                  if ($unsigned((($unsigned(reg2427) ?
                          (reg2579 * reg2828) : reg2783[(3'h4):(1'h0)]) ?
                      $signed(forvar2506[(4'hb):(2'h2)]) : reg2544[(4'hd):(4'h9)])))
                    begin
                      reg2878 <= (!$unsigned(((~|reg2617) >= ((8'h9f) ?
                          reg2819 : forvar2721))));
                      reg2879 <= reg2587;
                    end
                  else
                    begin
                      reg2878 <= forvar2694[(2'h2):(2'h2)];
                      reg2879 <= reg2790;
                    end
                  if ((((~forvar2442[(2'h2):(1'h1)]) & (^~forvar2656)) ?
                      ({reg2774[(2'h2):(2'h2)]} > ((^forvar2651) + (&reg2867))) : (8'hb0)))
                    begin
                      reg2880 <= (wire2514[(2'h3):(2'h2)] < (reg2441 && (reg2670[(1'h1):(1'h0)] ?
                          (forvar2666 ?
                              reg2824 : forvar2823) : $signed(reg2808))));
                    end
                  else
                    begin
                      reg2880 <= ($unsigned($unsigned(reg2815[(2'h2):(2'h2)])) ?
                          $unsigned((~|((8'h9f) & reg2555))) : $unsigned($signed($signed(reg2618))));
                    end
                  for (forvar2881 = (1'h0); (forvar2881 < (1'h1)); forvar2881 = (forvar2881 + (1'h1)))
                    begin
                      reg2882 <= ($signed((~^{reg2665})) <<< $signed((reg2761[(2'h2):(1'h1)] ?
                          (reg2746 ? reg2686 : (8'ha6)) : (reg2852 ?
                              reg2853 : forvar2693))));
                      reg2883 <= $unsigned({($signed(reg2579) ?
                              (reg2599 >> reg2481) : forvar2527[(4'hd):(4'hc)])});
                      reg2884 <= reg2659;
                      reg2885 <= $signed((~^reg2812[(2'h2):(1'h1)]));
                    end
                end
            end
          else
            begin
              reg2872 <= (-((reg2694[(1'h1):(1'h1)] ?
                  reg2755[(2'h2):(1'h1)] : (~^forvar2380)) ^~ reg2532[(3'h6):(2'h3)]));
            end
        end
      if (reg2522[(1'h0):(1'h0)])
        begin
          reg2886 <= ((forvar2552[(4'h8):(3'h6)] + {(reg2652 ~^ reg2705)}) ?
              $signed(forvar2785[(1'h0):(1'h0)]) : (((reg2568 ?
                      reg2588 : reg2483) - $unsigned(reg2861)) ?
                  {reg2481} : (forvar2381 >> reg2593[(2'h3):(1'h1)])));
          for (forvar2887 = (1'h0); (forvar2887 < (1'h1)); forvar2887 = (forvar2887 + (1'h1)))
            begin
              for (forvar2888 = (1'h0); (forvar2888 < (1'h0)); forvar2888 = (forvar2888 + (1'h1)))
                begin
                  if ((reg2718[(2'h3):(2'h3)] ?
                      (($unsigned(reg2681) ?
                              (~&forvar2872) : wire2514[(4'h8):(1'h0)]) ?
                          $unsigned(reg2599[(1'h0):(1'h0)]) : reg2582[(1'h1):(1'h0)]) : {$signed({(8'hba)})}))
                    begin
                      reg2889 <= (^$signed(forvar2545));
                    end
                  else
                    begin
                      reg2889 <= (^~$unsigned(reg2699));
                      reg2890 <= (reg2625 || $signed(((8'ha1) ?
                          reg2452 : $unsigned(reg2544))));
                      reg2891 <= {((reg2552[(1'h0):(1'h0)] ?
                                  $signed(reg2654) : (8'hb2)) ?
                              reg2517 : $unsigned($unsigned((8'ha9))))};
                    end
                end
            end
          for (forvar2892 = (1'h0); (forvar2892 < (2'h3)); forvar2892 = (forvar2892 + (1'h1)))
            begin
              reg2893 <= (reg2433 * $unsigned(((-reg2642) >= $unsigned((8'had)))));
              for (forvar2894 = (1'h0); (forvar2894 < (1'h1)); forvar2894 = (forvar2894 + (1'h1)))
                begin
                  for (forvar2895 = (1'h0); (forvar2895 < (1'h1)); forvar2895 = (forvar2895 + (1'h1)))
                    begin
                      reg2896 <= reg2843[(3'h5):(1'h1)];
                      reg2897 <= $signed(reg2857[(1'h0):(1'h0)]);
                      reg2898 <= {reg2619[(4'he):(4'h8)]};
                    end
                  reg2899 <= forvar2396;
                  for (forvar2900 = (1'h0); (forvar2900 < (1'h1)); forvar2900 = (forvar2900 + (1'h1)))
                    begin
                      reg2901 <= $signed(reg2674);
                      reg2902 <= (reg2481 + $signed($unsigned($unsigned(forvar2703))));
                    end
                  if ((^$unsigned($signed((reg2658 ?
                      forvar2651 : forvar2680)))))
                    begin
                      reg2903 <= (($signed((forvar2763 | reg2590)) ?
                          reg2463 : (reg2509[(3'h4):(2'h3)] ?
                              (~(8'hb6)) : $signed(reg2489))) | forvar2784[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg2903 <= $unsigned($unsigned($signed($unsigned((8'ha8)))));
                      reg2904 <= (|(forvar2536[(2'h2):(1'h1)] ?
                          $signed((!forvar2773)) : (!{(8'ha8)})));
                    end
                end
              for (forvar2905 = (1'h0); (forvar2905 < (2'h3)); forvar2905 = (forvar2905 + (1'h1)))
                begin
                  reg2906 <= (+$unsigned(reg2432[(3'h4):(1'h0)]));
                  for (forvar2907 = (1'h0); (forvar2907 < (1'h1)); forvar2907 = (forvar2907 + (1'h1)))
                    begin
                      reg2908 <= ({(8'hac)} == ((+$signed(reg2710)) ?
                          reg2849[(3'h4):(3'h4)] : reg2757[(1'h0):(1'h0)]));
                    end
                  for (forvar2909 = (1'h0); (forvar2909 < (2'h2)); forvar2909 = (forvar2909 + (1'h1)))
                    begin
                      reg2910 <= $unsigned($signed((reg2797 | {reg2844})));
                      reg2911 <= ((reg2814[(2'h2):(1'h1)] <<< ((+reg2552) ?
                          {wire2512} : forvar2716[(3'h4):(2'h2)])) | reg2801[(1'h0):(1'h0)]);
                      reg2912 <= reg2609[(2'h3):(2'h2)];
                    end
                end
            end
        end
      else
        begin
          if (forvar2435[(4'h9):(3'h7)])
            begin
              if ($unsigned($signed((reg2702 ^~ $signed(reg2859)))))
                begin
                  if (forvar2435)
                    begin
                      reg2886 <= $unsigned((^reg2791[(2'h3):(1'h0)]));
                      reg2887 <= (reg2843 ?
                          {reg2425[(4'h9):(3'h6)]} : (+((wire2377 ^ (8'haa)) << (reg2872 | reg2727))));
                      reg2888 <= ({$signed((forvar2473 ?
                              reg2561 : reg2495))} * {$unsigned({(8'hb0)})});
                      reg2889 <= forvar2799[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg2886 <= $unsigned($unsigned(forvar2694));
                    end
                  for (forvar2890 = (1'h0); (forvar2890 < (1'h1)); forvar2890 = (forvar2890 + (1'h1)))
                    begin
                      reg2891 <= {$unsigned(forvar2753[(2'h2):(1'h1)])};
                      reg2892 <= reg2677;
                      reg2893 <= (((^~{forvar2785}) ?
                          ($unsigned(reg2696) ?
                              $unsigned(forvar2892) : (8'ha2)) : ($signed((8'ha9)) | reg2537[(3'h6):(3'h4)])) < (^reg2508));
                    end
                end
              else
                begin
                  for (forvar2886 = (1'h0); (forvar2886 < (2'h3)); forvar2886 = (forvar2886 + (1'h1)))
                    begin
                      reg2887 <= (8'hb0);
                      reg2888 <= $signed(wire2378[(3'h4):(1'h1)]);
                      reg2889 <= $signed({$signed((^~forvar2784))});
                    end
                  for (forvar2890 = (1'h0); (forvar2890 < (1'h0)); forvar2890 = (forvar2890 + (1'h1)))
                    begin
                      reg2891 <= (reg2547 ?
                          (((^~reg2619) < (reg2879 ? forvar2601 : (8'ha1))) ?
                              reg2843[(3'h4):(2'h2)] : $signed($unsigned(reg2849))) : $signed((reg2711[(3'h4):(1'h0)] > (8'hba))));
                      reg2892 <= ((($signed(forvar2799) <= {wire2376}) ^~ (^{(8'hb9)})) ?
                          $unsigned(((8'ha9) ^~ reg2519[(2'h3):(2'h3)])) : (~&((|reg2430) != (reg2416 && forvar2379))));
                      reg2893 <= (~|(~&(forvar2593[(3'h5):(2'h3)] | reg2414[(4'h8):(1'h1)])));
                    end
                end
              for (forvar2894 = (1'h0); (forvar2894 < (1'h1)); forvar2894 = (forvar2894 + (1'h1)))
                begin
                  if ({$unsigned(reg2706[(3'h4):(3'h4)])})
                    begin
                      reg2895 <= $unsigned((~|{(^~reg2559)}));
                      reg2896 <= $unsigned(reg2648);
                      reg2897 <= forvar2394[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2895 <= {reg2552};
                      reg2896 <= reg2720;
                      reg2897 <= $signed((~|($signed(forvar2785) | {forvar2716})));
                    end
                  for (forvar2898 = (1'h0); (forvar2898 < (1'h0)); forvar2898 = (forvar2898 + (1'h1)))
                    begin
                      reg2899 <= $unsigned((~&$signed(reg2836[(3'h5):(3'h5)])));
                      reg2900 <= (forvar2629 ?
                          $unsigned(((reg2885 ? reg2635 : wire2511) ?
                              (+forvar2753) : $signed(reg2604))) : reg2807);
                    end
                end
            end
          else
            begin
              for (forvar2886 = (1'h0); (forvar2886 < (2'h2)); forvar2886 = (forvar2886 + (1'h1)))
                begin
                  for (forvar2887 = (1'h0); (forvar2887 < (2'h3)); forvar2887 = (forvar2887 + (1'h1)))
                    begin
                      reg2888 <= forvar2824[(2'h3):(1'h0)];
                      reg2889 <= forvar2611[(2'h2):(1'h1)];
                      reg2890 <= $unsigned($signed({$unsigned(reg2433)}));
                    end
                  if ($signed($signed($unsigned(reg2509[(3'h7):(1'h0)]))))
                    begin
                      reg2891 <= reg2659;
                      reg2892 <= (^~reg2561);
                      reg2893 <= (($unsigned((reg2777 > reg2707)) ?
                          (~|reg2599) : (&(reg2654 ?
                              reg2776 : wire2374))) <= reg2477);
                    end
                  else
                    begin
                      reg2891 <= (reg2756 >= forvar2409);
                      reg2892 <= ((8'hac) | $unsigned(reg2475));
                      reg2893 <= (^$signed($unsigned(((8'ha9) << reg2575))));
                    end
                  for (forvar2894 = (1'h0); (forvar2894 < (2'h2)); forvar2894 = (forvar2894 + (1'h1)))
                    begin
                      reg2895 <= (^(~^{reg2505[(1'h0):(1'h0)]}));
                      reg2896 <= (reg2595[(2'h2):(2'h2)] > (($signed(reg2555) ?
                              (8'haf) : reg2708[(1'h1):(1'h1)]) ?
                          ($signed(reg2727) || $unsigned(reg2717)) : (8'ha1)));
                      reg2897 <= ($signed(($unsigned(reg2732) ?
                              $unsigned(reg2559) : forvar2612)) ?
                          ($unsigned((^forvar2656)) <<< {$unsigned(forvar2527)}) : (8'hb8));
                    end
                  for (forvar2898 = (1'h0); (forvar2898 < (1'h0)); forvar2898 = (forvar2898 + (1'h1)))
                    begin
                      reg2899 <= ($unsigned(forvar2738[(2'h3):(1'h1)]) ?
                          {reg2686[(1'h1):(1'h1)]} : reg2637);
                      reg2900 <= reg2525[(3'h7):(1'h1)];
                      reg2901 <= reg2557[(3'h4):(3'h4)];
                      reg2902 <= ($signed(reg2812[(4'h9):(1'h1)]) >> $unsigned($unsigned($unsigned(reg2642))));
                    end
                end
            end
          for (forvar2903 = (1'h0); (forvar2903 < (1'h0)); forvar2903 = (forvar2903 + (1'h1)))
            begin
              reg2904 <= {(+{$signed(reg2618)})};
              for (forvar2905 = (1'h0); (forvar2905 < (1'h0)); forvar2905 = (forvar2905 + (1'h1)))
                begin
                  for (forvar2906 = (1'h0); (forvar2906 < (2'h3)); forvar2906 = (forvar2906 + (1'h1)))
                    begin
                      reg2907 <= $signed(forvar2601[(2'h3):(2'h2)]);
                      reg2908 <= forvar2401;
                    end
                  reg2909 <= (!reg2566[(2'h3):(1'h0)]);
                  reg2910 <= reg2579[(2'h2):(2'h2)];
                  if (forvar2702[(4'hc):(3'h4)])
                    begin
                      reg2911 <= reg2619;
                    end
                  else
                    begin
                      reg2911 <= $signed($unsigned($unsigned(forvar2756)));
                    end
                end
              for (forvar2912 = (1'h0); (forvar2912 < (2'h2)); forvar2912 = (forvar2912 + (1'h1)))
                begin
                  for (forvar2913 = (1'h0); (forvar2913 < (2'h2)); forvar2913 = (forvar2913 + (1'h1)))
                    begin
                      reg2914 <= ((|$unsigned({reg2483})) <= ($unsigned($signed((8'ha3))) ?
                          (wire2378[(2'h2):(1'h0)] ?
                              (reg2708 | forvar2821) : ((8'h9d) == forvar2824)) : (!reg2664)));
                      reg2915 <= $signed($unsigned($signed((reg2556 ?
                          reg2382 : forvar2703))));
                    end
                end
            end
        end
      reg2916 <= (wire2372[(3'h4):(3'h4)] ?
          $signed((forvar2616 + (~forvar2506))) : $unsigned($unsigned((+reg2533))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3117  (y, clk, wire3122, wire3121, wire3120, wire3119, wire3118);
  output wire [(32'ha0a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire3122;
  input wire [(4'hd):(1'h0)] wire3121;
  input wire [(4'he):(1'h0)] wire3120;
  input wire [(3'h4):(1'h0)] wire3119;
  input wire [(4'hd):(1'h0)] wire3118;
  reg signed [(3'h6):(1'h0)] reg3365 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3364 = (1'h0);
  reg [(4'he):(1'h0)] reg3363 = (1'h0);
  reg [(4'hc):(1'h0)] reg3362 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3361 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3360 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3357 = (1'h0);
  reg [(4'hc):(1'h0)] reg3353 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3350 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3345 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3342 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3338 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3359 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3358 = (1'h0);
  reg [(3'h5):(1'h0)] reg3357 = (1'h0);
  reg [(5'h10):(1'h0)] reg3356 = (1'h0);
  reg [(4'ha):(1'h0)] reg3355 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3354 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3353 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3352 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3351 = (1'h0);
  reg [(4'he):(1'h0)] reg3350 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3349 = (1'h0);
  reg [(3'h4):(1'h0)] reg3348 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3347 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3346 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3345 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3344 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3343 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3342 = (1'h0);
  reg [(4'hf):(1'h0)] reg3341 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3340 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3339 = (1'h0);
  reg [(4'ha):(1'h0)] reg3338 = (1'h0);
  reg [(4'hc):(1'h0)] reg3337 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3336 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3335 = (1'h0);
  reg [(4'h8):(1'h0)] reg3334 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3333 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3332 = (1'h0);
  reg [(4'hf):(1'h0)] reg3331 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3330 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3329 = (1'h0);
  reg [(4'h9):(1'h0)] reg3328 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3327 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3326 = (1'h0);
  reg [(2'h2):(1'h0)] reg3325 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3324 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3323 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3323 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3322 = (1'h0);
  reg [(3'h4):(1'h0)] reg3321 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3320 = (1'h0);
  reg [(3'h4):(1'h0)] reg3319 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3318 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3317 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3316 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3315 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3314 = (1'h0);
  reg [(3'h6):(1'h0)] reg3313 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3312 = (1'h0);
  reg [(4'hd):(1'h0)] reg3311 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3310 = (1'h0);
  reg [(3'h5):(1'h0)] reg3309 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3308 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3307 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3306 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3305 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3304 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3303 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3302 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3301 = (1'h0);
  reg [(4'hb):(1'h0)] reg3300 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3299 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3298 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3297 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3294 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3291 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3296 = (1'h0);
  reg [(2'h3):(1'h0)] reg3295 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3294 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3293 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3292 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3291 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3290 = (1'h0);
  reg [(3'h7):(1'h0)] reg3289 = (1'h0);
  reg [(4'h8):(1'h0)] reg3288 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3287 = (1'h0);
  reg [(4'h8):(1'h0)] reg3286 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3285 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3284 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3283 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3282 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire3281;
  reg [(5'h10):(1'h0)] reg3280 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3279 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3278 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3277 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3276 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3275 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3274 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3273 = (1'h0);
  reg [(2'h3):(1'h0)] reg3272 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3271 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3270 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3269 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3267 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3266 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3265 = (1'h0);
  reg [(4'he):(1'h0)] reg3264 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3258 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3263 = (1'h0);
  reg [(4'he):(1'h0)] forvar3262 = (1'h0);
  reg [(4'h9):(1'h0)] reg3261 = (1'h0);
  reg [(3'h6):(1'h0)] reg3260 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3259 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3258 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3255 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3253 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3252 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3249 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3245 = (1'h0);
  reg [(4'hd):(1'h0)] reg3257 = (1'h0);
  reg [(2'h3):(1'h0)] reg3256 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3255 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3254 = (1'h0);
  reg [(4'h8):(1'h0)] reg3253 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3252 = (1'h0);
  reg [(2'h3):(1'h0)] reg3251 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3250 = (1'h0);
  reg [(4'he):(1'h0)] reg3249 = (1'h0);
  reg [(3'h5):(1'h0)] reg3248 = (1'h0);
  reg [(3'h7):(1'h0)] reg3247 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3246 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3245 = (1'h0);
  reg [(4'h8):(1'h0)] reg3244 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3243 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3242 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3241 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3240 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3239 = (1'h0);
  reg [(4'he):(1'h0)] forvar3238 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3237 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3236 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3235 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3234 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3233 = (1'h0);
  reg [(3'h4):(1'h0)] reg3232 = (1'h0);
  reg [(2'h3):(1'h0)] reg3231 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3230 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3229 = (1'h0);
  reg [(3'h6):(1'h0)] reg3228 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3227 = (1'h0);
  reg [(5'h10):(1'h0)] reg3226 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3225 = (1'h0);
  reg [(2'h2):(1'h0)] reg3224 = (1'h0);
  reg [(4'hb):(1'h0)] reg3223 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3222 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3221 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3220 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3192 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3190 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3184 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3173 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3172 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3170 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3164 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3162 = (1'h0);
  reg [(4'hf):(1'h0)] reg3159 = (1'h0);
  reg [(3'h4):(1'h0)] reg3219 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3218 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3217 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3216 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3215 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3214 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3206 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3205 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3213 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3195 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3191 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3188 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3187 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3212 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3211 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3210 = (1'h0);
  reg [(4'hb):(1'h0)] reg3209 = (1'h0);
  reg [(4'hd):(1'h0)] reg3208 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3207 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3206 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3205 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3197 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3204 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3202 = (1'h0);
  reg [(3'h7):(1'h0)] reg3201 = (1'h0);
  reg [(3'h7):(1'h0)] reg3200 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3199 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3198 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3197 = (1'h0);
  reg [(4'hc):(1'h0)] reg3196 = (1'h0);
  reg [(5'h10):(1'h0)] reg3195 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3194 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3193 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3192 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3191 = (1'h0);
  reg [(4'h9):(1'h0)] reg3190 = (1'h0);
  reg [(5'h10):(1'h0)] reg3189 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3188 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3187 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3186 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3185 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3184 = (1'h0);
  reg [(4'hf):(1'h0)] reg3183 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3182 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3181 = (1'h0);
  reg [(4'ha):(1'h0)] reg3179 = (1'h0);
  reg [(2'h2):(1'h0)] reg3180 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3179 = (1'h0);
  reg [(4'hf):(1'h0)] reg3178 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3169 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3177 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3176 = (1'h0);
  reg [(2'h2):(1'h0)] reg3175 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3174 = (1'h0);
  reg [(3'h5):(1'h0)] reg3173 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3172 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3171 = (1'h0);
  reg [(3'h7):(1'h0)] reg3170 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3169 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3168 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3167 = (1'h0);
  reg [(4'he):(1'h0)] reg3166 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3165 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3164 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3163 = (1'h0);
  reg [(4'hf):(1'h0)] reg3162 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3161 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3157 = (1'h0);
  reg [(4'he):(1'h0)] reg3160 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3159 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3158 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3157 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3156 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3142 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3139 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3134 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3124 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3155 = (1'h0);
  reg [(3'h5):(1'h0)] reg3154 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3153 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3152 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3151 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3150 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3147 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3144 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3143 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3140 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3138 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3137 = (1'h0);
  reg [(3'h4):(1'h0)] reg3132 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3131 = (1'h0);
  reg [(4'ha):(1'h0)] reg3129 = (1'h0);
  reg [(3'h6):(1'h0)] reg3125 = (1'h0);
  reg [(3'h6):(1'h0)] reg3149 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3148 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3147 = (1'h0);
  reg [(4'hb):(1'h0)] reg3146 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3145 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3144 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3143 = (1'h0);
  reg [(3'h4):(1'h0)] reg3142 = (1'h0);
  reg [(4'ha):(1'h0)] reg3141 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3140 = (1'h0);
  reg [(4'hd):(1'h0)] reg3139 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3138 = (1'h0);
  reg [(5'h10):(1'h0)] reg3137 = (1'h0);
  reg [(5'h10):(1'h0)] reg3136 = (1'h0);
  reg [(3'h6):(1'h0)] reg3135 = (1'h0);
  reg [(3'h5):(1'h0)] reg3134 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3133 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3132 = (1'h0);
  reg [(4'hf):(1'h0)] reg3131 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3130 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3129 = (1'h0);
  reg [(3'h7):(1'h0)] reg3128 = (1'h0);
  reg [(4'he):(1'h0)] reg3127 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3126 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3125 = (1'h0);
  reg [(4'he):(1'h0)] reg3124 = (1'h0);
  reg [(3'h6):(1'h0)] reg3123 = (1'h0);
  assign y = {reg3365,
                 reg3364,
                 reg3363,
                 reg3362,
                 reg3361,
                 reg3360,
                 forvar3357,
                 reg3353,
                 forvar3350,
                 reg3345,
                 reg3342,
                 forvar3338,
                 reg3359,
                 reg3358,
                 reg3357,
                 reg3356,
                 reg3355,
                 reg3354,
                 forvar3353,
                 reg3352,
                 reg3351,
                 reg3350,
                 reg3349,
                 reg3348,
                 reg3347,
                 reg3346,
                 forvar3345,
                 reg3344,
                 reg3343,
                 forvar3342,
                 reg3341,
                 reg3340,
                 reg3339,
                 reg3338,
                 reg3337,
                 reg3336,
                 reg3335,
                 reg3334,
                 forvar3333,
                 forvar3332,
                 reg3331,
                 reg3330,
                 forvar3329,
                 reg3328,
                 reg3327,
                 reg3326,
                 reg3325,
                 reg3324,
                 forvar3323,
                 reg3323,
                 forvar3322,
                 reg3321,
                 reg3320,
                 reg3319,
                 reg3318,
                 forvar3317,
                 reg3316,
                 reg3315,
                 reg3314,
                 reg3313,
                 forvar3312,
                 reg3311,
                 forvar3310,
                 reg3309,
                 forvar3308,
                 forvar3307,
                 reg3306,
                 reg3305,
                 reg3304,
                 forvar3303,
                 reg3302,
                 reg3301,
                 reg3300,
                 reg3299,
                 forvar3298,
                 forvar3297,
                 reg3294,
                 forvar3291,
                 reg3296,
                 reg3295,
                 forvar3294,
                 reg3293,
                 reg3292,
                 reg3291,
                 forvar3290,
                 reg3289,
                 reg3288,
                 reg3287,
                 reg3286,
                 forvar3285,
                 forvar3284,
                 forvar3283,
                 reg3282,
                 wire3281,
                 reg3280,
                 reg3279,
                 reg3278,
                 forvar3277,
                 reg3276,
                 reg3275,
                 reg3274,
                 reg3273,
                 reg3272,
                 forvar3271,
                 reg3270,
                 reg3269,
                 reg3268,
                 reg3267,
                 forvar3266,
                 forvar3265,
                 reg3264,
                 forvar3258,
                 reg3263,
                 forvar3262,
                 reg3261,
                 reg3260,
                 reg3259,
                 reg3258,
                 reg3255,
                 forvar3253,
                 reg3252,
                 forvar3249,
                 forvar3245,
                 reg3257,
                 reg3256,
                 forvar3255,
                 reg3254,
                 reg3253,
                 forvar3252,
                 reg3251,
                 reg3250,
                 reg3249,
                 reg3248,
                 reg3247,
                 reg3246,
                 reg3245,
                 reg3244,
                 forvar3243,
                 reg3242,
                 reg3241,
                 reg3240,
                 reg3239,
                 forvar3238,
                 reg3237,
                 reg3236,
                 reg3235,
                 forvar3234,
                 reg3233,
                 reg3232,
                 reg3231,
                 reg3230,
                 forvar3229,
                 reg3228,
                 reg3227,
                 reg3226,
                 forvar3225,
                 reg3224,
                 reg3223,
                 forvar3222,
                 forvar3221,
                 forvar3220,
                 reg3192,
                 forvar3190,
                 forvar3184,
                 forvar3173,
                 forvar3172,
                 forvar3170,
                 reg3164,
                 forvar3162,
                 reg3159,
                 reg3219,
                 reg3218,
                 reg3217,
                 reg3216,
                 forvar3215,
                 forvar3214,
                 forvar3206,
                 reg3205,
                 reg3213,
                 forvar3195,
                 reg3191,
                 forvar3188,
                 forvar3187,
                 reg3212,
                 reg3211,
                 reg3210,
                 reg3209,
                 reg3208,
                 reg3207,
                 reg3206,
                 forvar3205,
                 forvar3197,
                 reg3204,
                 reg3203,
                 reg3202,
                 reg3201,
                 reg3200,
                 reg3199,
                 reg3198,
                 reg3197,
                 reg3196,
                 reg3195,
                 reg3194,
                 reg3193,
                 forvar3192,
                 forvar3191,
                 reg3190,
                 reg3189,
                 reg3188,
                 reg3187,
                 reg3186,
                 reg3185,
                 reg3184,
                 reg3183,
                 reg3182,
                 reg3181,
                 reg3179,
                 reg3180,
                 forvar3179,
                 reg3178,
                 reg3169,
                 reg3177,
                 reg3176,
                 reg3175,
                 reg3174,
                 reg3173,
                 reg3172,
                 reg3171,
                 reg3170,
                 forvar3169,
                 reg3168,
                 reg3167,
                 reg3166,
                 reg3165,
                 forvar3164,
                 reg3163,
                 reg3162,
                 reg3161,
                 reg3157,
                 reg3160,
                 forvar3159,
                 reg3158,
                 forvar3157,
                 forvar3156,
                 forvar3142,
                 forvar3139,
                 forvar3134,
                 forvar3124,
                 reg3155,
                 reg3154,
                 reg3153,
                 forvar3152,
                 reg3151,
                 reg3150,
                 reg3147,
                 reg3144,
                 reg3143,
                 reg3140,
                 forvar3138,
                 forvar3137,
                 reg3132,
                 forvar3131,
                 reg3129,
                 reg3125,
                 reg3149,
                 reg3148,
                 forvar3147,
                 reg3146,
                 reg3145,
                 forvar3144,
                 forvar3143,
                 reg3142,
                 reg3141,
                 forvar3140,
                 reg3139,
                 reg3138,
                 reg3137,
                 reg3136,
                 reg3135,
                 reg3134,
                 reg3133,
                 forvar3132,
                 reg3131,
                 reg3130,
                 forvar3129,
                 reg3128,
                 reg3127,
                 reg3126,
                 forvar3125,
                 reg3124,
                 reg3123,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg3123 <= ($signed(({wire3122} < wire3119)) <= wire3121);
      if (wire3120)
        begin
          reg3124 <= ($unsigned($unsigned((wire3121 ? (8'hb4) : (8'ha8)))) ?
              $unsigned($unsigned($signed(wire3122))) : ((8'haf) * {(wire3122 ?
                      wire3118 : wire3122)}));
          if (wire3118)
            begin
              if ((^$unsigned((8'ha0))))
                begin
                  for (forvar3125 = (1'h0); (forvar3125 < (2'h2)); forvar3125 = (forvar3125 + (1'h1)))
                    begin
                      reg3126 <= (~^wire3120[(2'h3):(1'h1)]);
                      reg3127 <= ((((~^wire3119) ^ $unsigned(wire3118)) ?
                              wire3121 : (wire3118 ?
                                  $unsigned(reg3123) : (8'haa))) ?
                          {($signed((8'hb2)) >= $signed(wire3118))} : $unsigned(wire3119[(1'h1):(1'h0)]));
                      reg3128 <= $unsigned((&$unsigned((+(8'ha0)))));
                    end
                end
              else
                begin
                  for (forvar3125 = (1'h0); (forvar3125 < (2'h2)); forvar3125 = (forvar3125 + (1'h1)))
                    begin
                      reg3126 <= {(8'hb6)};
                      reg3127 <= forvar3125;
                      reg3128 <= (^($unsigned((8'haa)) >> ($signed((8'h9c)) <<< reg3123)));
                    end
                  for (forvar3129 = (1'h0); (forvar3129 < (1'h0)); forvar3129 = (forvar3129 + (1'h1)))
                    begin
                      reg3130 <= $signed({((wire3122 | reg3127) ?
                              $unsigned(reg3126) : reg3123[(3'h4):(3'h4)])});
                      reg3131 <= $signed($signed(((!wire3118) ?
                          reg3126[(4'hc):(3'h5)] : wire3121[(4'h9):(3'h6)])));
                    end
                end
              if ($signed((reg3131 ? $signed($signed(reg3124)) : wire3122)))
                begin
                  for (forvar3132 = (1'h0); (forvar3132 < (2'h3)); forvar3132 = (forvar3132 + (1'h1)))
                    begin
                      reg3133 <= ((+(!$unsigned(wire3119))) != reg3124[(4'hc):(2'h2)]);
                      reg3134 <= wire3118[(4'hb):(3'h5)];
                      reg3135 <= ($unsigned($unsigned((reg3131 ?
                              reg3124 : reg3130))) ?
                          reg3124 : reg3128);
                    end
                  reg3136 <= $signed(forvar3129);
                  reg3137 <= (^~{forvar3129[(2'h2):(1'h1)]});
                end
              else
                begin
                  for (forvar3132 = (1'h0); (forvar3132 < (2'h2)); forvar3132 = (forvar3132 + (1'h1)))
                    begin
                      reg3133 <= ($signed($unsigned((8'hae))) == $unsigned(reg3126));
                      reg3134 <= $unsigned(reg3123[(1'h0):(1'h0)]);
                      reg3135 <= forvar3132[(2'h2):(2'h2)];
                      reg3136 <= ($unsigned(reg3133[(1'h0):(1'h0)]) ?
                          $unsigned({reg3126}) : $signed(wire3121[(4'hb):(3'h7)]));
                    end
                  if ((reg3130[(1'h1):(1'h1)] ?
                      (($signed(reg3124) ?
                              (reg3131 ?
                                  wire3121 : wire3121) : reg3126[(4'hb):(3'h6)]) ?
                          reg3133 : (forvar3125[(2'h3):(1'h1)] ?
                              reg3131 : wire3122)) : (reg3128 ?
                          $signed(reg3130) : $signed((~&reg3127)))))
                    begin
                      reg3137 <= $signed((^~(~reg3134[(2'h3):(1'h0)])));
                      reg3138 <= ((($signed(wire3118) <= $unsigned(reg3124)) ^~ reg3135) ?
                          reg3134[(1'h1):(1'h0)] : reg3133);
                    end
                  else
                    begin
                      reg3137 <= (~&wire3118);
                      reg3138 <= reg3138;
                      reg3139 <= $signed(($unsigned((reg3131 + forvar3129)) ^ wire3119[(1'h0):(1'h0)]));
                    end
                  for (forvar3140 = (1'h0); (forvar3140 < (2'h3)); forvar3140 = (forvar3140 + (1'h1)))
                    begin
                      reg3141 <= {(reg3123 ?
                              (&$unsigned((8'hb3))) : ($unsigned((8'hb2)) != (8'ha9)))};
                    end
                end
              reg3142 <= $unsigned(reg3138[(3'h7):(1'h0)]);
              for (forvar3143 = (1'h0); (forvar3143 < (1'h1)); forvar3143 = (forvar3143 + (1'h1)))
                begin
                  for (forvar3144 = (1'h0); (forvar3144 < (1'h1)); forvar3144 = (forvar3144 + (1'h1)))
                    begin
                      reg3145 <= (^$unsigned($signed($signed((8'ha6)))));
                      reg3146 <= $signed($unsigned(forvar3143));
                    end
                  for (forvar3147 = (1'h0); (forvar3147 < (1'h0)); forvar3147 = (forvar3147 + (1'h1)))
                    begin
                      reg3148 <= $unsigned($signed((~&(wire3120 ?
                          wire3122 : reg3141))));
                    end
                  reg3149 <= $signed(reg3148);
                end
            end
          else
            begin
              if ($unsigned($unsigned((~^reg3146))))
                begin
                  if (($unsigned(({(8'hae)} ?
                      {reg3126} : (8'hb8))) != $signed((((8'hb6) | (8'hb5)) ?
                      reg3146[(4'hb):(4'ha)] : (forvar3147 > wire3122)))))
                    begin
                      reg3125 <= ((!($unsigned(wire3118) > reg3126[(2'h3):(2'h3)])) * reg3126);
                      reg3126 <= $unsigned($signed((((8'hb8) ?
                          reg3138 : reg3146) && wire3122[(4'ha):(2'h2)])));
                      reg3127 <= wire3120[(3'h7):(1'h0)];
                    end
                  else
                    begin
                      reg3125 <= (~|(8'ha1));
                      reg3126 <= (reg3141[(3'h5):(3'h5)] || (^~{(~^reg3130)}));
                      reg3127 <= $signed($unsigned(reg3145[(3'h7):(3'h6)]));
                    end
                  if (reg3134[(3'h5):(3'h5)])
                    begin
                      reg3128 <= $unsigned((8'h9d));
                    end
                  else
                    begin
                      reg3128 <= (^~$signed((~|(&forvar3147))));
                      reg3129 <= forvar3143[(1'h0):(1'h0)];
                      reg3130 <= reg3141;
                    end
                  for (forvar3131 = (1'h0); (forvar3131 < (2'h3)); forvar3131 = (forvar3131 + (1'h1)))
                    begin
                      reg3132 <= wire3120[(4'h9):(1'h1)];
                      reg3133 <= (+wire3120);
                    end
                  reg3134 <= {reg3142};
                end
              else
                begin
                  for (forvar3125 = (1'h0); (forvar3125 < (1'h0)); forvar3125 = (forvar3125 + (1'h1)))
                    begin
                      reg3126 <= reg3141[(4'h9):(3'h5)];
                      reg3127 <= $signed((!(8'hb7)));
                      reg3128 <= wire3120[(2'h2):(1'h1)];
                      reg3129 <= (reg3142 ?
                          (^~($signed((8'hb0)) ?
                              (8'ha2) : $signed(reg3135))) : reg3146[(4'hb):(1'h0)]);
                    end
                  if ($signed(($unsigned({reg3125}) + (8'ha0))))
                    begin
                      reg3130 <= $signed((reg3138 ?
                          ((forvar3143 ?
                              reg3128 : (8'ha3)) << wire3120) : reg3138[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg3130 <= ($unsigned((^~reg3129)) & $unsigned(reg3146));
                      reg3131 <= $signed($unsigned($unsigned((reg3125 != reg3129))));
                    end
                  for (forvar3132 = (1'h0); (forvar3132 < (1'h0)); forvar3132 = (forvar3132 + (1'h1)))
                    begin
                      reg3133 <= $unsigned((((wire3122 + reg3130) && (reg3132 <<< reg3130)) && (~|(reg3138 ?
                          reg3138 : forvar3140))));
                      reg3134 <= {forvar3129};
                      reg3135 <= reg3131;
                      reg3136 <= {($unsigned((reg3128 != forvar3125)) | $signed((reg3138 > reg3128)))};
                    end
                end
              for (forvar3137 = (1'h0); (forvar3137 < (2'h2)); forvar3137 = (forvar3137 + (1'h1)))
                begin
                  for (forvar3138 = (1'h0); (forvar3138 < (1'h0)); forvar3138 = (forvar3138 + (1'h1)))
                    begin
                      reg3139 <= forvar3138;
                      reg3140 <= wire3120[(2'h2):(1'h1)];
                      reg3141 <= $unsigned($signed(((forvar3129 < reg3128) & (forvar3143 ?
                          (8'had) : wire3120))));
                      reg3142 <= $unsigned(reg3140[(3'h6):(1'h1)]);
                    end
                end
              reg3143 <= forvar3140;
              if (((8'ha6) ?
                  ($signed((reg3132 ? (8'hb4) : (8'ha8))) ?
                      $unsigned(reg3134) : (&{reg3145})) : forvar3144))
                begin
                  reg3144 <= {$signed((+(reg3145 ? reg3129 : reg3134)))};
                end
              else
                begin
                  if (reg3139[(3'h4):(2'h2)])
                    begin
                      reg3144 <= reg3138[(3'h6):(2'h3)];
                      reg3145 <= (-$unsigned(($unsigned(reg3135) * $signed(reg3143))));
                    end
                  else
                    begin
                      reg3144 <= reg3137;
                      reg3145 <= $signed(wire3122[(4'h8):(3'h4)]);
                      reg3146 <= ((|($unsigned(reg3129) ?
                              $unsigned(reg3143) : (reg3142 ?
                                  forvar3147 : forvar3137))) ?
                          reg3126[(3'h7):(1'h1)] : (~^$unsigned(reg3146)));
                      reg3147 <= reg3149[(3'h6):(2'h3)];
                    end
                  if (reg3130[(1'h0):(1'h0)])
                    begin
                      reg3148 <= (~forvar3144[(4'hf):(3'h6)]);
                      reg3149 <= (reg3124[(4'h8):(3'h5)] >= {$unsigned(((8'hb8) ?
                              reg3149 : reg3146))});
                      reg3150 <= reg3143;
                      reg3151 <= reg3133[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3148 <= forvar3132;
                      reg3149 <= (((wire3119[(1'h1):(1'h1)] + $signed(forvar3137)) && ($signed(reg3136) >= reg3146[(4'h8):(1'h0)])) ?
                          {(^{reg3134})} : $signed(((reg3126 - forvar3140) <= (8'hac))));
                      reg3150 <= reg3137[(4'h9):(1'h1)];
                    end
                  for (forvar3152 = (1'h0); (forvar3152 < (2'h2)); forvar3152 = (forvar3152 + (1'h1)))
                    begin
                      reg3153 <= $unsigned((reg3136 ?
                          $unsigned($signed(forvar3140)) : $unsigned((reg3124 >= reg3126))));
                      reg3154 <= reg3146;
                      reg3155 <= reg3143[(2'h3):(1'h0)];
                    end
                end
            end
        end
      else
        begin
          for (forvar3124 = (1'h0); (forvar3124 < (2'h2)); forvar3124 = (forvar3124 + (1'h1)))
            begin
              for (forvar3125 = (1'h0); (forvar3125 < (1'h0)); forvar3125 = (forvar3125 + (1'h1)))
                begin
                  if ($signed(({(wire3120 ? reg3139 : forvar3147)} ?
                      forvar3140[(3'h6):(1'h0)] : reg3127)))
                    begin
                      reg3126 <= (~|$signed((-(|reg3127))));
                      reg3127 <= $signed(($unsigned((^forvar3147)) ~^ $unsigned(reg3127[(1'h0):(1'h0)])));
                      reg3128 <= wire3119[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg3126 <= ($signed((+reg3145)) > reg3146);
                    end
                  for (forvar3129 = (1'h0); (forvar3129 < (2'h2)); forvar3129 = (forvar3129 + (1'h1)))
                    begin
                      reg3130 <= reg3141;
                      reg3131 <= (-$unsigned(reg3140));
                      reg3132 <= ($signed(reg3145) ^~ (($unsigned(reg3132) ?
                          (8'hac) : (8'hae)) + $unsigned(((8'hb2) ?
                          reg3146 : forvar3124))));
                      reg3133 <= forvar3132[(2'h2):(1'h0)];
                    end
                  for (forvar3134 = (1'h0); (forvar3134 < (1'h1)); forvar3134 = (forvar3134 + (1'h1)))
                    begin
                      reg3135 <= (-forvar3137);
                      reg3136 <= (({forvar3129[(2'h3):(1'h0)]} & forvar3143) == reg3142);
                      reg3137 <= forvar3152;
                      reg3138 <= reg3133;
                    end
                  for (forvar3139 = (1'h0); (forvar3139 < (1'h1)); forvar3139 = (forvar3139 + (1'h1)))
                    begin
                      reg3140 <= wire3118[(3'h5):(1'h0)];
                    end
                end
              reg3141 <= reg3149[(2'h2):(1'h1)];
              for (forvar3142 = (1'h0); (forvar3142 < (1'h0)); forvar3142 = (forvar3142 + (1'h1)))
                begin
                  reg3143 <= forvar3147;
                  reg3144 <= ((($signed(reg3146) < (|reg3148)) >>> forvar3140) ?
                      $signed(($unsigned(reg3124) ?
                          (reg3132 & reg3145) : reg3123[(2'h2):(1'h1)])) : $signed(reg3137));
                end
            end
          reg3145 <= $unsigned(forvar3139[(1'h0):(1'h0)]);
        end
      if ($signed($signed((~^(reg3123 <<< reg3129)))))
        begin
          for (forvar3156 = (1'h0); (forvar3156 < (1'h0)); forvar3156 = (forvar3156 + (1'h1)))
            begin
              if ($unsigned((|$unsigned($signed(forvar3140)))))
                begin
                  for (forvar3157 = (1'h0); (forvar3157 < (2'h3)); forvar3157 = (forvar3157 + (1'h1)))
                    begin
                      reg3158 <= $signed((+$signed($unsigned(reg3153))));
                    end
                  for (forvar3159 = (1'h0); (forvar3159 < (2'h2)); forvar3159 = (forvar3159 + (1'h1)))
                    begin
                      reg3160 <= $unsigned($unsigned(($signed(reg3135) ~^ $signed(reg3126))));
                    end
                end
              else
                begin
                  if ({(wire3119 << ($unsigned(reg3154) ?
                          forvar3147 : forvar3142[(3'h4):(2'h2)]))})
                    begin
                      reg3157 <= (($signed({reg3141}) ~^ reg3123[(2'h3):(2'h3)]) ?
                          $unsigned({((8'haa) == (8'ha7))}) : $unsigned($unsigned((reg3138 ?
                              wire3121 : (8'hb8)))));
                      reg3158 <= (($unsigned((^~reg3155)) * {(!reg3127)}) ^~ ($signed((forvar3147 << reg3127)) >= $unsigned(forvar3125)));
                    end
                  else
                    begin
                      reg3157 <= (~(~&reg3128));
                    end
                  for (forvar3159 = (1'h0); (forvar3159 < (2'h3)); forvar3159 = (forvar3159 + (1'h1)))
                    begin
                      reg3160 <= $signed((-(+$unsigned(reg3149))));
                      reg3161 <= $signed($unsigned(($signed(reg3150) ?
                          (|forvar3132) : $unsigned(reg3154))));
                      reg3162 <= ((&$signed(forvar3139[(2'h2):(1'h1)])) - (((!forvar3124) ?
                          forvar3132[(2'h2):(2'h2)] : $unsigned(reg3139)) <= ((reg3146 <= wire3118) || forvar3157[(2'h2):(2'h2)])));
                    end
                  reg3163 <= wire3118[(4'h9):(4'h9)];
                  for (forvar3164 = (1'h0); (forvar3164 < (2'h3)); forvar3164 = (forvar3164 + (1'h1)))
                    begin
                      reg3165 <= ({($signed((8'hba)) ?
                                  (^~(8'h9e)) : {reg3149})} ?
                          ((reg3129[(4'h9):(3'h5)] >>> reg3124) == $unsigned((~^wire3122))) : $unsigned(((~&forvar3157) ?
                              (&reg3134) : (-wire3122))));
                      reg3166 <= forvar3144[(3'h4):(3'h4)];
                      reg3167 <= (forvar3147[(2'h3):(1'h0)] >>> reg3129);
                    end
                end
              if ({(~|forvar3147[(3'h4):(3'h4)])})
                begin
                  reg3168 <= {(~^({wire3122} ?
                          $signed(reg3162) : (reg3135 & reg3158)))};
                  for (forvar3169 = (1'h0); (forvar3169 < (2'h2)); forvar3169 = (forvar3169 + (1'h1)))
                    begin
                      reg3170 <= (!(|forvar3134));
                      reg3171 <= (forvar3144[(3'h5):(3'h4)] ?
                          forvar3144[(3'h4):(1'h1)] : (&((!reg3137) != {forvar3139})));
                      reg3172 <= (reg3150 >= forvar3134);
                    end
                  if (((((reg3132 < reg3131) ^ $unsigned(reg3126)) ~^ ($signed(wire3119) ?
                          (forvar3144 ^ reg3170) : $unsigned(forvar3147))) ?
                      $signed(forvar3134) : wire3121[(1'h1):(1'h1)]))
                    begin
                      reg3173 <= (~forvar3156);
                    end
                  else
                    begin
                      reg3173 <= reg3123;
                      reg3174 <= forvar3131[(3'h4):(2'h3)];
                      reg3175 <= {(^reg3142[(1'h0):(1'h0)])};
                      reg3176 <= (+reg3155[(4'h9):(1'h0)]);
                    end
                  reg3177 <= (~|reg3172);
                end
              else
                begin
                  if (($unsigned(forvar3156[(3'h6):(3'h4)]) ^~ {((wire3119 <= reg3163) + (reg3172 >> reg3145))}))
                    begin
                      reg3168 <= forvar3143[(3'h7):(2'h3)];
                      reg3169 <= reg3142[(2'h3):(2'h2)];
                      reg3170 <= (($signed((reg3170 >>> forvar3156)) || (~|$unsigned(wire3118))) ?
                          reg3161[(1'h0):(1'h0)] : {reg3151[(3'h7):(3'h5)]});
                    end
                  else
                    begin
                      reg3168 <= (&(+(8'hb4)));
                      reg3169 <= $unsigned(reg3169[(3'h5):(1'h1)]);
                    end
                end
              reg3178 <= {(forvar3169 ? (~|$signed(reg3153)) : reg3158)};
            end
          if (reg3175[(1'h0):(1'h0)])
            begin
              if ((reg3142 ?
                  (~|reg3148[(3'h4):(2'h3)]) : $signed({(forvar3139 ?
                          reg3141 : reg3147)})))
                begin
                  for (forvar3179 = (1'h0); (forvar3179 < (1'h1)); forvar3179 = (forvar3179 + (1'h1)))
                    begin
                      reg3180 <= (forvar3142[(3'h4):(2'h3)] ?
                          (~{(reg3160 ?
                                  reg3150 : (8'ha2))}) : $signed($signed(reg3124[(2'h2):(2'h2)])));
                    end
                end
              else
                begin
                  if (forvar3131)
                    begin
                      reg3179 <= ((reg3135 ?
                              ((!forvar3139) ?
                                  (~^reg3137) : (reg3127 ?
                                      forvar3142 : reg3173)) : $signed(reg3160[(1'h0):(1'h0)])) ?
                          reg3180[(1'h1):(1'h1)] : (|($signed(reg3165) ?
                              (~&reg3157) : reg3132[(1'h0):(1'h0)])));
                      reg3180 <= ((reg3155 ?
                              reg3128[(2'h2):(1'h0)] : ((forvar3164 && forvar3132) ?
                                  $signed(forvar3132) : (reg3178 ?
                                      reg3142 : forvar3156))) ?
                          $unsigned($unsigned($signed(reg3145))) : $unsigned(reg3145[(1'h0):(1'h0)]));
                      reg3181 <= (-$signed($unsigned((|reg3140))));
                    end
                  else
                    begin
                      reg3179 <= {$signed($signed(reg3130[(1'h1):(1'h0)]))};
                      reg3180 <= $unsigned($signed($signed((~&reg3157))));
                      reg3181 <= $signed((!$signed((reg3124 ?
                          reg3171 : reg3142))));
                      reg3182 <= reg3124;
                    end
                  if (forvar3159[(4'ha):(1'h1)])
                    begin
                      reg3183 <= $unsigned($signed($unsigned(wire3121)));
                      reg3184 <= $unsigned((forvar3129 ?
                          (+(reg3167 == reg3172)) : {reg3127[(1'h1):(1'h1)]}));
                      reg3185 <= $signed((~|reg3168));
                      reg3186 <= reg3170;
                    end
                  else
                    begin
                      reg3183 <= (!((((8'h9e) >>> reg3144) + (~&(8'hb8))) ?
                          $unsigned((-(8'hba))) : wire3118));
                      reg3184 <= $unsigned((8'hae));
                    end
                  if ($signed({$signed(reg3124[(3'h6):(2'h2)])}))
                    begin
                      reg3187 <= (reg3185 | wire3120);
                      reg3188 <= ($signed($unsigned(((8'hb5) ?
                          wire3121 : reg3187))) - reg3169[(4'h9):(2'h2)]);
                      reg3189 <= ($signed((8'hb4)) ^~ reg3175[(1'h1):(1'h0)]);
                      reg3190 <= (!((~&reg3142) ^ reg3184[(4'he):(3'h5)]));
                    end
                  else
                    begin
                      reg3187 <= forvar3138;
                      reg3188 <= ((^$unsigned($signed(forvar3139))) >> reg3183[(4'ha):(4'h9)]);
                      reg3189 <= ((8'hb6) ? reg3126[(3'h5):(3'h4)] : reg3175);
                      reg3190 <= $unsigned({reg3133[(1'h1):(1'h1)]});
                    end
                end
              for (forvar3191 = (1'h0); (forvar3191 < (2'h3)); forvar3191 = (forvar3191 + (1'h1)))
                begin
                  for (forvar3192 = (1'h0); (forvar3192 < (2'h2)); forvar3192 = (forvar3192 + (1'h1)))
                    begin
                      reg3193 <= $unsigned({$signed(reg3145[(1'h1):(1'h0)])});
                      reg3194 <= {$unsigned($signed(reg3181))};
                      reg3195 <= ({(-reg3143[(2'h3):(1'h1)])} >>> $signed(reg3125[(3'h5):(2'h3)]));
                    end
                  reg3196 <= reg3190;
                end
              if (reg3151)
                begin
                  if ((8'hb7))
                    begin
                      reg3197 <= reg3194;
                      reg3198 <= forvar3144[(3'h6):(1'h1)];
                      reg3199 <= (!(8'hac));
                    end
                  else
                    begin
                      reg3197 <= (~&((~^{reg3187}) < (+reg3168)));
                      reg3198 <= (((8'ha9) > reg3171[(2'h2):(1'h1)]) ?
                          $signed((+{reg3166})) : $signed((~|{reg3158})));
                      reg3199 <= {reg3151};
                      reg3200 <= $unsigned(reg3157);
                    end
                  if ($signed((+(&$signed(reg3187)))))
                    begin
                      reg3201 <= (^~((forvar3138 ?
                          (reg3141 ~^ reg3155) : (forvar3137 & reg3127)) * reg3173[(2'h2):(1'h0)]));
                      reg3202 <= $unsigned((8'hb5));
                    end
                  else
                    begin
                      reg3201 <= reg3174[(3'h7):(1'h1)];
                      reg3202 <= (+(($signed((8'ha9)) ?
                              $signed((8'ha4)) : (forvar3156 ?
                                  (8'h9c) : reg3195)) ?
                          $unsigned((reg3181 ?
                              forvar3138 : reg3142)) : $unsigned({(8'ha7)})));
                      reg3203 <= (($signed(reg3183[(4'hb):(1'h1)]) && $signed((forvar3124 >= (8'haf)))) ?
                          reg3151 : (^reg3180));
                      reg3204 <= {$signed(forvar3191[(3'h6):(3'h4)])};
                    end
                end
              else
                begin
                  for (forvar3197 = (1'h0); (forvar3197 < (1'h0)); forvar3197 = (forvar3197 + (1'h1)))
                    begin
                      reg3198 <= ((8'ha0) || (reg3176 <<< reg3174[(3'h4):(1'h1)]));
                      reg3199 <= $signed({(8'h9e)});
                      reg3200 <= $unsigned((&$signed(reg3190)));
                    end
                  if ((8'ha8))
                    begin
                      reg3201 <= (-(reg3167 ? reg3124 : $signed(reg3151)));
                    end
                  else
                    begin
                      reg3201 <= $signed(forvar3152[(1'h1):(1'h1)]);
                      reg3202 <= ((^~{((8'ha4) && forvar3144)}) != reg3186);
                      reg3203 <= ($unsigned((~^$unsigned(reg3187))) >>> $signed((forvar3157[(2'h2):(2'h2)] && $signed(reg3151))));
                      reg3204 <= $unsigned((~(forvar3192 == reg3160[(4'h8):(1'h1)])));
                    end
                  for (forvar3205 = (1'h0); (forvar3205 < (2'h3)); forvar3205 = (forvar3205 + (1'h1)))
                    begin
                      reg3206 <= $signed((^~((reg3128 ? reg3198 : reg3203) ?
                          {reg3133} : $unsigned(wire3118))));
                      reg3207 <= (($unsigned($unsigned(forvar3157)) ?
                              ((forvar3156 ? forvar3152 : reg3125) ?
                                  ((8'ha2) << (8'hba)) : (+reg3197)) : ($signed(reg3158) ?
                                  (reg3131 ?
                                      (8'hb0) : (8'hb0)) : reg3158[(2'h2):(2'h2)])) ?
                          (((forvar3140 ^ reg3206) != {(8'ha7)}) ?
                              (|$signed((8'hb1))) : $unsigned(reg3168)) : reg3174[(4'h9):(4'h9)]);
                      reg3208 <= $signed(((|reg3130[(1'h1):(1'h1)]) < forvar3137));
                      reg3209 <= (((reg3157 + (reg3168 ^ reg3194)) ?
                              ($signed(forvar3159) ?
                                  (reg3149 ?
                                      forvar3197 : forvar3147) : (reg3206 ?
                                      reg3170 : forvar3138)) : $unsigned({reg3157})) ?
                          ($signed(reg3174[(4'h8):(3'h5)]) != ((~reg3125) ?
                              (8'hb3) : forvar3144[(3'h5):(3'h4)])) : (^$unsigned((~reg3157))));
                    end
                  if ($unsigned(reg3202))
                    begin
                      reg3210 <= reg3142[(2'h3):(2'h2)];
                      reg3211 <= $signed((^$signed(reg3132[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg3210 <= (~^((((8'hb5) <= reg3139) ^ (|reg3167)) ?
                          (reg3201[(3'h5):(1'h1)] | (|forvar3179)) : reg3127));
                      reg3211 <= (reg3193[(2'h2):(2'h2)] ^~ reg3129[(4'h8):(4'h8)]);
                      reg3212 <= ((~|forvar3132[(1'h1):(1'h0)]) ?
                          (~^($signed(forvar3169) ?
                              {(8'h9d)} : (8'hba))) : $signed((((8'hba) ?
                              reg3148 : reg3198) <<< reg3204)));
                    end
                end
            end
          else
            begin
              for (forvar3179 = (1'h0); (forvar3179 < (1'h1)); forvar3179 = (forvar3179 + (1'h1)))
                begin
                  if ((({$signed(reg3147)} ?
                          ((reg3173 + reg3169) > (^~reg3209)) : forvar3140[(1'h1):(1'h0)]) ?
                      reg3139[(4'h9):(3'h6)] : reg3183[(4'he):(3'h5)]))
                    begin
                      reg3180 <= ($signed((reg3188[(3'h4):(1'h1)] ?
                          $signed(reg3133) : (8'ha5))) ^~ forvar3157);
                      reg3181 <= $unsigned({$unsigned((+reg3133))});
                      reg3182 <= ((forvar3142 ?
                          $unsigned(forvar3132) : ((^~reg3125) & $unsigned(reg3132))) & reg3189);
                    end
                  else
                    begin
                      reg3180 <= ((forvar3144 ^ (8'ha7)) ?
                          ((^~(forvar3156 ?
                              reg3149 : reg3169)) && ((reg3174 ^~ reg3143) ?
                              $unsigned(reg3177) : reg3131)) : reg3165[(2'h2):(1'h1)]);
                      reg3181 <= wire3118[(4'h8):(3'h7)];
                      reg3182 <= $signed((($signed(forvar3191) ?
                              (forvar3124 ~^ reg3211) : $signed(forvar3125)) ?
                          reg3181[(3'h7):(3'h5)] : ((reg3133 >= reg3204) ?
                              $signed(reg3141) : (8'haf))));
                      reg3183 <= (reg3166 <<< ($signed(forvar3157[(1'h0):(1'h0)]) ?
                          ($signed(reg3189) * (reg3163 ?
                              (8'ha9) : (8'hb6))) : {$signed(reg3134)}));
                    end
                  if (reg3143[(3'h7):(3'h5)])
                    begin
                      reg3184 <= (($signed((reg3211 ? reg3203 : (8'hb5))) ?
                          $unsigned((reg3211 ?
                              reg3201 : reg3171)) : (-{forvar3164})) || {(~$signed(forvar3142))});
                      reg3185 <= reg3124;
                      reg3186 <= ($unsigned($unsigned(wire3119[(1'h1):(1'h1)])) && wire3122[(4'h9):(3'h5)]);
                    end
                  else
                    begin
                      reg3184 <= reg3136;
                    end
                end
              for (forvar3187 = (1'h0); (forvar3187 < (2'h2)); forvar3187 = (forvar3187 + (1'h1)))
                begin
                  for (forvar3188 = (1'h0); (forvar3188 < (1'h1)); forvar3188 = (forvar3188 + (1'h1)))
                    begin
                      reg3189 <= ($signed($unsigned($signed(reg3150))) ?
                          forvar3152 : $unsigned(($unsigned(reg3211) ?
                              (reg3143 ?
                                  reg3187 : reg3181) : (reg3197 >> forvar3138))));
                      reg3190 <= ((reg3169[(1'h0):(1'h0)] ?
                          $signed(reg3196[(4'hb):(1'h0)]) : {$unsigned(wire3120)}) ^~ $signed($unsigned((~&reg3147))));
                      reg3191 <= $signed((^~$signed($signed(reg3206))));
                    end
                  for (forvar3192 = (1'h0); (forvar3192 < (1'h1)); forvar3192 = (forvar3192 + (1'h1)))
                    begin
                      reg3193 <= ((({reg3162} ?
                                  (forvar3138 >> (8'h9c)) : {wire3119}) ?
                              reg3132 : (8'ha5)) ?
                          (forvar3138[(2'h2):(2'h2)] ?
                              (+reg3193) : reg3143[(3'h7):(3'h5)]) : ({(reg3125 & reg3186)} != $signed((^(8'ha3)))));
                      reg3194 <= $unsigned(((|(~|reg3181)) ?
                          (forvar3139 ?
                              ((8'ha7) || reg3161) : (~&reg3144)) : ((reg3210 ?
                                  forvar3132 : reg3165) ?
                              (-reg3161) : $signed(reg3129))));
                    end
                  for (forvar3195 = (1'h0); (forvar3195 < (2'h3)); forvar3195 = (forvar3195 + (1'h1)))
                    begin
                      reg3196 <= ((-(+$unsigned(reg3202))) ?
                          reg3202[(2'h2):(2'h2)] : (forvar3137 ?
                              (~&(^~(8'hb8))) : (~|{(8'hb6)})));
                      reg3197 <= (-($unsigned((~^reg3138)) ?
                          (~|reg3198) : {(forvar3124 + forvar3147)}));
                      reg3198 <= forvar3138;
                    end
                  if (((8'ha2) ?
                      (|reg3173) : ($unsigned($unsigned(reg3203)) ?
                          ($unsigned(reg3172) ?
                              (~|forvar3159) : $signed(reg3193)) : ({forvar3124} == (+reg3196)))))
                    begin
                      reg3199 <= reg3201[(3'h4):(1'h1)];
                      reg3200 <= $unsigned($unsigned($unsigned($unsigned(reg3201))));
                    end
                  else
                    begin
                      reg3199 <= $signed($unsigned({forvar3124}));
                      reg3200 <= reg3150;
                      reg3201 <= forvar3129;
                    end
                end
              if ((($signed(wire3121) ?
                      ($unsigned(forvar3164) ~^ (~reg3131)) : ($signed(reg3158) ~^ (reg3137 >>> forvar3138))) ?
                  (~|$signed((reg3179 ?
                      reg3123 : forvar3157))) : (reg3174 == ({reg3125} << $signed(reg3130)))))
                begin
                  if (reg3183)
                    begin
                      reg3202 <= (reg3195[(2'h2):(1'h0)] == reg3137);
                      reg3203 <= $unsigned(wire3118[(3'h5):(1'h0)]);
                      reg3204 <= {forvar3129};
                    end
                  else
                    begin
                      reg3202 <= reg3177;
                      reg3203 <= $signed(reg3125);
                    end
                  for (forvar3205 = (1'h0); (forvar3205 < (1'h1)); forvar3205 = (forvar3205 + (1'h1)))
                    begin
                      reg3206 <= reg3137[(2'h2):(2'h2)];
                      reg3207 <= (8'ha1);
                      reg3208 <= (8'hba);
                      reg3209 <= reg3133[(1'h0):(1'h0)];
                    end
                  if ((($unsigned((reg3187 > (8'ha5))) * (+{(8'h9c)})) ?
                      forvar3131[(2'h2):(1'h0)] : $signed($signed($unsigned(reg3200)))))
                    begin
                      reg3210 <= (((8'h9d) ~^ reg3202[(2'h2):(2'h2)]) ?
                          ((((8'hb5) ?
                              reg3171 : forvar3205) ^ (!(8'hb8))) ~^ $unsigned((reg3132 >= reg3191))) : ($unsigned((~^reg3203)) > reg3206[(3'h4):(2'h2)]));
                      reg3211 <= (^$unsigned($signed(reg3155[(3'h5):(1'h0)])));
                    end
                  else
                    begin
                      reg3210 <= reg3163[(2'h3):(2'h2)];
                      reg3211 <= $signed(reg3163);
                      reg3212 <= $signed({$unsigned((forvar3187 ?
                              reg3160 : forvar3147))});
                      reg3213 <= $signed((~reg3165));
                    end
                end
              else
                begin
                  if (reg3201)
                    begin
                      reg3202 <= reg3184[(1'h0):(1'h0)];
                      reg3203 <= (($unsigned((forvar3157 > reg3163)) ?
                          ((reg3144 ? (8'hb1) : reg3202) ?
                              ((8'hb5) <<< (8'hb9)) : reg3124) : (wire3121[(4'h9):(3'h4)] && $unsigned(reg3132))) == reg3154);
                      reg3204 <= $signed($signed(forvar3157[(2'h2):(1'h0)]));
                      reg3205 <= (reg3177 ?
                          forvar3147[(2'h3):(2'h3)] : forvar3124);
                    end
                  else
                    begin
                      reg3202 <= $unsigned(forvar3143[(3'h6):(3'h4)]);
                    end
                  for (forvar3206 = (1'h0); (forvar3206 < (1'h0)); forvar3206 = (forvar3206 + (1'h1)))
                    begin
                      reg3207 <= $unsigned({((reg3170 + forvar3131) ?
                              (8'h9e) : $signed(reg3144))});
                    end
                  reg3208 <= reg3161[(1'h1):(1'h0)];
                  if (($unsigned(({(8'hb9)} ?
                          reg3204[(1'h1):(1'h0)] : reg3196[(2'h2):(2'h2)])) ?
                      (^reg3133[(1'h0):(1'h0)]) : reg3138[(1'h0):(1'h0)]))
                    begin
                      reg3209 <= (($signed(reg3144) >= reg3193[(1'h1):(1'h0)]) + (-$unsigned($unsigned((8'h9e)))));
                      reg3210 <= reg3153;
                      reg3211 <= $unsigned((((&reg3182) ?
                          (8'hae) : $unsigned(reg3193)) ~^ ((8'hb0) ?
                          reg3143[(3'h5):(2'h3)] : reg3137)));
                      reg3212 <= reg3142[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg3209 <= $unsigned(reg3185);
                    end
                end
              for (forvar3214 = (1'h0); (forvar3214 < (2'h2)); forvar3214 = (forvar3214 + (1'h1)))
                begin
                  for (forvar3215 = (1'h0); (forvar3215 < (1'h1)); forvar3215 = (forvar3215 + (1'h1)))
                    begin
                      reg3216 <= (((|(-reg3209)) ?
                              $unsigned(forvar3147) : (forvar3140 == ((8'hac) ?
                                  reg3190 : reg3176))) ?
                          $unsigned(($signed(forvar3192) ?
                              reg3148[(4'ha):(1'h1)] : reg3149[(2'h2):(2'h2)])) : (8'ha5));
                      reg3217 <= reg3169;
                      reg3218 <= $unsigned(({(forvar3140 ?
                                  reg3146 : forvar3139)} ?
                          $unsigned({reg3175}) : {forvar3129[(4'ha):(4'ha)]}));
                      reg3219 <= reg3158;
                    end
                end
            end
        end
      else
        begin
          for (forvar3156 = (1'h0); (forvar3156 < (1'h1)); forvar3156 = (forvar3156 + (1'h1)))
            begin
              if ($signed($signed((~&{reg3178}))))
                begin
                  for (forvar3157 = (1'h0); (forvar3157 < (1'h0)); forvar3157 = (forvar3157 + (1'h1)))
                    begin
                      reg3158 <= (~|{{$unsigned(forvar3140)}});
                      reg3159 <= wire3120[(4'hb):(4'ha)];
                      reg3160 <= $unsigned(reg3182[(3'h4):(1'h1)]);
                      reg3161 <= $unsigned((((reg3136 - reg3148) || (reg3154 <= reg3198)) - (reg3184 * forvar3125[(1'h0):(1'h0)])));
                    end
                  for (forvar3162 = (1'h0); (forvar3162 < (1'h0)); forvar3162 = (forvar3162 + (1'h1)))
                    begin
                      reg3163 <= (((((8'haa) ?
                              reg3129 : reg3180) + (reg3193 | reg3138)) ?
                          reg3199[(1'h1):(1'h0)] : $signed($unsigned(reg3171))) + ($signed($signed(reg3200)) ?
                          reg3191[(3'h6):(3'h6)] : $unsigned($signed(forvar3132))));
                      reg3164 <= ((reg3204[(2'h3):(2'h2)] ?
                              ((forvar3169 ? forvar3143 : reg3137) ?
                                  $signed(reg3148) : (wire3121 ^ reg3142)) : reg3141[(1'h1):(1'h1)]) ?
                          $unsigned((reg3213[(4'h9):(1'h0)] ?
                              $signed(reg3208) : forvar3206[(1'h1):(1'h1)])) : (($signed(forvar3197) <<< {wire3118}) ~^ reg3135[(2'h3):(1'h0)]));
                      reg3165 <= forvar3143[(3'h5):(2'h3)];
                    end
                  if ($unsigned(((~&reg3209[(4'ha):(1'h1)]) <= (reg3200[(1'h1):(1'h1)] ?
                      (!reg3136) : {reg3208}))))
                    begin
                      reg3166 <= reg3157[(3'h5):(3'h5)];
                      reg3167 <= (!$unsigned((-forvar3197)));
                      reg3168 <= ((&((reg3219 - (8'hb1)) ?
                          ((8'hb2) ?
                              reg3172 : forvar3206) : $unsigned(reg3140))) >> $unsigned(wire3122[(4'hc):(2'h3)]));
                    end
                  else
                    begin
                      reg3166 <= (!forvar3124);
                    end
                end
              else
                begin
                  reg3157 <= ($signed((^~(8'ha5))) ?
                      $unsigned(forvar3134[(2'h2):(2'h2)]) : {$signed((reg3213 ?
                              reg3159 : reg3140))});
                  reg3158 <= ((!($unsigned(reg3132) ?
                          (~&reg3176) : $signed(reg3193))) ?
                      $unsigned((^~reg3193)) : {(~(reg3202 | (8'h9c)))});
                  for (forvar3159 = (1'h0); (forvar3159 < (2'h3)); forvar3159 = (forvar3159 + (1'h1)))
                    begin
                      reg3160 <= (reg3196 <= ((^~(forvar3138 >>> reg3218)) - $unsigned((reg3127 && reg3169))));
                    end
                  reg3161 <= reg3138[(2'h3):(2'h3)];
                end
            end
          for (forvar3169 = (1'h0); (forvar3169 < (1'h1)); forvar3169 = (forvar3169 + (1'h1)))
            begin
              for (forvar3170 = (1'h0); (forvar3170 < (2'h2)); forvar3170 = (forvar3170 + (1'h1)))
                begin
                  reg3171 <= $signed(forvar3191[(1'h1):(1'h1)]);
                end
              for (forvar3172 = (1'h0); (forvar3172 < (1'h1)); forvar3172 = (forvar3172 + (1'h1)))
                begin
                  for (forvar3173 = (1'h0); (forvar3173 < (1'h1)); forvar3173 = (forvar3173 + (1'h1)))
                    begin
                      reg3174 <= (!reg3208[(4'ha):(3'h4)]);
                      reg3175 <= ($signed({reg3183[(4'he):(4'hc)]}) ?
                          forvar3188[(1'h1):(1'h1)] : (~&($signed(forvar3131) ?
                              (8'had) : {(8'hac)})));
                      reg3176 <= (&$unsigned(reg3147[(2'h3):(2'h3)]));
                      reg3177 <= $signed((8'had));
                    end
                  if (reg3186)
                    begin
                      reg3178 <= ($signed(($unsigned((8'hb0)) ?
                              $signed(forvar3215) : $signed(wire3120))) ?
                          $signed($unsigned((reg3146 ?
                              reg3123 : forvar3195))) : ((((8'ha0) ?
                                      reg3155 : (8'h9f)) ?
                                  $signed((8'h9f)) : $signed(reg3185)) ?
                              reg3149[(2'h3):(1'h1)] : (reg3206 + reg3124)));
                      reg3179 <= wire3120[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3178 <= reg3217[(3'h4):(2'h3)];
                    end
                  if ($unsigned({forvar3144[(5'h10):(2'h2)]}))
                    begin
                      reg3180 <= reg3134;
                      reg3181 <= ($signed((~(!reg3197))) ?
                          $signed(((reg3123 | wire3120) & $signed((8'hab)))) : $signed(((reg3171 ?
                                  reg3124 : reg3123) ?
                              (^~(8'ha0)) : (forvar3137 | reg3137))));
                      reg3182 <= (~|$unsigned($signed((reg3136 == (8'h9c)))));
                      reg3183 <= (reg3167 >>> ($signed(forvar3187[(2'h2):(2'h2)]) - reg3149[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg3180 <= ((^~{reg3136[(4'ha):(2'h3)]}) ?
                          ((~|$signed(reg3142)) ?
                              forvar3134[(2'h2):(1'h0)] : ((^forvar3142) != (~reg3146))) : {($unsigned(reg3188) ?
                                  (reg3157 ? (8'h9d) : (8'hb5)) : (reg3160 ?
                                      reg3201 : forvar3125))});
                      reg3181 <= (~^(((forvar3156 || forvar3172) >= forvar3214) ?
                          $signed($unsigned(reg3154)) : $signed({reg3142})));
                    end
                  for (forvar3184 = (1'h0); (forvar3184 < (2'h3)); forvar3184 = (forvar3184 + (1'h1)))
                    begin
                      reg3185 <= reg3153[(4'he):(4'ha)];
                    end
                end
              reg3186 <= $unsigned({((8'hb3) ?
                      reg3182[(2'h2):(1'h1)] : forvar3172[(1'h0):(1'h0)])});
              if ($unsigned(reg3165[(2'h2):(2'h2)]))
                begin
                  if ((forvar3192 ?
                      $signed(((~|forvar3164) ?
                          reg3169[(4'ha):(4'ha)] : $signed(forvar3191))) : wire3121))
                    begin
                      reg3187 <= ($signed(forvar3147[(3'h5):(1'h0)]) <= $signed(reg3150[(3'h5):(1'h0)]));
                      reg3188 <= (~&wire3120[(1'h0):(1'h0)]);
                      reg3189 <= $unsigned($signed(reg3164[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg3187 <= {(!(forvar3214[(1'h0):(1'h0)] & (reg3133 ?
                              reg3138 : reg3194)))};
                    end
                  for (forvar3190 = (1'h0); (forvar3190 < (1'h1)); forvar3190 = (forvar3190 + (1'h1)))
                    begin
                      reg3191 <= $signed(reg3212);
                      reg3192 <= (reg3213 ?
                          $signed((forvar3173 >>> $signed(forvar3190))) : (^~(^{reg3206})));
                    end
                end
              else
                begin
                  for (forvar3187 = (1'h0); (forvar3187 < (1'h0)); forvar3187 = (forvar3187 + (1'h1)))
                    begin
                      reg3188 <= ((^~($signed(reg3146) ?
                              reg3167 : forvar3191[(3'h5):(3'h5)])) ?
                          forvar3138 : ($unsigned((8'hb8)) << (reg3212 ?
                              (!(8'hb9)) : $unsigned((8'haf)))));
                      reg3189 <= (8'hb8);
                    end
                end
            end
          reg3193 <= ($unsigned($unsigned((~forvar3188))) - {reg3167[(4'h9):(1'h0)]});
        end
      for (forvar3220 = (1'h0); (forvar3220 < (1'h1)); forvar3220 = (forvar3220 + (1'h1)))
        begin
          for (forvar3221 = (1'h0); (forvar3221 < (1'h0)); forvar3221 = (forvar3221 + (1'h1)))
            begin
              for (forvar3222 = (1'h0); (forvar3222 < (2'h2)); forvar3222 = (forvar3222 + (1'h1)))
                begin
                  reg3223 <= (^~(^~$unsigned(reg3195[(3'h6):(2'h2)])));
                  reg3224 <= $unsigned(reg3158);
                  for (forvar3225 = (1'h0); (forvar3225 < (2'h3)); forvar3225 = (forvar3225 + (1'h1)))
                    begin
                      reg3226 <= (-(~&forvar3157[(1'h0):(1'h0)]));
                      reg3227 <= (($signed($signed(forvar3124)) ?
                          reg3179 : (reg3146 ?
                              reg3136[(4'hf):(1'h1)] : reg3147)) <= $signed(($unsigned((8'haa)) ?
                          $signed(forvar3157) : $unsigned(forvar3169))));
                      reg3228 <= $signed({{(forvar3164 ?
                                  forvar3220 : reg3198)}});
                    end
                end
              for (forvar3229 = (1'h0); (forvar3229 < (2'h2)); forvar3229 = (forvar3229 + (1'h1)))
                begin
                  if (reg3153)
                    begin
                      reg3230 <= $signed($unsigned((reg3148[(1'h1):(1'h0)] <<< (reg3166 >= reg3189))));
                      reg3231 <= (forvar3206 ? $signed((8'h9e)) : reg3207);
                      reg3232 <= (+(~|(~|(~^forvar3139))));
                    end
                  else
                    begin
                      reg3230 <= $signed({$unsigned(((8'haa) ?
                              (8'ha8) : reg3161))});
                      reg3231 <= ($signed((!(reg3153 ?
                          reg3125 : forvar3132))) != ($signed($signed(reg3151)) ?
                          forvar3220 : $unsigned(((8'hb6) >= reg3172))));
                    end
                  reg3233 <= $unsigned(((^~reg3172) ?
                      reg3205[(1'h0):(1'h0)] : forvar3170));
                end
              if ((~^(8'hb1)))
                begin
                  for (forvar3234 = (1'h0); (forvar3234 < (1'h1)); forvar3234 = (forvar3234 + (1'h1)))
                    begin
                      reg3235 <= $signed(wire3121);
                    end
                  if ((reg3139 ?
                      (forvar3179 == ((+forvar3205) - reg3149[(2'h3):(2'h3)])) : forvar3191[(3'h6):(1'h0)]))
                    begin
                      reg3236 <= (reg3176[(2'h2):(1'h0)] ~^ {reg3187[(1'h1):(1'h0)]});
                      reg3237 <= reg3173[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg3236 <= forvar3234;
                      reg3237 <= $signed({((~^reg3124) >= (reg3145 ^~ (8'ha0)))});
                    end
                  for (forvar3238 = (1'h0); (forvar3238 < (1'h0)); forvar3238 = (forvar3238 + (1'h1)))
                    begin
                      reg3239 <= (((8'hb8) << reg3190) == ($signed(wire3120[(4'h8):(2'h2)]) ~^ (reg3185 == (^reg3218))));
                      reg3240 <= (reg3164[(3'h5):(2'h3)] ?
                          {$unsigned((~|reg3142))} : $signed(reg3204[(1'h1):(1'h0)]));
                      reg3241 <= $unsigned((~|{forvar3140[(3'h4):(3'h4)]}));
                      reg3242 <= reg3223;
                    end
                  for (forvar3243 = (1'h0); (forvar3243 < (1'h1)); forvar3243 = (forvar3243 + (1'h1)))
                    begin
                      reg3244 <= (reg3176 - forvar3225[(3'h6):(3'h4)]);
                    end
                end
              else
                begin
                  for (forvar3234 = (1'h0); (forvar3234 < (1'h1)); forvar3234 = (forvar3234 + (1'h1)))
                    begin
                      reg3235 <= (^{(|((8'haf) <<< forvar3190))});
                    end
                end
              if (({(~reg3232)} + reg3142))
                begin
                  if ((8'hb3))
                    begin
                      reg3245 <= ((forvar3179 ?
                          (~|((8'hab) < reg3237)) : ($unsigned(reg3163) <<< (reg3133 ?
                              reg3230 : (8'hb8)))) || (((-wire3121) >> (forvar3147 ?
                              reg3143 : forvar3221)) ?
                          ($unsigned(reg3235) ^~ (reg3191 ?
                              (8'hb5) : reg3175)) : $unsigned(reg3191[(1'h1):(1'h1)])));
                      reg3246 <= $signed((((+forvar3173) | (wire3122 ?
                              wire3122 : reg3128)) ?
                          {reg3203[(2'h3):(2'h3)]} : reg3193[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg3245 <= {{forvar3138}};
                      reg3246 <= forvar3159[(3'h4):(1'h1)];
                      reg3247 <= reg3129;
                    end
                  if (reg3141[(2'h3):(1'h1)])
                    begin
                      reg3248 <= (~&(($unsigned(forvar3170) ?
                          (-reg3194) : $signed(reg3246)) == ($unsigned(reg3228) == forvar3184[(2'h3):(1'h0)])));
                      reg3249 <= reg3159[(4'h9):(3'h5)];
                    end
                  else
                    begin
                      reg3248 <= reg3148;
                      reg3249 <= reg3195;
                      reg3250 <= {$unsigned($signed((forvar3220 ?
                              reg3163 : (8'hb0))))};
                      reg3251 <= $unsigned(reg3138[(2'h3):(2'h3)]);
                    end
                  for (forvar3252 = (1'h0); (forvar3252 < (1'h1)); forvar3252 = (forvar3252 + (1'h1)))
                    begin
                      reg3253 <= ($unsigned((~|(~^reg3125))) ?
                          forvar3169 : reg3143[(3'h4):(2'h3)]);
                      reg3254 <= {$signed(($unsigned(reg3168) & (reg3130 ?
                              forvar3143 : reg3213)))};
                    end
                  for (forvar3255 = (1'h0); (forvar3255 < (2'h2)); forvar3255 = (forvar3255 + (1'h1)))
                    begin
                      reg3256 <= reg3162;
                      reg3257 <= (~|(forvar3252 ?
                          $unsigned((~&reg3216)) : reg3247));
                    end
                end
              else
                begin
                  for (forvar3245 = (1'h0); (forvar3245 < (2'h3)); forvar3245 = (forvar3245 + (1'h1)))
                    begin
                      reg3246 <= {reg3176};
                      reg3247 <= (((|(8'h9f)) ^ ((reg3171 >= reg3173) ?
                              (^~reg3166) : reg3162[(4'hc):(4'h8)])) ?
                          $signed(((reg3197 | (8'hb6)) ?
                              forvar3188[(3'h7):(3'h4)] : {reg3127})) : ($unsigned(forvar3173) ?
                              {reg3201[(1'h1):(1'h1)]} : (wire3118[(2'h3):(1'h0)] ?
                                  {reg3245} : forvar3143)));
                      reg3248 <= reg3153[(4'hc):(3'h5)];
                    end
                  for (forvar3249 = (1'h0); (forvar3249 < (2'h3)); forvar3249 = (forvar3249 + (1'h1)))
                    begin
                      reg3250 <= ($signed((~&{reg3177})) ?
                          (!reg3134[(2'h2):(1'h1)]) : (($unsigned(forvar3205) * (8'ha9)) ?
                              ((8'hb4) ^ {reg3170}) : reg3180[(1'h0):(1'h0)]));
                      reg3251 <= ($signed(($signed(reg3226) <<< (forvar3159 <<< reg3145))) ?
                          (+((^~reg3205) >= (wire3118 ?
                              (8'hb8) : reg3242))) : (8'haf));
                      reg3252 <= reg3210;
                    end
                  for (forvar3253 = (1'h0); (forvar3253 < (2'h3)); forvar3253 = (forvar3253 + (1'h1)))
                    begin
                      reg3254 <= ($unsigned({reg3126}) ~^ reg3186);
                      reg3255 <= {(forvar3252 ?
                              $signed((forvar3156 != reg3169)) : {$signed(reg3161)})};
                      reg3256 <= $signed($signed(((reg3186 ?
                              (8'hb4) : reg3230) ?
                          (reg3166 + reg3251) : reg3257)));
                    end
                end
            end
          if ($unsigned({(~&$unsigned(reg3173))}))
            begin
              if (reg3159[(1'h0):(1'h0)])
                begin
                  if (reg3204[(3'h4):(3'h4)])
                    begin
                      reg3258 <= ($unsigned((forvar3252 ?
                          (reg3191 << reg3173) : $signed(reg3147))) > $signed($signed((|reg3177))));
                      reg3259 <= reg3163;
                      reg3260 <= {$unsigned($signed((~^(8'hae))))};
                      reg3261 <= (&$signed(reg3175));
                    end
                  else
                    begin
                      reg3258 <= (|reg3191);
                      reg3259 <= {((-{reg3181}) ? {{reg3158}} : {(~&reg3179)})};
                      reg3260 <= forvar3245[(1'h0):(1'h0)];
                    end
                  for (forvar3262 = (1'h0); (forvar3262 < (2'h2)); forvar3262 = (forvar3262 + (1'h1)))
                    begin
                      reg3263 <= $unsigned((reg3162[(4'ha):(3'h6)] ?
                          reg3252[(2'h2):(2'h2)] : (8'ha5)));
                    end
                end
              else
                begin
                  for (forvar3258 = (1'h0); (forvar3258 < (1'h1)); forvar3258 = (forvar3258 + (1'h1)))
                    begin
                      reg3259 <= $unsigned($unsigned(reg3261));
                      reg3260 <= $signed(reg3245[(4'h9):(4'h9)]);
                      reg3261 <= {$unsigned((~&(+reg3178)))};
                    end
                  for (forvar3262 = (1'h0); (forvar3262 < (1'h1)); forvar3262 = (forvar3262 + (1'h1)))
                    begin
                      reg3263 <= {($unsigned(forvar3159) != {$unsigned(reg3181)})};
                      reg3264 <= reg3205;
                    end
                end
              for (forvar3265 = (1'h0); (forvar3265 < (2'h3)); forvar3265 = (forvar3265 + (1'h1)))
                begin
                  for (forvar3266 = (1'h0); (forvar3266 < (2'h2)); forvar3266 = (forvar3266 + (1'h1)))
                    begin
                      reg3267 <= reg3241;
                      reg3268 <= (reg3204 >> (|$signed({forvar3172})));
                      reg3269 <= (reg3184[(4'hb):(1'h0)] ?
                          {$signed(reg3224[(2'h2):(2'h2)])} : ($signed($unsigned(forvar3164)) ?
                              {$signed(reg3203)} : (forvar3195[(1'h0):(1'h0)] | reg3198)));
                      reg3270 <= (forvar3252[(1'h0):(1'h0)] ?
                          (($unsigned((8'hb3)) * reg3123[(3'h6):(2'h3)]) ^ (forvar3197 ?
                              $signed(reg3160) : (forvar3129 ?
                                  forvar3265 : reg3175))) : (|reg3223[(3'h7):(3'h5)]));
                    end
                  for (forvar3271 = (1'h0); (forvar3271 < (1'h1)); forvar3271 = (forvar3271 + (1'h1)))
                    begin
                      reg3272 <= (({{reg3250}} ?
                              reg3208[(4'h9):(3'h6)] : reg3168[(1'h1):(1'h0)]) ?
                          ((8'ha1) & (|{(8'hab)})) : reg3167);
                      reg3273 <= forvar3139[(2'h2):(1'h1)];
                      reg3274 <= (reg3256 ?
                          $unsigned(forvar3253[(2'h2):(1'h1)]) : ($unsigned(forvar3245[(1'h0):(1'h0)]) ?
                              $unsigned((+(8'hb6))) : ((reg3206 ?
                                      forvar3262 : (8'ha1)) ?
                                  $signed(forvar3190) : ((8'hba) ?
                                      reg3256 : reg3197))));
                      reg3275 <= (reg3140[(4'h9):(4'h8)] ?
                          (~$unsigned(reg3203)) : ((8'had) >> {$signed(reg3128)}));
                    end
                  reg3276 <= $signed((~^((~^reg3176) ?
                      reg3236[(1'h1):(1'h0)] : (&reg3244))));
                end
              for (forvar3277 = (1'h0); (forvar3277 < (2'h3)); forvar3277 = (forvar3277 + (1'h1)))
                begin
                  if ($signed(($unsigned((reg3140 <<< forvar3140)) ?
                      ((-reg3255) ?
                          ((8'haa) << reg3202) : (~forvar3192)) : ($unsigned(reg3171) ?
                          reg3186[(3'h4):(1'h1)] : (~^reg3224)))))
                    begin
                      reg3278 <= ((($unsigned((8'ha8)) ?
                              {reg3207} : reg3180[(1'h1):(1'h1)]) && forvar3124[(3'h5):(1'h0)]) ?
                          reg3203 : $signed(reg3200[(3'h7):(3'h5)]));
                    end
                  else
                    begin
                      reg3278 <= (reg3217 ?
                          (~{(+forvar3152)}) : {(^(forvar3197 ?
                                  reg3224 : forvar3152))});
                    end
                end
            end
          else
            begin
              reg3258 <= (~|($signed(reg3192) < reg3194[(1'h1):(1'h1)]));
            end
        end
    end
  always
    @(posedge clk) begin
      reg3279 <= (~(8'ha2));
      reg3280 <= {wire3119};
    end
  assign wire3281 = (reg3185[(2'h3):(1'h0)] ? reg3125 : {forvar3188});
  always
    @(posedge clk) begin
      reg3282 <= forvar3157[(2'h2):(2'h2)];
      for (forvar3283 = (1'h0); (forvar3283 < (1'h1)); forvar3283 = (forvar3283 + (1'h1)))
        begin
          for (forvar3284 = (1'h0); (forvar3284 < (2'h3)); forvar3284 = (forvar3284 + (1'h1)))
            begin
              for (forvar3285 = (1'h0); (forvar3285 < (1'h0)); forvar3285 = (forvar3285 + (1'h1)))
                begin
                  if ($unsigned({($signed(forvar3262) + (reg3263 | reg3207))}))
                    begin
                      reg3286 <= {(8'h9c)};
                      reg3287 <= ((+$signed(reg3194[(1'h1):(1'h0)])) - forvar3271[(3'h4):(2'h2)]);
                      reg3288 <= $unsigned($signed(((~|(8'h9f)) - $unsigned(reg3146))));
                    end
                  else
                    begin
                      reg3286 <= $signed(reg3125[(3'h5):(2'h3)]);
                      reg3287 <= reg3181;
                      reg3288 <= reg3189[(3'h7):(2'h3)];
                      reg3289 <= reg3147[(4'hc):(3'h6)];
                    end
                end
            end
          for (forvar3290 = (1'h0); (forvar3290 < (2'h3)); forvar3290 = (forvar3290 + (1'h1)))
            begin
              if ((^reg3208[(4'hb):(3'h4)]))
                begin
                  if ((+(-((~^reg3195) ~^ ((8'ha0) <<< reg3202)))))
                    begin
                      reg3291 <= reg3201;
                    end
                  else
                    begin
                      reg3291 <= $signed($unsigned({reg3151}));
                      reg3292 <= (($signed($signed(reg3273)) >> (|$signed(reg3248))) ?
                          ($signed(reg3174[(4'h9):(1'h1)]) ?
                              ({forvar3206} ?
                                  $signed(wire3121) : $signed((8'ha4))) : $signed((reg3147 != reg3216))) : reg3180[(2'h2):(2'h2)]);
                      reg3293 <= (($signed((reg3255 ?
                              reg3191 : forvar3170)) - ({reg3195} ?
                              {(8'haf)} : {reg3148})) ?
                          (^{(forvar3195 > reg3141)}) : $unsigned(reg3174));
                    end
                  for (forvar3294 = (1'h0); (forvar3294 < (1'h1)); forvar3294 = (forvar3294 + (1'h1)))
                    begin
                      reg3295 <= $signed((~($unsigned(reg3268) ?
                          (reg3141 == reg3173) : (|(8'hba)))));
                    end
                  reg3296 <= (reg3254[(2'h3):(1'h1)] ?
                      reg3143[(3'h6):(2'h2)] : (reg3204 | $unsigned((&forvar3229))));
                end
              else
                begin
                  for (forvar3291 = (1'h0); (forvar3291 < (2'h3)); forvar3291 = (forvar3291 + (1'h1)))
                    begin
                      reg3292 <= $unsigned(($signed({reg3127}) ?
                          $unsigned($signed(forvar3229)) : $signed((reg3134 * forvar3190))));
                      reg3293 <= reg3206[(4'h8):(2'h2)];
                    end
                  if ((reg3143 ?
                      $unsigned({(reg3168 * reg3168)}) : $unsigned((~|(reg3130 ?
                          reg3223 : forvar3125)))))
                    begin
                      reg3294 <= (reg3264[(4'ha):(1'h0)] || $signed(reg3211));
                    end
                  else
                    begin
                      reg3294 <= wire3121;
                      reg3295 <= $signed((((8'haf) & {forvar3172}) ~^ (&$unsigned(reg3191))));
                    end
                end
              for (forvar3297 = (1'h0); (forvar3297 < (1'h0)); forvar3297 = (forvar3297 + (1'h1)))
                begin
                  for (forvar3298 = (1'h0); (forvar3298 < (1'h1)); forvar3298 = (forvar3298 + (1'h1)))
                    begin
                      reg3299 <= ((+((forvar3297 && forvar3220) ?
                          (reg3247 ? forvar3191 : wire3121) : (reg3247 ?
                              (8'hb0) : reg3178))) << reg3149[(3'h5):(2'h3)]);
                      reg3300 <= reg3223;
                      reg3301 <= reg3237[(3'h6):(3'h5)];
                      reg3302 <= $unsigned({(&reg3130)});
                    end
                  for (forvar3303 = (1'h0); (forvar3303 < (1'h0)); forvar3303 = (forvar3303 + (1'h1)))
                    begin
                      reg3304 <= reg3237;
                    end
                  reg3305 <= $signed($unsigned($signed((reg3194 ?
                      forvar3252 : (8'hab)))));
                end
              reg3306 <= $unsigned((+((&(8'ha9)) >= $unsigned(reg3155))));
            end
          for (forvar3307 = (1'h0); (forvar3307 < (1'h1)); forvar3307 = (forvar3307 + (1'h1)))
            begin
              for (forvar3308 = (1'h0); (forvar3308 < (2'h3)); forvar3308 = (forvar3308 + (1'h1)))
                begin
                  reg3309 <= (~|$signed(reg3293));
                end
              for (forvar3310 = (1'h0); (forvar3310 < (2'h2)); forvar3310 = (forvar3310 + (1'h1)))
                begin
                  reg3311 <= {$signed(($unsigned(forvar3140) ^ reg3147[(4'h9):(4'h9)]))};
                end
              for (forvar3312 = (1'h0); (forvar3312 < (2'h3)); forvar3312 = (forvar3312 + (1'h1)))
                begin
                  if (reg3253)
                    begin
                      reg3313 <= reg3181[(4'hd):(1'h0)];
                      reg3314 <= ((reg3129[(4'h8):(3'h7)] < $signed(forvar3238)) ?
                          (+$unsigned((8'ha7))) : {reg3224[(2'h2):(1'h1)]});
                      reg3315 <= (-{$unsigned((reg3153 <<< reg3264))});
                    end
                  else
                    begin
                      reg3313 <= forvar3238;
                      reg3314 <= (~&(&$unsigned(reg3314[(4'h9):(4'h9)])));
                      reg3315 <= (&{((8'hb4) ?
                              $signed((8'hb4)) : reg3263[(4'hb):(4'h9)])});
                      reg3316 <= (forvar3277 >= ((forvar3283 ?
                          reg3198 : (reg3185 | reg3274)) >> (&$signed(reg3239))));
                    end
                  for (forvar3317 = (1'h0); (forvar3317 < (2'h3)); forvar3317 = (forvar3317 + (1'h1)))
                    begin
                      reg3318 <= (~&forvar3143);
                    end
                  if ((~{(reg3276[(2'h3):(1'h1)] == (reg3149 ?
                          reg3179 : reg3252))}))
                    begin
                      reg3319 <= ($unsigned($unsigned($signed(reg3292))) || reg3250[(2'h3):(1'h1)]);
                      reg3320 <= {(~((reg3257 ^~ reg3199) <<< $unsigned(reg3299)))};
                      reg3321 <= reg3257;
                    end
                  else
                    begin
                      reg3319 <= ((((reg3142 >> reg3309) & (reg3142 ?
                                  forvar3290 : reg3184)) ?
                              reg3190[(3'h6):(3'h6)] : {reg3245[(3'h7):(3'h6)]}) ?
                          wire3120[(3'h5):(2'h2)] : reg3240[(2'h2):(1'h0)]);
                      reg3320 <= $unsigned($unsigned((!reg3131)));
                    end
                end
            end
        end
      if ({reg3193[(1'h1):(1'h1)]})
        begin
          for (forvar3322 = (1'h0); (forvar3322 < (2'h3)); forvar3322 = (forvar3322 + (1'h1)))
            begin
              reg3323 <= $signed(wire3122);
            end
        end
      else
        begin
          for (forvar3322 = (1'h0); (forvar3322 < (1'h0)); forvar3322 = (forvar3322 + (1'h1)))
            begin
              for (forvar3323 = (1'h0); (forvar3323 < (2'h3)); forvar3323 = (forvar3323 + (1'h1)))
                begin
                  if ($unsigned(forvar3144[(4'he):(4'h8)]))
                    begin
                      reg3324 <= $signed(($signed((reg3171 <= reg3279)) * forvar3308));
                      reg3325 <= {reg3233[(3'h5):(2'h2)]};
                      reg3326 <= (^(reg3210[(2'h2):(2'h2)] < (^~((8'hb5) ^ reg3240))));
                    end
                  else
                    begin
                      reg3324 <= (((~|{(8'ha5)}) ?
                          (~$unsigned((8'h9d))) : (8'hb6)) <<< $unsigned((~(&(8'hac)))));
                      reg3325 <= (|(forvar3262[(4'he):(3'h5)] ^~ ((!reg3319) >>> (reg3173 && reg3268))));
                      reg3326 <= (-$signed(reg3227));
                      reg3327 <= forvar3129;
                    end
                  reg3328 <= (!reg3228);
                end
            end
          for (forvar3329 = (1'h0); (forvar3329 < (2'h3)); forvar3329 = (forvar3329 + (1'h1)))
            begin
              reg3330 <= (($unsigned((reg3232 < reg3321)) ?
                      ((reg3202 ?
                          reg3207 : (8'ha2)) ^~ (forvar3159 && reg3274)) : reg3137) ?
                  (~&$unsigned(((8'hab) >> (8'hb0)))) : $signed($unsigned((^~forvar3329))));
              reg3331 <= $unsigned((-{$unsigned(reg3206)}));
            end
        end
      for (forvar3332 = (1'h0); (forvar3332 < (1'h1)); forvar3332 = (forvar3332 + (1'h1)))
        begin
          if ((~&forvar3147[(1'h0):(1'h0)]))
            begin
              if (forvar3156[(1'h0):(1'h0)])
                begin
                  for (forvar3333 = (1'h0); (forvar3333 < (1'h0)); forvar3333 = (forvar3333 + (1'h1)))
                    begin
                      reg3334 <= $unsigned(reg3313[(2'h3):(1'h0)]);
                      reg3335 <= forvar3157;
                      reg3336 <= $signed((~{forvar3249[(1'h1):(1'h0)]}));
                    end
                end
              else
                begin
                  for (forvar3333 = (1'h0); (forvar3333 < (1'h1)); forvar3333 = (forvar3333 + (1'h1)))
                    begin
                      reg3334 <= $signed(({{reg3264}} ?
                          (^~{reg3160}) : (8'h9f)));
                      reg3335 <= reg3199;
                      reg3336 <= (!(($signed(forvar3225) && (reg3325 ?
                              forvar3173 : (8'hba))) ?
                          $signed((reg3209 ^~ (8'hba))) : ((~^reg3247) >> $unsigned(forvar3310))));
                    end
                  if ((~^forvar3265))
                    begin
                      reg3337 <= $signed(reg3272);
                      reg3338 <= ($unsigned((reg3206[(3'h7):(2'h3)] ^~ reg3208[(4'h9):(4'h8)])) && (8'ha7));
                      reg3339 <= $signed(((!(8'hb6)) ?
                          (-(reg3208 ?
                              (8'hb3) : reg3269)) : $unsigned((forvar3142 ^~ forvar3192))));
                    end
                  else
                    begin
                      reg3337 <= (&$signed($unsigned((reg3324 ?
                          (8'hae) : reg3311))));
                      reg3338 <= $unsigned((((!forvar3329) ?
                              (-reg3195) : $signed(forvar3170)) ?
                          $signed((~&reg3230)) : forvar3205));
                    end
                  if ((reg3159[(4'h8):(3'h4)] >> $signed(reg3176[(1'h1):(1'h1)])))
                    begin
                      reg3340 <= reg3248[(2'h3):(2'h2)];
                      reg3341 <= $signed((((^reg3155) & forvar3297[(2'h2):(2'h2)]) ?
                          (8'hb9) : $unsigned(forvar3131[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg3340 <= ($unsigned(($signed(reg3184) | ((8'hb2) * reg3301))) < reg3201);
                    end
                end
              for (forvar3342 = (1'h0); (forvar3342 < (1'h1)); forvar3342 = (forvar3342 + (1'h1)))
                begin
                  reg3343 <= forvar3137[(4'h8):(2'h2)];
                  reg3344 <= (|(({reg3148} ?
                          (forvar3290 ? reg3245 : reg3135) : {reg3168}) ?
                      ((^reg3252) * reg3149[(1'h1):(1'h0)]) : (&(|reg3208))));
                  for (forvar3345 = (1'h0); (forvar3345 < (2'h3)); forvar3345 = (forvar3345 + (1'h1)))
                    begin
                      reg3346 <= $unsigned({reg3231});
                      reg3347 <= (~&((&(!reg3343)) >>> $signed((reg3192 ?
                          reg3137 : reg3154))));
                      reg3348 <= $unsigned((((forvar3284 >= reg3128) ?
                          reg3158 : ((8'ha2) ?
                              forvar3345 : reg3301)) & (reg3325[(1'h1):(1'h1)] <<< reg3219)));
                      reg3349 <= $signed((~&forvar3170));
                    end
                  if ($signed((reg3280 && forvar3134[(1'h0):(1'h0)])))
                    begin
                      reg3350 <= (($unsigned(reg3237) ?
                          $signed(((8'hb4) ?
                              forvar3222 : forvar3190)) : $signed((reg3319 ?
                              forvar3297 : forvar3188))) ~^ $unsigned(({(8'h9e)} >> (reg3203 ~^ reg3172))));
                      reg3351 <= ($unsigned($unsigned((reg3190 ?
                              reg3136 : reg3269))) ?
                          $signed(reg3213[(4'ha):(3'h7)]) : $unsigned($signed((forvar3225 ?
                              reg3142 : reg3179))));
                    end
                  else
                    begin
                      reg3350 <= (8'ha0);
                      reg3351 <= (8'ha1);
                    end
                end
              reg3352 <= $signed((forvar3169 ? forvar3187 : {(~^reg3275)}));
              for (forvar3353 = (1'h0); (forvar3353 < (2'h3)); forvar3353 = (forvar3353 + (1'h1)))
                begin
                  reg3354 <= {$unsigned({((8'ha4) ? reg3260 : (8'ha4))})};
                  if (reg3319)
                    begin
                      reg3355 <= (|reg3137[(4'ha):(3'h6)]);
                      reg3356 <= (~|$unsigned($signed((~^forvar3253))));
                      reg3357 <= (|($unsigned((^forvar3124)) << (!(reg3177 ?
                          (8'ha0) : reg3204))));
                    end
                  else
                    begin
                      reg3355 <= ($unsigned(reg3167[(4'he):(3'h7)]) >= ($unsigned($unsigned(reg3256)) ?
                          {(~&wire3121)} : $signed($signed(reg3140))));
                    end
                  if ((8'ha3))
                    begin
                      reg3358 <= ((8'hb4) | (^($signed(reg3232) ^~ $signed(reg3130))));
                    end
                  else
                    begin
                      reg3358 <= reg3251;
                    end
                  reg3359 <= reg3252;
                end
            end
          else
            begin
              for (forvar3333 = (1'h0); (forvar3333 < (1'h1)); forvar3333 = (forvar3333 + (1'h1)))
                begin
                  if ($unsigned(forvar3142[(2'h3):(1'h1)]))
                    begin
                      reg3334 <= (((!reg3314) <= ((reg3191 ?
                          forvar3312 : reg3170) >= reg3273)) <<< forvar3308[(3'h6):(3'h4)]);
                      reg3335 <= $unsigned($signed($unsigned($unsigned(forvar3312))));
                      reg3336 <= ({((^~reg3341) >>> {reg3288})} >> $unsigned(reg3208));
                      reg3337 <= ($signed(forvar3308[(3'h5):(3'h4)]) ?
                          (((~&forvar3156) ? $unsigned(reg3343) : reg3125) ?
                              reg3230 : $signed((reg3339 ?
                                  reg3193 : reg3193))) : $unsigned({{reg3244}}));
                    end
                  else
                    begin
                      reg3334 <= $signed((^(reg3301[(3'h4):(1'h1)] ?
                          $signed(reg3327) : forvar3221[(4'h8):(3'h4)])));
                    end
                  for (forvar3338 = (1'h0); (forvar3338 < (1'h1)); forvar3338 = (forvar3338 + (1'h1)))
                    begin
                      reg3339 <= ((^((reg3196 ? reg3133 : forvar3129) ?
                              $signed(reg3249) : ((8'hb2) ?
                                  reg3164 : reg3319))) ?
                          forvar3140 : ((-$unsigned(reg3195)) ?
                              forvar3284[(4'h8):(3'h6)] : {$signed((8'h9e))}));
                      reg3340 <= reg3227;
                      reg3341 <= (((&forvar3195) ^~ reg3130) ?
                          reg3144 : forvar3187);
                    end
                end
              if (((8'hb6) < (8'hab)))
                begin
                  if ((^~reg3198[(4'h8):(3'h6)]))
                    begin
                      reg3342 <= {$unsigned(forvar3222)};
                      reg3343 <= ({{(reg3305 ? reg3342 : forvar3147)}} ?
                          reg3136[(1'h0):(1'h0)] : (8'h9d));
                    end
                  else
                    begin
                      reg3342 <= ($signed(($unsigned(reg3161) - {reg3327})) || (|(-$signed((8'ha0)))));
                      reg3343 <= $signed((~|{(reg3264 ? reg3138 : reg3200)}));
                    end
                  reg3344 <= (($signed((reg3245 ? reg3305 : reg3166)) ?
                      reg3293 : forvar3308[(3'h6):(3'h4)]) ^ {{$unsigned(reg3288)}});
                end
              else
                begin
                  if ($signed(reg3325[(1'h1):(1'h0)]))
                    begin
                      reg3342 <= $signed({reg3257[(4'h8):(3'h4)]});
                      reg3343 <= (8'hae);
                    end
                  else
                    begin
                      reg3342 <= forvar3265;
                      reg3343 <= $signed(forvar3187[(4'hf):(3'h7)]);
                      reg3344 <= $signed(($signed((reg3202 ~^ reg3149)) && ($signed(reg3198) ?
                          (reg3313 ? reg3132 : reg3146) : (forvar3179 ?
                              forvar3285 : reg3258))));
                      reg3345 <= (^~reg3125[(3'h4):(2'h3)]);
                    end
                  if ((|{$signed($signed((8'hac)))}))
                    begin
                      reg3346 <= reg3208;
                      reg3347 <= reg3158[(2'h3):(2'h2)];
                      reg3348 <= forvar3322[(1'h1):(1'h1)];
                      reg3349 <= (($signed($unsigned(forvar3190)) ?
                              (-reg3301) : ($unsigned(reg3189) >> $unsigned(reg3128))) ?
                          reg3259[(2'h3):(2'h3)] : $unsigned($signed((reg3335 ?
                              reg3276 : reg3141))));
                    end
                  else
                    begin
                      reg3346 <= (reg3304 ?
                          reg3273[(1'h1):(1'h0)] : ($signed((&reg3249)) | ({wire3121} ~^ {reg3126})));
                      reg3347 <= {((reg3138[(3'h7):(3'h4)] ?
                              {forvar3195} : $unsigned(reg3157)) != reg3351)};
                      reg3348 <= $signed(($unsigned((8'h9f)) & ($signed(reg3346) ?
                          (+reg3154) : (reg3344 | forvar3134))));
                      reg3349 <= $unsigned($signed($unsigned((+reg3305))));
                    end
                  for (forvar3350 = (1'h0); (forvar3350 < (1'h0)); forvar3350 = (forvar3350 + (1'h1)))
                    begin
                      reg3351 <= (+$signed({$unsigned(reg3197)}));
                    end
                  if ((8'h9e))
                    begin
                      reg3352 <= (reg3163[(3'h4):(2'h3)] & {{(~&reg3261)}});
                      reg3353 <= {$unsigned(reg3339)};
                      reg3354 <= $unsigned(($unsigned($unsigned(reg3349)) < $signed((!reg3138))));
                    end
                  else
                    begin
                      reg3352 <= (8'ha7);
                      reg3353 <= ($unsigned($unsigned((reg3353 ?
                              forvar3188 : reg3244))) ?
                          $signed(reg3183[(4'ha):(4'ha)]) : $signed((reg3172[(3'h4):(3'h4)] * (forvar3350 ?
                              reg3181 : reg3223))));
                      reg3354 <= $unsigned((reg3184 ?
                          $signed({(8'ha5)}) : (^reg3204[(3'h4):(2'h3)])));
                      reg3355 <= $signed($signed(reg3235));
                    end
                end
              reg3356 <= forvar3303[(1'h1):(1'h1)];
              for (forvar3357 = (1'h0); (forvar3357 < (2'h2)); forvar3357 = (forvar3357 + (1'h1)))
                begin
                  reg3358 <= ({$unsigned((~^reg3253))} < (forvar3169[(2'h2):(1'h0)] * (forvar3125 != $signed(reg3248))));
                  if (reg3218[(1'h0):(1'h0)])
                    begin
                      reg3359 <= {$unsigned(reg3217)};
                      reg3360 <= (~|$unsigned($unsigned({reg3294})));
                      reg3361 <= forvar3243;
                    end
                  else
                    begin
                      reg3359 <= reg3309[(1'h0):(1'h0)];
                      reg3360 <= reg3207[(4'h9):(3'h7)];
                    end
                  if (reg3323[(2'h3):(2'h2)])
                    begin
                      reg3362 <= $unsigned($signed((~$signed(reg3276))));
                      reg3363 <= {$unsigned((reg3197[(1'h1):(1'h1)] & reg3306[(4'hc):(3'h5)]))};
                    end
                  else
                    begin
                      reg3362 <= (forvar3323[(2'h2):(2'h2)] ?
                          $unsigned({reg3191[(3'h5):(1'h1)]}) : {$signed((&reg3258))});
                      reg3363 <= {{((|reg3323) != $signed((8'ha8)))}};
                      reg3364 <= ($signed(forvar3262[(4'hb):(4'h8)]) <= (!$unsigned((-reg3189))));
                      reg3365 <= reg3180[(1'h0):(1'h0)];
                    end
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3769
#( parameter param4729 = (((((8'hb5) >>> (8'hb7)) >= ((8'hb6) <= (8'haf))) ? ((+(8'h9f)) - {(8'h9d)}) : (((8'hb7) != (8'ha6)) ? (8'hb4) : (!(8'ha4)))) ? ((((8'hb9) <= (8'ha4)) > (-(8'had))) ? {{(8'hb6)}} : ({(8'hb1)} ? ((8'hae) & (8'ha0)) : ((8'hb7) ^ (8'ha3)))) : (+(((8'hab) >> (8'hb4)) ? ((8'ha8) ? (8'ha2) : (8'haf)) : ((8'hb2) < (8'hb2))))) )
(y, clk, wire3773, wire3772, wire3771, wire3770);
  output wire [(32'hb6d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire3773;
  input wire signed [(4'h9):(1'h0)] wire3772;
  input wire signed [(5'h10):(1'h0)] wire3771;
  input wire [(4'h8):(1'h0)] wire3770;
  reg signed [(4'hf):(1'h0)] reg4728 = (1'h0);
  reg [(4'he):(1'h0)] reg4727 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4726 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4725 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4724 = (1'h0);
  reg [(3'h6):(1'h0)] reg4723 = (1'h0);
  reg [(4'h9):(1'h0)] reg4722 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4721 = (1'h0);
  reg [(4'hb):(1'h0)] reg4720 = (1'h0);
  reg [(5'h10):(1'h0)] reg4719 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4718 = (1'h0);
  reg [(3'h6):(1'h0)] reg4717 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4716 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4715 = (1'h0);
  reg [(4'he):(1'h0)] forvar4714 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4713 = (1'h0);
  reg [(4'hd):(1'h0)] reg4712 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4711 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4710 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4709 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4708 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4707 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4706 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4705 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4704 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4703 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4702 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4701 = (1'h0);
  reg [(4'he):(1'h0)] forvar4700 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4699 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4698 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4697 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4696 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4695 = (1'h0);
  reg [(2'h2):(1'h0)] reg4694 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4693 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4692 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4691 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4690 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4689 = (1'h0);
  reg [(4'he):(1'h0)] reg4688 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4687 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4686 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4685 = (1'h0);
  reg [(3'h7):(1'h0)] reg4684 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4683 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4682 = (1'h0);
  reg [(3'h7):(1'h0)] reg4681 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4680 = (1'h0);
  reg [(5'h10):(1'h0)] reg4679 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4678 = (1'h0);
  reg [(3'h7):(1'h0)] reg4677 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4676 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4675 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4674 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4673 = (1'h0);
  reg [(4'hc):(1'h0)] reg4672 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4671 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4670 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4663 = (1'h0);
  reg [(3'h5):(1'h0)] reg4669 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4668 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4667 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4666 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4665 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4664 = (1'h0);
  reg [(5'h10):(1'h0)] reg4663 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4662 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4661 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4660 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4659 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4658 = (1'h0);
  reg [(2'h3):(1'h0)] reg4657 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4656 = (1'h0);
  reg [(3'h4):(1'h0)] reg4655 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4654 = (1'h0);
  reg [(4'h8):(1'h0)] reg4653 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4652 = (1'h0);
  reg [(4'h8):(1'h0)] reg4651 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4650 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4649 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4648 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4647 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4646 = (1'h0);
  reg [(3'h7):(1'h0)] reg4645 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4644 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4643 = (1'h0);
  reg [(4'hd):(1'h0)] reg4642 = (1'h0);
  reg [(4'hd):(1'h0)] reg4641 = (1'h0);
  reg [(4'hf):(1'h0)] reg4640 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4639 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4638 = (1'h0);
  reg [(3'h5):(1'h0)] reg4637 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4636 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4635 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4625 = (1'h0);
  reg [(3'h6):(1'h0)] reg4624 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4621 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4634 = (1'h0);
  reg [(4'hd):(1'h0)] reg4633 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4632 = (1'h0);
  reg [(4'hc):(1'h0)] reg4631 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4630 = (1'h0);
  reg [(4'ha):(1'h0)] reg4629 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4628 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4627 = (1'h0);
  reg [(4'ha):(1'h0)] reg4626 = (1'h0);
  reg [(5'h10):(1'h0)] reg4625 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4624 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4623 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4622 = (1'h0);
  reg [(3'h6):(1'h0)] reg4621 = (1'h0);
  reg [(2'h2):(1'h0)] reg4620 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4619 = (1'h0);
  reg [(4'hc):(1'h0)] reg4618 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4617 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4614 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4611 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4610 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4607 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4604 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4593 = (1'h0);
  reg [(3'h5):(1'h0)] reg4609 = (1'h0);
  reg [(4'hc):(1'h0)] reg4606 = (1'h0);
  reg [(2'h2):(1'h0)] reg4605 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4603 = (1'h0);
  reg [(4'he):(1'h0)] forvar4602 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4600 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4597 = (1'h0);
  reg [(4'he):(1'h0)] forvar4596 = (1'h0);
  reg [(4'hb):(1'h0)] reg4594 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4592 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4616 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4615 = (1'h0);
  reg [(4'he):(1'h0)] reg4614 = (1'h0);
  reg [(4'hf):(1'h0)] reg4613 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4612 = (1'h0);
  reg [(4'hf):(1'h0)] reg4611 = (1'h0);
  reg [(4'hb):(1'h0)] reg4610 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4609 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4608 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4607 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4606 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4605 = (1'h0);
  reg [(2'h2):(1'h0)] reg4604 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4603 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4602 = (1'h0);
  reg [(5'h10):(1'h0)] reg4601 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4600 = (1'h0);
  reg [(4'ha):(1'h0)] reg4599 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4598 = (1'h0);
  reg [(4'hf):(1'h0)] reg4598 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4597 = (1'h0);
  reg [(4'hd):(1'h0)] reg4596 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4595 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4594 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4593 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4592 = (1'h0);
  reg [(4'h8):(1'h0)] reg4591 = (1'h0);
  reg [(4'ha):(1'h0)] reg4590 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4589 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4588 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire4587;
  reg [(2'h2):(1'h0)] reg4586 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4585 = (1'h0);
  reg [(4'hf):(1'h0)] reg4581 = (1'h0);
  reg [(3'h5):(1'h0)] reg4584 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4583 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4582 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4581 = (1'h0);
  reg [(2'h2):(1'h0)] reg4580 = (1'h0);
  reg [(3'h4):(1'h0)] reg4579 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4578 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4577 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4576 = (1'h0);
  reg [(3'h6):(1'h0)] reg4575 = (1'h0);
  reg [(3'h6):(1'h0)] reg4574 = (1'h0);
  reg [(4'h9):(1'h0)] reg4573 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4572 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4569 = (1'h0);
  reg [(2'h2):(1'h0)] reg4572 = (1'h0);
  reg [(4'hf):(1'h0)] reg4571 = (1'h0);
  reg [(4'hb):(1'h0)] reg4570 = (1'h0);
  reg [(4'hb):(1'h0)] reg4569 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4563 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4568 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4567 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4566 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4565 = (1'h0);
  reg [(4'hd):(1'h0)] reg4564 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4563 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4552 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4562 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4561 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4560 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4559 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4558 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4557 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4556 = (1'h0);
  reg [(2'h3):(1'h0)] reg4555 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4554 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4553 = (1'h0);
  reg [(3'h7):(1'h0)] reg4552 = (1'h0);
  reg [(4'hb):(1'h0)] reg4551 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4550 = (1'h0);
  reg [(4'he):(1'h0)] reg4549 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4548 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4547 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4546 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4545 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4544 = (1'h0);
  reg [(3'h4):(1'h0)] reg4543 = (1'h0);
  reg [(3'h5):(1'h0)] reg4542 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4541 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4540 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4539 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4538 = (1'h0);
  reg [(5'h10):(1'h0)] reg4537 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4536 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4536 = (1'h0);
  reg [(4'he):(1'h0)] reg4535 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4534 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4533 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4532 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4531 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4530 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4529 = (1'h0);
  reg [(2'h2):(1'h0)] reg4528 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4527 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4526 = (1'h0);
  reg [(4'h8):(1'h0)] reg4525 = (1'h0);
  reg [(3'h7):(1'h0)] reg4524 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4523 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4522 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4521 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4520 = (1'h0);
  reg [(4'hd):(1'h0)] reg4519 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4518 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4517 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4516 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4515 = (1'h0);
  reg [(4'hc):(1'h0)] reg4514 = (1'h0);
  reg [(5'h10):(1'h0)] reg4513 = (1'h0);
  reg [(4'hf):(1'h0)] reg4512 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4511 = (1'h0);
  reg [(4'h8):(1'h0)] reg4510 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4509 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4508 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4507 = (1'h0);
  reg [(4'hc):(1'h0)] reg4506 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4503 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4497 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4495 = (1'h0);
  reg [(3'h4):(1'h0)] reg4494 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4491 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4483 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4480 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4471 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4478 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4470 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4466 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4461 = (1'h0);
  reg [(4'hb):(1'h0)] reg4499 = (1'h0);
  reg [(4'ha):(1'h0)] reg4505 = (1'h0);
  reg [(4'hd):(1'h0)] reg4504 = (1'h0);
  reg [(4'h8):(1'h0)] reg4503 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4502 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4501 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4500 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4499 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4498 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4497 = (1'h0);
  reg [(3'h6):(1'h0)] reg4496 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4489 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4485 = (1'h0);
  reg [(4'hd):(1'h0)] reg4484 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4482 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4477 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4475 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4495 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4494 = (1'h0);
  reg [(3'h5):(1'h0)] reg4493 = (1'h0);
  reg [(4'hf):(1'h0)] reg4492 = (1'h0);
  reg [(3'h6):(1'h0)] reg4491 = (1'h0);
  reg [(5'h10):(1'h0)] reg4490 = (1'h0);
  reg [(3'h7):(1'h0)] reg4489 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4488 = (1'h0);
  reg [(2'h2):(1'h0)] reg4487 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4486 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4485 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4484 = (1'h0);
  reg [(4'he):(1'h0)] reg4483 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4482 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4481 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4480 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4479 = (1'h0);
  reg [(3'h6):(1'h0)] reg4478 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4477 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4476 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4475 = (1'h0);
  reg [(2'h2):(1'h0)] reg4474 = (1'h0);
  reg [(4'hf):(1'h0)] reg4473 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4472 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4471 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4470 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4469 = (1'h0);
  reg [(4'hd):(1'h0)] reg4468 = (1'h0);
  reg [(4'hf):(1'h0)] reg4467 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4466 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4465 = (1'h0);
  reg [(4'hb):(1'h0)] reg4464 = (1'h0);
  reg [(4'he):(1'h0)] reg4463 = (1'h0);
  reg [(4'hc):(1'h0)] reg4462 = (1'h0);
  reg [(2'h3):(1'h0)] reg4461 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4460 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4459 = (1'h0);
  wire [(4'hf):(1'h0)] wire4457;
  reg [(4'he):(1'h0)] reg3779 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire3778;
  wire signed [(4'h9):(1'h0)] wire3777;
  wire signed [(4'hf):(1'h0)] wire3776;
  wire signed [(4'hd):(1'h0)] wire3775;
  wire [(5'h10):(1'h0)] wire3774;
  assign y = {reg4728,
                 reg4727,
                 reg4726,
                 reg4725,
                 reg4724,
                 reg4723,
                 reg4722,
                 forvar4721,
                 reg4720,
                 reg4719,
                 reg4718,
                 reg4717,
                 reg4716,
                 reg4715,
                 forvar4714,
                 forvar4713,
                 reg4712,
                 reg4711,
                 reg4710,
                 forvar4709,
                 reg4708,
                 reg4707,
                 forvar4706,
                 forvar4705,
                 forvar4704,
                 reg4703,
                 forvar4702,
                 reg4701,
                 forvar4700,
                 reg4699,
                 reg4698,
                 reg4697,
                 reg4696,
                 forvar4695,
                 reg4694,
                 reg4693,
                 reg4692,
                 reg4691,
                 reg4690,
                 forvar4689,
                 reg4688,
                 forvar4687,
                 reg4686,
                 reg4685,
                 reg4684,
                 forvar4683,
                 reg4682,
                 reg4681,
                 reg4680,
                 reg4679,
                 forvar4678,
                 reg4677,
                 reg4676,
                 reg4675,
                 forvar4674,
                 reg4673,
                 reg4672,
                 forvar4671,
                 reg4670,
                 forvar4663,
                 reg4669,
                 reg4668,
                 forvar4667,
                 reg4666,
                 reg4665,
                 reg4664,
                 reg4663,
                 reg4662,
                 forvar4661,
                 forvar4660,
                 forvar4659,
                 forvar4658,
                 reg4657,
                 reg4656,
                 reg4655,
                 reg4654,
                 reg4653,
                 reg4652,
                 reg4651,
                 forvar4650,
                 forvar4649,
                 reg4648,
                 reg4647,
                 reg4646,
                 reg4645,
                 reg4644,
                 reg4643,
                 reg4642,
                 reg4641,
                 reg4640,
                 reg4639,
                 reg4638,
                 reg4637,
                 reg4636,
                 forvar4635,
                 forvar4625,
                 reg4624,
                 forvar4621,
                 reg4634,
                 reg4633,
                 reg4632,
                 reg4631,
                 reg4630,
                 reg4629,
                 reg4628,
                 reg4627,
                 reg4626,
                 reg4625,
                 forvar4624,
                 reg4623,
                 reg4622,
                 reg4621,
                 reg4620,
                 forvar4619,
                 reg4618,
                 reg4617,
                 forvar4614,
                 forvar4611,
                 forvar4610,
                 forvar4607,
                 forvar4604,
                 forvar4593,
                 reg4609,
                 reg4606,
                 reg4605,
                 forvar4603,
                 forvar4602,
                 reg4600,
                 forvar4597,
                 forvar4596,
                 reg4594,
                 reg4592,
                 reg4616,
                 reg4615,
                 reg4614,
                 reg4613,
                 reg4612,
                 reg4611,
                 reg4610,
                 forvar4609,
                 reg4608,
                 reg4607,
                 forvar4606,
                 forvar4605,
                 reg4604,
                 reg4603,
                 reg4602,
                 reg4601,
                 forvar4600,
                 reg4599,
                 forvar4598,
                 reg4598,
                 reg4597,
                 reg4596,
                 reg4595,
                 forvar4594,
                 reg4593,
                 forvar4592,
                 reg4591,
                 reg4590,
                 forvar4589,
                 forvar4588,
                 wire4587,
                 reg4586,
                 reg4585,
                 reg4581,
                 reg4584,
                 reg4583,
                 reg4582,
                 forvar4581,
                 reg4580,
                 reg4579,
                 reg4578,
                 reg4577,
                 reg4576,
                 reg4575,
                 reg4574,
                 reg4573,
                 forvar4572,
                 forvar4569,
                 reg4572,
                 reg4571,
                 reg4570,
                 reg4569,
                 forvar4563,
                 reg4568,
                 reg4567,
                 reg4566,
                 reg4565,
                 reg4564,
                 reg4563,
                 forvar4552,
                 reg4562,
                 reg4561,
                 reg4560,
                 reg4559,
                 reg4558,
                 forvar4557,
                 reg4556,
                 reg4555,
                 reg4554,
                 reg4553,
                 reg4552,
                 reg4551,
                 forvar4550,
                 reg4549,
                 reg4548,
                 reg4547,
                 forvar4546,
                 reg4545,
                 reg4544,
                 reg4543,
                 reg4542,
                 forvar4541,
                 reg4540,
                 forvar4539,
                 reg4538,
                 reg4537,
                 forvar4536,
                 reg4536,
                 reg4535,
                 forvar4534,
                 reg4533,
                 forvar4532,
                 forvar4531,
                 reg4530,
                 reg4529,
                 reg4528,
                 reg4527,
                 reg4526,
                 reg4525,
                 reg4524,
                 reg4523,
                 forvar4522,
                 forvar4521,
                 reg4520,
                 reg4519,
                 reg4518,
                 reg4517,
                 reg4516,
                 reg4515,
                 reg4514,
                 reg4513,
                 reg4512,
                 reg4511,
                 reg4510,
                 forvar4509,
                 forvar4508,
                 forvar4507,
                 reg4506,
                 forvar4503,
                 forvar4497,
                 forvar4495,
                 reg4494,
                 forvar4491,
                 forvar4483,
                 forvar4480,
                 forvar4471,
                 forvar4478,
                 reg4470,
                 forvar4466,
                 forvar4461,
                 reg4499,
                 reg4505,
                 reg4504,
                 reg4503,
                 reg4502,
                 reg4501,
                 reg4500,
                 forvar4499,
                 reg4498,
                 reg4497,
                 reg4496,
                 forvar4489,
                 forvar4485,
                 reg4484,
                 reg4482,
                 forvar4477,
                 forvar4475,
                 reg4495,
                 forvar4494,
                 reg4493,
                 reg4492,
                 reg4491,
                 reg4490,
                 reg4489,
                 reg4488,
                 reg4487,
                 reg4486,
                 reg4485,
                 forvar4484,
                 reg4483,
                 forvar4482,
                 reg4481,
                 reg4480,
                 reg4479,
                 reg4478,
                 forvar4476,
                 reg4477,
                 reg4476,
                 reg4475,
                 reg4474,
                 reg4473,
                 reg4472,
                 reg4471,
                 forvar4470,
                 reg4469,
                 reg4468,
                 reg4467,
                 reg4466,
                 reg4465,
                 reg4464,
                 reg4463,
                 reg4462,
                 reg4461,
                 forvar4460,
                 forvar4459,
                 wire4457,
                 reg3779,
                 wire3778,
                 wire3777,
                 wire3776,
                 wire3775,
                 wire3774,
                 (1'h0)};
  assign wire3774 = wire3772;
  assign wire3775 = $signed(wire3770);
  assign wire3776 = wire3772;
  assign wire3777 = $signed(wire3772);
  assign wire3778 = wire3775[(4'h8):(4'h8)];
  always
    @(posedge clk) begin
      reg3779 <= wire3771[(5'h10):(4'hd)];
    end
  module3780 modinst4458 (.wire3782(wire3770), .clk(clk), .wire3784(wire3772), .y(wire4457), .wire3781(wire3775), .wire3783(wire3778));
  always
    @(posedge clk) begin
      if (wire3770)
        begin
          for (forvar4459 = (1'h0); (forvar4459 < (2'h3)); forvar4459 = (forvar4459 + (1'h1)))
            begin
              for (forvar4460 = (1'h0); (forvar4460 < (2'h2)); forvar4460 = (forvar4460 + (1'h1)))
                begin
                  if (wire3770[(3'h6):(2'h2)])
                    begin
                      reg4461 <= (wire3770 ?
                          wire3774[(4'h9):(1'h0)] : $unsigned(($unsigned((8'hb1)) ?
                              $signed(wire3777) : forvar4460[(4'hb):(3'h7)])));
                      reg4462 <= {(((wire4457 ?
                                  (8'hb2) : reg3779) >>> (wire3773 ?
                                  wire3774 : forvar4459)) ?
                              {$unsigned(reg3779)} : ($signed(wire3771) ~^ wire3776))};
                    end
                  else
                    begin
                      reg4461 <= (-(~&$signed(wire3778)));
                      reg4462 <= ((~&wire3778) + $unsigned(reg3779[(3'h5):(2'h3)]));
                    end
                  if (((wire3778[(1'h0):(1'h0)] | ($signed((8'ha6)) ^~ {wire3778})) >= (reg4461 ?
                      (^~wire3773[(4'hc):(3'h4)]) : $signed((~&reg4462)))))
                    begin
                      reg4463 <= (~|($signed($unsigned(wire3771)) ?
                          {(forvar4459 + wire3771)} : wire3776[(3'h6):(2'h3)]));
                      reg4464 <= (8'hb0);
                    end
                  else
                    begin
                      reg4463 <= $unsigned((!wire3770[(3'h6):(1'h1)]));
                      reg4464 <= $unsigned($unsigned($signed($signed(wire3777))));
                      reg4465 <= (($signed($unsigned(wire3771)) >>> ((wire3770 ^~ wire3778) ?
                              (reg4463 == wire3776) : (~|wire3778))) ?
                          $unsigned(($signed(reg3779) & (wire3771 ?
                              wire4457 : wire3772))) : (~((^wire3773) - reg4461)));
                      reg4466 <= $signed($unsigned(($signed(reg3779) == $unsigned(wire3774))));
                    end
                  if ((^~(8'haa)))
                    begin
                      reg4467 <= (forvar4459 == $unsigned(forvar4460[(3'h5):(2'h2)]));
                      reg4468 <= (reg4464[(3'h5):(3'h5)] << $unsigned($unsigned($signed(wire3771))));
                      reg4469 <= (wire3777 ^~ $signed($unsigned({reg3779})));
                    end
                  else
                    begin
                      reg4467 <= (reg4466[(3'h7):(3'h5)] != {wire3771});
                    end
                  for (forvar4470 = (1'h0); (forvar4470 < (2'h3)); forvar4470 = (forvar4470 + (1'h1)))
                    begin
                      reg4471 <= wire3772[(1'h1):(1'h1)];
                      reg4472 <= {wire3776[(4'hc):(3'h6)]};
                      reg4473 <= (!$signed(((wire3774 > forvar4459) ?
                          (reg4468 > reg4461) : (forvar4470 ~^ forvar4459))));
                      reg4474 <= (~$signed($signed(wire3778)));
                    end
                end
            end
          if (reg4462)
            begin
              reg4475 <= ($unsigned({wire4457[(4'hb):(1'h1)]}) ?
                  $signed(wire3775[(4'hb):(3'h7)]) : (~&$signed(reg4469)));
              if ((|forvar4470[(2'h3):(1'h0)]))
                begin
                  if ((8'hb2))
                    begin
                      reg4476 <= {$unsigned(($unsigned((8'ha5)) ?
                              {forvar4460} : (wire3770 < (8'hb9))))};
                    end
                  else
                    begin
                      reg4476 <= $unsigned(((|(reg4472 ?
                          wire3778 : (8'h9d))) && $signed((reg3779 ?
                          forvar4470 : (8'hb6)))));
                      reg4477 <= reg4461[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar4476 = (1'h0); (forvar4476 < (2'h3)); forvar4476 = (forvar4476 + (1'h1)))
                    begin
                      reg4477 <= $unsigned(reg4473);
                      reg4478 <= $signed(wire3771[(1'h1):(1'h0)]);
                      reg4479 <= ((~reg4463[(3'h4):(1'h0)]) ?
                          (&$unsigned((wire4457 && wire3776))) : $signed({{reg4472}}));
                      reg4480 <= reg4475[(4'h8):(3'h4)];
                    end
                  reg4481 <= {$unsigned($signed(reg3779[(3'h7):(3'h4)]))};
                  for (forvar4482 = (1'h0); (forvar4482 < (1'h0)); forvar4482 = (forvar4482 + (1'h1)))
                    begin
                      reg4483 <= wire4457[(4'hc):(3'h6)];
                    end
                  for (forvar4484 = (1'h0); (forvar4484 < (2'h2)); forvar4484 = (forvar4484 + (1'h1)))
                    begin
                      reg4485 <= ((reg4481 >> (8'ha5)) ~^ $signed((!(-forvar4460))));
                      reg4486 <= ($signed(reg4465) & $unsigned((8'hb4)));
                      reg4487 <= ((((forvar4476 ? reg4474 : (8'hb5)) ?
                              (~forvar4484) : wire3777) ?
                          $unsigned((~reg4473)) : reg4466[(3'h4):(3'h4)]) & (!($signed(wire3774) >= (reg4476 ?
                          (8'hb8) : (8'hb1)))));
                    end
                end
              if (($signed((8'ha0)) != (((reg4477 ? wire3777 : reg4487) ?
                      $signed(wire3776) : (+wire3775)) ?
                  $signed({reg4461}) : ((reg4471 & (8'hb6)) - reg4478))))
                begin
                  if (((($signed(reg4465) ?
                      (!reg4473) : {reg4463}) || $signed($signed((8'hac)))) | ((reg4475 ~^ (forvar4460 ?
                      reg4463 : wire3772)) >= reg4478)))
                    begin
                      reg4488 <= $signed($unsigned(reg4479));
                    end
                  else
                    begin
                      reg4488 <= $signed(reg4479[(2'h3):(2'h2)]);
                      reg4489 <= ((($unsigned(reg4487) ?
                              $unsigned((8'hb4)) : $signed(reg4481)) ^ reg4476[(1'h0):(1'h0)]) ?
                          reg4467[(4'he):(2'h2)] : (reg4481[(4'h8):(2'h3)] ?
                              {(^~(8'hb6))} : $signed($unsigned(reg4469))));
                    end
                  if (reg4488)
                    begin
                      reg4490 <= {({(8'ha0)} ?
                              $signed(forvar4460) : (~reg4466[(2'h2):(1'h1)]))};
                      reg4491 <= (!({$unsigned(wire4457)} ?
                          $unsigned($unsigned(forvar4482)) : reg4468));
                      reg4492 <= reg4471[(2'h2):(1'h0)];
                      reg4493 <= {($unsigned(reg4491[(2'h3):(1'h0)]) ?
                              $signed((wire3772 ?
                                  reg4486 : reg4465)) : ($unsigned(reg4483) ?
                                  (~&reg4486) : (reg4473 ?
                                      forvar4476 : reg4463)))};
                    end
                  else
                    begin
                      reg4490 <= $unsigned(((|(+reg4472)) && {(wire3773 ^~ reg4486)}));
                      reg4491 <= (&(wire3772 >> reg4488[(2'h3):(1'h0)]));
                      reg4492 <= $signed((({reg4476} - (reg4469 ?
                          wire4457 : reg4488)) < (|(reg4468 >> reg4477))));
                    end
                  for (forvar4494 = (1'h0); (forvar4494 < (1'h0)); forvar4494 = (forvar4494 + (1'h1)))
                    begin
                      reg4495 <= $unsigned(reg4477[(3'h4):(1'h1)]);
                    end
                end
              else
                begin
                  if ((8'hb5))
                    begin
                      reg4488 <= $unsigned($signed($signed({reg4467})));
                    end
                  else
                    begin
                      reg4488 <= ((~^reg4490) >> {reg4486});
                      reg4489 <= (8'ha9);
                      reg4490 <= forvar4460[(3'h6):(3'h4)];
                    end
                end
            end
          else
            begin
              for (forvar4475 = (1'h0); (forvar4475 < (2'h3)); forvar4475 = (forvar4475 + (1'h1)))
                begin
                  reg4476 <= $signed($unsigned({(wire3771 <= wire3778)}));
                  for (forvar4477 = (1'h0); (forvar4477 < (1'h1)); forvar4477 = (forvar4477 + (1'h1)))
                    begin
                      reg4478 <= reg4469[(1'h0):(1'h0)];
                      reg4479 <= (wire3777[(1'h1):(1'h0)] ?
                          forvar4494[(1'h0):(1'h0)] : (~^({reg4475} ?
                              (forvar4475 ? wire3778 : reg4465) : (&reg4468))));
                      reg4480 <= $unsigned((~^$signed((forvar4459 * reg4485))));
                      reg4481 <= ({$signed($unsigned(reg4472))} >>> forvar4494);
                    end
                  if ((reg4475 == forvar4460[(1'h1):(1'h1)]))
                    begin
                      reg4482 <= (wire3774[(4'hb):(1'h0)] ?
                          $signed($unsigned((8'h9f))) : reg4480);
                    end
                  else
                    begin
                      reg4482 <= reg4478[(2'h3):(2'h3)];
                      reg4483 <= $unsigned(((reg4463[(4'ha):(4'h8)] ?
                          reg4481[(4'hb):(4'h8)] : (reg3779 != (8'had))) <= $unsigned({reg4467})));
                      reg4484 <= (reg4493 > {(|(&reg4473))});
                    end
                end
              for (forvar4485 = (1'h0); (forvar4485 < (2'h2)); forvar4485 = (forvar4485 + (1'h1)))
                begin
                  reg4486 <= {$unsigned(($signed(reg4490) | (|(8'hab))))};
                  reg4487 <= $unsigned(reg4489);
                  reg4488 <= wire3774;
                end
              for (forvar4489 = (1'h0); (forvar4489 < (1'h1)); forvar4489 = (forvar4489 + (1'h1)))
                begin
                  if ((-($unsigned((&reg4467)) | {(forvar4485 ?
                          wire3773 : (8'haa))})))
                    begin
                      reg4490 <= (wire3774[(2'h3):(2'h2)] << ((8'hb1) < reg4489));
                      reg4491 <= $signed(((^(wire3775 ?
                          reg4461 : wire3774)) < reg4488));
                      reg4492 <= $unsigned($unsigned($unsigned((8'ha4))));
                      reg4493 <= (~|{(forvar4470[(2'h2):(1'h1)] == $unsigned(reg4478))});
                    end
                  else
                    begin
                      reg4490 <= $unsigned($unsigned((8'haa)));
                      reg4491 <= $signed((~^{(^~forvar4484)}));
                      reg4492 <= reg3779[(2'h2):(1'h0)];
                    end
                  for (forvar4494 = (1'h0); (forvar4494 < (2'h2)); forvar4494 = (forvar4494 + (1'h1)))
                    begin
                      reg4495 <= (~&reg4481);
                      reg4496 <= (((+$unsigned(reg4479)) ?
                          $unsigned(forvar4476[(2'h3):(2'h2)]) : wire3774[(4'hb):(1'h1)]) ^~ $unsigned((~|reg4467[(4'hb):(1'h0)])));
                      reg4497 <= (reg4477 & ((8'ha9) >>> {(reg4492 && reg4490)}));
                    end
                  reg4498 <= $signed((reg4461[(2'h3):(1'h0)] ?
                      ({(8'hb8)} && ((8'h9c) | reg4479)) : ((reg4480 ?
                          (8'h9f) : wire3773) > $signed((8'hb2)))));
                end
              if (($signed(reg4466[(3'h6):(3'h4)]) ?
                  reg4487 : (!forvar4459[(3'h4):(2'h2)])))
                begin
                  for (forvar4499 = (1'h0); (forvar4499 < (2'h2)); forvar4499 = (forvar4499 + (1'h1)))
                    begin
                      reg4500 <= (^($signed((8'hb4)) == {(forvar4460 ?
                              forvar4477 : reg4481)}));
                      reg4501 <= reg4483;
                    end
                  if (((((forvar4499 <<< (8'hb4)) || (~(8'ha2))) ?
                          (+$signed((8'hb7))) : ($signed(reg4495) ?
                              reg4473[(3'h7):(2'h2)] : (reg4491 ?
                                  reg4474 : reg4462))) ?
                      reg4496[(1'h0):(1'h0)] : reg4467))
                    begin
                      reg4502 <= (8'ha7);
                      reg4503 <= reg4483;
                      reg4504 <= reg4490[(4'h8):(4'h8)];
                      reg4505 <= forvar4489;
                    end
                  else
                    begin
                      reg4502 <= wire3776;
                    end
                end
              else
                begin
                  if (reg4462[(1'h1):(1'h0)])
                    begin
                      reg4499 <= forvar4484;
                    end
                  else
                    begin
                      reg4499 <= (8'hac);
                      reg4500 <= reg4477;
                      reg4501 <= ((((forvar4476 <= (8'haf)) ?
                          (reg4482 >= (8'hb3)) : (reg4499 ?
                              (8'h9e) : reg4462)) >= (((8'hab) ^ reg3779) * $unsigned(reg4461))) & (($signed(reg4489) <= (8'hb6)) <<< (((8'ha3) ?
                              reg4491 : reg4504) ?
                          $signed(reg4471) : (wire3774 ? (8'hb2) : reg4503))));
                      reg4502 <= {reg4493};
                    end
                end
            end
        end
      else
        begin
          for (forvar4459 = (1'h0); (forvar4459 < (2'h2)); forvar4459 = (forvar4459 + (1'h1)))
            begin
              for (forvar4460 = (1'h0); (forvar4460 < (1'h1)); forvar4460 = (forvar4460 + (1'h1)))
                begin
                  for (forvar4461 = (1'h0); (forvar4461 < (2'h3)); forvar4461 = (forvar4461 + (1'h1)))
                    begin
                      reg4462 <= $signed(reg4471[(1'h1):(1'h1)]);
                      reg4463 <= (|wire3775);
                      reg4464 <= ((~($signed(wire3773) ?
                              {wire3777} : forvar4484[(3'h6):(3'h4)])) ?
                          {wire3771} : reg4475[(3'h4):(1'h1)]);
                      reg4465 <= $signed({{wire3772}});
                    end
                  for (forvar4466 = (1'h0); (forvar4466 < (1'h1)); forvar4466 = (forvar4466 + (1'h1)))
                    begin
                      reg4467 <= ($unsigned(((|reg4479) <<< $unsigned((8'hb2)))) | {(^$unsigned(reg4467))});
                      reg4468 <= {(~|(reg4463[(1'h1):(1'h1)] ?
                              $unsigned(forvar4489) : $signed(reg4493)))};
                      reg4469 <= ((wire3770[(1'h1):(1'h1)] ?
                              (+$signed(forvar4477)) : {(forvar4476 ?
                                      reg4491 : forvar4476)}) ?
                          $unsigned(($signed(forvar4459) >>> reg4495[(1'h1):(1'h1)])) : (~&$signed(forvar4466)));
                      reg4470 <= $signed(wire3778[(2'h3):(1'h1)]);
                    end
                end
              if ($unsigned((reg4496[(3'h4):(1'h1)] ?
                  $signed({wire3773}) : (-((8'hae) ? reg4495 : wire3773)))))
                begin
                  if ((($signed({wire3774}) ?
                          $unsigned(forvar4476) : (!reg4468)) ?
                      (~reg4500) : $unsigned((!$signed(reg4495)))))
                    begin
                      reg4471 <= reg4466;
                      reg4472 <= (~wire3776[(4'h8):(1'h0)]);
                      reg4473 <= (-(($unsigned(reg4482) <<< ((8'hb5) != reg4473)) ?
                          forvar4476[(2'h3):(1'h0)] : (^~(reg4500 ?
                              reg4482 : forvar4489))));
                      reg4474 <= (reg4488[(2'h3):(2'h3)] ?
                          (((&reg4465) * reg4500[(3'h7):(3'h6)]) ?
                              reg4488 : ($signed(forvar4475) ?
                                  (reg4466 >>> reg4469) : (!(8'h9f)))) : {(reg4490 <<< {(8'ha1)})});
                    end
                  else
                    begin
                      reg4471 <= $unsigned((forvar4476[(1'h1):(1'h0)] ?
                          ($signed(reg4476) ?
                              $unsigned(forvar4499) : forvar4485[(4'hc):(1'h0)]) : $signed(reg4464[(3'h4):(2'h2)])));
                    end
                  for (forvar4475 = (1'h0); (forvar4475 < (1'h1)); forvar4475 = (forvar4475 + (1'h1)))
                    begin
                      reg4476 <= {$signed(wire3776[(1'h0):(1'h0)])};
                      reg4477 <= (8'hb9);
                    end
                  for (forvar4478 = (1'h0); (forvar4478 < (2'h3)); forvar4478 = (forvar4478 + (1'h1)))
                    begin
                      reg4479 <= (wire3775 ?
                          (-($signed(reg4504) ?
                              $signed(forvar4484) : (8'h9c))) : $signed(($signed(reg4502) == $signed(wire3775))));
                    end
                  reg4480 <= reg4477[(1'h1):(1'h1)];
                end
              else
                begin
                  for (forvar4471 = (1'h0); (forvar4471 < (1'h1)); forvar4471 = (forvar4471 + (1'h1)))
                    begin
                      reg4472 <= ($signed($unsigned($signed((8'hac)))) >>> $unsigned($signed((wire3778 ?
                          reg4468 : reg4461))));
                      reg4473 <= {{(~^(reg4471 ? forvar4484 : reg4495))}};
                    end
                  if (reg4478)
                    begin
                      reg4474 <= (&((8'ha6) ~^ $signed(forvar4475)));
                      reg4475 <= (~|({(reg4479 ? forvar4460 : (8'hb1))} ?
                          forvar4471 : reg4485[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg4474 <= ({{reg4467}} ? $unsigned({reg4504}) : reg4490);
                      reg4475 <= ($signed(((reg4483 ?
                              forvar4477 : wire3778) < $signed(forvar4484))) ?
                          reg4491[(3'h6):(3'h5)] : $signed(($signed(reg4467) ?
                              (forvar4489 ~^ wire3778) : (reg4484 >>> reg4472))));
                    end
                  if ($unsigned($unsigned((reg4463 == (reg4504 == (8'hb5))))))
                    begin
                      reg4476 <= $signed(({wire3776[(3'h6):(3'h4)]} ?
                          forvar4477 : {(reg4469 ? (8'haf) : (8'hb2))}));
                      reg4477 <= forvar4485;
                      reg4478 <= (~forvar4460);
                      reg4479 <= $unsigned((((reg4504 ? reg4468 : reg4478) ?
                          (reg4481 != wire3778) : $signed(wire3777)) > ((reg4482 ?
                          wire4457 : forvar4470) >= $unsigned((8'hac)))));
                    end
                  else
                    begin
                      reg4476 <= $unsigned((~|{$unsigned(reg4472)}));
                      reg4477 <= $signed(($signed($unsigned((8'ha8))) ?
                          ((reg4466 ^~ reg4495) < {reg4481}) : (~&reg4461[(2'h3):(2'h2)])));
                      reg4478 <= (|$unsigned({(~&reg4467)}));
                    end
                  for (forvar4480 = (1'h0); (forvar4480 < (2'h3)); forvar4480 = (forvar4480 + (1'h1)))
                    begin
                      reg4481 <= (!forvar4480[(1'h0):(1'h0)]);
                      reg4482 <= (($signed($unsigned(reg4495)) ?
                          ((reg4495 ? reg4469 : forvar4471) ?
                              (forvar4475 ?
                                  reg4485 : reg4501) : (reg4476 < (8'ha3))) : ((^~reg4485) <= (&forvar4485))) << $signed(reg4489[(1'h0):(1'h0)]));
                    end
                end
              for (forvar4483 = (1'h0); (forvar4483 < (1'h0)); forvar4483 = (forvar4483 + (1'h1)))
                begin
                  for (forvar4484 = (1'h0); (forvar4484 < (2'h3)); forvar4484 = (forvar4484 + (1'h1)))
                    begin
                      reg4485 <= ((wire3777[(2'h3):(1'h0)] ?
                          ((forvar4489 == forvar4477) ?
                              reg4504 : reg4492[(4'hc):(4'hc)]) : reg4462) && (~^reg4490));
                      reg4486 <= wire3776[(1'h1):(1'h1)];
                      reg4487 <= $unsigned((!forvar4475[(1'h0):(1'h0)]));
                      reg4488 <= reg4466;
                    end
                  if ($signed(((-forvar4470) ?
                      reg4470 : $signed((^forvar4459)))))
                    begin
                      reg4489 <= (((~|{wire3771}) ^~ $signed($signed(wire3778))) ?
                          ($signed($unsigned(reg4480)) ?
                              $unsigned($signed(wire4457)) : (reg4461 + $signed(forvar4459))) : ((^~$signed((8'hb6))) << wire3770[(3'h4):(1'h1)]));
                      reg4490 <= reg4472[(4'hc):(1'h0)];
                    end
                  else
                    begin
                      reg4489 <= $unsigned({wire3775});
                    end
                  for (forvar4491 = (1'h0); (forvar4491 < (1'h0)); forvar4491 = (forvar4491 + (1'h1)))
                    begin
                      reg4492 <= {($signed($signed((8'hb1))) ?
                              reg4465[(3'h6):(3'h6)] : ({forvar4470} - (8'hab)))};
                      reg4493 <= $signed(forvar4459[(2'h2):(1'h1)]);
                      reg4494 <= (forvar4478[(3'h6):(2'h3)] >= $signed($unsigned((forvar4476 ?
                          reg4498 : reg4488))));
                    end
                end
            end
          for (forvar4495 = (1'h0); (forvar4495 < (2'h3)); forvar4495 = (forvar4495 + (1'h1)))
            begin
              if (reg4487)
                begin
                  reg4496 <= wire3775[(1'h0):(1'h0)];
                  if (((&$signed((&forvar4477))) ?
                      $unsigned(reg4490) : reg4495[(4'hb):(4'h8)]))
                    begin
                      reg4497 <= $unsigned(((reg4476 & $signed(reg4478)) ?
                          (!(forvar4480 <<< reg4498)) : reg4475[(4'h9):(4'h8)]));
                      reg4498 <= (^~{reg4500});
                      reg4499 <= ((reg4483[(4'hd):(2'h2)] ?
                              $unsigned(reg4501) : forvar4480) ?
                          (wire3776 + (reg4487[(1'h0):(1'h0)] ?
                              {forvar4485} : {(8'hb3)})) : $unsigned(reg3779));
                      reg4500 <= (($unsigned(wire3773) ?
                              ((forvar4478 ? reg4470 : reg4471) ?
                                  reg4492[(3'h7):(1'h1)] : reg4491) : ((wire3770 ?
                                      reg4490 : reg4500) ?
                                  $unsigned(reg4485) : $signed(reg4462))) ?
                          $signed($unsigned($signed(reg4471))) : $signed((8'hb7)));
                    end
                  else
                    begin
                      reg4497 <= reg4487[(2'h2):(1'h1)];
                      reg4498 <= forvar4489[(1'h1):(1'h0)];
                      reg4499 <= ($unsigned(($signed(forvar4476) ?
                          (forvar4478 ?
                              reg4489 : forvar4461) : forvar4475)) < ($signed((reg4465 ?
                              reg4470 : wire3771)) ?
                          (^forvar4480) : reg4483));
                      reg4500 <= (forvar4478[(2'h2):(1'h0)] ~^ (forvar4499 ?
                          $unsigned((~^reg4462)) : ($unsigned(reg4495) ?
                              $signed(reg4469) : (reg4492 >>> reg4498))));
                    end
                  if ((~|($unsigned(forvar4495) ?
                      wire3776 : $signed(forvar4478))))
                    begin
                      reg4501 <= (reg4487 <<< (^~(reg4474 ?
                          reg4482[(2'h3):(1'h1)] : forvar4485[(3'h5):(1'h0)])));
                      reg4502 <= (!{(&wire3775[(1'h1):(1'h1)])});
                    end
                  else
                    begin
                      reg4501 <= reg4484;
                      reg4502 <= {wire3774};
                    end
                end
              else
                begin
                  reg4496 <= (&$signed(reg4497[(4'h9):(3'h6)]));
                  for (forvar4497 = (1'h0); (forvar4497 < (1'h0)); forvar4497 = (forvar4497 + (1'h1)))
                    begin
                      reg4498 <= wire3776;
                      reg4499 <= reg4468[(4'ha):(4'ha)];
                      reg4500 <= (!reg4479);
                    end
                end
              for (forvar4503 = (1'h0); (forvar4503 < (2'h2)); forvar4503 = (forvar4503 + (1'h1)))
                begin
                  reg4504 <= ((+$unsigned($signed(wire3771))) * forvar4471[(2'h2):(2'h2)]);
                  reg4505 <= ((8'ha5) ? reg4481 : forvar4461);
                end
              reg4506 <= reg4486[(2'h3):(2'h2)];
            end
        end
      for (forvar4507 = (1'h0); (forvar4507 < (2'h3)); forvar4507 = (forvar4507 + (1'h1)))
        begin
          for (forvar4508 = (1'h0); (forvar4508 < (1'h0)); forvar4508 = (forvar4508 + (1'h1)))
            begin
              for (forvar4509 = (1'h0); (forvar4509 < (2'h3)); forvar4509 = (forvar4509 + (1'h1)))
                begin
                  if (forvar4507[(2'h2):(2'h2)])
                    begin
                      reg4510 <= forvar4471[(1'h0):(1'h0)];
                      reg4511 <= ((forvar4470 ^~ (wire4457 & (forvar4466 ?
                          (8'haa) : (8'ha3)))) ^~ reg4474[(1'h1):(1'h1)]);
                      reg4512 <= (^{reg4485[(1'h1):(1'h0)]});
                      reg4513 <= ({reg4484[(2'h3):(1'h0)]} | $signed(($unsigned(reg4494) ?
                          forvar4477[(1'h1):(1'h1)] : (8'ha4))));
                    end
                  else
                    begin
                      reg4510 <= reg4511;
                      reg4511 <= ($unsigned($signed($unsigned(reg4495))) ?
                          $signed($unsigned((8'hb0))) : $unsigned(((^~forvar4508) ^ reg4513[(4'h8):(1'h1)])));
                      reg4512 <= reg4479[(3'h6):(2'h3)];
                    end
                  if (wire3770[(2'h2):(1'h1)])
                    begin
                      reg4514 <= $signed((8'ha5));
                    end
                  else
                    begin
                      reg4514 <= $unsigned($signed($unsigned($unsigned(forvar4495))));
                      reg4515 <= ($unsigned(forvar4503[(3'h4):(1'h0)]) ?
                          $signed($signed($unsigned(reg4475))) : forvar4497);
                      reg4516 <= {$signed(reg4505)};
                    end
                  reg4517 <= (forvar4499 || wire3774);
                  if ((^~forvar4460[(4'h8):(3'h4)]))
                    begin
                      reg4518 <= $signed($unsigned($signed(reg4474[(2'h2):(1'h1)])));
                      reg4519 <= forvar4489;
                      reg4520 <= reg4504;
                    end
                  else
                    begin
                      reg4518 <= $unsigned((-(((8'hb0) ?
                          reg4510 : forvar4471) - (reg4506 ?
                          reg4489 : wire3772))));
                      reg4519 <= {$unsigned($signed({reg4466}))};
                    end
                end
              for (forvar4521 = (1'h0); (forvar4521 < (2'h3)); forvar4521 = (forvar4521 + (1'h1)))
                begin
                  for (forvar4522 = (1'h0); (forvar4522 < (1'h0)); forvar4522 = (forvar4522 + (1'h1)))
                    begin
                      reg4523 <= {$signed((reg4462 ?
                              forvar4460[(3'h6):(1'h1)] : ((8'haa) | (8'hae))))};
                      reg4524 <= ($unsigned(((reg4483 ? wire3773 : wire3771) ?
                          $unsigned((8'hae)) : forvar4475)) ^~ {(forvar4491[(1'h0):(1'h0)] == (reg4498 ?
                              reg4519 : wire3777))});
                    end
                  if ((reg4471 ? $unsigned(reg4486) : reg4475))
                    begin
                      reg4525 <= ((-($unsigned(reg4472) <<< $unsigned(reg4494))) < reg4471[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4525 <= (8'h9d);
                    end
                  if ((^~(&($unsigned(wire3777) ?
                      (reg4525 < reg4511) : reg4485[(2'h3):(1'h0)]))))
                    begin
                      reg4526 <= (~$signed(($unsigned(forvar4503) ~^ $signed((8'ha7)))));
                      reg4527 <= $signed(({$signed(reg4490)} ?
                          (~^$unsigned(wire3775)) : $signed((~^forvar4460))));
                      reg4528 <= $signed(reg4461);
                    end
                  else
                    begin
                      reg4526 <= $signed((+forvar4503));
                      reg4527 <= (((reg4510 >> $unsigned(reg4477)) ?
                          (8'ha0) : wire3775) ~^ {$signed((forvar4483 ?
                              reg4503 : forvar4491))});
                    end
                  if ($signed({((reg4467 << reg4468) || $unsigned(wire3772))}))
                    begin
                      reg4529 <= $unsigned($unsigned({{reg4515}}));
                    end
                  else
                    begin
                      reg4529 <= ((8'ha7) ?
                          $unsigned((^~$unsigned(reg4477))) : $unsigned(forvar4482[(1'h1):(1'h0)]));
                      reg4530 <= $unsigned((({forvar4480} < (8'hac)) ?
                          (^~reg4524[(2'h2):(1'h1)]) : (8'hba)));
                    end
                end
            end
        end
      for (forvar4531 = (1'h0); (forvar4531 < (2'h3)); forvar4531 = (forvar4531 + (1'h1)))
        begin
          for (forvar4532 = (1'h0); (forvar4532 < (1'h1)); forvar4532 = (forvar4532 + (1'h1)))
            begin
              if (((forvar4477 >> {(~&forvar4489)}) ?
                  reg4491 : $signed($unsigned($unsigned((8'hb8))))))
                begin
                  reg4533 <= {$signed($signed(forvar4470[(2'h2):(2'h2)]))};
                  for (forvar4534 = (1'h0); (forvar4534 < (1'h1)); forvar4534 = (forvar4534 + (1'h1)))
                    begin
                      reg4535 <= forvar4521;
                    end
                end
              else
                begin
                  reg4533 <= (!(-reg4470));
                end
              if (reg4493[(1'h1):(1'h1)])
                begin
                  reg4536 <= $unsigned((($signed((8'haf)) ?
                          ((8'h9f) ? reg4527 : reg4466) : (reg4470 ?
                              reg4464 : reg4514)) ?
                      (^~$unsigned(reg4505)) : (!(reg4492 ?
                          (8'hb6) : (8'hb6)))));
                end
              else
                begin
                  for (forvar4536 = (1'h0); (forvar4536 < (2'h3)); forvar4536 = (forvar4536 + (1'h1)))
                    begin
                      reg4537 <= wire3770[(3'h7):(3'h5)];
                    end
                  reg4538 <= {(~&$unsigned((^(8'hb0))))};
                  for (forvar4539 = (1'h0); (forvar4539 < (1'h1)); forvar4539 = (forvar4539 + (1'h1)))
                    begin
                      reg4540 <= {($unsigned($signed(reg4490)) >= $signed($signed(forvar4497)))};
                    end
                end
              if ($unsigned((~^reg4471)))
                begin
                  for (forvar4541 = (1'h0); (forvar4541 < (1'h0)); forvar4541 = (forvar4541 + (1'h1)))
                    begin
                      reg4542 <= ({(forvar4476 ?
                              ((8'ha3) ?
                                  reg4514 : forvar4536) : (wire3771 || (8'haf)))} <<< (~^$signed({(8'hba)})));
                      reg4543 <= ((~&(^(~&reg4528))) ?
                          $unsigned((+(!(8'hb3)))) : $unsigned(reg4538[(1'h1):(1'h1)]));
                      reg4544 <= reg4500[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar4541 = (1'h0); (forvar4541 < (1'h0)); forvar4541 = (forvar4541 + (1'h1)))
                    begin
                      reg4542 <= {$signed(((^~reg4514) ?
                              (reg4513 == reg4468) : (reg4493 * reg4470)))};
                      reg4543 <= (8'hb1);
                      reg4544 <= $signed((((forvar4507 ?
                              reg4471 : reg4538) < {reg4523}) ?
                          (^~{(8'ha4)}) : (^(&(8'ha3)))));
                      reg4545 <= reg4465;
                    end
                  for (forvar4546 = (1'h0); (forvar4546 < (2'h3)); forvar4546 = (forvar4546 + (1'h1)))
                    begin
                      reg4547 <= (|(|forvar4546[(4'hd):(1'h1)]));
                      reg4548 <= (reg4523 && (((~&forvar4539) ^ $unsigned((8'hb1))) >> $signed(reg4543)));
                    end
                  reg4549 <= reg4491[(2'h3):(2'h2)];
                end
            end
          for (forvar4550 = (1'h0); (forvar4550 < (2'h2)); forvar4550 = (forvar4550 + (1'h1)))
            begin
              if ((!reg4549[(2'h2):(1'h1)]))
                begin
                  if ($signed((wire3772[(4'h9):(4'h8)] ?
                      ($unsigned(reg4475) + reg4482) : $signed((reg4544 > reg4516)))))
                    begin
                      reg4551 <= ($signed(forvar4489) <= reg4517);
                      reg4552 <= $signed(reg4492);
                      reg4553 <= (~|{(8'hb8)});
                    end
                  else
                    begin
                      reg4551 <= {$signed((|{reg4540}))};
                      reg4552 <= (-wire3778[(1'h0):(1'h0)]);
                    end
                  if ($signed($signed(reg4482[(3'h4):(2'h3)])))
                    begin
                      reg4554 <= reg4464[(2'h2):(1'h1)];
                      reg4555 <= reg4542[(2'h3):(2'h3)];
                      reg4556 <= $unsigned($unsigned((reg4485 ?
                          reg3779 : $unsigned((8'hab)))));
                    end
                  else
                    begin
                      reg4554 <= (reg4491[(3'h5):(2'h2)] ?
                          (^reg4552) : (-$unsigned((reg4529 ?
                              reg4485 : reg4490))));
                    end
                  for (forvar4557 = (1'h0); (forvar4557 < (1'h1)); forvar4557 = (forvar4557 + (1'h1)))
                    begin
                      reg4558 <= {{({forvar4557} ?
                                  reg4464[(3'h7):(3'h6)] : (reg4525 ?
                                      reg4461 : wire3777))}};
                      reg4559 <= ($signed((~|(-reg4530))) == (+forvar4477));
                    end
                  if (reg4549)
                    begin
                      reg4560 <= reg4474;
                    end
                  else
                    begin
                      reg4560 <= (($signed($signed(reg4526)) <<< $signed(reg4496[(2'h2):(1'h0)])) >> $unsigned(forvar4531));
                      reg4561 <= reg4529;
                      reg4562 <= reg4513;
                    end
                end
              else
                begin
                  reg4551 <= ($unsigned((!reg4489[(3'h6):(3'h6)])) ?
                      ({(~&reg4551)} ?
                          ($signed(reg4510) ?
                              (~|(8'hb1)) : (^~forvar4541)) : $unsigned($signed(reg4472))) : reg4515[(4'hc):(2'h2)]);
                  for (forvar4552 = (1'h0); (forvar4552 < (2'h2)); forvar4552 = (forvar4552 + (1'h1)))
                    begin
                      reg4553 <= ((({forvar4521} ?
                              ((8'hb3) != reg4490) : reg4504[(4'hb):(2'h2)]) ^~ ((^~reg4486) ?
                              (~&forvar4482) : $unsigned(reg4472))) ?
                          {forvar4489[(1'h1):(1'h0)]} : $unsigned(((reg3779 ?
                                  forvar4539 : wire3776) ?
                              (^~reg4476) : (reg4552 < reg4503))));
                      reg4554 <= wire3773;
                      reg4555 <= ($unsigned((^$unsigned(reg4470))) * ((+(^reg4559)) ?
                          ({reg4551} ?
                              (^~reg4551) : (~|reg4483)) : $signed((reg4525 ?
                              forvar4532 : forvar4485))));
                      reg4556 <= ({wire3771} ?
                          (&$unsigned(reg4560)) : (+{reg4470}));
                    end
                end
              if ($unsigned(wire3774[(4'he):(2'h3)]))
                begin
                  if ((((reg4485[(1'h1):(1'h1)] == (reg4549 >= forvar4478)) ?
                          (+(8'ha5)) : forvar4476[(3'h4):(1'h1)]) ?
                      {{(reg4463 <= reg4496)}} : (!($unsigned(forvar4480) & $unsigned(reg4492)))))
                    begin
                      reg4563 <= reg4495[(4'h9):(1'h1)];
                      reg4564 <= reg4540[(4'h8):(2'h3)];
                    end
                  else
                    begin
                      reg4563 <= $signed($signed(reg4556[(2'h3):(1'h0)]));
                    end
                  reg4565 <= reg4484[(3'h6):(3'h6)];
                  if (wire3775)
                    begin
                      reg4566 <= $signed($signed(($signed(wire3777) <= (reg4563 ?
                          reg4528 : reg4518))));
                      reg4567 <= ($unsigned(((reg4538 ? reg4517 : reg4497) ?
                              (!reg4562) : $unsigned(reg4489))) ?
                          (($unsigned((8'h9c)) ? reg4549 : $signed(reg4558)) ?
                              $signed(forvar4503) : (wire4457 ?
                                  (reg4478 ?
                                      reg4558 : reg4493) : forvar4484[(4'h8):(3'h5)])) : reg4488[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg4566 <= $unsigned($signed($unsigned(forvar4461[(1'h0):(1'h0)])));
                      reg4567 <= {{forvar4478[(1'h0):(1'h0)]}};
                      reg4568 <= {((|(reg4504 ? forvar4461 : reg4479)) ?
                              $signed($signed(reg4525)) : $unsigned(reg4506))};
                    end
                end
              else
                begin
                  for (forvar4563 = (1'h0); (forvar4563 < (2'h2)); forvar4563 = (forvar4563 + (1'h1)))
                    begin
                      reg4564 <= reg4465[(2'h2):(1'h0)];
                      reg4565 <= (^~reg4484);
                    end
                  reg4566 <= ((^~$signed((reg4516 > reg4503))) ?
                      $signed((-$signed((8'hb7)))) : ({{reg4525}} < (|$unsigned(wire3773))));
                end
              if (({{((8'ha2) ?
                          reg4535 : reg4524)}} > $unsigned($unsigned((wire3776 ?
                  reg4548 : reg4558)))))
                begin
                  if ((({{forvar4536}} & ({reg4495} ?
                      reg4482 : $signed((8'h9c)))) + ($unsigned($signed(reg4526)) >= $signed(forvar4482[(2'h3):(1'h1)]))))
                    begin
                      reg4569 <= $signed(reg4526);
                      reg4570 <= ((~|(!(reg4474 <= forvar4541))) | wire3778[(1'h0):(1'h0)]);
                      reg4571 <= $signed($unsigned(reg4502));
                      reg4572 <= (~|$unsigned(forvar4491));
                    end
                  else
                    begin
                      reg4569 <= ($unsigned(reg4511[(1'h0):(1'h0)]) != wire3772[(3'h6):(2'h3)]);
                      reg4570 <= ($unsigned(reg4470[(3'h4):(2'h2)]) ?
                          $signed($signed(wire3775)) : (((8'hab) != (8'ha7)) ^~ forvar4563[(2'h2):(2'h2)]));
                      reg4571 <= $unsigned($signed((8'ha0)));
                    end
                end
              else
                begin
                  for (forvar4569 = (1'h0); (forvar4569 < (2'h3)); forvar4569 = (forvar4569 + (1'h1)))
                    begin
                      reg4570 <= reg4563[(3'h4):(1'h1)];
                      reg4571 <= ((reg4536[(3'h6):(1'h1)] ?
                          $signed((reg4484 || (8'hb2))) : ((reg4560 << reg4518) - (reg4475 | reg4469))) ^ ($signed({reg4555}) << reg4512[(2'h2):(1'h1)]));
                    end
                  for (forvar4572 = (1'h0); (forvar4572 < (1'h0)); forvar4572 = (forvar4572 + (1'h1)))
                    begin
                      reg4573 <= forvar4480;
                      reg4574 <= $unsigned(($signed(reg4492) ?
                          ((reg4504 ? reg4538 : reg4537) ?
                              reg4555[(2'h3):(2'h2)] : {reg4479}) : ($unsigned(forvar4484) <<< $signed(reg4471))));
                      reg4575 <= (-$signed($signed((reg4547 ^ reg4566))));
                      reg4576 <= reg4461;
                    end
                end
              if (forvar4532[(3'h4):(1'h0)])
                begin
                  if ($signed((($signed(forvar4509) + (forvar4503 ^ reg4530)) >>> (|{reg4512}))))
                    begin
                      reg4577 <= (~|($unsigned((forvar4478 >> reg4477)) ?
                          $unsigned(((8'ha6) || (8'h9c))) : (|((8'h9c) ?
                              reg4501 : reg4503))));
                      reg4578 <= {(~^reg4559[(2'h2):(2'h2)])};
                      reg4579 <= (+$signed(reg4469));
                    end
                  else
                    begin
                      reg4577 <= ((~|$unsigned((~|reg4547))) ?
                          (({reg4490} & $unsigned(reg4556)) ?
                              ($signed(forvar4499) * $signed(reg4524)) : (forvar4521[(4'h8):(1'h0)] ?
                                  reg4495 : reg4516)) : $signed(reg4575[(2'h2):(1'h1)]));
                      reg4578 <= (^~wire3777);
                      reg4579 <= (^{($signed(forvar4476) ~^ reg4552)});
                    end
                  reg4580 <= ((|(^(reg4491 ? reg4526 : reg4579))) * (reg4570 ?
                      (|(|reg4520)) : $signed($unsigned(wire3770))));
                  for (forvar4581 = (1'h0); (forvar4581 < (2'h3)); forvar4581 = (forvar4581 + (1'h1)))
                    begin
                      reg4582 <= $unsigned($signed(reg3779));
                      reg4583 <= {forvar4460};
                      reg4584 <= ($unsigned(reg4564[(1'h0):(1'h0)]) << $unsigned(($unsigned(forvar4572) > (reg4540 + reg4515))));
                    end
                end
              else
                begin
                  if ((reg4487 & $signed((&reg4543))))
                    begin
                      reg4577 <= forvar4460[(4'hb):(4'h8)];
                      reg4578 <= ($unsigned(($unsigned(reg4462) < {(8'had)})) ?
                          reg4526[(4'hf):(4'h8)] : (!((|(8'hba)) > (reg4485 ?
                              forvar4484 : wire4457))));
                      reg4579 <= reg4475;
                      reg4580 <= forvar4485[(4'hc):(1'h1)];
                    end
                  else
                    begin
                      reg4577 <= (~reg4568[(3'h5):(2'h2)]);
                      reg4578 <= ((reg4540 || (&(^~forvar4475))) ?
                          forvar4497[(2'h2):(2'h2)] : (reg4462[(4'ha):(4'ha)] * $unsigned($unsigned(forvar4508))));
                      reg4579 <= reg4512;
                    end
                  if (reg4552)
                    begin
                      reg4581 <= (^(&reg4478));
                      reg4582 <= $signed($unsigned(forvar4459));
                    end
                  else
                    begin
                      reg4581 <= $unsigned($unsigned($unsigned((8'h9e))));
                      reg4582 <= {{($signed(reg4549) <<< ((8'ha7) ?
                                  forvar4569 : (8'hb7)))}};
                    end
                  reg4583 <= (((&wire3771[(5'h10):(4'hb)]) || reg4566[(4'h9):(2'h2)]) & (forvar4466[(2'h2):(1'h0)] ^ $signed(reg4486[(2'h3):(1'h0)])));
                end
            end
          reg4585 <= reg4538;
        end
      reg4586 <= reg4468[(3'h4):(2'h2)];
    end
  assign wire4587 = wire3778[(3'h6):(1'h1)];
  always
    @(posedge clk) begin
      if ($unsigned(($signed(reg4471[(1'h0):(1'h0)]) ?
          (reg4578[(2'h2):(2'h2)] ~^ {reg4566}) : $unsigned(forvar4491[(3'h6):(3'h6)]))))
        begin
          for (forvar4588 = (1'h0); (forvar4588 < (2'h3)); forvar4588 = (forvar4588 + (1'h1)))
            begin
              for (forvar4589 = (1'h0); (forvar4589 < (1'h1)); forvar4589 = (forvar4589 + (1'h1)))
                begin
                  reg4590 <= $signed(reg4512[(1'h0):(1'h0)]);
                  reg4591 <= {({(~|(8'hba))} ?
                          (~^reg4466) : (^~reg4512[(4'ha):(1'h1)]))};
                  for (forvar4592 = (1'h0); (forvar4592 < (1'h0)); forvar4592 = (forvar4592 + (1'h1)))
                    begin
                      reg4593 <= ($unsigned(reg4576[(2'h2):(2'h2)]) ?
                          (&((forvar4476 > reg4463) ?
                              reg4554 : {reg4566})) : reg4524);
                    end
                end
              for (forvar4594 = (1'h0); (forvar4594 < (1'h1)); forvar4594 = (forvar4594 + (1'h1)))
                begin
                  reg4595 <= wire3778[(3'h6):(3'h6)];
                  reg4596 <= reg4475[(4'ha):(4'h9)];
                  reg4597 <= $signed((($unsigned((8'hb7)) > $signed(wire3773)) <<< $unsigned({(8'h9c)})));
                end
              if (((-((forvar4546 ? (8'hb3) : wire3771) ?
                      reg4486 : (~&forvar4466))) ?
                  (~|(|{reg4490})) : $unsigned((^~$unsigned(reg4468)))))
                begin
                  reg4598 <= (reg4497[(4'hc):(1'h0)] ?
                      $signed(reg4596) : $signed((~(reg4576 ?
                          reg4510 : (8'h9f)))));
                end
              else
                begin
                  for (forvar4598 = (1'h0); (forvar4598 < (1'h0)); forvar4598 = (forvar4598 + (1'h1)))
                    begin
                      reg4599 <= (8'hb9);
                    end
                  for (forvar4600 = (1'h0); (forvar4600 < (2'h2)); forvar4600 = (forvar4600 + (1'h1)))
                    begin
                      reg4601 <= (+$signed(reg4582[(2'h3):(2'h3)]));
                    end
                  if (($unsigned((&$signed(wire3772))) >= reg4559[(2'h2):(2'h2)]))
                    begin
                      reg4602 <= $signed(((reg4529 > reg4573) ?
                          ((reg4523 ?
                              (8'h9f) : reg4468) - wire4457[(2'h2):(1'h0)]) : reg4535[(4'hb):(3'h7)]));
                      reg4603 <= (^reg4584[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg4602 <= $signed({(reg4513[(4'hf):(3'h4)] ~^ reg4580[(1'h1):(1'h1)])});
                    end
                  reg4604 <= {(reg4493[(1'h0):(1'h0)] && $signed($signed((8'ha6))))};
                end
              for (forvar4605 = (1'h0); (forvar4605 < (2'h3)); forvar4605 = (forvar4605 + (1'h1)))
                begin
                  for (forvar4606 = (1'h0); (forvar4606 < (1'h1)); forvar4606 = (forvar4606 + (1'h1)))
                    begin
                      reg4607 <= $signed(reg4584);
                      reg4608 <= ({wire3770[(2'h2):(2'h2)]} ?
                          $unsigned(($signed(reg4553) < (^~wire3776))) : (^$unsigned($signed(wire3773))));
                    end
                  for (forvar4609 = (1'h0); (forvar4609 < (2'h2)); forvar4609 = (forvar4609 + (1'h1)))
                    begin
                      reg4610 <= reg4512;
                      reg4611 <= $unsigned((~({forvar4478} >> {forvar4546})));
                      reg4612 <= {(^wire3773[(3'h5):(1'h1)])};
                      reg4613 <= ($unsigned((~|$unsigned(reg4513))) | forvar4491[(2'h2):(1'h1)]);
                    end
                  if ({(forvar4460 ?
                          $signed(((8'ha3) >> reg4483)) : reg4582[(4'ha):(4'h9)])})
                    begin
                      reg4614 <= reg4567[(1'h1):(1'h0)];
                      reg4615 <= $signed(forvar4572[(4'ha):(1'h0)]);
                      reg4616 <= ($unsigned(reg4586) >= (!forvar4471[(3'h7):(1'h1)]));
                    end
                  else
                    begin
                      reg4614 <= (~|forvar4484[(3'h6):(2'h3)]);
                      reg4615 <= $unsigned($signed((-(-reg4556))));
                      reg4616 <= $signed((~&(^reg4513[(4'hd):(4'hb)])));
                    end
                end
            end
        end
      else
        begin
          if ($signed((|{(reg4545 - wire3774)})))
            begin
              for (forvar4588 = (1'h0); (forvar4588 < (1'h1)); forvar4588 = (forvar4588 + (1'h1)))
                begin
                  for (forvar4589 = (1'h0); (forvar4589 < (1'h1)); forvar4589 = (forvar4589 + (1'h1)))
                    begin
                      reg4590 <= ((~&({reg4501} ?
                          (reg4575 ?
                              reg4516 : reg4577) : reg4528[(1'h1):(1'h1)])) + reg4570);
                      reg4591 <= reg4502[(1'h1):(1'h1)];
                    end
                  if ($signed({reg4591[(3'h7):(1'h1)]}))
                    begin
                      reg4592 <= reg4510[(2'h2):(2'h2)];
                      reg4593 <= $unsigned({$signed(((8'hab) ?
                              reg4475 : (8'ha4)))});
                      reg4594 <= reg4463[(2'h3):(1'h0)];
                      reg4595 <= $unsigned((($unsigned(reg4535) && $unsigned(wire3771)) >> $signed((reg4542 ?
                          reg4607 : forvar4539))));
                    end
                  else
                    begin
                      reg4592 <= (&forvar4534[(3'h4):(3'h4)]);
                      reg4593 <= $signed(reg4520);
                      reg4594 <= (reg4462 && forvar4475);
                    end
                end
              for (forvar4596 = (1'h0); (forvar4596 < (2'h3)); forvar4596 = (forvar4596 + (1'h1)))
                begin
                  for (forvar4597 = (1'h0); (forvar4597 < (1'h0)); forvar4597 = (forvar4597 + (1'h1)))
                    begin
                      reg4598 <= ((^~($signed(wire3772) ^~ $unsigned((8'ha4)))) > (reg4538 - {(&reg4543)}));
                    end
                  if ((8'hb4))
                    begin
                      reg4599 <= ($signed(($signed(reg4471) - (~&reg4528))) * (reg4494 ^~ forvar4461));
                      reg4600 <= forvar4475[(4'h8):(2'h2)];
                    end
                  else
                    begin
                      reg4599 <= forvar4491[(3'h4):(2'h3)];
                    end
                end
              reg4601 <= ($unsigned(reg4492[(3'h6):(2'h3)]) ?
                  $signed((reg4471[(2'h3):(2'h3)] <<< ((8'h9c) ?
                      reg4490 : reg4613))) : (8'hb7));
              for (forvar4602 = (1'h0); (forvar4602 < (2'h2)); forvar4602 = (forvar4602 + (1'h1)))
                begin
                  for (forvar4603 = (1'h0); (forvar4603 < (1'h1)); forvar4603 = (forvar4603 + (1'h1)))
                    begin
                      reg4604 <= (~((reg4537 >>> (+reg4490)) ?
                          ((forvar4546 >= wire3771) ~^ forvar4597) : reg4603[(2'h2):(1'h1)]));
                      reg4605 <= (((8'hae) ?
                          ((reg4490 == reg4498) ?
                              (reg4575 ?
                                  reg4560 : forvar4482) : ((8'ha0) >>> (8'ha4))) : $unsigned($signed(reg4510))) == (reg4602[(4'h9):(4'h9)] != ($unsigned(reg4476) ?
                          (reg4491 <<< reg4466) : {reg4597})));
                      reg4606 <= {forvar4592};
                      reg4607 <= (8'ha6);
                    end
                  if ($unsigned($signed(((^(8'hba)) ^~ reg4558[(4'h8):(2'h2)]))))
                    begin
                      reg4608 <= $signed(reg4591);
                    end
                  else
                    begin
                      reg4608 <= reg4476;
                      reg4609 <= (forvar4483[(3'h4):(2'h2)] == (-reg4548[(1'h0):(1'h0)]));
                      reg4610 <= reg4568;
                    end
                end
            end
          else
            begin
              for (forvar4588 = (1'h0); (forvar4588 < (2'h3)); forvar4588 = (forvar4588 + (1'h1)))
                begin
                  for (forvar4589 = (1'h0); (forvar4589 < (1'h1)); forvar4589 = (forvar4589 + (1'h1)))
                    begin
                      reg4590 <= $unsigned(reg4523[(2'h3):(1'h1)]);
                      reg4591 <= ($signed(($signed(reg4599) < (reg4572 || reg4518))) - ($unsigned((!reg4566)) ~^ $signed($signed((8'hb2)))));
                      reg4592 <= $signed((reg4527[(3'h7):(1'h1)] ?
                          ($unsigned(reg4607) & (~|reg4514)) : {wire3773[(3'h4):(2'h2)]}));
                    end
                end
              for (forvar4593 = (1'h0); (forvar4593 < (2'h3)); forvar4593 = (forvar4593 + (1'h1)))
                begin
                  for (forvar4594 = (1'h0); (forvar4594 < (1'h0)); forvar4594 = (forvar4594 + (1'h1)))
                    begin
                      reg4595 <= reg4544;
                    end
                  for (forvar4596 = (1'h0); (forvar4596 < (1'h1)); forvar4596 = (forvar4596 + (1'h1)))
                    begin
                      reg4597 <= $unsigned({$signed($unsigned(reg4570))});
                      reg4598 <= reg4497;
                      reg4599 <= $unsigned(reg4593);
                    end
                end
              if ((~^$signed($unsigned((forvar4557 ? reg4600 : reg4591)))))
                begin
                  for (forvar4600 = (1'h0); (forvar4600 < (2'h2)); forvar4600 = (forvar4600 + (1'h1)))
                    begin
                      reg4601 <= (~^(reg4583 ?
                          $signed(reg4475) : $unsigned({reg4577})));
                      reg4602 <= ((($signed(reg4506) ?
                              (reg4499 << reg4462) : $signed(reg4573)) ?
                          ((forvar4499 >>> reg4584) ?
                              forvar4482[(3'h4):(1'h0)] : $unsigned(forvar4491)) : $unsigned((|wire3772))) << (|reg4615[(2'h3):(2'h2)]));
                      reg4603 <= reg4575;
                    end
                  for (forvar4604 = (1'h0); (forvar4604 < (2'h3)); forvar4604 = (forvar4604 + (1'h1)))
                    begin
                      reg4605 <= {$signed(reg4552[(3'h6):(3'h5)])};
                    end
                  if ($unsigned(reg4483[(3'h4):(2'h2)]))
                    begin
                      reg4606 <= (+($signed((forvar4507 ?
                              reg4577 : forvar4509)) ?
                          $unsigned({reg4476}) : reg4573));
                      reg4607 <= (8'hb8);
                      reg4608 <= ((reg4485[(2'h2):(1'h1)] != reg4610) ?
                          $signed($signed({forvar4597})) : ((~|$signed((8'hb0))) & forvar4460));
                    end
                  else
                    begin
                      reg4606 <= $signed({$signed((^~reg4605))});
                    end
                end
              else
                begin
                  reg4600 <= ((^$signed((forvar4589 ?
                      wire3778 : reg4484))) == reg4478[(2'h2):(1'h0)]);
                  if (($signed((~&forvar4569)) ?
                      (&reg4611) : (($signed(wire3774) == ((8'hb6) || reg4475)) ?
                          (reg4547 == $unsigned((8'hb7))) : ($unsigned(reg4598) ?
                              (8'hb5) : (reg4570 < reg4572)))))
                    begin
                      reg4601 <= ((forvar4546 ?
                              ((forvar4604 || reg4500) ?
                                  (-reg4602) : forvar4509[(1'h1):(1'h0)]) : reg4465) ?
                          $unsigned(((reg4526 ? (8'hba) : (8'hab)) ?
                              $unsigned((8'hab)) : (reg4562 ?
                                  reg4547 : reg4552))) : {reg4490[(1'h0):(1'h0)]});
                      reg4602 <= (&$unsigned($unsigned(forvar4598)));
                      reg4603 <= (&$unsigned((forvar4489 ?
                          $signed(reg4542) : $unsigned((8'hab)))));
                    end
                  else
                    begin
                      reg4601 <= reg4535[(3'h5):(1'h0)];
                      reg4602 <= $unsigned(reg4476[(1'h0):(1'h0)]);
                      reg4603 <= {forvar4541[(4'h8):(3'h7)]};
                      reg4604 <= (((reg4593[(4'hd):(4'hb)] <<< reg4499[(4'ha):(1'h0)]) ^ forvar4609) ?
                          (($unsigned(wire3778) ?
                              {reg4567} : reg4524) << $signed((forvar4497 ?
                              wire4587 : (8'ha5)))) : {(~^reg4569)});
                    end
                  for (forvar4605 = (1'h0); (forvar4605 < (2'h3)); forvar4605 = (forvar4605 + (1'h1)))
                    begin
                      reg4606 <= ($unsigned($unsigned((~^reg4575))) > $signed(reg4591));
                    end
                  for (forvar4607 = (1'h0); (forvar4607 < (1'h0)); forvar4607 = (forvar4607 + (1'h1)))
                    begin
                      reg4608 <= $signed((~&(forvar4572 & $signed(reg4519))));
                      reg4609 <= {(reg4515 || $signed(reg4523[(2'h2):(1'h0)]))};
                    end
                end
              for (forvar4610 = (1'h0); (forvar4610 < (1'h0)); forvar4610 = (forvar4610 + (1'h1)))
                begin
                  for (forvar4611 = (1'h0); (forvar4611 < (2'h2)); forvar4611 = (forvar4611 + (1'h1)))
                    begin
                      reg4612 <= ($signed($signed((reg4479 << reg4540))) == (reg4613[(4'h8):(3'h6)] ?
                          {reg4610} : reg4593));
                    end
                  reg4613 <= $unsigned(forvar4494[(3'h5):(2'h2)]);
                  for (forvar4614 = (1'h0); (forvar4614 < (2'h2)); forvar4614 = (forvar4614 + (1'h1)))
                    begin
                      reg4615 <= ($unsigned(forvar4466) ?
                          {(&$signed(reg4616))} : {(^(&(8'hba)))});
                      reg4616 <= wire4457;
                      reg4617 <= (|$unsigned(($signed((8'hba)) == (reg4543 <<< reg4466))));
                    end
                  reg4618 <= $signed(reg4513);
                end
            end
          for (forvar4619 = (1'h0); (forvar4619 < (2'h3)); forvar4619 = (forvar4619 + (1'h1)))
            begin
              if (({forvar4593} >= ($signed(reg4505) & $unsigned((forvar4572 >= (8'hb2))))))
                begin
                  if ((reg4553[(1'h0):(1'h0)] ?
                      ((forvar4594 ?
                          (~&reg4615) : $unsigned(reg4570)) < ($unsigned(reg4512) ?
                          (reg4516 <<< reg4560) : (!forvar4592))) : $signed((reg4473[(4'ha):(4'h9)] | $signed(forvar4539)))))
                    begin
                      reg4620 <= $signed(reg4564);
                      reg4621 <= forvar4491[(1'h0):(1'h0)];
                      reg4622 <= $signed({$signed((^reg4564))});
                      reg4623 <= ($signed($signed($signed(forvar4477))) ?
                          ((&reg4561[(4'h8):(3'h4)]) || (((8'ha9) >> reg4565) ?
                              forvar4602[(3'h7):(1'h1)] : $signed((8'hb6)))) : $unsigned((&$signed((8'ha7)))));
                    end
                  else
                    begin
                      reg4620 <= $unsigned({{reg4570[(3'h5):(2'h2)]}});
                      reg4621 <= ($unsigned(((forvar4484 ?
                              reg4471 : reg4462) != (^~reg4504))) ?
                          {$unsigned((~(8'hac)))} : reg4618[(2'h3):(1'h0)]);
                      reg4622 <= (|$signed(reg4567));
                    end
                  for (forvar4624 = (1'h0); (forvar4624 < (1'h0)); forvar4624 = (forvar4624 + (1'h1)))
                    begin
                      reg4625 <= reg4601[(3'h7):(3'h6)];
                      reg4626 <= forvar4569;
                    end
                  if ((forvar4624 ?
                      ((&reg4463) ^~ (reg4578 - (forvar4602 ?
                          forvar4460 : reg4495))) : $unsigned(forvar4598)))
                    begin
                      reg4627 <= reg4563;
                    end
                  else
                    begin
                      reg4627 <= forvar4557[(4'ha):(1'h0)];
                      reg4628 <= (-(-$signed(((8'hb7) ?
                          (8'ha9) : forvar4569))));
                      reg4629 <= (reg4567 | $signed($unsigned(wire4457[(4'hf):(4'hc)])));
                      reg4630 <= forvar4609[(1'h0):(1'h0)];
                    end
                  if ($signed(forvar4534[(4'h9):(3'h6)]))
                    begin
                      reg4631 <= reg4622;
                      reg4632 <= $unsigned($unsigned((reg4621 >>> $unsigned(reg4494))));
                      reg4633 <= ((forvar4536[(2'h3):(1'h1)] + (reg4560[(2'h2):(1'h0)] | forvar4522)) <<< forvar4604[(3'h6):(3'h5)]);
                      reg4634 <= ($unsigned((~^reg4575[(1'h1):(1'h0)])) ^ $unsigned((reg4466[(3'h7):(3'h7)] || forvar4461[(3'h5):(2'h2)])));
                    end
                  else
                    begin
                      reg4631 <= (($unsigned(reg4620[(2'h2):(2'h2)]) ?
                          forvar4594 : $signed((!reg4492))) != $unsigned(reg4548[(2'h3):(2'h3)]));
                      reg4632 <= wire3775[(4'hd):(4'hb)];
                      reg4633 <= reg4608[(4'h8):(1'h1)];
                      reg4634 <= (($unsigned((^~forvar4534)) ?
                              ((~reg4515) >> (reg4527 ^~ (8'hb9))) : ($unsigned(forvar4552) ?
                                  $signed(reg4626) : (forvar4489 ?
                                      forvar4588 : reg4495))) ?
                          reg4568[(3'h5):(1'h0)] : wire3774);
                    end
                end
              else
                begin
                  if ((^~$unsigned(forvar4508[(1'h0):(1'h0)])))
                    begin
                      reg4620 <= (($unsigned($unsigned(reg4566)) >= (~forvar4460)) ?
                          $unsigned(({reg4579} ?
                              reg4461 : {forvar4478})) : reg4562);
                    end
                  else
                    begin
                      reg4620 <= $unsigned(((~|reg4461[(2'h3):(2'h2)]) ?
                          ({forvar4563} ?
                              (forvar4541 ? (8'hb9) : reg4571) : (forvar4546 ?
                                  (8'hab) : reg4548)) : (+(reg4482 <<< (8'hab)))));
                    end
                  for (forvar4621 = (1'h0); (forvar4621 < (1'h1)); forvar4621 = (forvar4621 + (1'h1)))
                    begin
                      reg4622 <= {forvar4619[(1'h0):(1'h0)]};
                      reg4623 <= ((reg4577 * reg4503) << (~&$signed((&forvar4606))));
                      reg4624 <= (~&reg4479);
                    end
                  for (forvar4625 = (1'h0); (forvar4625 < (2'h2)); forvar4625 = (forvar4625 + (1'h1)))
                    begin
                      reg4626 <= ((|(~$signed(reg3779))) - $signed($signed(wire3773)));
                      reg4627 <= (|(reg4618[(1'h0):(1'h0)] <= (((8'ha9) ^ reg4538) ?
                          reg4602 : forvar4611)));
                    end
                end
              if (reg4535[(4'hb):(1'h1)])
                begin
                  for (forvar4635 = (1'h0); (forvar4635 < (2'h3)); forvar4635 = (forvar4635 + (1'h1)))
                    begin
                      reg4636 <= reg4602;
                    end
                end
              else
                begin
                  for (forvar4635 = (1'h0); (forvar4635 < (2'h2)); forvar4635 = (forvar4635 + (1'h1)))
                    begin
                      reg4636 <= {reg4499[(3'h4):(2'h3)]};
                      reg4637 <= forvar4508;
                      reg4638 <= $signed({$signed((+reg4489))});
                      reg4639 <= forvar4475;
                    end
                  if ((^reg4617))
                    begin
                      reg4640 <= ($unsigned($unsigned((reg4590 + reg4518))) ?
                          $signed(reg4516) : reg4514);
                      reg4641 <= ($signed((&(wire3775 ?
                          reg4479 : reg4468))) && reg4465);
                      reg4642 <= ($unsigned((!(reg4492 ?
                          reg4533 : reg4621))) == ({{reg4608}} << {reg4461}));
                      reg4643 <= forvar4609;
                    end
                  else
                    begin
                      reg4640 <= $signed(forvar4602);
                      reg4641 <= (+$unsigned({$signed(reg4564)}));
                      reg4642 <= $unsigned(reg4494[(3'h4):(2'h3)]);
                      reg4643 <= reg4493[(3'h4):(3'h4)];
                    end
                  reg4644 <= (~|(((!forvar4593) ?
                          (reg4476 ?
                              forvar4597 : reg4473) : (reg4573 < reg4552)) ?
                      reg4478 : {(~&wire3772)}));
                  if ((8'hb6))
                    begin
                      reg4645 <= ($unsigned(((forvar4609 ? (8'hb6) : reg4571) ?
                          (reg4503 ?
                              reg4638 : forvar4470) : wire3771)) + (({(8'ha5)} ?
                          {reg4556} : (reg4462 > reg4471)) >>> ((&(8'h9c)) ~^ $signed(reg4477))));
                      reg4646 <= wire3773[(3'h5):(1'h0)];
                      reg4647 <= (reg4555[(1'h0):(1'h0)] >> $unsigned({$unsigned(wire3778)}));
                      reg4648 <= $signed(((|$unsigned(reg4549)) ?
                          ((reg4601 ?
                              forvar4459 : reg4487) ^~ (reg4617 ^ reg4597)) : ({reg4519} <<< (-(8'hb5)))));
                    end
                  else
                    begin
                      reg4645 <= (($signed($unsigned(reg4491)) || ((8'h9c) ?
                              reg4604 : ((8'h9f) ? reg4636 : reg4561))) ?
                          (((reg4516 | reg4535) ?
                                  (reg4471 ?
                                      reg4554 : reg4511) : $signed((8'hba))) ?
                              (8'haa) : (((8'hb4) >= (8'h9f)) ?
                                  (reg4466 ?
                                      reg4520 : reg4543) : (~|reg4500))) : ($signed((forvar4508 ?
                                  (8'h9c) : reg4560)) ?
                              {reg4586} : $unsigned((reg4646 != forvar4495))));
                      reg4646 <= reg4502[(2'h3):(1'h1)];
                      reg4647 <= reg4603;
                      reg4648 <= ($signed($signed(reg4646[(1'h1):(1'h0)])) ?
                          forvar4508[(1'h1):(1'h1)] : (wire3778 && $signed(reg4487[(1'h0):(1'h0)])));
                    end
                end
              for (forvar4649 = (1'h0); (forvar4649 < (1'h0)); forvar4649 = (forvar4649 + (1'h1)))
                begin
                  for (forvar4650 = (1'h0); (forvar4650 < (1'h1)); forvar4650 = (forvar4650 + (1'h1)))
                    begin
                      reg4651 <= reg4462;
                      reg4652 <= forvar4624;
                    end
                  if ({($unsigned((8'hb2)) | (^~wire3770))})
                    begin
                      reg4653 <= reg4528;
                      reg4654 <= reg4628;
                      reg4655 <= (8'hb2);
                      reg4656 <= (^~forvar4522);
                    end
                  else
                    begin
                      reg4653 <= reg4602[(2'h2):(2'h2)];
                      reg4654 <= (8'hb5);
                    end
                end
            end
        end
      reg4657 <= $signed(($signed(forvar4614[(1'h1):(1'h1)]) ^ reg4505));
      for (forvar4658 = (1'h0); (forvar4658 < (1'h1)); forvar4658 = (forvar4658 + (1'h1)))
        begin
          for (forvar4659 = (1'h0); (forvar4659 < (1'h1)); forvar4659 = (forvar4659 + (1'h1)))
            begin
              for (forvar4660 = (1'h0); (forvar4660 < (2'h3)); forvar4660 = (forvar4660 + (1'h1)))
                begin
                  for (forvar4661 = (1'h0); (forvar4661 < (2'h2)); forvar4661 = (forvar4661 + (1'h1)))
                    begin
                      reg4662 <= (($unsigned((!forvar4497)) ?
                              $unsigned(forvar4594[(4'h8):(3'h4)]) : reg4471) ?
                          reg4560 : reg4500[(4'ha):(3'h7)]);
                    end
                end
              if ((((8'hb5) ~^ ((reg4464 ?
                  reg4633 : reg4655) <<< reg4501[(4'h9):(1'h0)])) <<< (~&reg4537)))
                begin
                  if ($unsigned($unsigned(((reg4510 ?
                      forvar4658 : forvar4593) >> (reg4642 && (8'haf))))))
                    begin
                      reg4663 <= ((+{(reg4570 != reg4483)}) ?
                          reg4629[(4'ha):(3'h4)] : $signed((~|reg4559)));
                      reg4664 <= (-reg4626[(3'h5):(3'h5)]);
                      reg4665 <= ({reg4523[(2'h3):(2'h2)]} ?
                          ((^(wire3778 ? reg4479 : reg4591)) ?
                              (^~{forvar4604}) : $signed(forvar4610)) : reg4514[(4'h9):(3'h5)]);
                      reg4666 <= (((reg4499[(3'h4):(1'h1)] ?
                              reg4652[(3'h4):(2'h2)] : forvar4600[(3'h4):(2'h2)]) ^~ ($signed(reg4547) ?
                              (reg4652 == forvar4659) : forvar4531)) ?
                          (~|{$signed(reg4470)}) : $unsigned(($unsigned(forvar4531) < (8'h9e))));
                    end
                  else
                    begin
                      reg4663 <= wire3778[(3'h5):(1'h1)];
                      reg4664 <= reg4492[(4'he):(4'h9)];
                      reg4665 <= $signed(((~^$unsigned(forvar4485)) == {reg4527[(2'h3):(1'h0)]}));
                    end
                  for (forvar4667 = (1'h0); (forvar4667 < (1'h1)); forvar4667 = (forvar4667 + (1'h1)))
                    begin
                      reg4668 <= forvar4470;
                      reg4669 <= reg4484[(4'h8):(3'h4)];
                    end
                end
              else
                begin
                  for (forvar4663 = (1'h0); (forvar4663 < (2'h3)); forvar4663 = (forvar4663 + (1'h1)))
                    begin
                      reg4664 <= $signed(forvar4546[(3'h7):(2'h2)]);
                      reg4665 <= reg4581[(4'hb):(4'h8)];
                      reg4666 <= ($unsigned((~forvar4604[(3'h4):(3'h4)])) ?
                          $unsigned((forvar4610 ?
                              (|reg4613) : ((8'ha5) >>> (8'hba)))) : $signed($unsigned({reg4524})));
                    end
                end
            end
          reg4670 <= reg4570[(2'h2):(2'h2)];
          if ($unsigned(($signed($unsigned(reg4526)) & (!wire3775))))
            begin
              for (forvar4671 = (1'h0); (forvar4671 < (1'h1)); forvar4671 = (forvar4671 + (1'h1)))
                begin
                  reg4672 <= (forvar4581 > ((reg4604[(1'h0):(1'h0)] >>> reg4484[(2'h3):(1'h1)]) * reg4492));
                  if ((!reg4607))
                    begin
                      reg4673 <= ((reg4488 ?
                              ((+reg4585) ?
                                  $unsigned(forvar4604) : (reg4503 >= forvar4485)) : $signed($signed(wire3775))) ?
                          forvar4667 : reg4629[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg4673 <= (+(reg4577[(4'h9):(2'h2)] ?
                          reg4490[(4'hf):(3'h6)] : (reg4593 ^~ $unsigned(reg4564))));
                    end
                end
              if ((forvar4541 ?
                  ((forvar4581 ?
                      (!reg4611) : reg4604) >> ((reg4556 || (8'ha2)) | $signed(reg4603))) : (reg4576 ~^ (^~(~|wire4587)))))
                begin
                  for (forvar4674 = (1'h0); (forvar4674 < (2'h2)); forvar4674 = (forvar4674 + (1'h1)))
                    begin
                      reg4675 <= $signed(forvar4650);
                      reg4676 <= forvar4497[(2'h3):(1'h0)];
                    end
                  reg4677 <= ((^(((8'h9c) - reg4566) || (forvar4485 == reg4566))) | forvar4572);
                  for (forvar4678 = (1'h0); (forvar4678 < (2'h3)); forvar4678 = (forvar4678 + (1'h1)))
                    begin
                      reg4679 <= (^~($signed((reg4524 ? reg4492 : reg4576)) ?
                          (((8'ha6) ?
                              forvar4614 : reg4536) << (^~(8'ha9))) : (&forvar4610)));
                      reg4680 <= {forvar4503};
                      reg4681 <= reg4549;
                      reg4682 <= forvar4521[(2'h2):(2'h2)];
                    end
                  for (forvar4683 = (1'h0); (forvar4683 < (2'h2)); forvar4683 = (forvar4683 + (1'h1)))
                    begin
                      reg4684 <= ((|$unsigned((reg4472 < reg4524))) != (!((reg4665 ?
                          reg4560 : reg4506) - reg4530[(4'h9):(1'h1)])));
                      reg4685 <= $signed($signed((!{reg4574})));
                      reg4686 <= (($unsigned(forvar4494) << $signed(forvar4531)) >>> (~^{(8'hb2)}));
                    end
                end
              else
                begin
                  for (forvar4674 = (1'h0); (forvar4674 < (2'h3)); forvar4674 = (forvar4674 + (1'h1)))
                    begin
                      reg4675 <= $signed(wire4457[(4'he):(4'hc)]);
                      reg4676 <= ((~(^$signed((8'h9e)))) >= reg4629[(2'h3):(2'h2)]);
                    end
                end
            end
          else
            begin
              for (forvar4671 = (1'h0); (forvar4671 < (2'h3)); forvar4671 = (forvar4671 + (1'h1)))
                begin
                  reg4672 <= ((~^((forvar4658 > reg4493) ?
                          $unsigned(reg4486) : (^forvar4658))) ?
                      reg4473 : $unsigned((+{wire3773})));
                end
            end
          for (forvar4687 = (1'h0); (forvar4687 < (1'h1)); forvar4687 = (forvar4687 + (1'h1)))
            begin
              reg4688 <= forvar4592[(1'h0):(1'h0)];
              for (forvar4689 = (1'h0); (forvar4689 < (1'h0)); forvar4689 = (forvar4689 + (1'h1)))
                begin
                  reg4690 <= $signed($unsigned($unsigned(reg4478[(1'h0):(1'h0)])));
                  if ($unsigned($signed(((forvar4689 ?
                      forvar4659 : reg4609) * (forvar4563 & reg4593)))))
                    begin
                      reg4691 <= ((reg4614[(4'hc):(2'h3)] + $signed((8'hb3))) ?
                          (~^(((8'had) - forvar4476) & (~&reg4476))) : $unsigned($unsigned($unsigned(forvar4532))));
                      reg4692 <= $signed(forvar4484[(3'h6):(1'h0)]);
                      reg4693 <= (-wire3773[(4'h9):(4'h9)]);
                    end
                  else
                    begin
                      reg4691 <= (&reg4504);
                    end
                  reg4694 <= {(8'ha5)};
                end
              if ((($signed({reg4516}) ?
                      ((+forvar4503) ~^ $signed((8'ha4))) : ($signed((8'ha5)) > (!reg4640))) ?
                  $unsigned($signed((^forvar4667))) : ($signed(reg4547[(3'h5):(1'h1)]) ?
                      reg4572[(2'h2):(1'h1)] : reg4479)))
                begin
                  for (forvar4695 = (1'h0); (forvar4695 < (1'h1)); forvar4695 = (forvar4695 + (1'h1)))
                    begin
                      reg4696 <= ($unsigned({$signed(reg4676)}) ?
                          (8'hae) : reg4641[(3'h6):(2'h2)]);
                      reg4697 <= $signed($unsigned((&(forvar4592 ?
                          reg4568 : reg4549))));
                      reg4698 <= forvar4460[(2'h2):(2'h2)];
                      reg4699 <= (~&reg4594);
                    end
                  for (forvar4700 = (1'h0); (forvar4700 < (2'h2)); forvar4700 = (forvar4700 + (1'h1)))
                    begin
                      reg4701 <= (reg4628[(1'h0):(1'h0)] ~^ $signed($signed((reg4485 ^~ (8'ha5)))));
                    end
                end
              else
                begin
                  for (forvar4695 = (1'h0); (forvar4695 < (1'h0)); forvar4695 = (forvar4695 + (1'h1)))
                    begin
                      reg4696 <= $signed(({reg4585[(2'h2):(1'h0)]} << reg4561));
                      reg4697 <= $unsigned(($unsigned($signed(reg4632)) ?
                          reg4607 : ($unsigned(forvar4611) ?
                              (forvar4624 || forvar4531) : reg4679[(4'hb):(2'h3)])));
                    end
                end
              for (forvar4702 = (1'h0); (forvar4702 < (2'h2)); forvar4702 = (forvar4702 + (1'h1)))
                begin
                  reg4703 <= (($unsigned($unsigned(reg4644)) ^~ reg4549) & $unsigned(reg4475[(4'hb):(1'h0)]));
                end
            end
        end
      for (forvar4704 = (1'h0); (forvar4704 < (1'h0)); forvar4704 = (forvar4704 + (1'h1)))
        begin
          for (forvar4705 = (1'h0); (forvar4705 < (2'h2)); forvar4705 = (forvar4705 + (1'h1)))
            begin
              if ({$unsigned((reg4698 <= (~^forvar4459)))})
                begin
                  for (forvar4706 = (1'h0); (forvar4706 < (2'h3)); forvar4706 = (forvar4706 + (1'h1)))
                    begin
                      reg4707 <= reg4471[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar4706 = (1'h0); (forvar4706 < (2'h3)); forvar4706 = (forvar4706 + (1'h1)))
                    begin
                      reg4707 <= (forvar4661 < reg4542);
                      reg4708 <= forvar4589;
                    end
                  for (forvar4709 = (1'h0); (forvar4709 < (2'h3)); forvar4709 = (forvar4709 + (1'h1)))
                    begin
                      reg4710 <= forvar4606[(3'h4):(2'h2)];
                      reg4711 <= forvar4689[(3'h7):(1'h1)];
                      reg4712 <= $signed(($unsigned((reg4646 ?
                          reg4685 : reg4542)) ~^ (reg4540 ?
                          reg4677[(3'h4):(2'h2)] : (reg4498 ?
                              forvar4659 : forvar4635))));
                    end
                end
              for (forvar4713 = (1'h0); (forvar4713 < (1'h0)); forvar4713 = (forvar4713 + (1'h1)))
                begin
                  for (forvar4714 = (1'h0); (forvar4714 < (2'h2)); forvar4714 = (forvar4714 + (1'h1)))
                    begin
                      reg4715 <= $signed((!(&(forvar4494 < reg4506))));
                      reg4716 <= ((((reg4554 ^~ forvar4619) ?
                          (reg4640 ?
                              reg4703 : reg4496) : {forvar4678}) >> ((forvar4606 ?
                              forvar4598 : reg4595) ?
                          $unsigned(reg4647) : {reg4644})) | (reg4641 <<< reg4582[(4'hc):(2'h2)]));
                    end
                  if (($signed(((forvar4702 - reg4562) ?
                          $unsigned(reg4591) : (forvar4614 ?
                              forvar4683 : reg4708))) ?
                      ($unsigned((8'ha1)) - $unsigned($signed(reg4655))) : forvar4667[(1'h1):(1'h1)]))
                    begin
                      reg4717 <= $unsigned((^reg4498[(3'h4):(2'h2)]));
                      reg4718 <= (-forvar4600[(2'h3):(1'h0)]);
                      reg4719 <= $signed(forvar4522);
                      reg4720 <= $signed({forvar4604[(2'h3):(1'h1)]});
                    end
                  else
                    begin
                      reg4717 <= ({(|(~|reg4574))} ~^ $signed(reg4581[(3'h6):(3'h5)]));
                    end
                  for (forvar4721 = (1'h0); (forvar4721 < (1'h0)); forvar4721 = (forvar4721 + (1'h1)))
                    begin
                      reg4722 <= reg4499[(2'h2):(1'h1)];
                      reg4723 <= $signed($unsigned((~$unsigned(forvar4489))));
                      reg4724 <= (8'hb9);
                      reg4725 <= ($unsigned($signed(forvar4594[(2'h3):(1'h0)])) ?
                          (&{$signed(reg4609)}) : forvar4494);
                    end
                  if (reg4563)
                    begin
                      reg4726 <= ($unsigned($signed($signed(reg4642))) == (-{$signed(forvar4593)}));
                    end
                  else
                    begin
                      reg4726 <= reg4592[(1'h0):(1'h0)];
                      reg4727 <= forvar4660[(4'ha):(3'h6)];
                      reg4728 <= reg4636;
                    end
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3780  (y, clk, wire3784, wire3783, wire3782, wire3781);
  output wire [(32'h11ec):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire3784;
  input wire [(3'h5):(1'h0)] wire3783;
  input wire signed [(3'h6):(1'h0)] wire3782;
  input wire [(4'hd):(1'h0)] wire3781;
  wire [(3'h5):(1'h0)] wire4456;
  reg signed [(5'h10):(1'h0)] reg4452 = (1'h0);
  reg [(2'h3):(1'h0)] reg4449 = (1'h0);
  reg [(3'h6):(1'h0)] reg4455 = (1'h0);
  reg [(4'hd):(1'h0)] reg4454 = (1'h0);
  reg [(4'hd):(1'h0)] reg4453 = (1'h0);
  reg [(4'he):(1'h0)] forvar4452 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4451 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4450 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4449 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4448 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4447 = (1'h0);
  reg [(3'h6):(1'h0)] reg4446 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4445 = (1'h0);
  reg [(4'hb):(1'h0)] reg4444 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4443 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4442 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4441 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4434 = (1'h0);
  reg [(4'hf):(1'h0)] reg4440 = (1'h0);
  reg [(3'h6):(1'h0)] reg4439 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4438 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4437 = (1'h0);
  reg [(3'h5):(1'h0)] reg4436 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4435 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4434 = (1'h0);
  reg [(4'h9):(1'h0)] reg4433 = (1'h0);
  reg [(4'hc):(1'h0)] reg4432 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4431 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4430 = (1'h0);
  reg [(4'he):(1'h0)] reg4429 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4428 = (1'h0);
  reg [(4'hb):(1'h0)] reg4422 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4420 = (1'h0);
  reg [(4'hd):(1'h0)] reg4428 = (1'h0);
  reg [(5'h10):(1'h0)] reg4427 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4426 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4425 = (1'h0);
  reg [(2'h3):(1'h0)] reg4424 = (1'h0);
  reg [(4'he):(1'h0)] reg4423 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4422 = (1'h0);
  reg [(4'hb):(1'h0)] reg4421 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4420 = (1'h0);
  reg [(4'hc):(1'h0)] reg4419 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4418 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4417 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4416 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4415 = (1'h0);
  reg [(3'h7):(1'h0)] reg4414 = (1'h0);
  reg [(2'h2):(1'h0)] reg4413 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4411 = (1'h0);
  reg [(4'hf):(1'h0)] reg4412 = (1'h0);
  reg [(2'h2):(1'h0)] reg4411 = (1'h0);
  reg [(4'ha):(1'h0)] reg4410 = (1'h0);
  reg [(4'hb):(1'h0)] reg4409 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4408 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4407 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4406 = (1'h0);
  reg [(4'he):(1'h0)] forvar4405 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4401 = (1'h0);
  reg [(5'h10):(1'h0)] reg4399 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4394 = (1'h0);
  reg [(4'hb):(1'h0)] reg4404 = (1'h0);
  reg [(4'hd):(1'h0)] reg4403 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4402 = (1'h0);
  reg [(2'h3):(1'h0)] reg4401 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4400 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4399 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4398 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4397 = (1'h0);
  reg [(2'h3):(1'h0)] reg4396 = (1'h0);
  reg [(5'h10):(1'h0)] reg4395 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4394 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4393 = (1'h0);
  reg [(4'h8):(1'h0)] reg4392 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4391 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4390 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4384 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4389 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4388 = (1'h0);
  reg [(4'h8):(1'h0)] reg4387 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4386 = (1'h0);
  reg [(4'he):(1'h0)] reg4385 = (1'h0);
  reg [(2'h3):(1'h0)] reg4384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4383 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4382 = (1'h0);
  reg [(4'hd):(1'h0)] reg4381 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4380 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4379 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4378 = (1'h0);
  reg [(3'h5):(1'h0)] reg4377 = (1'h0);
  reg [(2'h2):(1'h0)] reg4376 = (1'h0);
  reg [(4'hf):(1'h0)] reg4375 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4374 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4373 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4371 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4366 = (1'h0);
  reg [(5'h10):(1'h0)] reg4363 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4372 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4371 = (1'h0);
  reg [(2'h3):(1'h0)] reg4370 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4369 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4368 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4367 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4366 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4365 = (1'h0);
  reg [(4'hd):(1'h0)] reg4364 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4363 = (1'h0);
  reg [(4'h9):(1'h0)] reg4362 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4361 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4360 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4359 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4358 = (1'h0);
  reg [(3'h5):(1'h0)] reg4357 = (1'h0);
  reg [(3'h6):(1'h0)] reg4352 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4351 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4348 = (1'h0);
  reg [(4'hb):(1'h0)] reg4356 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4355 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4354 = (1'h0);
  reg [(3'h4):(1'h0)] reg4353 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4352 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4351 = (1'h0);
  reg [(4'hb):(1'h0)] reg4350 = (1'h0);
  reg [(3'h5):(1'h0)] reg4349 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4348 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4347 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4346 = (1'h0);
  reg [(4'h8):(1'h0)] reg4337 = (1'h0);
  reg [(4'ha):(1'h0)] reg4333 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4345 = (1'h0);
  reg [(4'hf):(1'h0)] reg4344 = (1'h0);
  reg [(2'h2):(1'h0)] reg4343 = (1'h0);
  reg [(2'h3):(1'h0)] reg4342 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4341 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4340 = (1'h0);
  reg [(4'hb):(1'h0)] reg4339 = (1'h0);
  reg [(4'ha):(1'h0)] reg4338 = (1'h0);
  reg [(4'he):(1'h0)] forvar4337 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4336 = (1'h0);
  reg [(4'hf):(1'h0)] reg4335 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4334 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4333 = (1'h0);
  reg [(4'hd):(1'h0)] reg4332 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4331 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4330 = (1'h0);
  reg [(2'h3):(1'h0)] reg4329 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4320 = (1'h0);
  reg [(4'hf):(1'h0)] reg4328 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4327 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4326 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4325 = (1'h0);
  reg [(4'hb):(1'h0)] reg4324 = (1'h0);
  reg [(4'hd):(1'h0)] reg4323 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4322 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4321 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4320 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4319 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4318 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4317 = (1'h0);
  reg [(4'he):(1'h0)] reg4316 = (1'h0);
  reg [(4'hf):(1'h0)] reg4315 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4314 = (1'h0);
  reg [(2'h2):(1'h0)] reg4313 = (1'h0);
  reg [(2'h3):(1'h0)] reg4312 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4311 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4310 = (1'h0);
  reg [(4'hd):(1'h0)] reg4309 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4308 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4307 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4306 = (1'h0);
  reg [(4'he):(1'h0)] reg4300 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4299 = (1'h0);
  reg [(2'h3):(1'h0)] reg4297 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4305 = (1'h0);
  reg [(4'hd):(1'h0)] reg4304 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4303 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4302 = (1'h0);
  reg [(3'h7):(1'h0)] reg4301 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4300 = (1'h0);
  reg [(3'h6):(1'h0)] reg4299 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4298 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4297 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4296 = (1'h0);
  reg [(4'h8):(1'h0)] reg4295 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4294 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4293 = (1'h0);
  reg [(4'ha):(1'h0)] reg4292 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4291 = (1'h0);
  reg [(5'h10):(1'h0)] reg4290 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4289 = (1'h0);
  reg [(4'h8):(1'h0)] reg4288 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4287 = (1'h0);
  reg [(2'h3):(1'h0)] reg4286 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4285 = (1'h0);
  reg [(5'h10):(1'h0)] reg4284 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4283 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4282 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4281 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4280 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4279 = (1'h0);
  reg [(2'h3):(1'h0)] reg4278 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4277 = (1'h0);
  reg [(2'h3):(1'h0)] reg4276 = (1'h0);
  reg [(4'h9):(1'h0)] reg4275 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4274 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4273 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4272 = (1'h0);
  reg [(4'hc):(1'h0)] reg4271 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4270 = (1'h0);
  reg [(3'h5):(1'h0)] reg4269 = (1'h0);
  reg [(4'hb):(1'h0)] reg4268 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4267 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4266 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4265 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4264 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4242 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4263 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4262 = (1'h0);
  reg [(4'hc):(1'h0)] reg4261 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4260 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4259 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4258 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4250 = (1'h0);
  reg [(3'h5):(1'h0)] reg4257 = (1'h0);
  reg [(4'h9):(1'h0)] reg4256 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4255 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4254 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4253 = (1'h0);
  reg [(4'hf):(1'h0)] reg4252 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4251 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4250 = (1'h0);
  reg [(5'h10):(1'h0)] reg4249 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4248 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4247 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4246 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4245 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4244 = (1'h0);
  reg [(4'ha):(1'h0)] reg4243 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4242 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4241 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4239 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4235 = (1'h0);
  reg [(3'h4):(1'h0)] reg4240 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4239 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4238 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4237 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4236 = (1'h0);
  reg [(2'h3):(1'h0)] reg4235 = (1'h0);
  reg [(4'hb):(1'h0)] reg4234 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4233 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4232 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4231 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4230 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4229 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4228 = (1'h0);
  reg [(4'h9):(1'h0)] reg4227 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4226 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4225 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4224 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4223 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4219 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4223 = (1'h0);
  reg [(4'ha):(1'h0)] reg4222 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4221 = (1'h0);
  reg [(4'hb):(1'h0)] reg4220 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4219 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4218 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4211 = (1'h0);
  reg [(4'he):(1'h0)] reg4210 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4208 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4206 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4217 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4216 = (1'h0);
  reg [(3'h7):(1'h0)] reg4215 = (1'h0);
  reg [(3'h4):(1'h0)] reg4214 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4213 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4212 = (1'h0);
  reg [(3'h5):(1'h0)] reg4211 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4210 = (1'h0);
  reg [(4'hb):(1'h0)] reg4209 = (1'h0);
  reg [(4'he):(1'h0)] reg4208 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4207 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4206 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4194 = (1'h0);
  reg [(3'h6):(1'h0)] reg4205 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4204 = (1'h0);
  reg [(4'hd):(1'h0)] reg4203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4202 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4201 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4200 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4199 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4198 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4197 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4196 = (1'h0);
  reg [(4'hd):(1'h0)] reg4195 = (1'h0);
  reg [(2'h2):(1'h0)] reg4194 = (1'h0);
  reg [(3'h6):(1'h0)] reg4193 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4192 = (1'h0);
  reg [(4'hb):(1'h0)] reg4191 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4190 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4189 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4188 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4187 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4186 = (1'h0);
  reg [(4'ha):(1'h0)] reg4185 = (1'h0);
  reg [(4'hf):(1'h0)] reg4184 = (1'h0);
  reg [(4'hb):(1'h0)] reg4183 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4182 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4181 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4180 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4179 = (1'h0);
  reg [(3'h5):(1'h0)] reg4178 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4177 = (1'h0);
  reg [(4'hd):(1'h0)] reg4176 = (1'h0);
  reg [(3'h7):(1'h0)] reg4175 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4174 = (1'h0);
  reg [(2'h2):(1'h0)] reg4173 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4172 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4171 = (1'h0);
  reg [(4'he):(1'h0)] reg4170 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4169 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4168 = (1'h0);
  reg [(4'ha):(1'h0)] reg4167 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4166 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4165 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4164 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4163 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4162 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4161 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4160 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4159 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4158 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4157 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4156 = (1'h0);
  wire [(2'h2):(1'h0)] wire4154;
  reg [(4'he):(1'h0)] reg3930 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3929 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3928 = (1'h0);
  reg [(3'h5):(1'h0)] reg3927 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3926 = (1'h0);
  reg [(4'h8):(1'h0)] reg3925 = (1'h0);
  reg [(4'hd):(1'h0)] reg3924 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3923 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3922 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3921 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3920 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3919 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3918 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3917 = (1'h0);
  reg [(4'h8):(1'h0)] reg3916 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3915 = (1'h0);
  reg [(5'h10):(1'h0)] reg3914 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3913 = (1'h0);
  reg [(3'h4):(1'h0)] reg3912 = (1'h0);
  reg [(5'h10):(1'h0)] reg3911 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3908 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3910 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3907 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3909 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3908 = (1'h0);
  reg [(4'hb):(1'h0)] reg3907 = (1'h0);
  reg [(3'h4):(1'h0)] reg3906 = (1'h0);
  reg [(4'he):(1'h0)] reg3905 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3904 = (1'h0);
  reg [(2'h2):(1'h0)] reg3903 = (1'h0);
  reg [(4'he):(1'h0)] reg3902 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3901 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3900 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3899 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3898 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3897 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3896 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3895 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3894 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3893 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3858 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3871 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3870 = (1'h0);
  reg [(4'hf):(1'h0)] reg3869 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3865 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3861 = (1'h0);
  reg [(2'h2):(1'h0)] reg3857 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3838 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3833 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3852 = (1'h0);
  reg [(4'h8):(1'h0)] reg3848 = (1'h0);
  reg [(4'ha):(1'h0)] reg3892 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3891 = (1'h0);
  reg [(4'ha):(1'h0)] reg3890 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3889 = (1'h0);
  reg [(3'h5):(1'h0)] reg3888 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3887 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3886 = (1'h0);
  reg [(3'h6):(1'h0)] reg3886 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3885 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3884 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3883 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3879 = (1'h0);
  reg [(3'h7):(1'h0)] reg3877 = (1'h0);
  reg [(4'h8):(1'h0)] reg3882 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3881 = (1'h0);
  reg [(3'h6):(1'h0)] reg3880 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3879 = (1'h0);
  reg [(4'h8):(1'h0)] reg3878 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3877 = (1'h0);
  reg [(3'h7):(1'h0)] reg3876 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3875 = (1'h0);
  reg [(3'h5):(1'h0)] reg3874 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3873 = (1'h0);
  reg [(4'h8):(1'h0)] reg3872 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3871 = (1'h0);
  reg [(3'h5):(1'h0)] reg3870 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3869 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3868 = (1'h0);
  reg [(3'h4):(1'h0)] reg3867 = (1'h0);
  reg [(4'hd):(1'h0)] reg3866 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3865 = (1'h0);
  reg [(3'h5):(1'h0)] reg3864 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3862 = (1'h0);
  reg [(2'h3):(1'h0)] reg3863 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3862 = (1'h0);
  reg [(2'h2):(1'h0)] reg3861 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3860 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3859 = (1'h0);
  reg [(4'ha):(1'h0)] reg3858 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3857 = (1'h0);
  reg [(4'hd):(1'h0)] reg3856 = (1'h0);
  reg [(4'h8):(1'h0)] reg3855 = (1'h0);
  reg [(4'he):(1'h0)] reg3854 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3849 = (1'h0);
  reg [(4'h8):(1'h0)] reg3853 = (1'h0);
  reg [(2'h2):(1'h0)] reg3852 = (1'h0);
  reg [(4'hf):(1'h0)] reg3851 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3850 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3849 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3848 = (1'h0);
  reg [(3'h4):(1'h0)] reg3847 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3846 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3843 = (1'h0);
  reg [(5'h10):(1'h0)] reg3841 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3840 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3837 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3845 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3844 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3843 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3842 = (1'h0);
  reg [(4'he):(1'h0)] forvar3841 = (1'h0);
  reg [(3'h4):(1'h0)] reg3840 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3836 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3834 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3832 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3839 = (1'h0);
  reg [(4'h8):(1'h0)] reg3838 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3837 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3836 = (1'h0);
  reg [(3'h6):(1'h0)] reg3835 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3834 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3833 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3832 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3831 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3830 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3829 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3828 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3827 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3826 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3825 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3824 = (1'h0);
  reg [(3'h7):(1'h0)] reg3823 = (1'h0);
  reg [(4'hd):(1'h0)] reg3822 = (1'h0);
  reg [(5'h10):(1'h0)] reg3821 = (1'h0);
  reg [(4'h8):(1'h0)] reg3820 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3819 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3818 = (1'h0);
  reg [(3'h5):(1'h0)] reg3787 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3786 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3785 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3817 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3816 = (1'h0);
  reg [(4'h9):(1'h0)] reg3815 = (1'h0);
  reg [(4'h9):(1'h0)] reg3814 = (1'h0);
  reg [(3'h5):(1'h0)] reg3813 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3812 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3811 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3810 = (1'h0);
  reg [(2'h3):(1'h0)] reg3809 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3808 = (1'h0);
  reg [(4'hf):(1'h0)] reg3807 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3806 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3805 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3804 = (1'h0);
  reg [(4'hb):(1'h0)] reg3803 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3802 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3801 = (1'h0);
  reg [(4'hb):(1'h0)] reg3800 = (1'h0);
  reg [(4'h8):(1'h0)] reg3799 = (1'h0);
  reg [(4'he):(1'h0)] reg3798 = (1'h0);
  reg [(4'he):(1'h0)] reg3797 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3796 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3795 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3794 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3793 = (1'h0);
  reg [(4'ha):(1'h0)] reg3792 = (1'h0);
  reg [(4'hf):(1'h0)] reg3791 = (1'h0);
  reg [(4'hb):(1'h0)] reg3790 = (1'h0);
  reg [(2'h3):(1'h0)] reg3789 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3788 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3787 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3786 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3785 = (1'h0);
  assign y = {wire4456,
                 reg4452,
                 reg4449,
                 reg4455,
                 reg4454,
                 reg4453,
                 forvar4452,
                 reg4451,
                 reg4450,
                 forvar4449,
                 forvar4448,
                 forvar4447,
                 reg4446,
                 forvar4445,
                 reg4444,
                 reg4443,
                 forvar4442,
                 reg4441,
                 reg4434,
                 reg4440,
                 reg4439,
                 reg4438,
                 reg4437,
                 reg4436,
                 reg4435,
                 forvar4434,
                 reg4433,
                 reg4432,
                 reg4431,
                 forvar4430,
                 reg4429,
                 forvar4428,
                 reg4422,
                 reg4420,
                 reg4428,
                 reg4427,
                 reg4426,
                 reg4425,
                 reg4424,
                 reg4423,
                 forvar4422,
                 reg4421,
                 forvar4420,
                 reg4419,
                 reg4418,
                 forvar4417,
                 reg4416,
                 forvar4415,
                 reg4414,
                 reg4413,
                 forvar4411,
                 reg4412,
                 reg4411,
                 reg4410,
                 reg4409,
                 reg4408,
                 reg4407,
                 forvar4406,
                 forvar4405,
                 forvar4401,
                 reg4399,
                 reg4394,
                 reg4404,
                 reg4403,
                 reg4402,
                 reg4401,
                 reg4400,
                 forvar4399,
                 reg4398,
                 reg4397,
                 reg4396,
                 reg4395,
                 forvar4394,
                 reg4393,
                 reg4392,
                 reg4391,
                 reg4390,
                 forvar4384,
                 reg4389,
                 reg4388,
                 reg4387,
                 reg4386,
                 reg4385,
                 reg4384,
                 reg4383,
                 forvar4382,
                 reg4381,
                 forvar4380,
                 reg4379,
                 reg4378,
                 reg4377,
                 reg4376,
                 reg4375,
                 forvar4374,
                 forvar4373,
                 reg4371,
                 reg4366,
                 reg4363,
                 reg4372,
                 forvar4371,
                 reg4370,
                 reg4369,
                 reg4368,
                 reg4367,
                 forvar4366,
                 reg4365,
                 reg4364,
                 forvar4363,
                 reg4362,
                 forvar4361,
                 forvar4360,
                 reg4359,
                 reg4358,
                 reg4357,
                 reg4352,
                 forvar4351,
                 forvar4348,
                 reg4356,
                 reg4355,
                 reg4354,
                 reg4353,
                 forvar4352,
                 reg4351,
                 reg4350,
                 reg4349,
                 reg4348,
                 reg4347,
                 forvar4346,
                 reg4337,
                 reg4333,
                 reg4345,
                 reg4344,
                 reg4343,
                 reg4342,
                 reg4341,
                 reg4340,
                 reg4339,
                 reg4338,
                 forvar4337,
                 reg4336,
                 reg4335,
                 reg4334,
                 forvar4333,
                 reg4332,
                 forvar4331,
                 forvar4330,
                 reg4329,
                 reg4320,
                 reg4328,
                 reg4327,
                 forvar4326,
                 reg4325,
                 reg4324,
                 reg4323,
                 reg4322,
                 reg4321,
                 forvar4320,
                 reg4319,
                 forvar4318,
                 forvar4317,
                 reg4316,
                 reg4315,
                 forvar4314,
                 reg4313,
                 reg4312,
                 reg4311,
                 reg4310,
                 reg4309,
                 reg4308,
                 reg4307,
                 reg4306,
                 reg4300,
                 forvar4299,
                 reg4297,
                 reg4305,
                 reg4304,
                 reg4303,
                 reg4302,
                 reg4301,
                 forvar4300,
                 reg4299,
                 forvar4298,
                 forvar4297,
                 forvar4296,
                 reg4295,
                 forvar4294,
                 reg4293,
                 reg4292,
                 forvar4291,
                 reg4290,
                 reg4289,
                 reg4288,
                 reg4287,
                 reg4286,
                 reg4285,
                 reg4284,
                 forvar4283,
                 reg4282,
                 reg4281,
                 reg4280,
                 forvar4279,
                 reg4278,
                 forvar4277,
                 reg4276,
                 reg4275,
                 forvar4274,
                 reg4273,
                 reg4272,
                 reg4271,
                 reg4270,
                 reg4269,
                 reg4268,
                 reg4267,
                 forvar4266,
                 forvar4265,
                 forvar4264,
                 reg4242,
                 reg4263,
                 forvar4262,
                 reg4261,
                 reg4260,
                 reg4259,
                 reg4258,
                 forvar4250,
                 reg4257,
                 reg4256,
                 reg4255,
                 reg4254,
                 forvar4253,
                 reg4252,
                 reg4251,
                 reg4250,
                 reg4249,
                 forvar4248,
                 reg4247,
                 reg4246,
                 forvar4245,
                 reg4244,
                 reg4243,
                 forvar4242,
                 forvar4241,
                 reg4239,
                 forvar4235,
                 reg4240,
                 forvar4239,
                 reg4238,
                 reg4237,
                 reg4236,
                 reg4235,
                 reg4234,
                 forvar4233,
                 forvar4232,
                 reg4231,
                 reg4230,
                 reg4229,
                 reg4228,
                 reg4227,
                 reg4226,
                 reg4225,
                 reg4224,
                 forvar4223,
                 reg4219,
                 reg4223,
                 reg4222,
                 reg4221,
                 reg4220,
                 forvar4219,
                 forvar4218,
                 forvar4211,
                 reg4210,
                 forvar4208,
                 reg4206,
                 reg4217,
                 reg4216,
                 reg4215,
                 reg4214,
                 reg4213,
                 reg4212,
                 reg4211,
                 forvar4210,
                 reg4209,
                 reg4208,
                 reg4207,
                 forvar4206,
                 forvar4194,
                 reg4205,
                 reg4204,
                 reg4203,
                 reg4202,
                 reg4201,
                 reg4200,
                 reg4199,
                 reg4198,
                 reg4197,
                 reg4196,
                 reg4195,
                 reg4194,
                 reg4193,
                 forvar4192,
                 reg4191,
                 reg4190,
                 reg4189,
                 reg4188,
                 forvar4187,
                 reg4186,
                 reg4185,
                 reg4184,
                 reg4183,
                 reg4182,
                 reg4181,
                 forvar4180,
                 forvar4179,
                 reg4178,
                 reg4177,
                 reg4176,
                 reg4175,
                 forvar4174,
                 reg4173,
                 reg4172,
                 forvar4171,
                 reg4170,
                 reg4169,
                 forvar4168,
                 reg4167,
                 reg4166,
                 forvar4165,
                 forvar4164,
                 forvar4163,
                 forvar4162,
                 reg4161,
                 reg4160,
                 forvar4159,
                 reg4158,
                 forvar4157,
                 forvar4156,
                 wire4154,
                 reg3930,
                 reg3929,
                 forvar3928,
                 reg3927,
                 reg3926,
                 reg3925,
                 reg3924,
                 reg3923,
                 reg3922,
                 reg3921,
                 forvar3920,
                 forvar3919,
                 reg3918,
                 reg3917,
                 reg3916,
                 forvar3915,
                 reg3914,
                 reg3913,
                 reg3912,
                 reg3911,
                 forvar3908,
                 reg3910,
                 forvar3907,
                 reg3909,
                 reg3908,
                 reg3907,
                 reg3906,
                 reg3905,
                 reg3904,
                 reg3903,
                 reg3902,
                 forvar3901,
                 reg3900,
                 reg3899,
                 reg3898,
                 reg3897,
                 reg3896,
                 reg3895,
                 forvar3894,
                 forvar3893,
                 forvar3858,
                 forvar3871,
                 forvar3870,
                 reg3869,
                 forvar3865,
                 forvar3861,
                 reg3857,
                 forvar3838,
                 forvar3833,
                 forvar3852,
                 reg3848,
                 reg3892,
                 reg3891,
                 reg3890,
                 forvar3889,
                 reg3888,
                 reg3887,
                 forvar3886,
                 reg3886,
                 reg3885,
                 forvar3884,
                 reg3883,
                 forvar3879,
                 reg3877,
                 reg3882,
                 reg3881,
                 reg3880,
                 reg3879,
                 reg3878,
                 forvar3877,
                 reg3876,
                 reg3875,
                 reg3874,
                 reg3873,
                 reg3872,
                 reg3871,
                 reg3870,
                 forvar3869,
                 reg3868,
                 reg3867,
                 reg3866,
                 reg3865,
                 reg3864,
                 reg3862,
                 reg3863,
                 forvar3862,
                 reg3861,
                 reg3860,
                 reg3859,
                 reg3858,
                 forvar3857,
                 reg3856,
                 reg3855,
                 reg3854,
                 forvar3849,
                 reg3853,
                 reg3852,
                 reg3851,
                 reg3850,
                 reg3849,
                 forvar3848,
                 reg3847,
                 reg3846,
                 forvar3843,
                 reg3841,
                 forvar3840,
                 forvar3837,
                 reg3845,
                 reg3844,
                 reg3843,
                 reg3842,
                 forvar3841,
                 reg3840,
                 forvar3836,
                 reg3834,
                 forvar3832,
                 reg3839,
                 reg3838,
                 reg3837,
                 reg3836,
                 reg3835,
                 forvar3834,
                 reg3833,
                 reg3832,
                 reg3831,
                 reg3830,
                 reg3829,
                 reg3828,
                 reg3827,
                 reg3826,
                 reg3825,
                 forvar3824,
                 reg3823,
                 reg3822,
                 reg3821,
                 reg3820,
                 reg3819,
                 forvar3818,
                 reg3787,
                 forvar3786,
                 forvar3785,
                 reg3817,
                 reg3816,
                 reg3815,
                 reg3814,
                 reg3813,
                 reg3812,
                 reg3811,
                 reg3810,
                 reg3809,
                 reg3808,
                 reg3807,
                 forvar3806,
                 reg3805,
                 reg3804,
                 reg3803,
                 reg3802,
                 reg3801,
                 reg3800,
                 reg3799,
                 reg3798,
                 reg3797,
                 reg3796,
                 forvar3795,
                 forvar3794,
                 reg3793,
                 reg3792,
                 reg3791,
                 reg3790,
                 reg3789,
                 reg3788,
                 forvar3787,
                 reg3786,
                 reg3785,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (((wire3784 != (~^(wire3783 ? (8'h9e) : wire3781))) ?
          $signed({(~|wire3781)}) : $unsigned(((~&(8'hb6)) > ((8'ha8) | (8'h9f))))))
        begin
          if (wire3781)
            begin
              reg3785 <= $signed(wire3782[(3'h6):(2'h3)]);
              if ($unsigned((((wire3781 ? (8'hb1) : wire3784) ?
                      wire3784[(3'h5):(2'h2)] : $signed(reg3785)) ?
                  $signed(((8'ha8) >> reg3785)) : (wire3781 > $signed(wire3781)))))
                begin
                  reg3786 <= (^~((~^(^wire3781)) && wire3784[(3'h5):(3'h4)]));
                  for (forvar3787 = (1'h0); (forvar3787 < (2'h3)); forvar3787 = (forvar3787 + (1'h1)))
                    begin
                      reg3788 <= (($unsigned((reg3786 ? wire3784 : wire3784)) ?
                              (~^$unsigned(reg3786)) : $signed($unsigned((8'had)))) ?
                          ($signed($signed(wire3782)) ?
                              wire3781 : wire3782[(3'h6):(3'h6)]) : (($signed(wire3782) ~^ wire3783[(3'h5):(3'h5)]) << {wire3782[(3'h4):(3'h4)]}));
                      reg3789 <= ({$signed((wire3783 ?
                              reg3786 : wire3782))} * (wire3781 ^ (^(~&wire3784))));
                      reg3790 <= ({$signed((8'hb8))} * ({$signed(reg3789)} ?
                          {reg3789} : $signed($signed(reg3788))));
                      reg3791 <= ((wire3781[(3'h5):(2'h2)] ?
                          (^~$signed(wire3783)) : (((8'ha0) ?
                              reg3785 : reg3790) - (reg3786 - wire3784))) >= $unsigned($unsigned((8'ha6))));
                    end
                  if ((((((8'ha2) - (8'ha7)) | (~|wire3782)) <= (+(reg3790 >= (8'hb7)))) ?
                      (^$unsigned(wire3782)) : ((-$unsigned(reg3789)) >= reg3786)))
                    begin
                      reg3792 <= ((^~((-(8'hb5)) >> (reg3790 >= (8'h9d)))) < (reg3785[(1'h0):(1'h0)] ?
                          $signed((reg3785 ?
                              reg3785 : (8'ha7))) : (|{reg3789})));
                      reg3793 <= (($signed((wire3783 ^ reg3790)) * wire3781[(4'hc):(1'h0)]) ?
                          (wire3784[(1'h0):(1'h0)] ?
                              reg3790[(3'h7):(2'h2)] : $signed($signed(forvar3787))) : reg3788);
                    end
                  else
                    begin
                      reg3792 <= $signed({($signed(reg3791) ^ (wire3783 ~^ (8'h9d)))});
                    end
                end
              else
                begin
                  reg3786 <= reg3785[(1'h0):(1'h0)];
                  for (forvar3787 = (1'h0); (forvar3787 < (1'h0)); forvar3787 = (forvar3787 + (1'h1)))
                    begin
                      reg3788 <= (-wire3784);
                    end
                  if ($signed((&(~^{wire3784}))))
                    begin
                      reg3789 <= reg3790;
                    end
                  else
                    begin
                      reg3789 <= (((~^((8'hb3) != wire3781)) >> ((reg3785 ^ reg3788) ?
                          {reg3786} : forvar3787[(1'h0):(1'h0)])) ~^ $unsigned((~wire3782)));
                      reg3790 <= {(~|((reg3785 * reg3788) >>> $signed(reg3790)))};
                    end
                end
              for (forvar3794 = (1'h0); (forvar3794 < (2'h2)); forvar3794 = (forvar3794 + (1'h1)))
                begin
                  for (forvar3795 = (1'h0); (forvar3795 < (2'h3)); forvar3795 = (forvar3795 + (1'h1)))
                    begin
                      reg3796 <= reg3789;
                      reg3797 <= $unsigned((reg3792 ?
                          reg3791[(4'ha):(3'h6)] : $unsigned((~&forvar3787))));
                      reg3798 <= ((($unsigned(reg3788) ?
                                  forvar3787[(1'h1):(1'h0)] : {forvar3794}) ?
                              (reg3797[(1'h0):(1'h0)] ?
                                  (8'haa) : {(8'h9e)}) : ((-reg3790) != (|wire3781))) ?
                          ({$unsigned(reg3786)} < reg3792[(2'h3):(1'h1)]) : $signed((!reg3786)));
                    end
                  if ((((^$signed(wire3784)) ~^ $signed((forvar3787 + forvar3795))) ?
                      $unsigned((+(^~(8'hb7)))) : {$signed($unsigned(reg3786))}))
                    begin
                      reg3799 <= reg3785;
                      reg3800 <= $unsigned($signed($unsigned(wire3782[(2'h3):(2'h3)])));
                      reg3801 <= $signed((reg3800[(4'h9):(3'h4)] ?
                          reg3793 : forvar3787));
                      reg3802 <= $unsigned((forvar3795[(3'h5):(1'h1)] ?
                          (&reg3796[(2'h3):(1'h0)]) : (^$unsigned(reg3800))));
                    end
                  else
                    begin
                      reg3799 <= $signed(((8'hac) ?
                          $unsigned((reg3785 + reg3793)) : (reg3792 ?
                              reg3786[(2'h3):(1'h1)] : (^~reg3793))));
                      reg3800 <= ({$unsigned((~&reg3802))} ?
                          ($unsigned(reg3801[(2'h2):(1'h1)]) ?
                              (+(^~reg3789)) : ($signed(reg3790) == $signed(reg3791))) : $unsigned($unsigned($signed((8'haa)))));
                      reg3801 <= $unsigned({forvar3787});
                      reg3802 <= reg3796;
                    end
                  if (reg3785[(2'h3):(2'h3)])
                    begin
                      reg3803 <= (-reg3789[(2'h2):(1'h0)]);
                      reg3804 <= ($unsigned($signed((reg3786 ?
                          reg3799 : reg3792))) <= $unsigned(((&(8'ha1)) ?
                          $unsigned((8'ha4)) : $unsigned((8'hb7)))));
                      reg3805 <= ((~&((reg3791 ? reg3789 : reg3793) ?
                          $unsigned(reg3792) : (!wire3781))) != (reg3792[(3'h4):(2'h3)] << reg3799));
                    end
                  else
                    begin
                      reg3803 <= {reg3803[(3'h5):(1'h1)]};
                      reg3804 <= ((reg3799[(1'h1):(1'h1)] + (wire3784 ?
                          (reg3805 ?
                              reg3804 : wire3783) : $unsigned(reg3791))) != {((&(8'haf)) ?
                              {reg3790} : wire3781[(3'h6):(3'h6)])});
                    end
                end
              if ($signed((&wire3781)))
                begin
                  for (forvar3806 = (1'h0); (forvar3806 < (2'h2)); forvar3806 = (forvar3806 + (1'h1)))
                    begin
                      reg3807 <= reg3793;
                      reg3808 <= $signed($unsigned($unsigned(((8'hb1) ?
                          reg3789 : reg3805))));
                      reg3809 <= (reg3807 - (+$unsigned($unsigned(forvar3795))));
                    end
                  if (reg3805[(2'h2):(1'h1)])
                    begin
                      reg3810 <= forvar3806;
                      reg3811 <= wire3783;
                      reg3812 <= reg3791[(4'hc):(2'h2)];
                      reg3813 <= reg3808;
                    end
                  else
                    begin
                      reg3810 <= ((reg3797[(4'he):(3'h7)] * (-reg3802[(3'h6):(3'h5)])) <<< (&(8'ha2)));
                      reg3811 <= (reg3807 + (reg3813 != ($unsigned((8'hb7)) >> wire3783)));
                      reg3812 <= $unsigned((&(+reg3793)));
                      reg3813 <= ({((reg3800 && reg3785) >> {(8'haf)})} ?
                          (reg3812 ?
                              (reg3788 ?
                                  (~forvar3795) : (8'haf)) : (&{(8'ha7)})) : $signed((~&reg3805[(2'h2):(2'h2)])));
                    end
                  if ($unsigned({($unsigned((8'ha7)) ?
                          $signed((8'hb4)) : (reg3809 >= reg3788))}))
                    begin
                      reg3814 <= reg3812[(2'h2):(2'h2)];
                      reg3815 <= $signed($signed(reg3807[(4'ha):(4'h9)]));
                      reg3816 <= reg3804[(1'h1):(1'h0)];
                      reg3817 <= ((reg3808[(4'hc):(4'hb)] ?
                              (8'hb4) : (&reg3816[(3'h5):(1'h1)])) ?
                          ({reg3808[(3'h4):(1'h0)]} ~^ $signed((|wire3783))) : reg3796);
                    end
                  else
                    begin
                      reg3814 <= reg3812;
                      reg3815 <= ($unsigned((~^(reg3815 ?
                          forvar3787 : reg3788))) && (({wire3782} >= (|(8'ha6))) - $unsigned($signed(reg3792))));
                      reg3816 <= (~&{$signed((~^reg3791))});
                    end
                end
              else
                begin
                  for (forvar3806 = (1'h0); (forvar3806 < (2'h2)); forvar3806 = (forvar3806 + (1'h1)))
                    begin
                      reg3807 <= $unsigned((&{(reg3813 ? reg3790 : reg3812)}));
                    end
                  if (($unsigned((reg3817[(3'h7):(3'h5)] ?
                      (&reg3791) : $unsigned(wire3782))) == (^~{(reg3809 ?
                          reg3807 : reg3792)})))
                    begin
                      reg3808 <= (&$signed(($signed(reg3813) ?
                          (forvar3806 | reg3800) : forvar3806)));
                      reg3809 <= reg3785[(2'h3):(1'h1)];
                      reg3810 <= $unsigned(((^$signed(forvar3787)) < (~^$signed(forvar3806))));
                    end
                  else
                    begin
                      reg3808 <= reg3802;
                      reg3809 <= reg3786[(3'h7):(1'h1)];
                      reg3810 <= wire3782[(2'h3):(1'h0)];
                      reg3811 <= (reg3815 == (~^(reg3808[(4'he):(4'hd)] <= $signed(reg3814))));
                    end
                end
            end
          else
            begin
              for (forvar3785 = (1'h0); (forvar3785 < (2'h3)); forvar3785 = (forvar3785 + (1'h1)))
                begin
                  for (forvar3786 = (1'h0); (forvar3786 < (2'h2)); forvar3786 = (forvar3786 + (1'h1)))
                    begin
                      reg3787 <= ($signed(reg3811) ?
                          {(~^reg3793[(1'h0):(1'h0)])} : {(wire3782[(1'h0):(1'h0)] ^~ $unsigned(wire3781))});
                    end
                end
            end
          for (forvar3818 = (1'h0); (forvar3818 < (2'h3)); forvar3818 = (forvar3818 + (1'h1)))
            begin
              reg3819 <= {($signed((|reg3796)) - $signed((wire3781 ?
                      (8'h9c) : reg3788)))};
              if ($unsigned(reg3819[(1'h0):(1'h0)]))
                begin
                  reg3820 <= $unsigned({reg3787});
                end
              else
                begin
                  if (reg3809[(2'h2):(1'h0)])
                    begin
                      reg3820 <= $unsigned(((|reg3786[(3'h7):(2'h3)]) ?
                          $unsigned((reg3810 - reg3814)) : {{(8'hb9)}}));
                      reg3821 <= (-(8'hb8));
                    end
                  else
                    begin
                      reg3820 <= $signed(({{reg3817}} > reg3815[(3'h5):(2'h2)]));
                      reg3821 <= reg3808[(4'he):(4'ha)];
                      reg3822 <= ($signed((reg3809[(1'h1):(1'h1)] ?
                          (reg3788 > wire3781) : $unsigned(reg3801))) || ((~(forvar3787 <<< reg3787)) <= reg3817));
                      reg3823 <= (~^reg3807);
                    end
                  for (forvar3824 = (1'h0); (forvar3824 < (1'h1)); forvar3824 = (forvar3824 + (1'h1)))
                    begin
                      reg3825 <= forvar3818;
                      reg3826 <= reg3816;
                      reg3827 <= reg3799[(1'h1):(1'h0)];
                    end
                  if ((8'ha6))
                    begin
                      reg3828 <= (reg3804[(1'h1):(1'h0)] ?
                          ({(+reg3790)} ?
                              $unsigned(reg3817) : reg3785) : (((^reg3812) ?
                                  (!(8'had)) : $unsigned(reg3793)) ?
                              ($unsigned(reg3796) ?
                                  (~&(8'haf)) : (-reg3826)) : (|(~^reg3790))));
                      reg3829 <= reg3803;
                      reg3830 <= $signed($unsigned($unsigned(forvar3824)));
                    end
                  else
                    begin
                      reg3828 <= (|reg3822);
                      reg3829 <= reg3785;
                    end
                  if ((~^$unsigned((reg3823[(3'h5):(2'h2)] | (forvar3794 != reg3797)))))
                    begin
                      reg3831 <= wire3783;
                    end
                  else
                    begin
                      reg3831 <= (8'hb6);
                    end
                end
            end
        end
      else
        begin
          reg3785 <= ($signed($signed(((8'ha6) ^ reg3789))) ?
              forvar3794[(4'hb):(4'hb)] : reg3810[(4'h8):(3'h7)]);
        end
      if ({forvar3818[(3'h5):(2'h3)]})
        begin
          if (reg3813[(3'h5):(3'h4)])
            begin
              if (($signed((|(wire3781 <<< reg3828))) ?
                  reg3798[(3'h6):(2'h2)] : $signed((8'hab))))
                begin
                  reg3832 <= {forvar3818};
                  reg3833 <= ($signed((~^$signed(reg3826))) ?
                      reg3827[(1'h1):(1'h0)] : (|(reg3799 ?
                          (reg3810 ? reg3828 : reg3797) : $unsigned(reg3821))));
                  for (forvar3834 = (1'h0); (forvar3834 < (1'h0)); forvar3834 = (forvar3834 + (1'h1)))
                    begin
                      reg3835 <= $signed((~&((reg3800 + forvar3785) ~^ $signed(reg3786))));
                      reg3836 <= ((~$signed(((8'hba) ? reg3815 : (8'hb0)))) ?
                          $signed(($signed(reg3786) >= $signed(reg3820))) : {wire3782[(2'h2):(1'h0)]});
                      reg3837 <= (8'ha4);
                    end
                  if ($unsigned((~^reg3790[(3'h7):(1'h1)])))
                    begin
                      reg3838 <= (reg3815 * reg3803[(1'h0):(1'h0)]);
                      reg3839 <= (reg3793[(1'h0):(1'h0)] ^~ ($unsigned($unsigned(reg3797)) >>> (+{reg3832})));
                    end
                  else
                    begin
                      reg3838 <= $unsigned($unsigned((~^$unsigned(reg3839))));
                      reg3839 <= reg3821[(4'hc):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar3832 = (1'h0); (forvar3832 < (1'h0)); forvar3832 = (forvar3832 + (1'h1)))
                    begin
                      reg3833 <= (+(((~forvar3794) ?
                              reg3789 : $unsigned(reg3822)) ?
                          $signed($unsigned(forvar3786)) : reg3796[(2'h3):(1'h0)]));
                      reg3834 <= reg3822;
                    end
                  reg3835 <= (~^(8'h9e));
                  for (forvar3836 = (1'h0); (forvar3836 < (1'h0)); forvar3836 = (forvar3836 + (1'h1)))
                    begin
                      reg3837 <= reg3826[(4'h8):(3'h5)];
                      reg3838 <= $signed($signed($unsigned(reg3792[(2'h2):(2'h2)])));
                      reg3839 <= $unsigned((^(&(-wire3783))));
                      reg3840 <= $signed({((reg3797 ?
                              wire3781 : reg3833) >> (^reg3829))});
                    end
                  for (forvar3841 = (1'h0); (forvar3841 < (1'h1)); forvar3841 = (forvar3841 + (1'h1)))
                    begin
                      reg3842 <= (reg3786[(1'h0):(1'h0)] + wire3781);
                      reg3843 <= forvar3824;
                      reg3844 <= ((~^((reg3836 != reg3785) ?
                              reg3791[(3'h4):(2'h3)] : (reg3819 ?
                                  reg3812 : reg3798))) ?
                          (($unsigned(reg3837) ?
                                  (8'hb7) : wire3783[(2'h2):(1'h1)]) ?
                              ($unsigned(reg3787) ^ (reg3800 >> reg3826)) : ((reg3816 ?
                                  (8'hae) : reg3833) >>> reg3842)) : reg3837[(4'hb):(2'h2)]);
                      reg3845 <= reg3835;
                    end
                end
            end
          else
            begin
              if ($unsigned(($signed((~&forvar3832)) ?
                  $unsigned((+reg3835)) : (reg3796[(1'h1):(1'h1)] <<< {forvar3806}))))
                begin
                  if (((reg3787 - reg3832) ?
                      $signed(reg3809) : reg3811[(4'ha):(3'h7)]))
                    begin
                      reg3832 <= $unsigned(forvar3786);
                      reg3833 <= ({$unsigned($unsigned(reg3804))} ?
                          forvar3818[(3'h7):(1'h1)] : (((+reg3843) ?
                              reg3802[(3'h7):(3'h5)] : (^reg3802)) && $signed(((8'ha1) & reg3811))));
                      reg3834 <= ($signed(wire3784[(2'h2):(1'h0)]) ?
                          ($signed((reg3801 <= reg3801)) ?
                              (~&$unsigned(reg3844)) : (reg3797 ?
                                  $unsigned(reg3812) : (8'hb4))) : $signed((|forvar3836[(3'h5):(3'h5)])));
                    end
                  else
                    begin
                      reg3832 <= forvar3832;
                      reg3833 <= wire3784;
                    end
                  reg3835 <= forvar3785;
                  reg3836 <= ((reg3791[(3'h4):(2'h2)] >> reg3843) ?
                      $signed(({wire3782} - $signed(reg3820))) : $unsigned($unsigned($signed(reg3803))));
                end
              else
                begin
                  for (forvar3832 = (1'h0); (forvar3832 < (2'h3)); forvar3832 = (forvar3832 + (1'h1)))
                    begin
                      reg3833 <= (({$signed(reg3789)} - $unsigned((!reg3821))) || $unsigned(reg3811[(4'ha):(3'h5)]));
                      reg3834 <= reg3790[(4'h9):(4'h9)];
                      reg3835 <= $signed(((8'hb1) && $unsigned((reg3813 ^ reg3811))));
                      reg3836 <= (~^$unsigned((((8'hac) > reg3822) >>> $unsigned((8'h9f)))));
                    end
                  for (forvar3837 = (1'h0); (forvar3837 < (2'h3)); forvar3837 = (forvar3837 + (1'h1)))
                    begin
                      reg3838 <= $signed((~^(&(~^reg3835))));
                      reg3839 <= reg3787[(2'h3):(1'h0)];
                    end
                end
              if ((|(~|(8'ha0))))
                begin
                  for (forvar3840 = (1'h0); (forvar3840 < (2'h3)); forvar3840 = (forvar3840 + (1'h1)))
                    begin
                      reg3841 <= $signed(reg3817[(3'h6):(2'h2)]);
                      reg3842 <= (reg3789[(1'h1):(1'h1)] ?
                          (~$signed({reg3792})) : wire3781[(4'ha):(4'h9)]);
                    end
                  for (forvar3843 = (1'h0); (forvar3843 < (2'h3)); forvar3843 = (forvar3843 + (1'h1)))
                    begin
                      reg3844 <= (+reg3841[(1'h0):(1'h0)]);
                    end
                  if (reg3791)
                    begin
                      reg3845 <= $signed((^$unsigned((^reg3820))));
                    end
                  else
                    begin
                      reg3845 <= $signed(($signed($unsigned((8'h9d))) ?
                          $signed(forvar3840) : {reg3830[(2'h2):(1'h0)]}));
                      reg3846 <= reg3821[(4'hc):(3'h6)];
                      reg3847 <= $signed($signed((-(reg3809 | reg3820))));
                    end
                end
              else
                begin
                  for (forvar3840 = (1'h0); (forvar3840 < (1'h1)); forvar3840 = (forvar3840 + (1'h1)))
                    begin
                      reg3841 <= $unsigned(reg3835[(2'h3):(2'h3)]);
                      reg3842 <= $signed(reg3827);
                    end
                  if (reg3804[(2'h3):(2'h3)])
                    begin
                      reg3843 <= reg3837[(3'h5):(3'h5)];
                      reg3844 <= ((!((reg3800 ? reg3797 : (8'ha5)) ?
                              (&(8'h9e)) : forvar3837[(1'h1):(1'h1)])) ?
                          ((!reg3846) << $signed({wire3783})) : $unsigned($signed(((8'hba) ?
                              reg3841 : (8'hae)))));
                    end
                  else
                    begin
                      reg3843 <= ($signed({$signed((8'hba))}) ?
                          (~^$signed($signed(reg3844))) : $signed((reg3803[(1'h0):(1'h0)] ?
                              reg3846[(3'h7):(2'h2)] : reg3801)));
                    end
                end
            end
          if (reg3827)
            begin
              for (forvar3848 = (1'h0); (forvar3848 < (2'h2)); forvar3848 = (forvar3848 + (1'h1)))
                begin
                  if (reg3822[(4'hd):(4'h9)])
                    begin
                      reg3849 <= (-{$signed(reg3805)});
                    end
                  else
                    begin
                      reg3849 <= {$signed((8'hb2))};
                    end
                  if (reg3802[(3'h4):(2'h2)])
                    begin
                      reg3850 <= (8'ha1);
                      reg3851 <= $signed(forvar3837[(1'h1):(1'h1)]);
                      reg3852 <= ({reg3827[(3'h7):(3'h6)]} ?
                          forvar3786 : reg3829);
                    end
                  else
                    begin
                      reg3850 <= (^~((8'ha1) && (((8'h9c) > forvar3837) ?
                          reg3841 : (reg3850 ? (8'hb3) : (8'hb2)))));
                      reg3851 <= $signed(reg3813[(2'h3):(2'h2)]);
                      reg3852 <= $unsigned($unsigned($signed(forvar3834)));
                      reg3853 <= (&(8'ha8));
                    end
                end
            end
          else
            begin
              for (forvar3848 = (1'h0); (forvar3848 < (1'h1)); forvar3848 = (forvar3848 + (1'h1)))
                begin
                  for (forvar3849 = (1'h0); (forvar3849 < (2'h2)); forvar3849 = (forvar3849 + (1'h1)))
                    begin
                      reg3850 <= $unsigned(reg3802[(1'h0):(1'h0)]);
                      reg3851 <= $signed((-wire3782));
                      reg3852 <= $signed(reg3840);
                      reg3853 <= ((((reg3821 | reg3852) ^ $signed(forvar3794)) ?
                              $unsigned((~&reg3827)) : $unsigned((reg3822 ?
                                  reg3793 : (8'hba)))) ?
                          (+$unsigned($unsigned(forvar3787))) : $signed($signed(wire3784[(1'h1):(1'h0)])));
                    end
                  if (({($signed((8'ha6)) > (reg3825 & (8'hba)))} <= reg3845))
                    begin
                      reg3854 <= {$signed({(reg3835 ? reg3787 : (8'haf))})};
                    end
                  else
                    begin
                      reg3854 <= $unsigned((forvar3806[(2'h2):(1'h1)] << reg3809));
                      reg3855 <= (8'ha5);
                      reg3856 <= forvar3824;
                    end
                  for (forvar3857 = (1'h0); (forvar3857 < (1'h1)); forvar3857 = (forvar3857 + (1'h1)))
                    begin
                      reg3858 <= (($signed((^reg3831)) ?
                          {forvar3824} : $signed(reg3856)) > wire3781[(1'h1):(1'h0)]);
                      reg3859 <= reg3810;
                      reg3860 <= reg3816[(3'h5):(1'h0)];
                      reg3861 <= (|$signed((~&((8'h9e) == reg3792))));
                    end
                end
              if ({$unsigned((reg3815 < (reg3796 ~^ wire3783)))})
                begin
                  for (forvar3862 = (1'h0); (forvar3862 < (2'h2)); forvar3862 = (forvar3862 + (1'h1)))
                    begin
                      reg3863 <= $signed($signed((!$unsigned(reg3838))));
                    end
                end
              else
                begin
                  if ({{(~^(forvar3787 ? reg3821 : reg3844))}})
                    begin
                      reg3862 <= $unsigned(({(~&reg3854)} && $unsigned($signed(reg3855))));
                      reg3863 <= ({reg3849} + ({$signed(reg3807)} ?
                          (~$unsigned(forvar3834)) : $unsigned({reg3803})));
                      reg3864 <= $signed($unsigned((|(~&(8'hb8)))));
                    end
                  else
                    begin
                      reg3862 <= reg3862[(3'h5):(2'h3)];
                      reg3863 <= ($signed($signed(forvar3818[(4'hc):(2'h3)])) > (~^($unsigned(reg3788) <= (forvar3849 ?
                          forvar3786 : reg3861))));
                      reg3864 <= (8'hb5);
                    end
                  if ((8'h9c))
                    begin
                      reg3865 <= {forvar3785};
                      reg3866 <= {(~|(&reg3800[(4'h8):(3'h5)]))};
                      reg3867 <= wire3782;
                      reg3868 <= $unsigned({(8'ha4)});
                    end
                  else
                    begin
                      reg3865 <= wire3782;
                      reg3866 <= reg3823;
                    end
                  for (forvar3869 = (1'h0); (forvar3869 < (1'h1)); forvar3869 = (forvar3869 + (1'h1)))
                    begin
                      reg3870 <= reg3864[(3'h5):(2'h3)];
                      reg3871 <= reg3817;
                      reg3872 <= $signed(((&{reg3786}) ?
                          {$signed(reg3867)} : $unsigned(((8'ha6) && (8'haf)))));
                      reg3873 <= ({($signed(forvar3857) ?
                              forvar3794[(1'h1):(1'h0)] : (8'hb9))} & $unsigned({(reg3837 <<< forvar3794)}));
                    end
                  if ((forvar3824 ?
                      ((+reg3831) ^ ($unsigned((8'ha8)) ?
                          $signed((8'ha1)) : {reg3856})) : ($signed(reg3790[(3'h7):(3'h5)]) << ({reg3853} ?
                          $unsigned(reg3837) : $signed(reg3808)))))
                    begin
                      reg3874 <= ((~|($unsigned(reg3820) ?
                              $unsigned(reg3799) : $signed(reg3864))) ?
                          $signed((+(|reg3821))) : {(+((8'hae) ?
                                  reg3822 : (8'ha1)))});
                      reg3875 <= $unsigned((!reg3864));
                      reg3876 <= $unsigned($signed($unsigned({forvar3857})));
                    end
                  else
                    begin
                      reg3874 <= ((~^forvar3832[(4'hb):(4'hb)]) ?
                          {($unsigned(reg3793) >= $unsigned(reg3845))} : (&forvar3869));
                      reg3875 <= ((((~&(8'ha5)) ^~ {reg3801}) ?
                              ($signed(reg3807) >> ((8'hb9) ?
                                  reg3866 : reg3842)) : $unsigned((forvar3832 ?
                                  reg3856 : (8'hb1)))) ?
                          ($signed((reg3789 >>> (8'ha9))) + (+(forvar3862 == reg3855))) : $unsigned($signed((reg3852 ^ reg3813))));
                      reg3876 <= reg3870[(1'h1):(1'h1)];
                    end
                end
              if ({(-forvar3795[(1'h0):(1'h0)])})
                begin
                  for (forvar3877 = (1'h0); (forvar3877 < (1'h0)); forvar3877 = (forvar3877 + (1'h1)))
                    begin
                      reg3878 <= ((($signed(reg3812) ?
                          (wire3782 >> (8'ha3)) : reg3796) >= $signed({reg3851})) >= $signed(((reg3785 ?
                              forvar3832 : forvar3841) ?
                          $signed(reg3799) : $signed(reg3813))));
                      reg3879 <= (~|({$signed((8'ha0))} << {$signed(reg3861)}));
                    end
                  if ((~|$signed($unsigned($unsigned(reg3813)))))
                    begin
                      reg3880 <= $signed(wire3784[(3'h6):(1'h1)]);
                      reg3881 <= reg3791;
                      reg3882 <= ((~|$signed($unsigned((8'ha9)))) > ((((8'hb7) ?
                          reg3871 : reg3870) < ((8'hae) < reg3874)) >= ((|forvar3849) ?
                          ((8'ha8) ?
                              forvar3785 : reg3831) : (reg3825 == reg3812))));
                    end
                  else
                    begin
                      reg3880 <= (+(8'h9d));
                      reg3881 <= $unsigned(reg3850[(4'hf):(2'h2)]);
                      reg3882 <= ((^(8'hb2)) << $signed(forvar3787));
                    end
                end
              else
                begin
                  if ({forvar3840})
                    begin
                      reg3877 <= wire3783;
                    end
                  else
                    begin
                      reg3877 <= reg3789;
                    end
                  reg3878 <= (8'h9d);
                  for (forvar3879 = (1'h0); (forvar3879 < (1'h0)); forvar3879 = (forvar3879 + (1'h1)))
                    begin
                      reg3880 <= $unsigned($unsigned($unsigned((~&reg3808))));
                      reg3881 <= $signed({reg3841});
                      reg3882 <= reg3877;
                    end
                  reg3883 <= reg3845;
                end
              if (({$unsigned({reg3829})} ?
                  reg3845[(4'hb):(1'h1)] : $unsigned(reg3785)))
                begin
                  for (forvar3884 = (1'h0); (forvar3884 < (1'h0)); forvar3884 = (forvar3884 + (1'h1)))
                    begin
                      reg3885 <= (reg3863 ?
                          $unsigned(($unsigned((8'hba)) * {forvar3787})) : reg3850[(3'h4):(1'h1)]);
                      reg3886 <= ((|$signed((8'hb4))) < reg3835[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar3884 = (1'h0); (forvar3884 < (1'h0)); forvar3884 = (forvar3884 + (1'h1)))
                    begin
                      reg3885 <= {reg3829};
                    end
                  for (forvar3886 = (1'h0); (forvar3886 < (2'h3)); forvar3886 = (forvar3886 + (1'h1)))
                    begin
                      reg3887 <= reg3821;
                      reg3888 <= reg3829;
                    end
                  for (forvar3889 = (1'h0); (forvar3889 < (1'h0)); forvar3889 = (forvar3889 + (1'h1)))
                    begin
                      reg3890 <= $unsigned((forvar3836[(2'h2):(1'h1)] ?
                          reg3868 : reg3817));
                      reg3891 <= (~&$signed((+(reg3868 < reg3827))));
                      reg3892 <= $unsigned($unsigned((reg3839[(3'h5):(1'h0)] < reg3855[(3'h4):(1'h1)])));
                    end
                end
            end
        end
      else
        begin
          reg3832 <= (~$signed((~|(reg3861 < reg3888))));
          if (((($unsigned(reg3833) ?
              reg3858[(2'h3):(1'h0)] : forvar3857) << $signed((reg3799 >> reg3820))) - forvar3787))
            begin
              if (reg3861)
                begin
                  reg3833 <= $unsigned($unsigned(($signed((8'hab)) ?
                      $signed(reg3862) : $signed(reg3874))));
                  reg3834 <= {($signed((~&(8'ha3))) <<< ((8'hab) ?
                          ((8'haf) ? reg3880 : reg3788) : (&reg3867)))};
                end
              else
                begin
                  if ({($signed((~^reg3863)) ?
                          (reg3832 ?
                              {reg3842} : reg3802[(1'h0):(1'h0)]) : ($unsigned(reg3883) ?
                              (reg3823 | reg3800) : forvar3818[(3'h6):(3'h5)]))})
                    begin
                      reg3833 <= forvar3834[(4'hc):(3'h4)];
                    end
                  else
                    begin
                      reg3833 <= (~|$signed(reg3822[(1'h1):(1'h1)]));
                      reg3834 <= (reg3800[(2'h2):(2'h2)] * ({(reg3835 ?
                              reg3880 : reg3847)} > (~(8'ha8))));
                      reg3835 <= $signed($unsigned((((8'ha2) ?
                          reg3813 : reg3862) && (~reg3828))));
                    end
                  if (reg3858)
                    begin
                      reg3836 <= (~|$unsigned((-reg3867)));
                      reg3837 <= $unsigned({forvar3889});
                      reg3838 <= (reg3837 & (^~$signed(reg3812[(4'hc):(4'hb)])));
                      reg3839 <= reg3807[(4'ha):(4'ha)];
                    end
                  else
                    begin
                      reg3836 <= $unsigned(($signed((forvar3884 ?
                          reg3823 : reg3834)) > {((8'ha4) ?
                              reg3788 : reg3868)}));
                      reg3837 <= (forvar3889[(4'ha):(4'h9)] ?
                          (reg3802[(3'h5):(3'h5)] ?
                              (forvar3795[(1'h0):(1'h0)] <<< (forvar3877 ~^ reg3833)) : forvar3787) : reg3831[(4'h8):(3'h7)]);
                      reg3838 <= $unsigned((~&(&reg3786)));
                      reg3839 <= $signed((reg3843[(3'h7):(3'h5)] | $unsigned(((8'ha7) - reg3809))));
                    end
                  if ((8'hae))
                    begin
                      reg3840 <= ((~&(forvar3824[(1'h0):(1'h0)] ?
                              $signed(forvar3857) : forvar3841[(4'hc):(2'h2)])) ?
                          wire3783[(3'h5):(2'h2)] : ({((8'hae) ^~ reg3822)} ?
                              reg3849[(2'h3):(1'h0)] : ($signed(reg3861) ?
                                  $unsigned(reg3879) : reg3819[(2'h3):(1'h0)])));
                      reg3841 <= $unsigned(reg3832[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg3840 <= ((forvar3832[(2'h3):(1'h1)] & $unsigned((reg3819 ?
                              reg3868 : reg3813))) ?
                          (8'h9e) : $unsigned((~^$unsigned(reg3888))));
                      reg3841 <= $unsigned($signed(reg3825[(3'h4):(2'h2)]));
                      reg3842 <= {(8'hba)};
                      reg3843 <= $unsigned($unsigned($signed((reg3820 ?
                          forvar3836 : (8'h9d)))));
                    end
                end
              reg3844 <= $unsigned(reg3844[(2'h3):(2'h2)]);
              if ((&reg3865))
                begin
                  if (({((^reg3836) ?
                              (forvar3869 ?
                                  wire3781 : wire3784) : $signed(reg3888))} ?
                      reg3791[(3'h4):(1'h0)] : reg3845))
                    begin
                      reg3845 <= (8'h9c);
                      reg3846 <= (($signed({reg3793}) ?
                              reg3785[(3'h4):(3'h4)] : (reg3842 ?
                                  (~&reg3873) : reg3859[(2'h3):(1'h1)])) ?
                          (($signed((8'h9e)) ?
                                  (reg3853 ?
                                      reg3810 : reg3880) : $signed(reg3863)) ?
                              $unsigned(reg3858) : (forvar3818[(4'h9):(3'h4)] ?
                                  reg3798[(3'h6):(1'h1)] : (reg3803 * forvar3849))) : wire3784);
                      reg3847 <= (8'ha2);
                    end
                  else
                    begin
                      reg3845 <= (forvar3785[(4'h8):(3'h7)] ?
                          (reg3877 && $unsigned((forvar3837 == reg3822))) : ((8'hb4) ?
                              ($signed(reg3861) ?
                                  reg3858[(3'h6):(3'h5)] : (^~reg3885)) : reg3891[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  if (reg3816)
                    begin
                      reg3845 <= forvar3869[(4'h9):(4'h8)];
                      reg3846 <= ($unsigned($signed(reg3880)) & $unsigned((8'h9f)));
                    end
                  else
                    begin
                      reg3845 <= $unsigned((((wire3784 | reg3874) ?
                              $signed(reg3827) : (reg3832 ^ reg3874)) ?
                          (+forvar3836[(2'h3):(2'h3)]) : reg3891));
                      reg3846 <= reg3840;
                      reg3847 <= $unsigned(((~$signed(reg3888)) ?
                          ($signed((8'hae)) || $unsigned((8'hae))) : $unsigned($signed(reg3785))));
                    end
                  if (reg3872)
                    begin
                      reg3848 <= $signed((~$unsigned((^reg3822))));
                      reg3849 <= reg3829;
                      reg3850 <= reg3835;
                      reg3851 <= reg3791;
                    end
                  else
                    begin
                      reg3848 <= (8'hb8);
                      reg3849 <= {(8'ha6)};
                      reg3850 <= forvar3824;
                    end
                  for (forvar3852 = (1'h0); (forvar3852 < (2'h2)); forvar3852 = (forvar3852 + (1'h1)))
                    begin
                      reg3853 <= ($unsigned($unsigned(reg3833)) ?
                          ($unsigned({forvar3879}) ?
                              $unsigned(forvar3848[(4'h9):(1'h1)]) : $unsigned({reg3881})) : reg3842[(3'h4):(2'h2)]);
                      reg3854 <= (|(|reg3809));
                      reg3855 <= reg3863[(1'h0):(1'h0)];
                      reg3856 <= (forvar3862[(3'h6):(1'h0)] + (reg3871 <= reg3866[(3'h5):(3'h4)]));
                    end
                end
            end
          else
            begin
              for (forvar3833 = (1'h0); (forvar3833 < (1'h1)); forvar3833 = (forvar3833 + (1'h1)))
                begin
                  if ($unsigned((($unsigned(forvar3857) >> reg3813[(1'h1):(1'h0)]) ?
                      reg3851[(3'h7):(3'h7)] : reg3883[(4'h8):(1'h0)])))
                    begin
                      reg3834 <= (reg3798[(3'h5):(3'h5)] ? reg3847 : reg3820);
                      reg3835 <= $signed(((reg3891 ?
                          $unsigned(reg3817) : (&reg3844)) && {forvar3834[(4'ha):(2'h2)]}));
                    end
                  else
                    begin
                      reg3834 <= reg3885;
                      reg3835 <= {reg3811};
                      reg3836 <= reg3814;
                    end
                  reg3837 <= reg3849;
                  for (forvar3838 = (1'h0); (forvar3838 < (2'h3)); forvar3838 = (forvar3838 + (1'h1)))
                    begin
                      reg3839 <= {$signed($signed($signed(reg3808)))};
                      reg3840 <= (reg3876 == $unsigned(reg3833));
                      reg3841 <= (forvar3787[(4'h8):(3'h5)] ~^ $signed($unsigned(reg3870)));
                      reg3842 <= reg3845;
                    end
                end
            end
          if (((forvar3884 ?
              $signed($signed(reg3871)) : forvar3824[(4'h8):(4'h8)]) ^~ $signed($signed(reg3827[(4'h8):(3'h4)]))))
            begin
              if ({$unsigned(reg3787[(3'h5):(3'h4)])})
                begin
                  reg3857 <= ((~|reg3805[(3'h4):(2'h2)]) - $signed($signed(reg3851[(3'h6):(1'h0)])));
                  if ({reg3821})
                    begin
                      reg3858 <= reg3827;
                    end
                  else
                    begin
                      reg3858 <= (forvar3877[(5'h10):(3'h5)] > {wire3783[(2'h3):(2'h3)]});
                      reg3859 <= reg3828[(3'h4):(1'h0)];
                    end
                end
              else
                begin
                  if ((reg3802[(4'ha):(1'h0)] * (+(~$unsigned(reg3851)))))
                    begin
                      reg3857 <= ((^{reg3853[(2'h3):(1'h0)]}) ?
                          $unsigned({(reg3790 || wire3782)}) : (&(!forvar3862)));
                      reg3858 <= reg3886;
                      reg3859 <= $signed((~reg3808[(1'h0):(1'h0)]));
                      reg3860 <= (8'hb6);
                    end
                  else
                    begin
                      reg3857 <= (({{(8'ha3)}} ?
                          {$unsigned(reg3814)} : (^$unsigned(reg3826))) ~^ (($unsigned(forvar3806) ?
                              $unsigned(forvar3869) : $signed(reg3796)) ?
                          {((8'hb6) ?
                                  reg3823 : reg3847)} : $unsigned($unsigned(reg3865))));
                      reg3858 <= ((-reg3860) * (|forvar3852));
                    end
                  for (forvar3861 = (1'h0); (forvar3861 < (2'h2)); forvar3861 = (forvar3861 + (1'h1)))
                    begin
                      reg3862 <= reg3891[(1'h1):(1'h0)];
                      reg3863 <= ((($unsigned(reg3868) ?
                                  (reg3851 ~^ wire3783) : reg3838[(3'h4):(2'h3)]) ?
                              (|wire3782) : (8'ha9)) ?
                          $signed($signed($unsigned(reg3885))) : {($unsigned(reg3802) >= (!reg3862))});
                      reg3864 <= reg3822;
                    end
                  for (forvar3865 = (1'h0); (forvar3865 < (2'h3)); forvar3865 = (forvar3865 + (1'h1)))
                    begin
                      reg3866 <= {$unsigned(((forvar3886 > reg3832) ?
                              (reg3878 ?
                                  reg3885 : forvar3832) : reg3788[(3'h6):(1'h1)]))};
                      reg3867 <= (^~(~|((reg3850 ^~ reg3861) ?
                          (reg3841 ?
                              forvar3879 : reg3851) : $signed(reg3882))));
                      reg3868 <= $unsigned((+reg3873));
                      reg3869 <= ($unsigned($unsigned((reg3853 ^~ reg3850))) ?
                          $signed(reg3827) : $signed($unsigned((8'hb1))));
                    end
                end
              for (forvar3870 = (1'h0); (forvar3870 < (2'h3)); forvar3870 = (forvar3870 + (1'h1)))
                begin
                  for (forvar3871 = (1'h0); (forvar3871 < (2'h3)); forvar3871 = (forvar3871 + (1'h1)))
                    begin
                      reg3872 <= (!reg3812[(2'h3):(1'h0)]);
                      reg3873 <= (8'ha1);
                    end
                  if (reg3793)
                    begin
                      reg3874 <= (-({$unsigned(forvar3836)} ?
                          (~^(reg3885 ?
                              forvar3794 : reg3822)) : $signed((reg3797 == forvar3879))));
                      reg3875 <= {(($unsigned(reg3825) ?
                                  (reg3888 ?
                                      (8'h9f) : forvar3836) : (^~reg3885)) ?
                              $signed(reg3796) : (~|$signed(forvar3879)))};
                    end
                  else
                    begin
                      reg3874 <= reg3883;
                      reg3875 <= $signed({(|$unsigned(reg3890))});
                      reg3876 <= ({reg3872[(2'h2):(1'h0)]} >= reg3869);
                    end
                end
            end
          else
            begin
              for (forvar3857 = (1'h0); (forvar3857 < (2'h3)); forvar3857 = (forvar3857 + (1'h1)))
                begin
                  for (forvar3858 = (1'h0); (forvar3858 < (2'h3)); forvar3858 = (forvar3858 + (1'h1)))
                    begin
                      reg3859 <= {reg3802};
                    end
                  reg3860 <= reg3856[(3'h4):(2'h3)];
                  if ((~|reg3838))
                    begin
                      reg3861 <= ((((!reg3833) ^ (~^reg3834)) << (^~(reg3841 ?
                          forvar3879 : reg3787))) | reg3811);
                    end
                  else
                    begin
                      reg3861 <= (reg3847[(2'h2):(1'h0)] != reg3843);
                    end
                  reg3862 <= $unsigned((-reg3877));
                end
            end
        end
      for (forvar3893 = (1'h0); (forvar3893 < (1'h1)); forvar3893 = (forvar3893 + (1'h1)))
        begin
          for (forvar3894 = (1'h0); (forvar3894 < (1'h1)); forvar3894 = (forvar3894 + (1'h1)))
            begin
              if ((8'hb2))
                begin
                  if (reg3877)
                    begin
                      reg3895 <= forvar3849[(1'h0):(1'h0)];
                      reg3896 <= ($unsigned($unsigned(reg3864)) ?
                          $signed($unsigned($unsigned(reg3848))) : {forvar3862});
                    end
                  else
                    begin
                      reg3895 <= $signed(reg3830[(2'h2):(1'h0)]);
                      reg3896 <= reg3813[(2'h3):(1'h0)];
                    end
                  if (reg3869)
                    begin
                      reg3897 <= ($signed(reg3891) == (((reg3863 ~^ forvar3848) ?
                          {forvar3877} : wire3782[(1'h0):(1'h0)]) && (reg3843[(2'h3):(2'h2)] ?
                          $unsigned(reg3847) : reg3881)));
                    end
                  else
                    begin
                      reg3897 <= (((~&$signed(forvar3840)) ?
                          reg3827 : $signed(reg3800)) ~^ (^~(!((8'ha4) ~^ reg3881))));
                      reg3898 <= ((reg3844[(2'h2):(2'h2)] < (~^reg3854[(4'ha):(4'h9)])) ?
                          forvar3841 : (($unsigned(reg3809) >>> $signed(forvar3818)) ?
                              (~(8'h9d)) : $signed($signed(reg3812))));
                      reg3899 <= (((^(forvar3849 ? forvar3894 : reg3887)) ?
                              (+(^~reg3843)) : reg3804) ?
                          (((+(8'hb4)) - $unsigned(reg3832)) ?
                              $unsigned((reg3887 >>> (8'hb9))) : reg3812) : {(~^$unsigned(reg3843))});
                      reg3900 <= $unsigned(reg3854);
                    end
                  for (forvar3901 = (1'h0); (forvar3901 < (1'h0)); forvar3901 = (forvar3901 + (1'h1)))
                    begin
                      reg3902 <= reg3786;
                      reg3903 <= reg3797;
                      reg3904 <= ((~&reg3899) <<< $signed($unsigned((~|reg3872))));
                      reg3905 <= $signed(forvar3862[(2'h3):(1'h0)]);
                    end
                  reg3906 <= $signed(reg3865);
                end
              else
                begin
                  reg3895 <= $signed($signed($signed((forvar3877 << reg3813))));
                end
            end
          if ({$unsigned((^~reg3791[(4'h9):(3'h4)]))})
            begin
              if (forvar3857[(3'h5):(3'h4)])
                begin
                  reg3907 <= reg3815;
                  if (reg3836)
                    begin
                      reg3908 <= ({(^~$signed(forvar3886))} >> (($unsigned(reg3882) && reg3886[(3'h6):(3'h5)]) ?
                          reg3873 : (8'hb8)));
                      reg3909 <= reg3836[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg3908 <= reg3902[(2'h2):(1'h0)];
                      reg3909 <= $signed($signed(reg3862[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar3907 = (1'h0); (forvar3907 < (1'h0)); forvar3907 = (forvar3907 + (1'h1)))
                    begin
                      reg3908 <= {((8'ha1) > reg3870)};
                      reg3909 <= {reg3803};
                      reg3910 <= forvar3795[(2'h3):(2'h2)];
                    end
                end
            end
          else
            begin
              reg3907 <= reg3804;
              for (forvar3908 = (1'h0); (forvar3908 < (2'h3)); forvar3908 = (forvar3908 + (1'h1)))
                begin
                  if ($unsigned((((reg3873 && (8'haa)) ?
                      {reg3859} : (reg3831 ?
                          reg3789 : forvar3787)) & $signed(wire3781[(2'h3):(1'h1)]))))
                    begin
                      reg3909 <= (reg3846[(2'h3):(2'h3)] ?
                          (~^$signed(((8'hac) ?
                              reg3850 : reg3899))) : (reg3825[(1'h0):(1'h0)] ?
                              $signed(reg3879[(4'ha):(3'h5)]) : reg3892[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg3909 <= $unsigned((!((forvar3832 ?
                          reg3853 : reg3881) - (forvar3834 & forvar3901))));
                      reg3910 <= reg3908[(4'hb):(1'h0)];
                      reg3911 <= $unsigned(({(forvar3852 >>> (8'haf))} - $unsigned((~|(8'h9f)))));
                      reg3912 <= $signed(reg3831);
                    end
                  reg3913 <= ((~&reg3904[(1'h0):(1'h0)]) < $unsigned(($unsigned(reg3840) >>> $unsigned((8'hb9)))));
                  reg3914 <= ($signed($signed((forvar3785 ?
                      reg3865 : forvar3795))) || (^~forvar3865[(1'h1):(1'h1)]));
                  for (forvar3915 = (1'h0); (forvar3915 < (2'h2)); forvar3915 = (forvar3915 + (1'h1)))
                    begin
                      reg3916 <= (~&$unsigned(($signed((8'hb3)) * $signed(reg3825))));
                      reg3917 <= reg3850[(4'hb):(3'h4)];
                    end
                end
              reg3918 <= ({((reg3917 << forvar3879) ?
                          reg3877[(2'h2):(2'h2)] : reg3859)} ?
                  $signed($signed($unsigned(forvar3787))) : (forvar3862 == $unsigned($unsigned((8'ha1)))));
              for (forvar3919 = (1'h0); (forvar3919 < (2'h3)); forvar3919 = (forvar3919 + (1'h1)))
                begin
                  for (forvar3920 = (1'h0); (forvar3920 < (1'h0)); forvar3920 = (forvar3920 + (1'h1)))
                    begin
                      reg3921 <= $unsigned(reg3803);
                      reg3922 <= reg3861[(1'h1):(1'h0)];
                      reg3923 <= $unsigned(reg3911[(4'hd):(3'h4)]);
                      reg3924 <= (({$unsigned(forvar3840)} ?
                          $signed(reg3910[(1'h0):(1'h0)]) : (reg3837 ?
                              (reg3810 ?
                                  reg3800 : forvar3806) : (^reg3888))) >> reg3916);
                    end
                  if ((~&$signed(((reg3828 ? reg3917 : reg3923) ?
                      (&reg3874) : (reg3866 ? (8'haa) : reg3912)))))
                    begin
                      reg3925 <= (reg3872 <<< $signed(((forvar3871 & reg3910) ?
                          $signed(reg3864) : reg3843[(1'h1):(1'h0)])));
                      reg3926 <= $signed($unsigned(forvar3818[(4'ha):(1'h1)]));
                    end
                  else
                    begin
                      reg3925 <= $signed(reg3909[(1'h1):(1'h0)]);
                      reg3926 <= reg3878[(2'h3):(1'h1)];
                      reg3927 <= {reg3863};
                    end
                  for (forvar3928 = (1'h0); (forvar3928 < (1'h0)); forvar3928 = (forvar3928 + (1'h1)))
                    begin
                      reg3929 <= (~|reg3786[(3'h6):(3'h5)]);
                      reg3930 <= (8'haf);
                    end
                end
            end
        end
    end
  module3931 modinst4155 (.clk(clk), .wire3932(wire3781), .wire3933(forvar3869), .y(wire4154), .wire3934(reg3906), .wire3935(reg3825));
  always
    @(posedge clk) begin
      for (forvar4156 = (1'h0); (forvar4156 < (2'h2)); forvar4156 = (forvar4156 + (1'h1)))
        begin
          for (forvar4157 = (1'h0); (forvar4157 < (2'h3)); forvar4157 = (forvar4157 + (1'h1)))
            begin
              reg4158 <= {(reg3877 <= $signed(forvar3838[(3'h4):(3'h4)]))};
              for (forvar4159 = (1'h0); (forvar4159 < (1'h0)); forvar4159 = (forvar4159 + (1'h1)))
                begin
                  if (($unsigned(forvar3832) >= ($signed(reg3803) ?
                      $unsigned((reg3874 > reg3895)) : (reg3828 & (~|reg3918)))))
                    begin
                      reg4160 <= reg3876;
                      reg4161 <= $signed((+$unsigned((reg3858 * reg3909))));
                    end
                  else
                    begin
                      reg4160 <= (((forvar3928 && reg3883) < (|(reg3828 - reg3834))) ?
                          ((reg3860[(3'h7):(3'h5)] ?
                              (reg3923 < (8'hb0)) : {forvar3893}) >= ((forvar3908 * reg3883) ?
                              (reg3844 <<< reg3865) : ((8'hba) ?
                                  (8'hb7) : reg3791))) : ($signed({(8'hba)}) <<< (((8'h9f) | reg3927) - (forvar3861 <= reg3847))));
                    end
                end
            end
        end
      for (forvar4162 = (1'h0); (forvar4162 < (2'h2)); forvar4162 = (forvar4162 + (1'h1)))
        begin
          for (forvar4163 = (1'h0); (forvar4163 < (1'h0)); forvar4163 = (forvar4163 + (1'h1)))
            begin
              for (forvar4164 = (1'h0); (forvar4164 < (2'h2)); forvar4164 = (forvar4164 + (1'h1)))
                begin
                  for (forvar4165 = (1'h0); (forvar4165 < (2'h2)); forvar4165 = (forvar4165 + (1'h1)))
                    begin
                      reg4166 <= reg3876[(3'h6):(3'h4)];
                      reg4167 <= (wire3784 >> forvar3928[(1'h0):(1'h0)]);
                    end
                  for (forvar4168 = (1'h0); (forvar4168 < (1'h0)); forvar4168 = (forvar4168 + (1'h1)))
                    begin
                      reg4169 <= (8'hac);
                      reg4170 <= {($unsigned((~|forvar3833)) ?
                              reg3905[(4'hd):(4'hc)] : forvar3785)};
                    end
                  for (forvar4171 = (1'h0); (forvar4171 < (2'h2)); forvar4171 = (forvar4171 + (1'h1)))
                    begin
                      reg4172 <= $unsigned(forvar3908);
                      reg4173 <= forvar3907[(4'he):(4'ha)];
                    end
                  for (forvar4174 = (1'h0); (forvar4174 < (1'h0)); forvar4174 = (forvar4174 + (1'h1)))
                    begin
                      reg4175 <= $unsigned($signed($signed((~&reg3899))));
                      reg4176 <= {$unsigned(reg3912)};
                      reg4177 <= $unsigned({(+$signed(reg3899))});
                      reg4178 <= $unsigned(reg3830);
                    end
                end
              for (forvar4179 = (1'h0); (forvar4179 < (2'h2)); forvar4179 = (forvar4179 + (1'h1)))
                begin
                  for (forvar4180 = (1'h0); (forvar4180 < (1'h0)); forvar4180 = (forvar4180 + (1'h1)))
                    begin
                      reg4181 <= reg3788[(1'h1):(1'h1)];
                      reg4182 <= reg3825[(2'h3):(2'h3)];
                      reg4183 <= reg3816;
                    end
                  if (((!$signed((reg3826 ?
                      reg3887 : forvar3862))) - $signed($unsigned((forvar3861 ?
                      reg3839 : reg3905)))))
                    begin
                      reg4184 <= ($unsigned(((reg3917 ?
                          reg3872 : reg3890) ^~ (-forvar3824))) >= ((~|(8'hab)) >>> (reg3860[(3'h5):(1'h0)] <= (~|reg3804))));
                    end
                  else
                    begin
                      reg4184 <= (reg3902 != $unsigned((reg3797 ?
                          {reg3855} : (forvar3838 ? reg3827 : reg3926))));
                      reg4185 <= ((((8'hb4) - forvar4180) ?
                          forvar3869[(2'h3):(1'h1)] : reg3883) << $signed((reg3853[(3'h7):(1'h1)] ?
                          ((8'ha9) || reg3872) : $unsigned(forvar3861))));
                      reg4186 <= reg3814[(4'h8):(3'h5)];
                    end
                  for (forvar4187 = (1'h0); (forvar4187 < (2'h2)); forvar4187 = (forvar4187 + (1'h1)))
                    begin
                      reg4188 <= (forvar3915 < $signed(($signed(reg3878) >> $unsigned(reg3830))));
                      reg4189 <= {(~^((forvar4164 ?
                              reg3825 : forvar3818) < $signed((8'hb4))))};
                      reg4190 <= forvar3852;
                    end
                  reg4191 <= $signed(((~|reg3883[(4'ha):(4'ha)]) * ((reg4169 ?
                          (8'ha8) : reg3905) ?
                      (reg3871 ? (8'ha2) : forvar4164) : (reg3798 ?
                          reg3927 : forvar3834))));
                end
              if (forvar4174[(3'h6):(2'h3)])
                begin
                  for (forvar4192 = (1'h0); (forvar4192 < (1'h1)); forvar4192 = (forvar4192 + (1'h1)))
                    begin
                      reg4193 <= forvar4171[(1'h1):(1'h1)];
                      reg4194 <= reg3872[(3'h4):(2'h3)];
                      reg4195 <= ((((~|(8'ha5)) ?
                                  forvar3928[(1'h0):(1'h0)] : (reg3885 | (8'ha6))) ?
                              $unsigned(reg4190[(1'h1):(1'h1)]) : forvar3919[(2'h3):(1'h1)]) ?
                          (~|$unsigned(reg3912[(1'h0):(1'h0)])) : ((reg3851 | $unsigned(reg3873)) << {{forvar3838}}));
                      reg4196 <= ($unsigned(reg3879) ?
                          ($unsigned((reg3812 >>> wire4154)) ^ (!reg3846)) : reg3828[(4'hd):(3'h6)]);
                    end
                  reg4197 <= reg3847;
                  if ((reg3822[(4'h8):(4'h8)] ?
                      $unsigned($unsigned((8'h9e))) : reg3866))
                    begin
                      reg4198 <= $unsigned($unsigned(reg3849[(1'h0):(1'h0)]));
                      reg4199 <= (^~wire3783[(1'h0):(1'h0)]);
                      reg4200 <= $unsigned(forvar3865[(1'h0):(1'h0)]);
                      reg4201 <= {(~reg3848[(3'h5):(2'h3)])};
                    end
                  else
                    begin
                      reg4198 <= $unsigned((|(|{(8'hb9)})));
                      reg4199 <= $unsigned((($signed(reg3907) ?
                              {forvar4165} : forvar3869[(3'h4):(1'h1)]) ?
                          $signed((^forvar4168)) : ($unsigned(reg3921) <<< (^forvar3915))));
                    end
                  if (forvar3886)
                    begin
                      reg4202 <= ($signed((~&$unsigned(reg4196))) << $signed(({forvar3852} ?
                          $unsigned(reg3791) : forvar4163)));
                    end
                  else
                    begin
                      reg4202 <= reg3822[(1'h0):(1'h0)];
                      reg4203 <= (!$unsigned((~(~^reg3909))));
                      reg4204 <= (+(+($unsigned((8'hb5)) ^~ (reg4200 ?
                          reg3882 : reg3897))));
                      reg4205 <= (!reg3819[(2'h3):(2'h3)]);
                    end
                end
              else
                begin
                  for (forvar4192 = (1'h0); (forvar4192 < (1'h1)); forvar4192 = (forvar4192 + (1'h1)))
                    begin
                      reg4193 <= $signed(reg3923);
                    end
                  for (forvar4194 = (1'h0); (forvar4194 < (2'h2)); forvar4194 = (forvar4194 + (1'h1)))
                    begin
                      reg4195 <= reg3786[(2'h3):(1'h1)];
                      reg4196 <= $unsigned($unsigned($signed($signed(reg3854))));
                      reg4197 <= (reg3838[(3'h7):(3'h6)] >>> {$signed((reg3871 ?
                              reg3877 : reg3797))});
                      reg4198 <= ($signed((reg4186 <<< reg3856[(3'h5):(3'h4)])) & {$unsigned($signed(reg4201))});
                    end
                  reg4199 <= $unsigned(forvar3852);
                end
              if ((reg3858[(3'h6):(3'h6)] ?
                  reg3923[(4'ha):(3'h5)] : (!($signed(reg3807) || reg4170))))
                begin
                  for (forvar4206 = (1'h0); (forvar4206 < (1'h0)); forvar4206 = (forvar4206 + (1'h1)))
                    begin
                      reg4207 <= ($signed({reg3913[(2'h3):(1'h1)]}) > reg3859[(1'h1):(1'h1)]);
                      reg4208 <= $signed((^~$unsigned(reg3839)));
                      reg4209 <= (^(+reg3913[(3'h7):(1'h0)]));
                    end
                  for (forvar4210 = (1'h0); (forvar4210 < (1'h1)); forvar4210 = (forvar4210 + (1'h1)))
                    begin
                      reg4211 <= reg3877[(1'h1):(1'h0)];
                      reg4212 <= $unsigned((reg3887 ?
                          (reg4177[(3'h6):(1'h0)] && (reg4182 + forvar3857)) : forvar4159));
                    end
                  reg4213 <= ($unsigned({$unsigned(reg4182)}) ?
                      $signed(((forvar3865 ? forvar3907 : forvar3837) ?
                          $signed(reg3918) : reg3921[(2'h2):(2'h2)])) : {$unsigned(reg3832)});
                  if (((~&($signed(forvar4168) * (~forvar4157))) ?
                      $unsigned($signed(reg3837)) : reg4211[(1'h1):(1'h0)]))
                    begin
                      reg4214 <= forvar3786[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg4214 <= (((~|reg4209) != (~^reg3821)) < $unsigned(($signed(forvar3908) >= (-reg3886))));
                      reg4215 <= $unsigned({$unsigned($signed(reg4183))});
                      reg4216 <= $unsigned((forvar4210[(2'h2):(1'h0)] ?
                          $unsigned($unsigned((8'ha7))) : {$unsigned(reg3808)}));
                      reg4217 <= (8'hac);
                    end
                end
              else
                begin
                  reg4206 <= $unsigned($signed(((forvar4179 ?
                          reg3815 : forvar4206) ?
                      (reg3851 ^~ reg3892) : $signed(reg4197))));
                  reg4207 <= $unsigned(forvar3836);
                  for (forvar4208 = (1'h0); (forvar4208 < (1'h0)); forvar4208 = (forvar4208 + (1'h1)))
                    begin
                      reg4209 <= ($unsigned(forvar3838[(4'h8):(1'h0)]) ?
                          forvar3901 : reg4197[(3'h4):(2'h2)]);
                      reg4210 <= (forvar3838[(4'ha):(3'h4)] * (reg3815 ?
                          $signed($signed(reg3876)) : reg3926[(1'h0):(1'h0)]));
                    end
                  for (forvar4211 = (1'h0); (forvar4211 < (1'h1)); forvar4211 = (forvar4211 + (1'h1)))
                    begin
                      reg4212 <= (^~(&reg3792));
                    end
                end
            end
          for (forvar4218 = (1'h0); (forvar4218 < (1'h1)); forvar4218 = (forvar4218 + (1'h1)))
            begin
              if (((+((reg3853 != reg3907) ?
                  {reg4191} : $unsigned(reg3846))) < ({$unsigned(reg4206)} * (reg3908[(4'h9):(3'h5)] ^~ $unsigned(reg4170)))))
                begin
                  for (forvar4219 = (1'h0); (forvar4219 < (2'h3)); forvar4219 = (forvar4219 + (1'h1)))
                    begin
                      reg4220 <= (reg4200 >>> ($unsigned((^reg3847)) ?
                          reg4161 : forvar4180));
                      reg4221 <= $signed(reg3845);
                      reg4222 <= {reg3882[(1'h0):(1'h0)]};
                      reg4223 <= $unsigned((forvar3836[(1'h1):(1'h0)] ?
                          reg4185 : $unsigned((|reg4203))));
                    end
                end
              else
                begin
                  if (((!($signed(reg4181) ?
                      $unsigned((8'had)) : forvar4219[(3'h4):(1'h1)])) >> $unsigned({(reg3789 ?
                          reg3899 : reg4160)})))
                    begin
                      reg4219 <= reg4212[(1'h0):(1'h0)];
                      reg4220 <= reg3905;
                    end
                  else
                    begin
                      reg4219 <= reg4188;
                      reg4220 <= $signed((reg3826[(3'h6):(1'h1)] > $signed((reg3809 <= reg3869))));
                      reg4221 <= (reg3853 ?
                          (reg4216[(3'h4):(1'h1)] ?
                              {(reg4216 >= reg3790)} : $unsigned($unsigned(reg4207))) : forvar3843);
                      reg4222 <= $signed(($signed((reg3850 + reg3845)) << (wire3784[(3'h4):(1'h1)] ?
                          (~&reg3862) : (reg4223 * forvar4187))));
                    end
                  for (forvar4223 = (1'h0); (forvar4223 < (1'h1)); forvar4223 = (forvar4223 + (1'h1)))
                    begin
                      reg4224 <= (!{reg4207[(4'hc):(4'hb)]});
                      reg4225 <= reg3793[(3'h5):(3'h5)];
                    end
                  if (((!($signed(reg3861) * $unsigned(reg4221))) >> ($signed($unsigned(reg3913)) ?
                      $unsigned({reg4169}) : forvar3871[(1'h1):(1'h0)])))
                    begin
                      reg4226 <= {($signed(forvar3871[(2'h2):(1'h1)]) == ($signed(reg4184) ?
                              (|reg3886) : (forvar4223 ? reg3837 : reg3815)))};
                      reg4227 <= ((^~(reg3819[(1'h0):(1'h0)] ~^ $signed(reg3929))) ?
                          (-((forvar3928 >>> forvar3795) ?
                              (reg4206 ?
                                  forvar3832 : forvar4218) : wire4154[(1'h0):(1'h0)])) : reg3880);
                      reg4228 <= reg3796[(1'h0):(1'h0)];
                      reg4229 <= (-(((+reg3827) ? $signed(reg3878) : (8'hb5)) ?
                          ($unsigned(reg4211) ?
                              (reg4216 << reg4197) : (reg4167 ?
                                  reg3831 : reg3905)) : forvar3834[(4'hb):(4'h8)]));
                    end
                  else
                    begin
                      reg4226 <= $signed((~|$unsigned(forvar3889)));
                    end
                end
              reg4230 <= $unsigned(forvar4210[(1'h1):(1'h1)]);
              reg4231 <= $signed(($signed(forvar4187) ?
                  reg4177[(4'h9):(2'h2)] : forvar4206));
            end
          for (forvar4232 = (1'h0); (forvar4232 < (1'h0)); forvar4232 = (forvar4232 + (1'h1)))
            begin
              for (forvar4233 = (1'h0); (forvar4233 < (2'h3)); forvar4233 = (forvar4233 + (1'h1)))
                begin
                  reg4234 <= $signed($signed((reg3921 + $unsigned(reg4188))));
                end
              if ($signed(((reg3924[(3'h7):(1'h1)] ^~ $signed(reg4204)) ^ $signed(reg3814))))
                begin
                  if ((!(~|(^~(reg4158 ? forvar3787 : reg4170)))))
                    begin
                      reg4235 <= $unsigned((8'hb9));
                    end
                  else
                    begin
                      reg4235 <= (($unsigned((^reg4212)) ?
                          ($signed(forvar4192) ?
                              $signed(reg3888) : $signed(reg4223)) : reg3792[(3'h7):(1'h1)]) ^~ $signed(((|forvar3857) <<< (reg3838 ^ reg3842))));
                      reg4236 <= reg3800;
                      reg4237 <= (reg4221[(4'h8):(1'h0)] * reg3788);
                      reg4238 <= reg3821;
                    end
                  for (forvar4239 = (1'h0); (forvar4239 < (1'h0)); forvar4239 = (forvar4239 + (1'h1)))
                    begin
                      reg4240 <= $unsigned(({reg4207[(4'hb):(4'h9)]} <= {$unsigned(reg3929)}));
                    end
                end
              else
                begin
                  for (forvar4235 = (1'h0); (forvar4235 < (2'h3)); forvar4235 = (forvar4235 + (1'h1)))
                    begin
                      reg4236 <= (forvar3837 << $unsigned($unsigned({reg4211})));
                    end
                  if ($unsigned(forvar3879[(1'h1):(1'h1)]))
                    begin
                      reg4237 <= (reg3815 || ($signed($unsigned(reg3844)) ?
                          {$unsigned(reg3927)} : forvar3871[(1'h1):(1'h0)]));
                      reg4238 <= ($signed(reg4170[(3'h7):(3'h7)]) ?
                          (~^(8'hb4)) : ($signed((-forvar4187)) ?
                              $unsigned({forvar3833}) : $signed((reg3822 ?
                                  forvar3806 : reg4221))));
                      reg4239 <= forvar3870[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg4237 <= forvar4164;
                      reg4238 <= $signed(reg4197[(4'h8):(3'h7)]);
                    end
                end
            end
          if ($unsigned({reg3880[(3'h5):(3'h4)]}))
            begin
              for (forvar4241 = (1'h0); (forvar4241 < (1'h1)); forvar4241 = (forvar4241 + (1'h1)))
                begin
                  for (forvar4242 = (1'h0); (forvar4242 < (1'h0)); forvar4242 = (forvar4242 + (1'h1)))
                    begin
                      reg4243 <= $signed((^~(((8'h9d) & reg3848) != $signed(reg4199))));
                    end
                  reg4244 <= $unsigned(reg3925[(1'h1):(1'h1)]);
                  for (forvar4245 = (1'h0); (forvar4245 < (1'h0)); forvar4245 = (forvar4245 + (1'h1)))
                    begin
                      reg4246 <= reg3871[(1'h1):(1'h1)];
                      reg4247 <= {(reg4208[(4'ha):(1'h1)] ?
                              ((-forvar3865) ?
                                  reg4217[(3'h5):(3'h4)] : (forvar3893 ?
                                      wire3784 : (8'ha7))) : reg3895[(2'h2):(1'h1)])};
                    end
                  for (forvar4248 = (1'h0); (forvar4248 < (2'h2)); forvar4248 = (forvar4248 + (1'h1)))
                    begin
                      reg4249 <= (-(|{{wire3783}}));
                    end
                end
              if (reg3914[(4'h9):(3'h7)])
                begin
                  if ($unsigned(forvar4241))
                    begin
                      reg4250 <= (reg3816 ~^ ((-(8'hb1)) ?
                          reg4181 : ($unsigned(reg3823) ?
                              {reg4230} : $unsigned(forvar4164))));
                      reg4251 <= reg4243[(1'h0):(1'h0)];
                      reg4252 <= ({{((8'ha6) ~^ reg3834)}} + ($signed(reg3903[(1'h1):(1'h0)]) ^~ $unsigned($unsigned((8'haa)))));
                    end
                  else
                    begin
                      reg4250 <= reg4219;
                      reg4251 <= reg3830;
                    end
                  for (forvar4253 = (1'h0); (forvar4253 < (1'h1)); forvar4253 = (forvar4253 + (1'h1)))
                    begin
                      reg4254 <= ($unsigned($signed({reg4213})) ?
                          reg4223[(2'h2):(2'h2)] : {$unsigned({reg3839})});
                      reg4255 <= $unsigned($unsigned(($signed(reg3930) + $signed((8'hb4)))));
                      reg4256 <= reg3786;
                    end
                  reg4257 <= (((+{forvar4233}) ?
                          (+(reg3876 ?
                              (8'hba) : (8'hb0))) : $unsigned((~reg4189))) ?
                      $unsigned($signed((reg3790 & reg3812))) : $signed(reg4234[(4'h9):(3'h5)]));
                end
              else
                begin
                  for (forvar4250 = (1'h0); (forvar4250 < (1'h0)); forvar4250 = (forvar4250 + (1'h1)))
                    begin
                      reg4251 <= reg4229;
                      reg4252 <= forvar4210[(2'h3):(2'h2)];
                    end
                  for (forvar4253 = (1'h0); (forvar4253 < (1'h0)); forvar4253 = (forvar4253 + (1'h1)))
                    begin
                      reg4254 <= reg4198;
                      reg4255 <= {(~^(((8'ha0) ^~ reg3858) ?
                              (forvar3894 ? reg3797 : reg4223) : (-reg3887)))};
                      reg4256 <= ((reg3811 ?
                              $signed((+forvar4245)) : $unsigned(forvar3901[(3'h6):(3'h5)])) ?
                          (((8'ha1) << $unsigned(reg3791)) ?
                              (!(forvar4168 >>> reg3842)) : $signed($unsigned(reg4256))) : $unsigned(forvar3838[(4'hc):(3'h4)]));
                    end
                  if (((-($unsigned((8'hb9)) ?
                      $signed(reg3792) : (~|forvar3824))) || $unsigned($unsigned(reg3804[(1'h0):(1'h0)]))))
                    begin
                      reg4257 <= forvar4159;
                      reg4258 <= ((reg3911 ?
                              {(reg3885 || (8'hb6))} : ({(8'h9d)} ?
                                  (reg3848 || forvar4233) : ((8'hb1) ?
                                      reg4224 : forvar4242))) ?
                          reg3869 : $signed((~((8'haf) | reg4191))));
                      reg4259 <= (~&(!$signed($unsigned(reg4184))));
                    end
                  else
                    begin
                      reg4257 <= forvar4206[(2'h3):(1'h0)];
                      reg4258 <= reg3786[(2'h3):(1'h1)];
                      reg4259 <= {((reg3925 * (-forvar3870)) ?
                              $signed($signed(reg3823)) : reg4207[(4'h8):(3'h6)])};
                      reg4260 <= $unsigned($signed((forvar4248 ?
                          $unsigned(reg3929) : $unsigned(forvar3848))));
                    end
                end
              reg4261 <= forvar4156[(4'h9):(4'h9)];
              for (forvar4262 = (1'h0); (forvar4262 < (2'h3)); forvar4262 = (forvar4262 + (1'h1)))
                begin
                  reg4263 <= forvar4218[(4'h8):(3'h7)];
                end
            end
          else
            begin
              for (forvar4241 = (1'h0); (forvar4241 < (2'h2)); forvar4241 = (forvar4241 + (1'h1)))
                begin
                  reg4242 <= $unsigned(reg3857[(1'h1):(1'h0)]);
                end
            end
        end
      for (forvar4264 = (1'h0); (forvar4264 < (2'h3)); forvar4264 = (forvar4264 + (1'h1)))
        begin
          for (forvar4265 = (1'h0); (forvar4265 < (2'h3)); forvar4265 = (forvar4265 + (1'h1)))
            begin
              for (forvar4266 = (1'h0); (forvar4266 < (1'h1)); forvar4266 = (forvar4266 + (1'h1)))
                begin
                  if ($unsigned((($signed(reg4259) ^~ (forvar4248 + reg4183)) ?
                      {(|reg3786)} : $signed($signed(forvar4157)))))
                    begin
                      reg4267 <= (^~$unsigned(reg3867));
                    end
                  else
                    begin
                      reg4267 <= $signed({$signed($signed((8'hb7)))});
                      reg4268 <= forvar3858[(3'h5):(1'h1)];
                      reg4269 <= reg3861[(1'h0):(1'h0)];
                    end
                  if ($signed($unsigned(reg4216[(4'hd):(3'h5)])))
                    begin
                      reg4270 <= ((reg3826 + reg4234) ?
                          $unsigned(reg4158[(1'h0):(1'h0)]) : $unsigned(reg4197));
                    end
                  else
                    begin
                      reg4270 <= (((((8'haf) >= forvar3908) ?
                              $signed(reg3808) : $signed(forvar3838)) >> $unsigned((|reg4190))) ?
                          {forvar4253} : $signed((reg4259 ?
                              (~^reg3792) : (reg4167 == reg3810))));
                      reg4271 <= {($unsigned(forvar3884[(4'h9):(3'h6)]) ?
                              ((~&reg3831) + $signed(reg4182)) : reg4203[(3'h4):(2'h3)])};
                      reg4272 <= $unsigned($signed($unsigned(reg3819[(1'h0):(1'h0)])));
                      reg4273 <= ((reg3908[(4'h8):(1'h0)] ?
                              ((reg3924 ?
                                  reg3926 : (8'hb4)) == (8'hb5)) : reg3844[(4'h8):(1'h0)]) ?
                          {forvar4187[(1'h1):(1'h1)]} : (forvar4192[(2'h2):(2'h2)] ?
                              {{reg4226}} : reg4226));
                    end
                  for (forvar4274 = (1'h0); (forvar4274 < (2'h3)); forvar4274 = (forvar4274 + (1'h1)))
                    begin
                      reg4275 <= forvar4239[(3'h4):(2'h2)];
                      reg4276 <= $unsigned($signed($unsigned(((8'hac) ?
                          reg3868 : reg4197))));
                    end
                  for (forvar4277 = (1'h0); (forvar4277 < (1'h1)); forvar4277 = (forvar4277 + (1'h1)))
                    begin
                      reg4278 <= $signed(reg3842);
                    end
                end
              for (forvar4279 = (1'h0); (forvar4279 < (1'h0)); forvar4279 = (forvar4279 + (1'h1)))
                begin
                  if (reg3892[(3'h5):(1'h1)])
                    begin
                      reg4280 <= $unsigned($signed(forvar3848[(1'h0):(1'h0)]));
                      reg4281 <= ($unsigned(reg3875) >>> $unsigned(reg4255));
                    end
                  else
                    begin
                      reg4280 <= {{(&(~&reg3902))}};
                    end
                end
              if ((~($unsigned(reg4189) && reg4183[(4'h8):(2'h2)])))
                begin
                  reg4282 <= (8'hb5);
                  for (forvar4283 = (1'h0); (forvar4283 < (1'h1)); forvar4283 = (forvar4283 + (1'h1)))
                    begin
                      reg4284 <= $signed($signed($unsigned((forvar3806 ?
                          reg3897 : reg3888))));
                      reg4285 <= (+$unsigned(($signed((8'haa)) >> {reg3787})));
                      reg4286 <= ($unsigned($signed((|forvar4279))) ?
                          reg3895[(4'h9):(3'h6)] : reg4200);
                    end
                  if ($signed($signed(reg3864[(3'h4):(3'h4)])))
                    begin
                      reg4287 <= reg3845;
                    end
                  else
                    begin
                      reg4287 <= $signed({(-forvar3785)});
                      reg4288 <= {{($unsigned(reg4196) >= (|reg3925))}};
                      reg4289 <= $unsigned(((8'hb9) ^ (~|$unsigned(reg4191))));
                      reg4290 <= reg4222[(3'h4):(1'h0)];
                    end
                  for (forvar4291 = (1'h0); (forvar4291 < (1'h1)); forvar4291 = (forvar4291 + (1'h1)))
                    begin
                      reg4292 <= ($unsigned($unsigned((reg4209 + reg4194))) | forvar3886[(2'h2):(1'h1)]);
                      reg4293 <= forvar3889;
                    end
                end
              else
                begin
                  reg4282 <= (wire4154 ?
                      (((forvar4274 ?
                          reg4238 : reg4221) <= $unsigned((8'hae))) * ((forvar4253 ?
                          reg4166 : reg3886) != reg4276)) : (^reg4201[(2'h2):(1'h1)]));
                  for (forvar4283 = (1'h0); (forvar4283 < (1'h1)); forvar4283 = (forvar4283 + (1'h1)))
                    begin
                      reg4284 <= $signed($signed($unsigned((reg3880 ?
                          reg4214 : reg3849))));
                      reg4285 <= $signed((forvar4194[(4'h8):(2'h3)] >>> forvar3857));
                      reg4286 <= {$signed(($signed(reg3807) < $signed(reg4270)))};
                    end
                  if ((-$signed($unsigned((+(8'hae))))))
                    begin
                      reg4287 <= reg3912;
                    end
                  else
                    begin
                      reg4287 <= forvar4262[(1'h0):(1'h0)];
                    end
                end
              for (forvar4294 = (1'h0); (forvar4294 < (1'h1)); forvar4294 = (forvar4294 + (1'h1)))
                begin
                  reg4295 <= reg3916;
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar4296 = (1'h0); (forvar4296 < (2'h2)); forvar4296 = (forvar4296 + (1'h1)))
        begin
          if ((reg3891 ? reg4292 : $signed($unsigned(reg4240))))
            begin
              for (forvar4297 = (1'h0); (forvar4297 < (1'h0)); forvar4297 = (forvar4297 + (1'h1)))
                begin
                  for (forvar4298 = (1'h0); (forvar4298 < (1'h0)); forvar4298 = (forvar4298 + (1'h1)))
                    begin
                      reg4299 <= ((reg3831 >= {(~|reg3836)}) ?
                          forvar4297 : ((8'ha5) ?
                              (reg4254 ?
                                  {reg4292} : (8'hab)) : {((8'h9f) >> forvar3806)}));
                    end
                  for (forvar4300 = (1'h0); (forvar4300 < (1'h0)); forvar4300 = (forvar4300 + (1'h1)))
                    begin
                      reg4301 <= $signed((!(reg4292 ?
                          (+reg4189) : $signed((8'hb4)))));
                    end
                  if (reg4278)
                    begin
                      reg4302 <= reg3862;
                      reg4303 <= (((~(reg4220 == reg4278)) ?
                          reg4284 : (((8'hb9) <= reg3831) >> $unsigned((8'ha3)))) >>> reg4158);
                      reg4304 <= (((reg3888 | (reg3792 ?
                          reg4175 : forvar3852)) >= ((&(8'hb4)) ?
                          $unsigned(forvar3901) : (~(8'hb3)))) & (($unsigned(reg4239) != $unsigned(reg3854)) << ($signed(reg4207) > $signed(reg4254))));
                    end
                  else
                    begin
                      reg4302 <= ((($unsigned(forvar4164) ?
                                  (^~forvar3907) : $unsigned(reg3863)) ?
                              $signed(((8'hb5) ?
                                  forvar3886 : (8'h9c))) : $unsigned((-reg3796))) ?
                          forvar3824[(2'h3):(1'h1)] : (((forvar4279 <<< reg3926) <= reg3832) ?
                              (reg4215 > (reg3905 ^~ forvar4157)) : ((+reg3810) <= $signed(reg3834))));
                      reg4303 <= ($signed(forvar4279[(2'h3):(1'h1)]) ~^ reg4254[(4'hf):(3'h4)]);
                      reg4304 <= (|(~^(|reg4235[(1'h1):(1'h0)])));
                      reg4305 <= forvar4164[(1'h1):(1'h0)];
                    end
                end
            end
          else
            begin
              reg4297 <= reg4182[(4'h8):(3'h4)];
              for (forvar4298 = (1'h0); (forvar4298 < (1'h1)); forvar4298 = (forvar4298 + (1'h1)))
                begin
                  for (forvar4299 = (1'h0); (forvar4299 < (1'h0)); forvar4299 = (forvar4299 + (1'h1)))
                    begin
                      reg4300 <= ({$signed($unsigned(reg4203))} ?
                          reg4288 : (+((reg3896 ?
                              reg4260 : reg3927) ^ reg3835)));
                      reg4301 <= forvar4241;
                      reg4302 <= ((reg4191[(1'h0):(1'h0)] == $unsigned((~forvar4171))) ?
                          reg4234[(3'h4):(3'h4)] : reg3929[(1'h1):(1'h0)]);
                    end
                  if ((forvar3884 ?
                      reg3798 : $unsigned((reg3805[(1'h1):(1'h0)] ?
                          $signed(reg4217) : $signed(forvar4223)))))
                    begin
                      reg4303 <= reg4214[(2'h3):(2'h2)];
                      reg4304 <= (&{{((8'h9c) ? reg3930 : forvar3877)}});
                      reg4305 <= ({reg3899[(4'hc):(2'h3)]} << reg4263);
                    end
                  else
                    begin
                      reg4303 <= (^$signed({reg4285}));
                      reg4304 <= reg3851;
                      reg4305 <= $signed(($signed((reg4239 == reg4182)) ?
                          $unsigned((~|forvar4242)) : $signed($signed(reg3801))));
                      reg4306 <= (forvar3840[(3'h5):(2'h2)] == ({reg3852} <= $signed({forvar4233})));
                    end
                end
              if (($unsigned(reg4209) > (forvar3865 ?
                  reg4254[(1'h0):(1'h0)] : reg4237)))
                begin
                  reg4307 <= reg4183[(2'h2):(1'h1)];
                  reg4308 <= forvar3919[(3'h5):(2'h3)];
                  if (({($signed(reg3852) + ((8'h9d) ?
                          forvar3848 : (8'ha3)))} || (({(8'h9e)} <= (8'hb9)) >>> reg3847[(1'h0):(1'h0)])))
                    begin
                      reg4309 <= ($signed({{reg4197}}) ?
                          reg3848[(3'h4):(1'h1)] : (^(((8'ha9) << reg4194) < $signed((8'hab)))));
                      reg4310 <= (forvar4283[(1'h1):(1'h0)] && {(&forvar3833)});
                      reg4311 <= reg4210[(4'ha):(2'h2)];
                    end
                  else
                    begin
                      reg4309 <= reg4297[(1'h0):(1'h0)];
                      reg4310 <= ($unsigned($signed($unsigned(reg4231))) ?
                          $unsigned($unsigned({reg3807})) : reg4235[(1'h0):(1'h0)]);
                    end
                  reg4312 <= ($unsigned($signed(reg3905)) >>> reg3823[(3'h6):(3'h5)]);
                end
              else
                begin
                  if (((((reg4308 ?
                      reg4243 : reg3926) >= {reg4221}) << forvar4208) ^~ (^~(reg4242 ?
                      (reg3861 ? reg3867 : reg3852) : $unsigned(reg3908)))))
                    begin
                      reg4307 <= $signed({reg3857});
                      reg4308 <= $signed(forvar4235);
                      reg4309 <= (((reg3856 ? (+reg3896) : forvar4264) ?
                          $signed($signed(reg4237)) : ((|reg3848) ?
                              reg4204 : (reg3812 ?
                                  forvar3786 : reg4280))) && reg4276);
                    end
                  else
                    begin
                      reg4307 <= $signed($signed(reg3876[(3'h5):(1'h1)]));
                      reg4308 <= (reg4259[(2'h3):(1'h0)] & $signed(((reg3819 ?
                              reg3790 : forvar3834) ?
                          $unsigned(reg3883) : reg3837[(2'h2):(2'h2)])));
                    end
                  if (($unsigned(((8'ha7) << $signed((8'haf)))) ^~ ($signed($signed((8'hb1))) ?
                      reg3879 : (+$signed(reg4234)))))
                    begin
                      reg4310 <= forvar4165[(1'h0):(1'h0)];
                      reg4311 <= (({reg4230} ^ (8'hb3)) < $signed(($signed(forvar4180) != (~&reg4247))));
                      reg4312 <= {reg4222};
                    end
                  else
                    begin
                      reg4310 <= reg4198[(3'h4):(2'h2)];
                      reg4311 <= ($signed((reg3852[(1'h1):(1'h1)] ^ $signed((8'hb7)))) ?
                          (~^(((8'hae) >>> reg4255) ?
                              {(8'hab)} : $unsigned(reg4244))) : (-$signed($signed(reg4175))));
                      reg4312 <= {forvar4245};
                      reg4313 <= reg4184;
                    end
                  for (forvar4314 = (1'h0); (forvar4314 < (2'h3)); forvar4314 = (forvar4314 + (1'h1)))
                    begin
                      reg4315 <= $signed(forvar4233[(2'h3):(1'h1)]);
                      reg4316 <= $unsigned(reg3819);
                    end
                end
            end
        end
      for (forvar4317 = (1'h0); (forvar4317 < (1'h0)); forvar4317 = (forvar4317 + (1'h1)))
        begin
          if ($signed($signed(((^(8'hab)) ?
              reg4306[(2'h3):(1'h1)] : (forvar4168 != reg4199)))))
            begin
              for (forvar4318 = (1'h0); (forvar4318 < (2'h3)); forvar4318 = (forvar4318 + (1'h1)))
                begin
                  reg4319 <= (reg4209[(1'h1):(1'h0)] >= ((|{forvar4219}) ?
                      reg4185[(1'h1):(1'h1)] : (reg3854[(3'h4):(1'h0)] ?
                          ((8'ha0) ?
                              reg4299 : reg4300) : (reg4206 || reg4235))));
                  for (forvar4320 = (1'h0); (forvar4320 < (2'h2)); forvar4320 = (forvar4320 + (1'h1)))
                    begin
                      reg4321 <= (8'ha6);
                      reg4322 <= {$signed((reg3808 == ((8'ha8) ?
                              reg4186 : (8'ha6))))};
                      reg4323 <= $unsigned(reg4200);
                      reg4324 <= {$unsigned(((forvar4156 > reg4290) ?
                              $unsigned(reg4207) : $signed((8'hab))))};
                    end
                  reg4325 <= (-(^~reg3872));
                  for (forvar4326 = (1'h0); (forvar4326 < (1'h1)); forvar4326 = (forvar4326 + (1'h1)))
                    begin
                      reg4327 <= $unsigned((^~(-$signed((8'ha1)))));
                      reg4328 <= ((|$unsigned($unsigned(reg3925))) ?
                          ({(forvar3928 ? reg3896 : (8'hb6))} ?
                              ((~|reg3929) > (reg3903 ?
                                  reg4196 : forvar4156)) : (reg4231 ?
                                  {reg4290} : reg4229)) : ({$signed(forvar4223)} - ({reg4250} + (forvar3879 < reg4194))));
                    end
                end
            end
          else
            begin
              for (forvar4318 = (1'h0); (forvar4318 < (2'h3)); forvar4318 = (forvar4318 + (1'h1)))
                begin
                  if (($unsigned((8'hb7)) >= (forvar3785 > (&reg4177[(1'h0):(1'h0)]))))
                    begin
                      reg4319 <= reg3883[(2'h2):(1'h1)];
                      reg4320 <= reg4236;
                      reg4321 <= ((&reg4243[(2'h2):(2'h2)]) || $unsigned($unsigned(reg3841)));
                      reg4322 <= (forvar3865[(1'h1):(1'h1)] - (((reg3909 << (8'hb7)) ?
                              (-forvar4168) : (~forvar4192)) ?
                          {(reg3848 ?
                                  reg3870 : reg4227)} : $signed($signed(forvar4218))));
                    end
                  else
                    begin
                      reg4319 <= (forvar4223 ?
                          $signed({$signed(reg4182)}) : $unsigned((!reg3845[(4'hb):(1'h0)])));
                      reg4320 <= (^$unsigned(((!reg4208) & (reg4185 - reg3871))));
                    end
                  reg4323 <= $signed((~($signed(reg4286) + forvar3907[(4'hf):(2'h2)])));
                end
              reg4324 <= ($unsigned($unsigned({reg3927})) == reg3800[(1'h0):(1'h0)]);
            end
          reg4329 <= (+(+$unsigned($unsigned(reg3916))));
        end
      for (forvar4330 = (1'h0); (forvar4330 < (1'h1)); forvar4330 = (forvar4330 + (1'h1)))
        begin
          for (forvar4331 = (1'h0); (forvar4331 < (1'h0)); forvar4331 = (forvar4331 + (1'h1)))
            begin
              if ($signed($signed((&(forvar3824 && reg4323)))))
                begin
                  reg4332 <= {((^~(~forvar4208)) && (reg4309[(1'h0):(1'h0)] ?
                          (reg3831 >> reg4225) : (reg3800 ?
                              reg3922 : reg4205)))};
                  for (forvar4333 = (1'h0); (forvar4333 < (2'h2)); forvar4333 = (forvar4333 + (1'h1)))
                    begin
                      reg4334 <= (-reg3927);
                      reg4335 <= $signed($signed((^~(8'hb2))));
                      reg4336 <= $signed((($unsigned(reg3822) ?
                              (^~reg3891) : (forvar3919 ? reg4214 : (8'hba))) ?
                          $unsigned($unsigned(forvar4165)) : (-(reg4186 ?
                              reg3879 : reg3865))));
                    end
                  for (forvar4337 = (1'h0); (forvar4337 < (1'h1)); forvar4337 = (forvar4337 + (1'h1)))
                    begin
                      reg4338 <= reg3927;
                      reg4339 <= (!reg4254);
                      reg4340 <= $signed({reg3820});
                      reg4341 <= $signed(reg3918);
                    end
                  if (($unsigned({forvar4296}) != ($unsigned((forvar4331 ?
                      reg3921 : reg4235)) <<< reg3791[(2'h3):(2'h2)])))
                    begin
                      reg4342 <= forvar4245;
                      reg4343 <= ((~^(reg4256 ?
                          $signed(reg4280) : $unsigned(forvar4274))) ~^ reg3885);
                      reg4344 <= $unsigned(($unsigned($unsigned(forvar3889)) >= reg4263));
                      reg4345 <= (^reg3913);
                    end
                  else
                    begin
                      reg4342 <= (((reg3888[(2'h2):(1'h1)] ?
                              (forvar3858 ?
                                  reg4315 : forvar4333) : (reg3842 | reg4204)) ?
                          (+$signed(reg3904)) : $signed(forvar4265[(1'h1):(1'h0)])) << ($signed($unsigned(forvar4210)) == ((reg3811 >= reg3850) != (~^forvar3886))));
                      reg4343 <= {($unsigned(reg4186) & (~^$signed(reg4286)))};
                      reg4344 <= reg3803;
                      reg4345 <= {(({reg4292} || reg3822[(4'hd):(4'h8)]) | reg3812[(4'h9):(4'h8)])};
                    end
                end
              else
                begin
                  if ((reg4228 ?
                      {((&reg3807) ?
                              (~|(8'h9f)) : (reg3929 - reg4261))} : (^$signed(reg3790[(1'h1):(1'h0)]))))
                    begin
                      reg4332 <= (!$unsigned(reg4210[(3'h5):(2'h2)]));
                    end
                  else
                    begin
                      reg4332 <= (8'ha0);
                    end
                  if ((reg4212 ? reg3854[(4'h9):(2'h2)] : reg4278))
                    begin
                      reg4333 <= forvar4235;
                      reg4334 <= reg4268;
                    end
                  else
                    begin
                      reg4333 <= $unsigned($unsigned(((&reg4161) ?
                          (reg3841 ? (8'hb3) : forvar4162) : reg3848)));
                      reg4334 <= (reg3831 - reg3853[(1'h1):(1'h0)]);
                      reg4335 <= $signed({reg4332[(3'h4):(3'h4)]});
                      reg4336 <= {reg4191[(4'hb):(4'ha)]};
                    end
                  if (((~^$unsigned(reg4300)) ?
                      reg3842 : {$signed((~|reg4205))}))
                    begin
                      reg4337 <= $unsigned($signed($signed((reg3786 >>> reg3897))));
                      reg4338 <= reg3838[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg4337 <= ($signed((reg4210[(4'hc):(3'h7)] ?
                          (forvar4219 <<< reg4160) : $signed((8'ha9)))) ~^ (&(~^$unsigned(reg4276))));
                      reg4338 <= {$unsigned((|(forvar4320 >> forvar4250)))};
                    end
                end
            end
          if ({{(~&reg4193[(1'h1):(1'h0)])}})
            begin
              for (forvar4346 = (1'h0); (forvar4346 < (1'h1)); forvar4346 = (forvar4346 + (1'h1)))
                begin
                  if (((((forvar4179 <= (8'hb6)) ?
                          $unsigned((8'hb0)) : $signed(reg4324)) >>> (reg3850 << (~&forvar4210))) ?
                      (~($unsigned(reg3817) > ((8'h9e) ?
                          reg3853 : reg4189))) : forvar3840[(1'h0):(1'h0)]))
                    begin
                      reg4347 <= $unsigned((((reg3796 < reg3796) ?
                          (+reg4210) : (^forvar4346)) > reg3785));
                      reg4348 <= reg3860;
                      reg4349 <= $unsigned((reg4268 ?
                          $signed($unsigned(reg3918)) : (!$signed(reg4269))));
                    end
                  else
                    begin
                      reg4347 <= reg3866;
                      reg4348 <= reg4275[(2'h2):(1'h0)];
                      reg4349 <= {$signed($signed($signed(reg3926)))};
                      reg4350 <= forvar4245[(3'h4):(1'h0)];
                    end
                  if ((reg3807[(2'h2):(1'h1)] ~^ forvar4162[(3'h7):(3'h6)]))
                    begin
                      reg4351 <= reg3838[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg4351 <= ($signed(($unsigned(reg4226) && (reg4334 > forvar4171))) ?
                          reg4234 : ((-{reg3826}) ?
                              $signed((forvar4314 + (8'ha2))) : ((~^reg3789) ?
                                  (|(8'hb1)) : reg4243[(4'h8):(1'h0)])));
                    end
                  for (forvar4352 = (1'h0); (forvar4352 < (1'h0)); forvar4352 = (forvar4352 + (1'h1)))
                    begin
                      reg4353 <= forvar3886;
                      reg4354 <= reg4216;
                      reg4355 <= ((~|forvar4266[(4'h8):(1'h1)]) ?
                          forvar3908 : reg4257[(2'h3):(2'h2)]);
                      reg4356 <= ($unsigned($unsigned($unsigned(reg3891))) >> (^~$signed((reg3918 & reg4227))));
                    end
                end
            end
          else
            begin
              if ($unsigned($signed(($signed((8'hb0)) ?
                  (~^reg4356) : $signed(reg4282)))))
                begin
                  for (forvar4346 = (1'h0); (forvar4346 < (2'h3)); forvar4346 = (forvar4346 + (1'h1)))
                    begin
                      reg4347 <= ((reg4276[(1'h0):(1'h0)] ?
                              ((reg3785 > reg4195) - forvar4279[(4'h8):(3'h5)]) : ((reg4176 ?
                                      reg4293 : (8'haf)) ?
                                  $unsigned(reg3881) : reg4205)) ?
                          (+reg3902) : (^~reg3849[(5'h10):(3'h6)]));
                    end
                  for (forvar4348 = (1'h0); (forvar4348 < (1'h1)); forvar4348 = (forvar4348 + (1'h1)))
                    begin
                      reg4349 <= $signed(forvar4219[(3'h4):(1'h1)]);
                      reg4350 <= {reg3843};
                    end
                  for (forvar4351 = (1'h0); (forvar4351 < (1'h0)); forvar4351 = (forvar4351 + (1'h1)))
                    begin
                      reg4352 <= ((((reg4348 ? forvar4233 : (8'ha3)) ?
                                  forvar3843 : (!reg4252)) ?
                              forvar4235[(1'h1):(1'h0)] : (8'ha9)) ?
                          $unsigned({forvar4298[(2'h3):(1'h0)]}) : $signed(($signed(reg4186) ?
                              (reg3930 != forvar4262) : reg4325[(3'h6):(3'h6)])));
                      reg4353 <= $signed(reg3853);
                      reg4354 <= reg4250;
                    end
                  if (reg3923[(3'h6):(3'h6)])
                    begin
                      reg4355 <= reg4238;
                    end
                  else
                    begin
                      reg4355 <= reg4286[(1'h1):(1'h0)];
                      reg4356 <= forvar3832;
                      reg4357 <= (~|$signed({forvar4297}));
                      reg4358 <= reg3906[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar4346 = (1'h0); (forvar4346 < (2'h3)); forvar4346 = (forvar4346 + (1'h1)))
                    begin
                      reg4347 <= $signed(($unsigned($unsigned(reg4244)) > $signed($signed(reg3836))));
                      reg4348 <= reg4258;
                      reg4349 <= (-$signed((~|(-reg4308))));
                      reg4350 <= reg3851;
                    end
                end
              reg4359 <= $signed(((!reg3817[(4'hc):(3'h6)]) ?
                  reg4284 : reg3867));
            end
          for (forvar4360 = (1'h0); (forvar4360 < (2'h2)); forvar4360 = (forvar4360 + (1'h1)))
            begin
              if (forvar4219[(3'h7):(3'h5)])
                begin
                  for (forvar4361 = (1'h0); (forvar4361 < (2'h3)); forvar4361 = (forvar4361 + (1'h1)))
                    begin
                      reg4362 <= (8'ha5);
                    end
                  for (forvar4363 = (1'h0); (forvar4363 < (1'h0)); forvar4363 = (forvar4363 + (1'h1)))
                    begin
                      reg4364 <= reg4282;
                      reg4365 <= forvar3871;
                    end
                  for (forvar4366 = (1'h0); (forvar4366 < (1'h1)); forvar4366 = (forvar4366 + (1'h1)))
                    begin
                      reg4367 <= {$unsigned({$signed(reg4271)})};
                      reg4368 <= ({(-$signed(reg4348))} * $signed((|$unsigned(forvar4326))));
                      reg4369 <= reg4334[(3'h4):(2'h3)];
                      reg4370 <= $signed(reg4182[(2'h2):(1'h0)]);
                    end
                  for (forvar4371 = (1'h0); (forvar4371 < (2'h2)); forvar4371 = (forvar4371 + (1'h1)))
                    begin
                      reg4372 <= {(forvar3858 >> forvar4294[(3'h6):(3'h4)])};
                    end
                end
              else
                begin
                  for (forvar4361 = (1'h0); (forvar4361 < (2'h3)); forvar4361 = (forvar4361 + (1'h1)))
                    begin
                      reg4362 <= (forvar3862[(4'hb):(4'hb)] ?
                          reg4261 : (^{$unsigned((8'hba))}));
                      reg4363 <= reg4254[(4'he):(4'ha)];
                      reg4364 <= {$signed(forvar4371[(4'h8):(2'h3)])};
                      reg4365 <= $unsigned((~reg3812));
                    end
                  if ((!(!($unsigned(forvar3785) <= (forvar4211 ?
                      forvar4250 : reg3924)))))
                    begin
                      reg4366 <= (forvar4168[(1'h1):(1'h1)] >= forvar4233[(4'hb):(3'h4)]);
                      reg4367 <= reg4351[(2'h2):(2'h2)];
                      reg4368 <= reg4213[(4'h9):(3'h4)];
                    end
                  else
                    begin
                      reg4366 <= ((|$signed((reg4247 * reg3908))) ?
                          ((^~((8'ha4) >= reg4323)) && forvar4371) : (reg4367[(4'h8):(1'h1)] ?
                              (~|$signed(reg4172)) : $unsigned($unsigned(reg3871))));
                      reg4367 <= (8'ha0);
                      reg4368 <= {($unsigned($unsigned(reg4282)) ?
                              (reg4227[(1'h0):(1'h0)] ?
                                  {reg4292} : ((8'hb7) + reg4242)) : ({reg3841} < (reg3908 ?
                                  reg4343 : forvar4241)))};
                      reg4369 <= forvar4283;
                    end
                  reg4370 <= forvar4168;
                  if ({reg4329[(1'h0):(1'h0)]})
                    begin
                      reg4371 <= ((~^reg4186[(2'h2):(1'h1)]) >>> $signed(($unsigned((8'h9d)) ?
                          (reg4249 ? reg3839 : reg3793) : (&forvar4291))));
                      reg4372 <= $unsigned((8'hab));
                    end
                  else
                    begin
                      reg4371 <= $unsigned((^reg4176));
                    end
                end
              for (forvar4373 = (1'h0); (forvar4373 < (1'h1)); forvar4373 = (forvar4373 + (1'h1)))
                begin
                  for (forvar4374 = (1'h0); (forvar4374 < (2'h2)); forvar4374 = (forvar4374 + (1'h1)))
                    begin
                      reg4375 <= ((^$unsigned(reg4365[(3'h6):(3'h4)])) || (((reg4206 ?
                          forvar4242 : reg4319) > $unsigned((8'had))) && reg4160));
                      reg4376 <= forvar3785;
                      reg4377 <= {$unsigned($signed((reg3827 ?
                              reg4303 : reg4345)))};
                      reg4378 <= (&(+$signed((~|reg3857))));
                    end
                  reg4379 <= reg3800[(4'hb):(3'h4)];
                  for (forvar4380 = (1'h0); (forvar4380 < (2'h3)); forvar4380 = (forvar4380 + (1'h1)))
                    begin
                      reg4381 <= (~|forvar3849);
                    end
                  for (forvar4382 = (1'h0); (forvar4382 < (2'h3)); forvar4382 = (forvar4382 + (1'h1)))
                    begin
                      reg4383 <= $signed(($unsigned((forvar4331 <= reg3895)) ?
                          (reg4281[(1'h1):(1'h1)] ?
                              (reg3864 * (8'ha7)) : $unsigned(reg3908)) : $signed(forvar4179[(1'h0):(1'h0)])));
                    end
                end
              if (reg3808[(4'ha):(2'h3)])
                begin
                  reg4384 <= forvar3806[(3'h4):(2'h3)];
                  if (reg4254[(2'h2):(2'h2)])
                    begin
                      reg4385 <= {($signed(((8'hb2) - reg4190)) ?
                              (((8'haa) ? forvar3787 : forvar4208) ?
                                  reg3908[(2'h2):(1'h0)] : (~|forvar4331)) : reg4205)};
                    end
                  else
                    begin
                      reg4385 <= (reg4161 * ({reg4356} + $unsigned((reg4275 ^~ forvar3920))));
                      reg4386 <= $unsigned(reg4286);
                    end
                  if ((^~(^~(-{reg4189}))))
                    begin
                      reg4387 <= $unsigned((({reg4228} ?
                          (^~(8'hab)) : $signed(reg3807)) << (^~(forvar3865 && reg3793))));
                      reg4388 <= forvar4211;
                      reg4389 <= reg4347;
                    end
                  else
                    begin
                      reg4387 <= (8'haa);
                      reg4388 <= $unsigned(((8'haf) ?
                          reg4307 : (reg3875 ?
                              reg4200[(1'h0):(1'h0)] : $unsigned(forvar4374))));
                      reg4389 <= $unsigned({$signed((8'hb6))});
                    end
                end
              else
                begin
                  for (forvar4384 = (1'h0); (forvar4384 < (1'h1)); forvar4384 = (forvar4384 + (1'h1)))
                    begin
                      reg4385 <= forvar3852[(1'h0):(1'h0)];
                      reg4386 <= reg4328[(4'hd):(4'hb)];
                      reg4387 <= $unsigned($signed($unsigned(reg3895[(1'h0):(1'h0)])));
                      reg4388 <= ($signed(reg3903[(1'h1):(1'h1)]) << $signed(($signed(reg4166) * forvar4180[(2'h2):(2'h2)])));
                    end
                  reg4389 <= $signed((&({(8'hab)} <= $signed((8'ha5)))));
                  if ($unsigned(($unsigned((reg4313 ^ reg4320)) > {(!forvar4235)})))
                    begin
                      reg4390 <= ($unsigned({$signed((8'hab))}) + (!{(forvar4366 ?
                              (8'hb8) : (8'ha3))}));
                      reg4391 <= $unsigned($unsigned(reg4250));
                      reg4392 <= ((~(forvar4330 ?
                              (^~reg4320) : reg4235[(1'h0):(1'h0)])) ?
                          ($signed(reg4276[(1'h0):(1'h0)]) ?
                              {$unsigned(reg4225)} : $unsigned($unsigned(forvar3871))) : $unsigned({$signed(reg4210)}));
                      reg4393 <= $signed((forvar3787[(3'h6):(1'h1)] + reg4344[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg4390 <= (forvar4348 != $signed(($unsigned(reg3821) ?
                          $signed(reg4249) : forvar3849[(3'h5):(2'h2)])));
                      reg4391 <= $signed(({$signed(reg4259)} ?
                          ($signed(forvar4235) <= (-reg3830)) : $unsigned(((8'h9d) - forvar4239))));
                      reg4392 <= reg4243;
                    end
                end
              if ($signed((-$unsigned(forvar4317[(2'h3):(1'h0)]))))
                begin
                  for (forvar4394 = (1'h0); (forvar4394 < (2'h3)); forvar4394 = (forvar4394 + (1'h1)))
                    begin
                      reg4395 <= (reg3882[(1'h0):(1'h0)] >> {$unsigned((|reg4252))});
                      reg4396 <= (reg4282 ? forvar4296 : reg4269);
                      reg4397 <= $unsigned($unsigned(forvar4235));
                      reg4398 <= reg4222[(3'h4):(2'h2)];
                    end
                  for (forvar4399 = (1'h0); (forvar4399 < (2'h2)); forvar4399 = (forvar4399 + (1'h1)))
                    begin
                      reg4400 <= $signed($signed($unsigned(reg4365)));
                      reg4401 <= $signed(((forvar4194[(4'hb):(4'h9)] && $signed(reg3912)) && (8'hb4)));
                      reg4402 <= ($unsigned(forvar3920) ?
                          {reg4191[(3'h4):(2'h3)]} : ($unsigned(forvar4331) ?
                              ({reg3791} >= forvar4314[(1'h0):(1'h0)]) : (~|$unsigned(reg4333))));
                    end
                  if ((reg4234 ^~ (reg3840[(3'h4):(1'h1)] <<< ((-forvar4235) | forvar4346))))
                    begin
                      reg4403 <= reg4311[(4'h8):(3'h6)];
                      reg4404 <= ($unsigned($unsigned((~|reg4288))) >> forvar4211);
                    end
                  else
                    begin
                      reg4403 <= ($unsigned(reg4392) ?
                          {reg3914[(1'h0):(1'h0)]} : reg4400);
                    end
                end
              else
                begin
                  if (reg3799)
                    begin
                      reg4394 <= (({reg4286} < reg4242) << $unsigned((^{reg3854})));
                      reg4395 <= (reg3886 ? reg3887 : reg4392[(1'h0):(1'h0)]);
                      reg4396 <= {reg4282};
                      reg4397 <= {$signed(((reg3817 ?
                              reg4227 : (8'h9f)) >>> (~reg3859)))};
                    end
                  else
                    begin
                      reg4394 <= $unsigned(((8'hb5) ?
                          $unsigned((forvar3785 << reg4257)) : (^(~^reg4325))));
                    end
                  reg4398 <= {(reg4172[(3'h4):(2'h3)] && $signed(((8'ha0) > reg4214)))};
                  if ({{$unsigned(reg3908)}})
                    begin
                      reg4399 <= reg3900;
                      reg4400 <= reg4301;
                    end
                  else
                    begin
                      reg4399 <= $signed((forvar4232 + (~|(reg3835 ?
                          reg4379 : reg3877))));
                    end
                  for (forvar4401 = (1'h0); (forvar4401 < (2'h3)); forvar4401 = (forvar4401 + (1'h1)))
                    begin
                      reg4402 <= reg4222;
                      reg4403 <= ($unsigned(reg4392) ?
                          $signed(($unsigned(forvar4384) >>> ((8'h9d) << reg4207))) : (8'hba));
                      reg4404 <= forvar4218;
                    end
                end
            end
          for (forvar4405 = (1'h0); (forvar4405 < (2'h3)); forvar4405 = (forvar4405 + (1'h1)))
            begin
              if (reg4251[(1'h0):(1'h0)])
                begin
                  for (forvar4406 = (1'h0); (forvar4406 < (1'h1)); forvar4406 = (forvar4406 + (1'h1)))
                    begin
                      reg4407 <= (&reg4297);
                      reg4408 <= $signed((((+forvar3893) > ((8'hab) <<< forvar4165)) ?
                          (|(reg4311 ?
                              reg4336 : reg4188)) : forvar4192[(1'h0):(1'h0)]));
                      reg4409 <= (-$unsigned({{reg3829}}));
                    end
                  if (wire3781)
                    begin
                      reg4410 <= $unsigned(reg4175);
                      reg4411 <= (forvar3862 ?
                          reg4354[(1'h0):(1'h0)] : ($signed($signed(reg4214)) == $unsigned(reg4349)));
                    end
                  else
                    begin
                      reg4410 <= reg3814[(1'h0):(1'h0)];
                      reg4411 <= (+(reg4392 - (~&{reg3880})));
                      reg4412 <= (+($signed($signed((8'hb1))) & (reg4371 ?
                          forvar4250 : (reg4394 ? reg4269 : (8'h9e)))));
                    end
                end
              else
                begin
                  for (forvar4406 = (1'h0); (forvar4406 < (1'h0)); forvar4406 = (forvar4406 + (1'h1)))
                    begin
                      reg4407 <= forvar4192[(3'h6):(3'h5)];
                      reg4408 <= reg4410[(2'h2):(1'h1)];
                      reg4409 <= (~^(~reg4249[(4'hb):(4'ha)]));
                      reg4410 <= reg4400;
                    end
                  for (forvar4411 = (1'h0); (forvar4411 < (2'h3)); forvar4411 = (forvar4411 + (1'h1)))
                    begin
                      reg4412 <= ((reg4385[(4'hc):(3'h6)] > $unsigned($unsigned((8'h9d)))) + forvar4394[(1'h0):(1'h0)]);
                      reg4413 <= reg4409[(3'h6):(3'h6)];
                      reg4414 <= (8'h9f);
                    end
                  for (forvar4415 = (1'h0); (forvar4415 < (2'h3)); forvar4415 = (forvar4415 + (1'h1)))
                    begin
                      reg4416 <= reg4203;
                    end
                  for (forvar4417 = (1'h0); (forvar4417 < (1'h1)); forvar4417 = (forvar4417 + (1'h1)))
                    begin
                      reg4418 <= (~&$unsigned(((+reg4372) >= (reg3877 << reg3887))));
                      reg4419 <= (~$unsigned(forvar4232));
                    end
                end
              if ((($unsigned({reg4200}) ?
                      reg3838[(3'h6):(1'h1)] : reg4247[(2'h3):(1'h1)]) ?
                  (reg4237 ? reg3855[(3'h6):(3'h6)] : reg3866) : wire4154))
                begin
                  for (forvar4420 = (1'h0); (forvar4420 < (2'h3)); forvar4420 = (forvar4420 + (1'h1)))
                    begin
                      reg4421 <= reg3887;
                    end
                  for (forvar4422 = (1'h0); (forvar4422 < (2'h2)); forvar4422 = (forvar4422 + (1'h1)))
                    begin
                      reg4423 <= reg3857[(1'h1):(1'h0)];
                      reg4424 <= (^~(~|$unsigned({reg3860})));
                      reg4425 <= $signed($signed($unsigned(reg4301[(3'h6):(2'h2)])));
                      reg4426 <= $unsigned($unsigned(reg3841[(1'h0):(1'h0)]));
                    end
                  if (reg4418[(1'h1):(1'h0)])
                    begin
                      reg4427 <= reg3886[(3'h4):(1'h0)];
                      reg4428 <= reg4395;
                    end
                  else
                    begin
                      reg4427 <= {(reg4425[(3'h6):(1'h0)] ?
                              ({reg4421} ?
                                  $unsigned(reg3836) : $signed(reg3905)) : (^~reg4304))};
                      reg4428 <= ($unsigned((reg3826[(1'h0):(1'h0)] ?
                              (reg4377 ?
                                  (8'ha3) : forvar4187) : $signed(reg4208))) ?
                          $unsigned((-reg4195)) : reg3846);
                    end
                end
              else
                begin
                  if ($unsigned(reg4178))
                    begin
                      reg4420 <= reg3842[(4'hf):(1'h1)];
                    end
                  else
                    begin
                      reg4420 <= $unsigned(({(forvar4405 ?
                              forvar4299 : reg4366)} > $unsigned((~^reg4421))));
                      reg4421 <= (((~(forvar4235 ?
                          forvar3920 : forvar4174)) & $unsigned((reg3796 << reg4321))) >= reg4414[(3'h4):(2'h3)]);
                      reg4422 <= (~|reg4293);
                      reg4423 <= (|$unsigned(reg4418[(4'h9):(4'h9)]));
                    end
                  if ((($unsigned($unsigned(reg4339)) ?
                          ((reg4402 ? (8'hb4) : reg3916) ?
                              forvar4300[(1'h1):(1'h0)] : (forvar4380 ?
                                  reg3791 : reg3898)) : $signed(reg4160)) ?
                      (+(|reg4352[(3'h6):(2'h3)])) : $unsigned(reg4289)))
                    begin
                      reg4424 <= forvar3806;
                    end
                  else
                    begin
                      reg4424 <= forvar3879;
                      reg4425 <= (!reg4202);
                      reg4426 <= (reg4242[(4'ha):(1'h0)] ?
                          (($unsigned(reg3887) ?
                              reg3878 : $unsigned(reg4345)) <= $unsigned({reg4196})) : forvar4174[(3'h6):(3'h4)]);
                      reg4427 <= forvar4171;
                    end
                  for (forvar4428 = (1'h0); (forvar4428 < (1'h0)); forvar4428 = (forvar4428 + (1'h1)))
                    begin
                      reg4429 <= reg3851;
                    end
                end
              for (forvar4430 = (1'h0); (forvar4430 < (1'h0)); forvar4430 = (forvar4430 + (1'h1)))
                begin
                  reg4431 <= $signed($signed($signed($unsigned(reg3801))));
                  if ({(reg3825 ?
                          (reg3869[(3'h5):(2'h3)] ?
                              {reg3885} : {forvar4363}) : reg3841[(1'h0):(1'h0)])})
                    begin
                      reg4432 <= $unsigned($signed({reg3816[(2'h2):(2'h2)]}));
                      reg4433 <= ((^(reg3816 ?
                              (reg4210 && reg3905) : (forvar4337 >> reg4412))) ?
                          reg3918 : reg3859[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg4432 <= $unsigned(($unsigned((reg4398 >> reg3798)) ^ {reg3799}));
                      reg4433 <= (forvar4417[(2'h2):(1'h0)] >>> (~{(~^reg3896)}));
                    end
                end
              if ({$signed({(&forvar4223)})})
                begin
                  for (forvar4434 = (1'h0); (forvar4434 < (2'h2)); forvar4434 = (forvar4434 + (1'h1)))
                    begin
                      reg4435 <= ((reg4166 ?
                          (^{(8'ha1)}) : forvar3871) ^ $signed(reg3790[(2'h3):(2'h3)]));
                      reg4436 <= {(|$unsigned(reg4433[(4'h9):(3'h4)]))};
                    end
                  if ($signed($signed((forvar4405 >= (forvar3894 ?
                      forvar4265 : forvar4422)))))
                    begin
                      reg4437 <= ({reg4353} <= reg4205);
                      reg4438 <= ((reg4321[(3'h7):(2'h3)] ?
                          (-(wire4154 + reg4383)) : {reg3914[(3'h7):(3'h7)]}) > reg4216[(2'h2):(1'h1)]);
                      reg4439 <= reg3810[(3'h4):(1'h1)];
                      reg4440 <= ($signed(reg3905[(2'h3):(2'h3)]) << ((reg4185[(1'h0):(1'h0)] ?
                          (forvar4394 ?
                              forvar4163 : forvar4262) : reg4356) > (reg3799[(4'h8):(3'h4)] ^ $unsigned((8'haa)))));
                    end
                  else
                    begin
                      reg4437 <= (($signed(forvar3834) != ($signed((8'h9d)) > $unsigned((8'h9d)))) ^~ (($signed(reg4220) ?
                          $signed(reg4439) : $signed(reg3837)) >> (~(8'h9f))));
                      reg4438 <= reg4257;
                      reg4439 <= ($unsigned(($signed(forvar3785) ~^ forvar3915[(3'h6):(3'h6)])) <<< (+forvar4274));
                      reg4440 <= $unsigned((~&(~&reg4234[(4'hb):(4'h9)])));
                    end
                end
              else
                begin
                  if ($unsigned(reg4190))
                    begin
                      reg4434 <= (^~reg3800);
                      reg4435 <= {forvar3837[(1'h1):(1'h1)]};
                      reg4436 <= reg4304;
                    end
                  else
                    begin
                      reg4434 <= (~(({reg4297} <= (reg3900 ?
                          reg4353 : forvar4401)) << forvar3894));
                      reg4435 <= (($unsigned($signed(reg4203)) <<< $unsigned((forvar4241 ?
                              forvar3928 : reg3927))) ?
                          reg4341 : ($unsigned((^forvar4262)) ?
                              (-$unsigned((8'hb4))) : reg4172));
                      reg4436 <= $unsigned((forvar3879[(4'h8):(3'h7)] == reg4313[(1'h1):(1'h0)]));
                      reg4437 <= $signed($signed(forvar4219));
                    end
                  if (reg4349[(1'h1):(1'h0)])
                    begin
                      reg4438 <= (^~(reg4357 || ((reg4249 && reg4197) >> {(8'h9d)})));
                      reg4439 <= $signed((((^reg3913) ?
                          reg4403[(4'hb):(3'h7)] : reg3786[(1'h1):(1'h1)]) >= (8'ha7)));
                      reg4440 <= (&(-(8'hac)));
                    end
                  else
                    begin
                      reg4438 <= (reg4339 | reg3864[(2'h2):(1'h1)]);
                      reg4439 <= $unsigned(reg4178);
                      reg4440 <= ((|((wire3781 ?
                              (8'h9c) : reg4424) ~^ (+(8'ha8)))) ?
                          ($unsigned({forvar4283}) ?
                              reg3878 : (|(8'ha4))) : reg4271);
                      reg4441 <= forvar4380;
                    end
                  for (forvar4442 = (1'h0); (forvar4442 < (1'h0)); forvar4442 = (forvar4442 + (1'h1)))
                    begin
                      reg4443 <= (+($unsigned($unsigned(forvar4299)) ?
                          $signed((8'h9f)) : (&$signed(reg4203))));
                      reg4444 <= $signed((~&reg4229[(4'hd):(4'h8)]));
                    end
                  for (forvar4445 = (1'h0); (forvar4445 < (1'h1)); forvar4445 = (forvar4445 + (1'h1)))
                    begin
                      reg4446 <= $signed((^~(forvar4283 <= $unsigned(reg4228))));
                    end
                end
            end
        end
      for (forvar4447 = (1'h0); (forvar4447 < (2'h3)); forvar4447 = (forvar4447 + (1'h1)))
        begin
          for (forvar4448 = (1'h0); (forvar4448 < (1'h0)); forvar4448 = (forvar4448 + (1'h1)))
            begin
              if (reg3874[(1'h1):(1'h1)])
                begin
                  for (forvar4449 = (1'h0); (forvar4449 < (1'h0)); forvar4449 = (forvar4449 + (1'h1)))
                    begin
                      reg4450 <= $signed($unsigned($unsigned((8'hba))));
                      reg4451 <= {reg4322};
                    end
                  for (forvar4452 = (1'h0); (forvar4452 < (1'h1)); forvar4452 = (forvar4452 + (1'h1)))
                    begin
                      reg4453 <= $signed((($signed(reg4170) ?
                              (forvar4235 || reg3817) : $unsigned((8'hab))) ?
                          ($signed(forvar3795) ?
                              reg4325[(3'h6):(1'h0)] : (reg4172 ?
                                  (8'haf) : reg4420)) : $signed((reg4403 >> reg4324))));
                    end
                  if ({(-$unsigned(((8'h9d) ^~ forvar4206)))})
                    begin
                      reg4454 <= reg3923;
                      reg4455 <= $unsigned({(&(~reg4234))});
                    end
                  else
                    begin
                      reg4454 <= (8'hac);
                    end
                end
              else
                begin
                  if ((reg4429 ?
                      ($signed((|reg4328)) ?
                          forvar4411[(2'h2):(2'h2)] : (8'ha8)) : (({forvar4382} ?
                          reg4200[(3'h6):(3'h4)] : reg4375) >> {$signed(reg4401)})))
                    begin
                      reg4449 <= (~$signed(($signed(reg3885) < (reg4437 ^ forvar3920))));
                      reg4450 <= reg4439;
                    end
                  else
                    begin
                      reg4449 <= (+$unsigned($signed((forvar4384 ?
                          reg4372 : (8'hb3)))));
                    end
                  if (((^~(~(~reg4390))) ?
                      $unsigned({(~&reg3890)}) : $signed(forvar4242)))
                    begin
                      reg4451 <= reg4349[(3'h5):(3'h5)];
                      reg4452 <= (!forvar4380);
                      reg4453 <= reg4244;
                      reg4454 <= ($signed(($signed(forvar4384) >= $unsigned(reg4353))) ?
                          $signed(reg4341[(3'h5):(2'h2)]) : reg4349);
                    end
                  else
                    begin
                      reg4451 <= (~reg3897[(4'h9):(2'h2)]);
                    end
                end
            end
        end
    end
  assign wire4456 = (8'hb0);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3931
#( parameter param4153 = (&(-(((8'hb3) ? (8'hb6) : (8'hac)) ? ((8'h9c) ? (8'h9f) : (8'ha0)) : ((8'haa) ~^ (8'ha5))))) )
(y, clk, wire3935, wire3934, wire3933, wire3932);
  output wire [(32'h89b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire3935;
  input wire [(2'h3):(1'h0)] wire3934;
  input wire [(4'hd):(1'h0)] wire3933;
  input wire [(2'h3):(1'h0)] wire3932;
  wire signed [(4'hc):(1'h0)] wire4152;
  wire [(3'h6):(1'h0)] wire4151;
  wire [(3'h5):(1'h0)] wire4150;
  wire signed [(4'he):(1'h0)] wire4149;
  reg [(4'hf):(1'h0)] reg4148 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4147 = (1'h0);
  reg [(2'h3):(1'h0)] reg4146 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4145 = (1'h0);
  reg [(3'h5):(1'h0)] reg4144 = (1'h0);
  reg [(3'h7):(1'h0)] reg4143 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4142 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4141 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4140 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4139 = (1'h0);
  reg [(2'h3):(1'h0)] reg4138 = (1'h0);
  reg [(3'h7):(1'h0)] reg4137 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4136 = (1'h0);
  reg [(4'h9):(1'h0)] reg4135 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4134 = (1'h0);
  reg [(4'ha):(1'h0)] reg4133 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4131 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4127 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4123 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4122 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4120 = (1'h0);
  reg [(4'hd):(1'h0)] reg4132 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4131 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4130 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4129 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4128 = (1'h0);
  reg [(4'ha):(1'h0)] reg4127 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4126 = (1'h0);
  reg [(4'ha):(1'h0)] reg4125 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4124 = (1'h0);
  reg [(3'h5):(1'h0)] reg4123 = (1'h0);
  reg [(3'h6):(1'h0)] reg4122 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4121 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4120 = (1'h0);
  reg [(4'he):(1'h0)] reg4119 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4118 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4117 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4116 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4115 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4114 = (1'h0);
  reg [(3'h5):(1'h0)] reg4113 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4112 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4111 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4110 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4109 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4108 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4107 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4106 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4105 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4104 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4103 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4102 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4101 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4098 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4094 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4092 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4100 = (1'h0);
  reg [(3'h6):(1'h0)] reg4097 = (1'h0);
  reg [(3'h4):(1'h0)] reg4096 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4095 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4093 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4091 = (1'h0);
  reg [(2'h2):(1'h0)] reg4089 = (1'h0);
  reg [(3'h4):(1'h0)] reg4083 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4082 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4081 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4099 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4098 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4097 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4096 = (1'h0);
  reg [(4'hb):(1'h0)] reg4095 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4094 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4093 = (1'h0);
  reg [(5'h10):(1'h0)] reg4092 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4091 = (1'h0);
  reg [(4'hd):(1'h0)] reg4090 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4089 = (1'h0);
  reg [(3'h7):(1'h0)] reg4088 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4087 = (1'h0);
  reg [(5'h10):(1'h0)] reg4086 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4085 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4084 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4083 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4082 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4081 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4080 = (1'h0);
  reg [(4'hd):(1'h0)] reg4079 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4078 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4077 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4076 = (1'h0);
  reg [(4'h8):(1'h0)] reg4075 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4074 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4073 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4072 = (1'h0);
  reg [(4'hd):(1'h0)] reg4071 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4070 = (1'h0);
  reg [(4'ha):(1'h0)] reg4069 = (1'h0);
  reg [(4'he):(1'h0)] reg4068 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4067 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4064 = (1'h0);
  reg [(3'h6):(1'h0)] reg4066 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4065 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4064 = (1'h0);
  reg [(3'h5):(1'h0)] reg4063 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4062 = (1'h0);
  reg [(4'h9):(1'h0)] reg4061 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4060 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4059 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4058 = (1'h0);
  reg [(4'hf):(1'h0)] reg4057 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4056 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4055 = (1'h0);
  reg [(4'h8):(1'h0)] reg4048 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4054 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4053 = (1'h0);
  reg [(5'h10):(1'h0)] reg4052 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4051 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4050 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4049 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4048 = (1'h0);
  reg [(5'h10):(1'h0)] reg4047 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4046 = (1'h0);
  reg [(2'h3):(1'h0)] reg4045 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4044 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4043 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4042 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4041 = (1'h0);
  reg [(4'he):(1'h0)] reg4040 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4039 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4038 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4037 = (1'h0);
  reg [(3'h7):(1'h0)] reg4036 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4035 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4034 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4033 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4032 = (1'h0);
  reg [(3'h5):(1'h0)] reg4031 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4030 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4029 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4028 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4026 = (1'h0);
  reg [(4'ha):(1'h0)] reg4029 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4028 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4027 = (1'h0);
  reg [(4'he):(1'h0)] reg4023 = (1'h0);
  reg [(5'h10):(1'h0)] reg4022 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4026 = (1'h0);
  reg [(4'he):(1'h0)] reg4025 = (1'h0);
  reg [(5'h10):(1'h0)] reg4024 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4023 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4022 = (1'h0);
  reg [(4'ha):(1'h0)] reg4021 = (1'h0);
  reg [(4'hd):(1'h0)] reg4020 = (1'h0);
  reg [(5'h10):(1'h0)] reg4019 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4018 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4017 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4016 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4015 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4014 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4013 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4012 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4011 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4010 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3978 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3977 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3975 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3973 = (1'h0);
  reg [(4'hb):(1'h0)] reg4009 = (1'h0);
  reg [(4'hf):(1'h0)] reg4008 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4007 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4006 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4005 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4004 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4003 = (1'h0);
  reg [(4'hb):(1'h0)] reg4002 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4001 = (1'h0);
  reg [(4'he):(1'h0)] reg4000 = (1'h0);
  reg [(2'h3):(1'h0)] reg3999 = (1'h0);
  reg [(3'h6):(1'h0)] reg3998 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3997 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3996 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3995 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3994 = (1'h0);
  reg [(4'he):(1'h0)] reg3993 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3992 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3991 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3990 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3989 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3988 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3987 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3986 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3985 = (1'h0);
  reg [(5'h10):(1'h0)] reg3984 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3983 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3982 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3981 = (1'h0);
  reg [(3'h5):(1'h0)] reg3980 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3979 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3978 = (1'h0);
  reg [(3'h5):(1'h0)] reg3977 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3976 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3975 = (1'h0);
  reg [(3'h6):(1'h0)] reg3974 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3973 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3972 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3971 = (1'h0);
  reg [(3'h7):(1'h0)] reg3971 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3970 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3969 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3968 = (1'h0);
  reg [(4'hb):(1'h0)] reg3967 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3966 = (1'h0);
  reg [(5'h10):(1'h0)] reg3965 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3964 = (1'h0);
  reg [(4'hf):(1'h0)] reg3963 = (1'h0);
  reg [(2'h3):(1'h0)] reg3962 = (1'h0);
  reg [(4'ha):(1'h0)] reg3961 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3960 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3959 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3957 = (1'h0);
  reg [(4'he):(1'h0)] reg3952 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3958 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3957 = (1'h0);
  reg [(3'h6):(1'h0)] reg3956 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3955 = (1'h0);
  reg [(2'h3):(1'h0)] reg3954 = (1'h0);
  reg [(2'h3):(1'h0)] reg3953 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3952 = (1'h0);
  reg [(4'he):(1'h0)] reg3951 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3950 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3949 = (1'h0);
  reg [(4'h8):(1'h0)] reg3948 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3947 = (1'h0);
  reg [(4'hf):(1'h0)] reg3946 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3945 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3944 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3943 = (1'h0);
  reg [(2'h3):(1'h0)] reg3943 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3942 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3941 = (1'h0);
  wire [(2'h2):(1'h0)] wire3940;
  reg signed [(3'h4):(1'h0)] reg3939 = (1'h0);
  reg [(3'h6):(1'h0)] reg3938 = (1'h0);
  wire [(4'h8):(1'h0)] wire3937;
  wire [(3'h6):(1'h0)] wire3936;
  assign y = {wire4152,
                 wire4151,
                 wire4150,
                 wire4149,
                 reg4148,
                 forvar4147,
                 reg4146,
                 reg4145,
                 reg4144,
                 reg4143,
                 reg4142,
                 forvar4141,
                 forvar4140,
                 forvar4139,
                 reg4138,
                 reg4137,
                 forvar4136,
                 reg4135,
                 reg4134,
                 reg4133,
                 forvar4131,
                 forvar4127,
                 forvar4123,
                 forvar4122,
                 reg4120,
                 reg4132,
                 reg4131,
                 reg4130,
                 reg4129,
                 reg4128,
                 reg4127,
                 reg4126,
                 reg4125,
                 reg4124,
                 reg4123,
                 reg4122,
                 reg4121,
                 forvar4120,
                 reg4119,
                 reg4118,
                 reg4117,
                 forvar4116,
                 forvar4115,
                 forvar4114,
                 reg4113,
                 reg4112,
                 reg4111,
                 reg4110,
                 forvar4109,
                 forvar4108,
                 reg4107,
                 reg4106,
                 forvar4105,
                 forvar4104,
                 reg4103,
                 forvar4102,
                 reg4101,
                 forvar4098,
                 reg4094,
                 forvar4092,
                 reg4100,
                 reg4097,
                 reg4096,
                 forvar4095,
                 reg4093,
                 forvar4091,
                 reg4089,
                 reg4083,
                 reg4082,
                 forvar4081,
                 reg4099,
                 reg4098,
                 forvar4097,
                 forvar4096,
                 reg4095,
                 forvar4094,
                 forvar4093,
                 reg4092,
                 reg4091,
                 reg4090,
                 forvar4089,
                 reg4088,
                 reg4087,
                 reg4086,
                 reg4085,
                 reg4084,
                 forvar4083,
                 forvar4082,
                 reg4081,
                 reg4080,
                 reg4079,
                 reg4078,
                 forvar4077,
                 reg4076,
                 reg4075,
                 reg4074,
                 reg4073,
                 forvar4072,
                 reg4071,
                 reg4070,
                 reg4069,
                 reg4068,
                 forvar4067,
                 reg4064,
                 reg4066,
                 reg4065,
                 forvar4064,
                 reg4063,
                 reg4062,
                 reg4061,
                 forvar4060,
                 reg4059,
                 reg4058,
                 reg4057,
                 reg4056,
                 forvar4055,
                 reg4048,
                 reg4054,
                 reg4053,
                 reg4052,
                 reg4051,
                 reg4050,
                 reg4049,
                 forvar4048,
                 reg4047,
                 reg4046,
                 reg4045,
                 forvar4044,
                 reg4043,
                 reg4042,
                 forvar4041,
                 reg4040,
                 forvar4039,
                 forvar4038,
                 reg4037,
                 reg4036,
                 reg4035,
                 reg4034,
                 forvar4033,
                 forvar4032,
                 reg4031,
                 reg4030,
                 forvar4029,
                 reg4028,
                 forvar4026,
                 reg4029,
                 forvar4028,
                 reg4027,
                 reg4023,
                 reg4022,
                 reg4026,
                 reg4025,
                 reg4024,
                 forvar4023,
                 forvar4022,
                 reg4021,
                 reg4020,
                 reg4019,
                 reg4018,
                 forvar4017,
                 reg4016,
                 reg4015,
                 reg4014,
                 reg4013,
                 forvar4012,
                 forvar4011,
                 forvar4010,
                 reg3978,
                 forvar3977,
                 forvar3975,
                 reg3973,
                 reg4009,
                 reg4008,
                 forvar4007,
                 forvar4006,
                 reg4005,
                 reg4004,
                 reg4003,
                 reg4002,
                 forvar4001,
                 reg4000,
                 reg3999,
                 reg3998,
                 forvar3997,
                 reg3996,
                 forvar3995,
                 reg3994,
                 reg3993,
                 forvar3992,
                 reg3991,
                 reg3990,
                 forvar3989,
                 reg3988,
                 reg3987,
                 forvar3986,
                 forvar3985,
                 reg3984,
                 reg3983,
                 reg3982,
                 forvar3981,
                 reg3980,
                 reg3979,
                 forvar3978,
                 reg3977,
                 reg3976,
                 reg3975,
                 reg3974,
                 forvar3973,
                 reg3972,
                 forvar3971,
                 reg3971,
                 reg3970,
                 reg3969,
                 forvar3968,
                 reg3967,
                 reg3966,
                 reg3965,
                 reg3964,
                 reg3963,
                 reg3962,
                 reg3961,
                 forvar3960,
                 forvar3959,
                 forvar3957,
                 reg3952,
                 reg3958,
                 reg3957,
                 reg3956,
                 reg3955,
                 reg3954,
                 reg3953,
                 forvar3952,
                 reg3951,
                 reg3950,
                 reg3949,
                 reg3948,
                 reg3947,
                 reg3946,
                 forvar3945,
                 reg3944,
                 forvar3943,
                 reg3943,
                 forvar3942,
                 forvar3941,
                 wire3940,
                 reg3939,
                 reg3938,
                 wire3937,
                 wire3936,
                 (1'h0)};
  assign wire3936 = $signed($unsigned($signed((wire3932 | wire3934))));
  assign wire3937 = wire3936;
  always
    @(posedge clk) begin
      reg3938 <= $unsigned(wire3934[(1'h0):(1'h0)]);
      reg3939 <= wire3937[(3'h5):(1'h1)];
    end
  assign wire3940 = (wire3933[(4'hb):(2'h3)] || $unsigned(reg3939[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      for (forvar3941 = (1'h0); (forvar3941 < (2'h3)); forvar3941 = (forvar3941 + (1'h1)))
        begin
          for (forvar3942 = (1'h0); (forvar3942 < (1'h0)); forvar3942 = (forvar3942 + (1'h1)))
            begin
              if ((8'hb6))
                begin
                  if ({forvar3942[(3'h5):(3'h4)]})
                    begin
                      reg3943 <= $signed($signed(($signed(forvar3941) >= reg3939)));
                    end
                  else
                    begin
                      reg3943 <= (((^(wire3940 | wire3935)) ?
                              $unsigned($unsigned(forvar3941)) : reg3943) ?
                          $signed(wire3933[(1'h0):(1'h0)]) : ((-(reg3938 ?
                                  (8'h9e) : wire3940)) ?
                              (+$unsigned(wire3940)) : wire3932));
                    end
                end
              else
                begin
                  for (forvar3943 = (1'h0); (forvar3943 < (1'h1)); forvar3943 = (forvar3943 + (1'h1)))
                    begin
                      reg3944 <= ((|forvar3942) ?
                          (~&$unsigned(reg3939)) : wire3934);
                    end
                  for (forvar3945 = (1'h0); (forvar3945 < (2'h3)); forvar3945 = (forvar3945 + (1'h1)))
                    begin
                      reg3946 <= wire3936[(3'h4):(1'h0)];
                      reg3947 <= {(!{$signed(reg3943)})};
                      reg3948 <= (wire3940[(1'h0):(1'h0)] | reg3938[(3'h4):(2'h3)]);
                    end
                end
            end
          reg3949 <= ((^~$unsigned((~&reg3938))) & $signed(reg3946[(1'h1):(1'h1)]));
        end
      if ((~^$unsigned({{forvar3941}})))
        begin
          reg3950 <= ((~|wire3935) ~^ reg3939);
          if ({forvar3942})
            begin
              reg3951 <= $unsigned(reg3939);
              if (({reg3946[(3'h5):(2'h2)]} ?
                  (^(reg3951 ?
                      (wire3934 < forvar3941) : reg3943[(2'h2):(1'h1)])) : reg3949[(4'hc):(4'h9)]))
                begin
                  for (forvar3952 = (1'h0); (forvar3952 < (1'h1)); forvar3952 = (forvar3952 + (1'h1)))
                    begin
                      reg3953 <= (~^(8'ha2));
                    end
                  reg3954 <= wire3933;
                  if ((^~{(reg3949 < (reg3943 < forvar3941))}))
                    begin
                      reg3955 <= $signed(wire3932);
                      reg3956 <= {wire3933};
                      reg3957 <= (($signed($signed(wire3940)) ?
                              (forvar3943[(1'h0):(1'h0)] ^ (reg3948 & reg3948)) : reg3948) ?
                          $signed((^~(wire3936 ^~ reg3950))) : wire3934);
                      reg3958 <= (|(reg3946 ?
                          forvar3952[(3'h4):(1'h1)] : ((reg3947 < wire3937) - reg3953[(2'h2):(2'h2)])));
                    end
                  else
                    begin
                      reg3955 <= reg3949;
                      reg3956 <= (~((&reg3948[(3'h6):(1'h0)]) < reg3949));
                      reg3957 <= ((^$signed(forvar3945[(3'h5):(2'h2)])) <= ($signed($unsigned(wire3933)) ?
                          (wire3933 + {wire3934}) : ((^reg3950) << reg3958)));
                      reg3958 <= (^((((8'hb7) ?
                          (8'hab) : reg3955) || $signed(forvar3942)) + $unsigned({reg3953})));
                    end
                end
              else
                begin
                  for (forvar3952 = (1'h0); (forvar3952 < (2'h3)); forvar3952 = (forvar3952 + (1'h1)))
                    begin
                      reg3953 <= (((^~(&reg3956)) ? (8'h9f) : (-(^wire3940))) ?
                          $unsigned($signed($signed(reg3938))) : $unsigned(((&(8'h9f)) ?
                              (reg3956 ~^ wire3936) : $signed(wire3933))));
                      reg3954 <= $signed({reg3944[(4'hb):(4'ha)]});
                      reg3955 <= reg3950;
                      reg3956 <= ($unsigned(((~^forvar3942) >= (reg3950 ?
                          (8'hb7) : reg3947))) >= {(reg3954 ?
                              reg3955[(4'ha):(3'h6)] : (wire3937 ?
                                  reg3946 : reg3953))});
                    end
                  reg3957 <= {wire3936[(3'h5):(2'h3)]};
                end
            end
          else
            begin
              if ($unsigned(wire3933[(4'ha):(4'h9)]))
                begin
                  reg3951 <= ($signed(reg3949) ?
                      $signed(((reg3951 ?
                          reg3951 : (8'ha8)) <<< (forvar3945 >> wire3936))) : $unsigned($unsigned((|reg3939))));
                  if ((^$signed((forvar3952[(3'h5):(3'h4)] ?
                      $unsigned(wire3933) : (reg3939 ~^ forvar3943)))))
                    begin
                      reg3952 <= $signed(reg3955);
                    end
                  else
                    begin
                      reg3952 <= $signed($unsigned(((reg3948 != forvar3945) | (wire3933 ?
                          wire3934 : reg3955))));
                    end
                  if (reg3953[(2'h2):(2'h2)])
                    begin
                      reg3953 <= wire3934[(1'h0):(1'h0)];
                      reg3954 <= (forvar3952[(2'h2):(2'h2)] ?
                          (&reg3949[(4'hc):(2'h2)]) : (~&(reg3953[(1'h0):(1'h0)] ?
                              (forvar3941 ?
                                  reg3957 : wire3932) : (~|reg3950))));
                    end
                  else
                    begin
                      reg3953 <= $signed(reg3943);
                      reg3954 <= (~|forvar3943);
                      reg3955 <= $signed(reg3943[(1'h0):(1'h0)]);
                      reg3956 <= (8'hba);
                    end
                  for (forvar3957 = (1'h0); (forvar3957 < (1'h0)); forvar3957 = (forvar3957 + (1'h1)))
                    begin
                      reg3958 <= (^(~|(forvar3952 ?
                          {reg3954} : $unsigned((8'ha2)))));
                    end
                end
              else
                begin
                  if ((~(8'h9f)))
                    begin
                      reg3951 <= (forvar3943 ^ $signed((~|(reg3952 <= forvar3941))));
                    end
                  else
                    begin
                      reg3951 <= $unsigned(((8'ha7) ?
                          (!wire3932) : ((8'had) ?
                              reg3951[(2'h2):(1'h1)] : (^~forvar3941))));
                      reg3952 <= $unsigned($unsigned(reg3954[(1'h1):(1'h0)]));
                      reg3953 <= ((forvar3952 ?
                          $signed(((8'had) + reg3946)) : (8'hb0)) >= ({$signed(forvar3941)} ?
                          ({reg3947} ?
                              (!reg3955) : (wire3932 ?
                                  wire3935 : forvar3957)) : {(8'hb8)}));
                      reg3954 <= (reg3956[(2'h2):(1'h1)] ?
                          {({forvar3943} ?
                                  $unsigned((8'hab)) : ((8'ha1) ?
                                      wire3935 : wire3933))} : (($signed(reg3943) ?
                              $signed((8'ha6)) : forvar3943) <<< forvar3957[(4'h9):(3'h5)]));
                    end
                end
              for (forvar3959 = (1'h0); (forvar3959 < (1'h1)); forvar3959 = (forvar3959 + (1'h1)))
                begin
                  for (forvar3960 = (1'h0); (forvar3960 < (1'h1)); forvar3960 = (forvar3960 + (1'h1)))
                    begin
                      reg3961 <= wire3935[(2'h3):(2'h2)];
                      reg3962 <= $unsigned((8'hb5));
                      reg3963 <= (!({(forvar3942 ?
                              (8'hb5) : reg3951)} - (|$signed(wire3932))));
                    end
                  if ((&($signed(reg3948) ? reg3957 : (&reg3943))))
                    begin
                      reg3964 <= $unsigned((((reg3963 ?
                          wire3937 : (8'hb0)) - $signed(reg3955)) < (reg3943 ?
                          {(8'hb2)} : reg3961)));
                    end
                  else
                    begin
                      reg3964 <= reg3954;
                      reg3965 <= reg3939[(2'h2):(1'h1)];
                    end
                  if (($signed({$signed(reg3961)}) ?
                      (|(forvar3941[(2'h3):(2'h2)] ?
                          (reg3951 ~^ (8'hb2)) : (reg3954 ?
                              wire3937 : wire3937))) : $unsigned(reg3955[(4'ha):(4'h8)])))
                    begin
                      reg3966 <= $unsigned(reg3961);
                      reg3967 <= $unsigned($signed($unsigned($unsigned(reg3938))));
                    end
                  else
                    begin
                      reg3966 <= ($signed((-forvar3943)) << reg3947[(2'h3):(2'h3)]);
                      reg3967 <= (^~(|$signed(wire3932[(1'h1):(1'h1)])));
                    end
                  for (forvar3968 = (1'h0); (forvar3968 < (1'h0)); forvar3968 = (forvar3968 + (1'h1)))
                    begin
                      reg3969 <= $unsigned($unsigned(($unsigned(wire3932) ?
                          {reg3947} : $signed(reg3961))));
                      reg3970 <= $unsigned($signed({(reg3961 ?
                              reg3946 : reg3939)}));
                    end
                end
            end
        end
      else
        begin
          reg3950 <= {$signed(wire3934)};
        end
      if ((reg3964 < $unsigned($signed($signed((8'ha1))))))
        begin
          reg3971 <= $signed((&$unsigned(reg3954)));
        end
      else
        begin
          if (reg3948[(4'h8):(4'h8)])
            begin
              for (forvar3971 = (1'h0); (forvar3971 < (2'h2)); forvar3971 = (forvar3971 + (1'h1)))
                begin
                  reg3972 <= reg3957;
                  for (forvar3973 = (1'h0); (forvar3973 < (2'h3)); forvar3973 = (forvar3973 + (1'h1)))
                    begin
                      reg3974 <= (reg3953 ?
                          {wire3940[(2'h2):(2'h2)]} : (((+reg3952) ?
                                  $signed(forvar3943) : $unsigned(reg3967)) ?
                              reg3958 : (&reg3939)));
                      reg3975 <= $signed((&(|$unsigned(reg3944))));
                      reg3976 <= $unsigned((forvar3952 << (reg3961[(3'h6):(3'h5)] == (forvar3943 & reg3950))));
                      reg3977 <= $signed(reg3938[(3'h6):(3'h4)]);
                    end
                  for (forvar3978 = (1'h0); (forvar3978 < (1'h1)); forvar3978 = (forvar3978 + (1'h1)))
                    begin
                      reg3979 <= (8'ha9);
                      reg3980 <= forvar3968;
                    end
                  for (forvar3981 = (1'h0); (forvar3981 < (1'h0)); forvar3981 = (forvar3981 + (1'h1)))
                    begin
                      reg3982 <= $unsigned((&forvar3973));
                      reg3983 <= ({($signed(reg3982) <<< $signed((8'hb8)))} ?
                          (+(^~$signed(reg3976))) : ((reg3963 ?
                              $signed(reg3976) : reg3946) - (~&{(8'ha3)})));
                      reg3984 <= (+reg3976);
                    end
                end
              for (forvar3985 = (1'h0); (forvar3985 < (2'h2)); forvar3985 = (forvar3985 + (1'h1)))
                begin
                  for (forvar3986 = (1'h0); (forvar3986 < (2'h2)); forvar3986 = (forvar3986 + (1'h1)))
                    begin
                      reg3987 <= $unsigned($unsigned(($signed(reg3939) ?
                          (reg3955 || reg3979) : forvar3968)));
                    end
                  reg3988 <= (((reg3964 ?
                          wire3933 : ((8'ha8) ? forvar3978 : reg3982)) ?
                      {(reg3969 ?
                              reg3949 : reg3972)} : reg3948[(1'h1):(1'h0)]) ~^ {$unsigned((reg3961 ?
                          reg3982 : (8'haa)))});
                  for (forvar3989 = (1'h0); (forvar3989 < (1'h0)); forvar3989 = (forvar3989 + (1'h1)))
                    begin
                      reg3990 <= reg3987[(2'h2):(2'h2)];
                      reg3991 <= wire3940;
                    end
                end
              for (forvar3992 = (1'h0); (forvar3992 < (1'h0)); forvar3992 = (forvar3992 + (1'h1)))
                begin
                  if ($unsigned(($unsigned((reg3938 ?
                      reg3947 : reg3967)) > ((reg3971 ^~ (8'ha7)) & $signed(reg3991)))))
                    begin
                      reg3993 <= ((($signed(reg3975) && $signed(reg3977)) ?
                          ($signed(forvar3973) ~^ (8'hab)) : $signed(reg3943)) >> $signed($signed($signed(reg3956))));
                      reg3994 <= (8'h9e);
                    end
                  else
                    begin
                      reg3993 <= ($unsigned(reg3994[(2'h2):(2'h2)]) >> (reg3962[(1'h1):(1'h1)] ?
                          forvar3952 : (~^(~&wire3932))));
                      reg3994 <= (({((8'haf) << forvar3971)} >>> reg3950) ?
                          (reg3987[(1'h0):(1'h0)] ?
                              wire3932 : ($unsigned(reg3965) ^~ $unsigned(reg3969))) : $unsigned(((+(8'hb4)) > forvar3945[(1'h0):(1'h0)])));
                    end
                  for (forvar3995 = (1'h0); (forvar3995 < (2'h2)); forvar3995 = (forvar3995 + (1'h1)))
                    begin
                      reg3996 <= wire3934;
                    end
                  for (forvar3997 = (1'h0); (forvar3997 < (1'h1)); forvar3997 = (forvar3997 + (1'h1)))
                    begin
                      reg3998 <= forvar3968[(3'h7):(2'h3)];
                      reg3999 <= (~&forvar3943);
                      reg4000 <= reg3966[(1'h1):(1'h0)];
                    end
                  for (forvar4001 = (1'h0); (forvar4001 < (2'h2)); forvar4001 = (forvar4001 + (1'h1)))
                    begin
                      reg4002 <= reg3971;
                      reg4003 <= {forvar3992};
                      reg4004 <= (wire3933 ?
                          reg3955 : (+((reg3961 ? reg3949 : reg3987) ?
                              $signed(reg3951) : (reg3970 << reg4000))));
                      reg4005 <= (+$unsigned($unsigned((8'hac))));
                    end
                end
              for (forvar4006 = (1'h0); (forvar4006 < (1'h0)); forvar4006 = (forvar4006 + (1'h1)))
                begin
                  for (forvar4007 = (1'h0); (forvar4007 < (2'h3)); forvar4007 = (forvar4007 + (1'h1)))
                    begin
                      reg4008 <= reg3955[(4'h9):(4'h9)];
                      reg4009 <= forvar3943;
                    end
                end
            end
          else
            begin
              for (forvar3971 = (1'h0); (forvar3971 < (1'h1)); forvar3971 = (forvar3971 + (1'h1)))
                begin
                  if ((-reg3971[(3'h7):(1'h1)]))
                    begin
                      reg3972 <= reg3984;
                      reg3973 <= {(&(8'ha8))};
                    end
                  else
                    begin
                      reg3972 <= ($signed(forvar3997) ?
                          $signed((8'ha1)) : (reg3972 >>> {$unsigned(forvar3945)}));
                      reg3973 <= (!$unsigned(wire3940));
                      reg3974 <= forvar3981[(1'h0):(1'h0)];
                    end
                end
              for (forvar3975 = (1'h0); (forvar3975 < (1'h0)); forvar3975 = (forvar3975 + (1'h1)))
                begin
                  if ((~&((~&(~&reg3957)) ^~ $signed($signed(reg3977)))))
                    begin
                      reg3976 <= ($signed({reg3939}) <<< (~&($signed(reg3999) ?
                          (reg3994 <<< forvar3960) : (~reg3953))));
                    end
                  else
                    begin
                      reg3976 <= (reg3943[(1'h0):(1'h0)] | reg3951[(4'hd):(2'h3)]);
                    end
                  for (forvar3977 = (1'h0); (forvar3977 < (1'h1)); forvar3977 = (forvar3977 + (1'h1)))
                    begin
                      reg3978 <= ((|(~$signed((8'ha5)))) + ((8'ha5) ?
                          ({forvar3941} ?
                              $unsigned(reg3987) : $signed(reg3964)) : reg3946[(4'hc):(4'ha)]));
                    end
                  reg3979 <= $signed((!reg3946));
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar4010 = (1'h0); (forvar4010 < (2'h2)); forvar4010 = (forvar4010 + (1'h1)))
        begin
          for (forvar4011 = (1'h0); (forvar4011 < (2'h2)); forvar4011 = (forvar4011 + (1'h1)))
            begin
              for (forvar4012 = (1'h0); (forvar4012 < (2'h2)); forvar4012 = (forvar4012 + (1'h1)))
                begin
                  if ((forvar3992[(4'hb):(3'h5)] ?
                      (($signed(forvar4010) < (^reg3953)) ?
                          reg3954[(2'h3):(1'h0)] : $signed({forvar3978})) : (+{{(8'hb4)}})))
                    begin
                      reg4013 <= $unsigned(reg3999);
                      reg4014 <= (&(-(|(reg4005 ? reg3969 : reg3953))));
                      reg4015 <= reg3975;
                      reg4016 <= $signed((-wire3934[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg4013 <= $signed(forvar4001[(2'h3):(2'h2)]);
                    end
                  for (forvar4017 = (1'h0); (forvar4017 < (2'h2)); forvar4017 = (forvar4017 + (1'h1)))
                    begin
                      reg4018 <= (~reg4009);
                      reg4019 <= (^(($unsigned(reg3991) ?
                          reg3947 : $signed(forvar4007)) != (+{reg3973})));
                      reg4020 <= ($signed($unsigned((^~reg3953))) - ($signed((8'hae)) * $unsigned({reg3969})));
                    end
                end
              reg4021 <= (8'hb9);
            end
          if ((forvar4017 ?
              (((reg3996 ? forvar3960 : (8'ha7)) ?
                  reg4020[(4'h9):(2'h3)] : (reg4003 - wire3935)) != reg3951) : (($unsigned(reg3987) ?
                  {reg3947} : $signed(reg3991)) && (~^(reg3993 ?
                  forvar4001 : wire3940)))))
            begin
              for (forvar4022 = (1'h0); (forvar4022 < (2'h2)); forvar4022 = (forvar4022 + (1'h1)))
                begin
                  for (forvar4023 = (1'h0); (forvar4023 < (2'h3)); forvar4023 = (forvar4023 + (1'h1)))
                    begin
                      reg4024 <= $unsigned((((~(8'hb1)) ?
                          {(8'h9d)} : (forvar4017 ?
                              reg4008 : (8'hac))) >> ($signed(reg3938) ?
                          $signed((8'hb5)) : {reg3957})));
                      reg4025 <= $signed((^~reg4013));
                      reg4026 <= ($signed(wire3933) ?
                          reg4003[(2'h3):(2'h2)] : ($signed($unsigned(forvar3960)) ?
                              reg3993[(3'h7):(3'h5)] : ($unsigned(reg4002) <<< (reg3954 ?
                                  reg4008 : (8'hb9)))));
                    end
                end
            end
          else
            begin
              if (reg4025[(4'h9):(4'h9)])
                begin
                  if (reg4019)
                    begin
                      reg4022 <= (($unsigned({reg3965}) ?
                          $signed((8'ha2)) : (8'hae)) ^ $signed({(~^reg3950)}));
                    end
                  else
                    begin
                      reg4022 <= ((^((reg3952 ?
                          reg3951 : reg3972) <<< (|reg4026))) <<< (8'ha4));
                      reg4023 <= (reg3987[(1'h1):(1'h0)] < reg3962);
                      reg4024 <= forvar3992;
                    end
                  if (reg3978)
                    begin
                      reg4025 <= reg3952;
                      reg4026 <= $signed(((8'hae) ?
                          forvar4007[(1'h1):(1'h1)] : ((reg3961 ^~ reg3951) ?
                              (^reg4015) : reg3977)));
                      reg4027 <= ((~^(|{reg3949})) != $signed($unsigned(reg4026)));
                    end
                  else
                    begin
                      reg4025 <= forvar3959;
                    end
                  for (forvar4028 = (1'h0); (forvar4028 < (1'h1)); forvar4028 = (forvar4028 + (1'h1)))
                    begin
                      reg4029 <= forvar3952;
                    end
                end
              else
                begin
                  if ($signed(reg4014))
                    begin
                      reg4022 <= wire3933;
                    end
                  else
                    begin
                      reg4022 <= $signed(reg3948);
                      reg4023 <= wire3934;
                      reg4024 <= reg3994;
                      reg4025 <= forvar3989;
                    end
                  for (forvar4026 = (1'h0); (forvar4026 < (1'h0)); forvar4026 = (forvar4026 + (1'h1)))
                    begin
                      reg4027 <= (($signed((reg3962 & reg3980)) ?
                          $signed((reg4020 ?
                              reg3961 : forvar3971)) : (reg4000[(2'h3):(1'h1)] ?
                              reg3950 : $signed(reg3998))) && (&wire3936));
                      reg4028 <= (reg4015 >> (($signed(forvar3957) | reg4005) && (&$unsigned(reg3990))));
                    end
                  for (forvar4029 = (1'h0); (forvar4029 < (2'h2)); forvar4029 = (forvar4029 + (1'h1)))
                    begin
                      reg4030 <= {reg3943[(1'h0):(1'h0)]};
                      reg4031 <= $signed((~^reg3962[(2'h2):(1'h0)]));
                    end
                end
              for (forvar4032 = (1'h0); (forvar4032 < (2'h3)); forvar4032 = (forvar4032 + (1'h1)))
                begin
                  for (forvar4033 = (1'h0); (forvar4033 < (2'h3)); forvar4033 = (forvar4033 + (1'h1)))
                    begin
                      reg4034 <= (!($unsigned($signed(forvar4032)) ~^ $unsigned($unsigned(wire3935))));
                      reg4035 <= $unsigned((~^(!(forvar3973 ?
                          reg3996 : forvar3952))));
                      reg4036 <= (((-(reg4008 ?
                              reg3953 : reg4003)) || ($unsigned(forvar4017) ?
                              $signed(forvar4023) : (forvar3978 << reg3970))) ?
                          ($signed((reg3999 ~^ reg3999)) | forvar3975) : (reg3991 ?
                              (((8'hb1) ?
                                  forvar3981 : forvar3957) ~^ (reg4008 & reg3999)) : reg3946));
                      reg4037 <= reg3980;
                    end
                end
            end
          for (forvar4038 = (1'h0); (forvar4038 < (2'h3)); forvar4038 = (forvar4038 + (1'h1)))
            begin
              for (forvar4039 = (1'h0); (forvar4039 < (2'h3)); forvar4039 = (forvar4039 + (1'h1)))
                begin
                  reg4040 <= {$unsigned(reg4036[(3'h7):(1'h1)])};
                  for (forvar4041 = (1'h0); (forvar4041 < (2'h3)); forvar4041 = (forvar4041 + (1'h1)))
                    begin
                      reg4042 <= reg3984[(2'h3):(1'h1)];
                      reg4043 <= (~|$unsigned(reg4030));
                    end
                  for (forvar4044 = (1'h0); (forvar4044 < (2'h2)); forvar4044 = (forvar4044 + (1'h1)))
                    begin
                      reg4045 <= $unsigned((-(~forvar3992[(3'h6):(1'h0)])));
                    end
                end
              if ({{(((8'h9e) ? reg3962 : (8'h9f)) >> reg4018)}})
                begin
                  reg4046 <= ({$signed($signed(forvar3971))} <<< (forvar3992 * ((^wire3940) ?
                      (|reg3954) : {reg4019})));
                  reg4047 <= reg4045[(2'h3):(1'h1)];
                  for (forvar4048 = (1'h0); (forvar4048 < (1'h0)); forvar4048 = (forvar4048 + (1'h1)))
                    begin
                      reg4049 <= (8'ha3);
                      reg4050 <= $signed((~^($signed(reg3946) ?
                          $unsigned(forvar3943) : forvar4011[(2'h2):(1'h0)])));
                      reg4051 <= $unsigned(reg4005[(1'h0):(1'h0)]);
                    end
                  if ($unsigned($unsigned((^~(&(8'hb7))))))
                    begin
                      reg4052 <= $unsigned(forvar3960);
                      reg4053 <= (($signed(((8'h9e) == reg3965)) < (|{forvar3943})) == (~forvar3989[(1'h1):(1'h1)]));
                      reg4054 <= (~|({(~&forvar4001)} ?
                          ($unsigned((8'h9f)) ?
                              (reg4024 >>> (8'ha8)) : (reg4000 ?
                                  reg4034 : reg4023)) : {(reg3974 <= forvar4038)}));
                    end
                  else
                    begin
                      reg4052 <= reg3967[(4'h8):(3'h4)];
                      reg4053 <= (8'hb4);
                      reg4054 <= $unsigned(reg3973);
                    end
                end
              else
                begin
                  reg4046 <= (|(8'h9f));
                  if ((|(&$signed({reg3977}))))
                    begin
                      reg4047 <= $unsigned((^forvar3968[(3'h7):(2'h3)]));
                      reg4048 <= $signed(($signed((|reg3944)) ?
                          $unsigned(((8'ha9) ?
                              forvar3975 : reg3961)) : reg3964[(2'h3):(1'h0)]));
                      reg4049 <= $unsigned(forvar3995[(3'h7):(1'h0)]);
                    end
                  else
                    begin
                      reg4047 <= reg4049;
                      reg4048 <= {$unsigned((8'hab))};
                    end
                  reg4050 <= $signed(reg3980);
                end
            end
          for (forvar4055 = (1'h0); (forvar4055 < (1'h1)); forvar4055 = (forvar4055 + (1'h1)))
            begin
              if (reg3961)
                begin
                  if ($signed({$unsigned(forvar3959[(4'ha):(3'h6)])}))
                    begin
                      reg4056 <= (~&{((|forvar4033) ?
                              ((8'ha1) | forvar3973) : $unsigned(reg3955))});
                      reg4057 <= (^~(($unsigned(reg3976) - (+wire3940)) >= $unsigned($unsigned(reg4036))));
                      reg4058 <= (+($unsigned($signed(forvar3957)) ?
                          ((reg3954 >= reg3983) ?
                              (reg3973 != reg3983) : wire3937) : $signed((reg4024 ?
                              reg3939 : reg4040))));
                      reg4059 <= (($unsigned({forvar3973}) ?
                          (forvar4012 ?
                              (reg3939 ?
                                  forvar4017 : reg4019) : (!forvar3957)) : $unsigned(reg4002[(3'h4):(1'h1)])) - $signed($signed((~|reg3979))));
                    end
                  else
                    begin
                      reg4056 <= reg4022[(3'h7):(3'h7)];
                      reg4057 <= $unsigned($unsigned(reg3949[(1'h1):(1'h1)]));
                    end
                  for (forvar4060 = (1'h0); (forvar4060 < (2'h2)); forvar4060 = (forvar4060 + (1'h1)))
                    begin
                      reg4061 <= (^~reg4003[(2'h3):(2'h3)]);
                      reg4062 <= (reg3977 ?
                          (~&reg3993[(3'h7):(1'h1)]) : (reg3999[(2'h3):(1'h1)] ?
                              reg4061 : ((reg3990 ?
                                  reg4023 : reg4056) > (8'hb9))));
                    end
                  reg4063 <= $unsigned((&($signed(forvar4028) <= $unsigned(reg3978))));
                  for (forvar4064 = (1'h0); (forvar4064 < (2'h2)); forvar4064 = (forvar4064 + (1'h1)))
                    begin
                      reg4065 <= {forvar4006};
                      reg4066 <= reg3993;
                    end
                end
              else
                begin
                  if ((reg4002 - reg4037))
                    begin
                      reg4056 <= {(~reg4009)};
                    end
                  else
                    begin
                      reg4056 <= $signed(reg4002[(3'h7):(1'h1)]);
                      reg4057 <= (!(~|$signed((reg3974 ?
                          forvar4041 : reg3956))));
                      reg4058 <= (~|(reg4048[(4'h8):(2'h2)] ?
                          $signed((reg3980 >>> (8'h9e))) : ((reg4016 ?
                              reg4004 : forvar4041) < forvar3977)));
                      reg4059 <= (reg3979[(4'h9):(1'h1)] ?
                          (reg3983[(1'h1):(1'h0)] & $signed(reg4005)) : ($signed((reg4031 != reg4024)) ?
                              (^reg3980[(1'h1):(1'h1)]) : $signed((~|reg3991))));
                    end
                  for (forvar4060 = (1'h0); (forvar4060 < (2'h2)); forvar4060 = (forvar4060 + (1'h1)))
                    begin
                      reg4061 <= reg3955;
                      reg4062 <= reg3943[(2'h3):(2'h2)];
                      reg4063 <= (~&($unsigned($signed(forvar4038)) ?
                          forvar3992[(4'h9):(4'h8)] : ($unsigned(reg4037) ?
                              (+forvar3943) : (~^forvar3959))));
                    end
                  reg4064 <= reg4023[(4'h8):(3'h7)];
                  reg4065 <= ({($unsigned((8'ha7)) ?
                          reg3967[(3'h4):(2'h3)] : forvar3945[(1'h1):(1'h0)])} <= $signed(((reg4047 ?
                      wire3936 : (8'hb1)) << reg4036[(1'h1):(1'h1)])));
                end
              if (({$unsigned({forvar4001})} ? reg4058 : {reg4052}))
                begin
                  for (forvar4067 = (1'h0); (forvar4067 < (1'h1)); forvar4067 = (forvar4067 + (1'h1)))
                    begin
                      reg4068 <= ($signed($signed(reg3957)) ?
                          ($signed((+reg4013)) ?
                              (forvar4067 > $unsigned(reg4053)) : {(forvar3952 & reg3971)}) : forvar3981[(1'h0):(1'h0)]);
                      reg4069 <= ({$unsigned((&forvar4060))} * reg3961[(2'h2):(1'h1)]);
                      reg4070 <= (8'ha3);
                      reg4071 <= ((+$signed(forvar4023[(1'h1):(1'h0)])) > (((reg4023 == reg4026) ?
                          {reg3953} : (~^forvar4022)) > $unsigned($signed(forvar4017))));
                    end
                  for (forvar4072 = (1'h0); (forvar4072 < (2'h2)); forvar4072 = (forvar4072 + (1'h1)))
                    begin
                      reg4073 <= $signed((reg4002[(4'hb):(4'hb)] << (reg3947[(2'h3):(2'h2)] >> reg4018)));
                      reg4074 <= wire3932;
                      reg4075 <= $signed($signed((forvar3957[(2'h2):(1'h0)] * reg4013)));
                      reg4076 <= $signed((((reg4065 * forvar4012) ?
                          (reg4015 > reg3987) : reg3949[(2'h3):(1'h1)]) * (reg3991[(3'h6):(2'h3)] <= $signed(reg3947))));
                    end
                end
              else
                begin
                  for (forvar4067 = (1'h0); (forvar4067 < (2'h2)); forvar4067 = (forvar4067 + (1'h1)))
                    begin
                      reg4068 <= forvar4010[(2'h3):(2'h2)];
                      reg4069 <= {$unsigned(reg3971[(3'h4):(2'h2)])};
                    end
                end
              for (forvar4077 = (1'h0); (forvar4077 < (1'h1)); forvar4077 = (forvar4077 + (1'h1)))
                begin
                  if (((!((-reg4048) ? {forvar3941} : (~&forvar3941))) ?
                      reg4028 : reg4057))
                    begin
                      reg4078 <= ((!(forvar3952[(2'h2):(2'h2)] ^~ (reg3983 ?
                          reg4063 : reg4026))) != reg4021);
                    end
                  else
                    begin
                      reg4078 <= (($unsigned($unsigned(reg3955)) | ((~&(8'hb9)) ?
                          reg3944[(4'hc):(1'h1)] : $unsigned(forvar3986))) <<< ($signed($signed((8'ha3))) ?
                          reg3947[(2'h3):(1'h1)] : ($signed(reg4047) - (reg4018 | reg3975))));
                      reg4079 <= $unsigned(forvar4064[(4'h9):(3'h4)]);
                    end
                end
            end
        end
      reg4080 <= $signed(({(~^reg4022)} >>> reg3973[(4'h8):(4'h8)]));
    end
  always
    @(posedge clk) begin
      if ((8'hb6))
        begin
          reg4081 <= (-$signed(reg3983));
          for (forvar4082 = (1'h0); (forvar4082 < (2'h2)); forvar4082 = (forvar4082 + (1'h1)))
            begin
              for (forvar4083 = (1'h0); (forvar4083 < (2'h3)); forvar4083 = (forvar4083 + (1'h1)))
                begin
                  if (((reg3996[(3'h4):(3'h4)] | {forvar4067}) ?
                      forvar4012 : reg4061))
                    begin
                      reg4084 <= reg4053[(3'h7):(3'h4)];
                    end
                  else
                    begin
                      reg4084 <= (forvar4032 ?
                          $signed((^~$unsigned(forvar4039))) : forvar4001[(1'h0):(1'h0)]);
                    end
                  if ($unsigned((reg4029 ?
                      ((8'hb2) ?
                          reg4000 : forvar4072[(2'h2):(1'h0)]) : $unsigned((wire3935 ?
                          reg3962 : wire3936)))))
                    begin
                      reg4085 <= ((^~reg4043) ?
                          ($signed($signed(reg4036)) ?
                              reg4066[(3'h4):(2'h3)] : (|(|reg3963))) : reg4076[(4'ha):(4'h9)]);
                      reg4086 <= (^{({(8'ha3)} ?
                              $unsigned(forvar4048) : (~|forvar4012))});
                      reg4087 <= ($signed((-(~|reg4048))) ?
                          ((reg3983 ?
                                  $unsigned(reg3973) : reg4042[(2'h3):(1'h1)]) ?
                              reg3999 : (^~$signed(reg3972))) : {((reg3991 == reg4046) && $signed(wire3934))});
                      reg4088 <= reg4081;
                    end
                  else
                    begin
                      reg4085 <= {$signed(((!reg4070) ?
                              $signed(forvar3971) : $unsigned(forvar4026)))};
                    end
                  for (forvar4089 = (1'h0); (forvar4089 < (1'h1)); forvar4089 = (forvar4089 + (1'h1)))
                    begin
                      reg4090 <= $unsigned((reg4009 ?
                          reg3952[(4'hc):(2'h3)] : (~&forvar3968)));
                      reg4091 <= (&reg4075[(1'h1):(1'h0)]);
                      reg4092 <= (+(~^reg4025));
                    end
                end
              for (forvar4093 = (1'h0); (forvar4093 < (1'h1)); forvar4093 = (forvar4093 + (1'h1)))
                begin
                  for (forvar4094 = (1'h0); (forvar4094 < (1'h1)); forvar4094 = (forvar4094 + (1'h1)))
                    begin
                      reg4095 <= $signed($unsigned($signed($unsigned((8'ha4)))));
                    end
                end
            end
          for (forvar4096 = (1'h0); (forvar4096 < (2'h3)); forvar4096 = (forvar4096 + (1'h1)))
            begin
              for (forvar4097 = (1'h0); (forvar4097 < (1'h0)); forvar4097 = (forvar4097 + (1'h1)))
                begin
                  reg4098 <= forvar3945[(4'h9):(4'h8)];
                end
            end
          reg4099 <= ((~^reg3996[(3'h5):(1'h0)]) ? reg4065 : (8'ha6));
        end
      else
        begin
          if (($unsigned(reg4028[(1'h1):(1'h1)]) ?
              $signed(forvar3975) : (~((reg3984 + forvar3968) << (reg4068 ^~ reg4050)))))
            begin
              if ((~^(reg3973 ? {$signed((8'ha6))} : forvar4006)))
                begin
                  for (forvar4081 = (1'h0); (forvar4081 < (2'h2)); forvar4081 = (forvar4081 + (1'h1)))
                    begin
                      reg4082 <= $unsigned(reg4074);
                      reg4083 <= {(((reg3991 && (8'hab)) + (reg4003 ?
                              (8'haf) : reg3993)) ^ reg4079[(4'ha):(1'h0)])};
                      reg4084 <= forvar3941[(2'h3):(1'h0)];
                      reg4085 <= reg4059[(4'ha):(3'h5)];
                    end
                  if (reg3972[(3'h5):(2'h2)])
                    begin
                      reg4086 <= forvar4089;
                      reg4087 <= $unsigned((reg4073[(3'h5):(1'h1)] ?
                          ({forvar4026} ?
                              (forvar4082 ?
                                  reg3946 : reg4036) : ((8'ha8) < reg4058)) : ((!reg3983) ?
                              (8'ha8) : $signed(reg3998))));
                      reg4088 <= (+reg3947[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg4086 <= $unsigned((+((reg4058 == (8'hb3)) ?
                          (reg4013 ? reg4065 : reg4070) : (~|reg4046))));
                      reg4087 <= $unsigned(reg4076[(4'he):(4'h9)]);
                    end
                  if ((~^(~|(+(+reg4063)))))
                    begin
                      reg4089 <= (-(forvar4011 && (^~(reg3952 ?
                          reg4076 : forvar4077))));
                      reg4090 <= forvar3941[(4'h9):(1'h1)];
                    end
                  else
                    begin
                      reg4089 <= $signed($signed(reg3950[(4'ha):(3'h6)]));
                      reg4090 <= (~reg3969);
                    end
                  for (forvar4091 = (1'h0); (forvar4091 < (2'h2)); forvar4091 = (forvar4091 + (1'h1)))
                    begin
                      reg4092 <= ($signed({(~^reg3994)}) ?
                          $signed((reg3962 ?
                              reg4009 : $signed(reg3970))) : $unsigned($signed(reg4083)));
                    end
                end
              else
                begin
                  for (forvar4081 = (1'h0); (forvar4081 < (2'h3)); forvar4081 = (forvar4081 + (1'h1)))
                    begin
                      reg4082 <= $signed($signed($signed((^reg4046))));
                      reg4083 <= (reg4091 && {forvar4033[(4'h8):(3'h4)]});
                      reg4084 <= ($unsigned(forvar4044) ?
                          $unsigned(forvar4029[(3'h4):(1'h1)]) : (reg4009 ?
                              $unsigned((~&(8'hb8))) : {$unsigned(reg4013)}));
                    end
                end
              reg4093 <= $signed({{(forvar4038 >= reg4009)}});
              for (forvar4094 = (1'h0); (forvar4094 < (2'h2)); forvar4094 = (forvar4094 + (1'h1)))
                begin
                  for (forvar4095 = (1'h0); (forvar4095 < (1'h1)); forvar4095 = (forvar4095 + (1'h1)))
                    begin
                      reg4096 <= {forvar4048};
                      reg4097 <= ($signed(({forvar4017} ?
                              $signed(forvar4083) : (reg4089 >> reg3957))) ?
                          (8'hb0) : reg4009[(1'h1):(1'h0)]);
                      reg4098 <= $unsigned((~($unsigned(reg4075) ?
                          (forvar3959 ? reg4013 : reg4049) : {forvar3975})));
                      reg4099 <= (|$unsigned(((~&reg4088) ?
                          $unsigned(reg4063) : {reg4068})));
                    end
                end
              reg4100 <= ($unsigned(((^~reg4061) ?
                  reg4058[(4'hc):(4'h8)] : reg3961)) ^~ reg4049);
            end
          else
            begin
              if ($unsigned(((8'h9e) >>> $signed((forvar3941 ?
                  forvar4029 : reg4020)))))
                begin
                  for (forvar4081 = (1'h0); (forvar4081 < (2'h2)); forvar4081 = (forvar4081 + (1'h1)))
                    begin
                      reg4082 <= (8'hb8);
                      reg4083 <= reg3987[(1'h0):(1'h0)];
                      reg4084 <= {(reg4054[(3'h6):(3'h4)] << forvar4097)};
                      reg4085 <= ((8'ha0) | forvar3968[(3'h5):(3'h5)]);
                    end
                end
              else
                begin
                  if (((({reg4081} && reg4068) | (~reg3954)) < $signed(((8'hab) == reg3958))))
                    begin
                      reg4081 <= (forvar4023[(1'h0):(1'h0)] ?
                          $unsigned(reg3954) : (forvar4055 ?
                              ($signed(forvar4022) > $signed(reg3961)) : {(reg4074 ?
                                      reg3963 : (8'h9e))}));
                      reg4082 <= wire3933[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg4081 <= $unsigned($signed((8'ha5)));
                      reg4082 <= forvar4095[(3'h5):(3'h5)];
                      reg4083 <= $signed(reg3964[(3'h7):(3'h5)]);
                    end
                  if (reg4004[(2'h3):(1'h0)])
                    begin
                      reg4084 <= reg4004[(3'h4):(1'h0)];
                      reg4085 <= reg3955[(4'ha):(2'h2)];
                    end
                  else
                    begin
                      reg4084 <= (reg4016[(3'h5):(2'h3)] ?
                          reg3947 : $signed((-(~reg4015))));
                      reg4085 <= forvar4033[(2'h2):(1'h1)];
                      reg4086 <= reg3947;
                      reg4087 <= reg4085;
                    end
                  if ($unsigned($signed(reg3996)))
                    begin
                      reg4088 <= (!reg4009[(4'hb):(4'ha)]);
                      reg4089 <= $signed((~|$unsigned($unsigned((8'hb3)))));
                    end
                  else
                    begin
                      reg4088 <= reg3955[(1'h0):(1'h0)];
                      reg4089 <= (~|$unsigned(wire3933));
                      reg4090 <= wire3935[(1'h1):(1'h0)];
                      reg4091 <= reg4089[(1'h1):(1'h0)];
                    end
                end
              for (forvar4092 = (1'h0); (forvar4092 < (1'h1)); forvar4092 = (forvar4092 + (1'h1)))
                begin
                  for (forvar4093 = (1'h0); (forvar4093 < (2'h3)); forvar4093 = (forvar4093 + (1'h1)))
                    begin
                      reg4094 <= $signed($unsigned((+reg4097[(1'h0):(1'h0)])));
                      reg4095 <= $signed(((!(reg3961 ? reg4052 : reg3975)) ?
                          reg4016[(3'h6):(3'h4)] : ((!reg3971) >> (reg3955 ?
                              reg3976 : (8'hb9)))));
                      reg4096 <= ($signed(wire3933[(4'hd):(4'ha)]) ?
                          $unsigned(reg4009[(3'h5):(1'h0)]) : reg4052[(4'hc):(3'h7)]);
                      reg4097 <= reg4099;
                    end
                  for (forvar4098 = (1'h0); (forvar4098 < (1'h0)); forvar4098 = (forvar4098 + (1'h1)))
                    begin
                      reg4099 <= reg4090[(4'hd):(2'h2)];
                      reg4100 <= (8'hab);
                    end
                  reg4101 <= {{((^forvar3960) ? reg4085 : (!reg4047))}};
                  for (forvar4102 = (1'h0); (forvar4102 < (2'h3)); forvar4102 = (forvar4102 + (1'h1)))
                    begin
                      reg4103 <= (8'ha8);
                    end
                end
              for (forvar4104 = (1'h0); (forvar4104 < (1'h1)); forvar4104 = (forvar4104 + (1'h1)))
                begin
                  for (forvar4105 = (1'h0); (forvar4105 < (2'h2)); forvar4105 = (forvar4105 + (1'h1)))
                    begin
                      reg4106 <= reg4016[(2'h3):(2'h2)];
                      reg4107 <= $unsigned($signed({$signed(reg3943)}));
                    end
                end
              for (forvar4108 = (1'h0); (forvar4108 < (1'h0)); forvar4108 = (forvar4108 + (1'h1)))
                begin
                  for (forvar4109 = (1'h0); (forvar4109 < (2'h2)); forvar4109 = (forvar4109 + (1'h1)))
                    begin
                      reg4110 <= $signed({$signed(forvar4055)});
                    end
                  if (((~^(8'hab)) ?
                      (~|forvar4010[(2'h3):(1'h1)]) : $signed((8'ha1))))
                    begin
                      reg4111 <= reg4016;
                      reg4112 <= (^reg3998[(3'h4):(2'h3)]);
                      reg4113 <= wire3932;
                    end
                  else
                    begin
                      reg4111 <= {$signed({reg4015})};
                      reg4112 <= reg4059;
                      reg4113 <= {reg3991[(1'h0):(1'h0)]};
                    end
                end
            end
          for (forvar4114 = (1'h0); (forvar4114 < (2'h3)); forvar4114 = (forvar4114 + (1'h1)))
            begin
              for (forvar4115 = (1'h0); (forvar4115 < (1'h1)); forvar4115 = (forvar4115 + (1'h1)))
                begin
                  for (forvar4116 = (1'h0); (forvar4116 < (2'h3)); forvar4116 = (forvar4116 + (1'h1)))
                    begin
                      reg4117 <= (((-$unsigned(reg4029)) & {(forvar4089 ?
                                  reg3952 : reg4113)}) ?
                          {reg4025} : forvar4044);
                      reg4118 <= $unsigned(((^$signed(forvar3941)) ?
                          (~|reg3949[(4'ha):(1'h1)]) : forvar4104[(3'h5):(3'h5)]));
                      reg4119 <= (^reg4084[(1'h0):(1'h0)]);
                    end
                end
            end
          if ($unsigned(reg3939[(2'h2):(1'h1)]))
            begin
              for (forvar4120 = (1'h0); (forvar4120 < (2'h2)); forvar4120 = (forvar4120 + (1'h1)))
                begin
                  if ($unsigned($unsigned(reg4052[(5'h10):(4'he)])))
                    begin
                      reg4121 <= (reg4005 ?
                          (8'haf) : ($signed((forvar3959 == reg4056)) || (|(forvar4083 != reg4019))));
                    end
                  else
                    begin
                      reg4121 <= reg3990;
                      reg4122 <= reg3961;
                      reg4123 <= $unsigned((8'h9e));
                      reg4124 <= ((~|((reg4101 * reg3971) || (forvar3992 == forvar3960))) ^~ (8'hb3));
                    end
                  if (reg3954)
                    begin
                      reg4125 <= $signed((^~{forvar3986[(4'hc):(1'h1)]}));
                    end
                  else
                    begin
                      reg4125 <= (reg4089 || reg4119);
                      reg4126 <= reg3967[(3'h4):(3'h4)];
                      reg4127 <= reg4079[(3'h6):(3'h4)];
                    end
                  if ($signed($unsigned({(~^reg3972)})))
                    begin
                      reg4128 <= {(reg4034[(1'h0):(1'h0)] <<< (-reg4027))};
                      reg4129 <= (8'ha5);
                      reg4130 <= (8'hab);
                      reg4131 <= (~|reg4020[(4'hd):(4'hb)]);
                    end
                  else
                    begin
                      reg4128 <= $unsigned(($unsigned($signed((8'hb0))) == reg4005[(4'h8):(3'h7)]));
                      reg4129 <= ((^{wire3937[(2'h3):(1'h0)]}) ?
                          $unsigned((~(~&reg4078))) : $signed($signed($unsigned(wire3937))));
                      reg4130 <= $signed(forvar4102);
                    end
                end
              reg4132 <= forvar4022;
            end
          else
            begin
              reg4120 <= $unsigned((8'hb4));
              reg4121 <= $signed((($signed((8'ha5)) ?
                  $unsigned(reg4013) : $signed(reg4093)) ~^ $signed(forvar3985[(2'h2):(1'h0)])));
              for (forvar4122 = (1'h0); (forvar4122 < (1'h1)); forvar4122 = (forvar4122 + (1'h1)))
                begin
                  for (forvar4123 = (1'h0); (forvar4123 < (2'h3)); forvar4123 = (forvar4123 + (1'h1)))
                    begin
                      reg4124 <= ($unsigned(forvar4120[(3'h5):(3'h4)]) ?
                          ((reg3964[(3'h6):(3'h5)] * (|reg3946)) ?
                              ((+reg4075) << reg4022) : ((reg3991 ?
                                  reg3947 : reg4078) > forvar3968[(4'hd):(1'h1)])) : (forvar4017[(4'h8):(3'h6)] ?
                              reg4118[(4'hc):(2'h2)] : forvar4029[(1'h1):(1'h1)]));
                      reg4125 <= ((+(forvar4026[(1'h0):(1'h0)] ?
                              (reg4098 ?
                                  reg4031 : forvar4120) : reg4016[(1'h1):(1'h1)])) ?
                          $unsigned((8'hb4)) : $signed($unsigned((reg4107 ?
                              reg4113 : reg4128))));
                      reg4126 <= $signed(forvar4072);
                    end
                  for (forvar4127 = (1'h0); (forvar4127 < (1'h0)); forvar4127 = (forvar4127 + (1'h1)))
                    begin
                      reg4128 <= (reg3955 ?
                          ({(8'hb9)} << ((reg3976 ?
                              reg4126 : reg4013) & forvar4010[(2'h2):(1'h1)])) : ((~^((8'hb1) | reg4092)) ?
                              forvar4108 : (reg3965[(4'he):(4'hd)] ?
                                  (-(8'hb7)) : $signed(reg3984))));
                      reg4129 <= ((reg4126 ?
                          reg4037 : reg3956) <= (forvar4048[(3'h6):(3'h5)] && ($signed(forvar3945) ?
                          reg4128 : {reg4025})));
                      reg4130 <= (~|forvar4127);
                    end
                  for (forvar4131 = (1'h0); (forvar4131 < (2'h3)); forvar4131 = (forvar4131 + (1'h1)))
                    begin
                      reg4132 <= forvar3973[(4'h8):(2'h2)];
                      reg4133 <= ((8'h9c) ?
                          reg3998[(3'h4):(1'h1)] : (((reg4106 >>> reg4054) ?
                                  wire3935[(1'h1):(1'h0)] : (reg3950 > reg3983)) ?
                              (!forvar4114) : {reg4113[(2'h2):(1'h1)]}));
                      reg4134 <= (forvar4011[(3'h4):(2'h3)] ?
                          ($unsigned($signed(reg3980)) - forvar4115[(1'h1):(1'h0)]) : $signed(((8'hba) && (~(8'hb9)))));
                      reg4135 <= $signed((~|$signed(reg3944)));
                    end
                end
              for (forvar4136 = (1'h0); (forvar4136 < (1'h0)); forvar4136 = (forvar4136 + (1'h1)))
                begin
                  if ({(reg4122[(3'h4):(2'h3)] ?
                          reg4084 : $unsigned(forvar4032[(3'h7):(1'h0)]))})
                    begin
                      reg4137 <= (|(8'h9e));
                    end
                  else
                    begin
                      reg4137 <= $unsigned(reg4123[(2'h3):(2'h2)]);
                      reg4138 <= {($signed($unsigned((8'ha0))) + (((8'ha2) >> forvar4096) | $signed(forvar4098)))};
                    end
                end
            end
          for (forvar4139 = (1'h0); (forvar4139 < (1'h1)); forvar4139 = (forvar4139 + (1'h1)))
            begin
              for (forvar4140 = (1'h0); (forvar4140 < (2'h3)); forvar4140 = (forvar4140 + (1'h1)))
                begin
                  for (forvar4141 = (1'h0); (forvar4141 < (1'h1)); forvar4141 = (forvar4141 + (1'h1)))
                    begin
                      reg4142 <= reg4078[(1'h0):(1'h0)];
                      reg4143 <= reg3994[(2'h2):(2'h2)];
                      reg4144 <= (forvar3971[(4'hc):(4'h9)] ?
                          $signed({forvar4023}) : {forvar3957[(3'h5):(2'h3)]});
                    end
                end
              reg4145 <= (~&((reg4059 * reg4129) ?
                  $signed(((8'hb1) ? reg4014 : forvar4001)) : reg3996));
              reg4146 <= (reg4066[(2'h3):(2'h3)] ?
                  (!(forvar3968[(4'h9):(4'h9)] ?
                      reg4074 : (8'hac))) : (&($signed(reg4085) ^ {reg4080})));
              for (forvar4147 = (1'h0); (forvar4147 < (2'h2)); forvar4147 = (forvar4147 + (1'h1)))
                begin
                  reg4148 <= ((-(~|$unsigned(reg3990))) ~^ ((reg3979[(4'ha):(2'h2)] + $unsigned(reg3999)) < $unsigned((reg3950 != reg4133))));
                end
            end
        end
    end
  assign wire4149 = forvar3968;
  assign wire4150 = ($unsigned((-forvar4048)) ?
                        (&($unsigned(forvar4114) ?
                            reg4051[(3'h5):(2'h3)] : (reg4048 ?
                                reg4037 : (8'hae)))) : {forvar4092});
  assign wire4151 = ($unsigned(reg3996[(2'h2):(2'h2)]) | (((~&reg4094) ?
                        reg4143[(3'h4):(2'h3)] : reg4124) == reg3988[(3'h5):(2'h3)]));
  assign wire4152 = (((|{reg3943}) > (-forvar4089[(3'h6):(1'h0)])) - (^~(&(reg3938 * forvar4127))));
endmodule