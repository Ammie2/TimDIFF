(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [32'b00000000000000000000001001101111:32'b00000000000000000000000000000000] y;
  input wire [1'b10:1'b10] clk;
  input wire [4'b10101110:1'b10] wire0;
  input wire [5'b0001110101:1'b00] wire1;
  input wire signed [5'b0001110101:1'b00] wire2;
  input wire [5'b1111010100:1'b00] wire3;
  reg [5'b0101010011:1'b10] reg324 = (1'h0);
  reg [4'b10101110:1'b10] reg323 = (1'h0);
  reg [2'b1011:1'b00] reg322 = (1'h0);
  reg [4'b11111000:1'b00] reg321 = (1'h0);
  reg [2'b1011:1'b00] reg320 = (1'h0);
  wire [4'b00101011:1'b00] wire273;
  wire [5'b1000110000:1'b0] wire4;
  wire signed [5'b0001110101:1'b00] wire74;
  wire [4'b01001111:1'b10] wire271;
  wire signed [5'b1111010100:1'b00] wire275;
  reg signed [5'b1111010100:1'b00] reg276 = (1'h0);
  reg signed [2'b1011:1'b00] reg277 = (1'h0);
  reg signed [3'b000101:1'b00] reg278 = (1'h0);
  reg [4'b00101011:1'b00] reg279 = (1'h0);
  reg signed [5'b0001110101:1'b00] reg280 = (1'h0);
  reg [5'b1110001:1'b10] reg281 = (1'h0);
  reg signed [3'b001111:1'b00] reg282 = (1'h0);
  reg [5'b1110001:1'b10] reg283 = (1'h0);
  reg signed [4'b11111000:1'b00] reg284 = (1'h0);
  reg [4'b11011001:1'b10] reg285 = (1'h0);
  reg signed [5'b0001010010:1'b10] reg286 = (1'h0);
  reg [3'b001111:1'b00] reg287 = (1'h0);
  reg signed [4'b11111000:1'b00] reg288 = (1'h0);
  reg [5'b1110001:1'b10] reg289 = (1'h0);
  reg signed [4'b10001101:1'b10] reg290 = (1'h0);
  reg signed [5'b0001110101:1'b00] reg291 = (1'h0);
  reg signed [5'b1110001:1'b10] reg292 = (1'h0);
  reg [3'b000101:1'b00] reg293 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg294 = (1'h0);
  reg signed [3'b000110:1'b00] reg295 = (1'h0);
  reg signed [5'b0001010010:1'b10] reg296 = (1'h0);
  reg signed [2'b010:1'b10] reg297 = (1'h0);
  reg [4'b00101011:1'b00] reg298 = (1'h0);
  reg signed [4'b11011001:1'b10] reg299 = (1'h0);
  reg [5'b1110001:1'b10] reg300 = (1'h0);
  reg [5'b1111010100:1'b00] reg301 = (1'h0);
  reg [4'b10001101:1'b10] reg302 = (1'h0);
  reg [3'b000110:1'b00] reg303 = (1'h0);
  reg [4'b10001101:1'b10] reg304 = (1'h0);
  reg [5'b0001110101:1'b00] reg305 = (1'h0);
  reg [2'b010:1'b10] reg306 = (1'h0);
  reg signed [2'b1011:1'b00] reg307 = (1'h0);
  reg [4'b00101011:1'b00] reg308 = (1'h0);
  reg [3'b001111:1'b00] reg309 = (1'h0);
  reg signed [5'b1110001:1'b10] reg310 = (1'h0);
  wire signed [4'b10101110:1'b10] wire311;
  wire signed [3'b000110:1'b00] wire312;
  wire [5'b1000110000:1'b0] wire313;
  wire signed [2'b010:1'b10] wire314;
  wire signed [5'b0101010011:1'b10] wire315;
  wire signed [2'b010:1'b10] wire316;
  wire signed [4'b00101011:1'b00] wire317;
  wire [2'b1011:1'b00] wire318;
  assign y = {reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 wire273,
                 wire4,
                 wire74,
                 wire271,
                 wire275,
                 reg276,
                 reg277,
                 reg278,
                 reg279,
                 reg280,
                 reg281,
                 reg282,
                 reg283,
                 reg284,
                 reg285,
                 reg286,
                 reg287,
                 reg288,
                 reg289,
                 reg290,
                 reg291,
                 reg292,
                 reg293,
                 reg294,
                 reg295,
                 reg296,
                 reg297,
                 reg298,
                 reg299,
                 reg300,
                 reg301,
                 reg302,
                 reg303,
                 reg304,
                 reg305,
                 reg306,
                 reg307,
                 reg308,
                 reg309,
                 reg310,
                 wire311,
                 wire312,
                 wire313,
                 wire314,
                 wire315,
                 wire316,
                 wire317,
                 wire318,
                 (1'h0)};
  assign wire4 = (^~wire0);
  module5 modinst75 (wire74, clk, wire2, wire3, wire1, wire0);
  module76 modinst272 (wire271, clk, wire3, wire0, wire2, wire74, wire4);
  module76 modinst274 (.wire80(wire271), .wire81(wire2), .wire78(wire1), .wire79(wire74), .clk(clk), .wire77(wire4), .y(wire273));
  assign wire275 = ((wire273 ?
                       (!wire74) : (+(~^((8'ha7) >>> wire2)))) ~^ (-wire271));
  always
    @(posedge clk) begin
      if (($unsigned(wire0) ^~ wire275))
        begin
          reg276 <= (~(($unsigned((!(8'ha7))) >= $signed((wire0 != wire275))) >= $unsigned((8'hb9))));
          reg277 <= $unsigned($unsigned(((^wire2) ~^ wire3)));
          reg278 <= wire2;
          reg279 <= ($signed((8'hb5)) ^ (wire0 <= $signed(({reg278} ~^ $unsigned(reg276)))));
        end
      else
        begin
          if ((wire275 && (wire0 ?
              (~wire3) : $unsigned(wire275[3'b101110:3'b011110]))))
            begin
              reg276 <= reg279[1'b11:1'b00];
              reg277 <= $signed($unsigned($unsigned({wire0[4'b10111101:4'b00001011],
                  ((8'hbf) | wire0)})));
              reg278 <= wire2;
            end
          else
            begin
              reg276 <= ((~(reg277 ?
                  $signed({reg278, reg276}) : ((wire74 ?
                      (8'ha2) : reg278) <= (wire275 + (8'hb3))))) + $unsigned({((wire275 <<< reg277) == wire3),
                  (wire4 << {(7'h41)})}));
            end
          if (wire2[1'b01:1'b11])
            begin
              reg279 <= $signed($signed(((wire275 ? wire0 : $signed(reg276)) ?
                  wire3[3'b000101:2'b0111] : $signed(wire2))));
              reg280 <= wire74;
              reg281 <= (&($unsigned($unsigned(wire271[2'b1111:1'b11])) && $unsigned(reg276[1'b10:1'b10])));
              reg282 <= $unsigned(((reg281[2'b1011:1'b00] ?
                      wire4 : (^(reg279 ~^ wire1))) ?
                  $signed(wire1[3'b101110:3'b011110]) : {(~&(~reg279)),
                      $signed($signed(wire0))}));
              reg283 <= (~|reg282[2'b0111:2'b10]);
            end
          else
            begin
              reg279 <= {$unsigned($unsigned($signed(wire4))),
                  $unsigned($signed(((8'h9c) ?
                      ((8'hb2) ? wire74 : wire271) : reg281)))};
              reg280 <= (!wire273);
              reg281 <= $unsigned({$unsigned(((wire74 == (8'hbc)) * (8'haf)))});
              reg282 <= $unsigned(reg278);
            end
          reg284 <= wire74;
          if (($signed((!wire74[2'b1110:2'b0110])) ?
              (|($signed((reg282 ^~ reg279)) ?
                  reg283[2'b010:1'b10] : $unsigned(wire2[1'b10:1'b10]))) : {($unsigned(wire271) ?
                      $unsigned($signed(wire74)) : $unsigned($signed(wire3))),
                  (~(^{wire275}))}))
            begin
              reg285 <= ((-wire0[3'b000101:1'b00]) >> (reg282[1'b01:1'b11] ?
                  $signed(reg283[4'b00001101:4'b00101100]) : $signed((wire74[4'b11001011:4'b10101011] + (reg279 - wire0)))));
            end
          else
            begin
              reg285 <= $signed(((^~wire3) >> $unsigned(reg276)));
            end
          reg286 <= {($unsigned((8'ha5)) ~^ $unsigned(reg282[1'b11:1'b00])),
              {wire74[1'b01:1'b11]}};
        end
      if ($signed(reg285))
        begin
          if (reg284[2'b1110:2'b0110])
            begin
              reg287 <= (~wire0);
              reg288 <= $signed($unsigned($signed(reg283)));
            end
          else
            begin
              reg287 <= (8'h9c);
              reg288 <= reg277;
              reg289 <= ((reg281 < (~&{reg282[3'b001100:3'b001100], (~reg285)})) ?
                  wire4[4'b00111111:4'b00011101] : wire1[3'b110101:1'b11]);
            end
        end
      else
        begin
          if ((wire3 >= wire273))
            begin
              reg287 <= (~|$signed((wire2 ?
                  (~|$unsigned(reg279)) : (reg277 < (~|reg278)))));
              reg288 <= (&reg281[3'b000101:2'b0111]);
              reg289 <= $signed((($signed((wire74 ? wire1 : reg287)) ?
                      ($unsigned(wire1) ?
                          (wire2 < reg285) : ((8'hbf) ?
                              wire1 : (8'hb9))) : ((&wire2) - (wire2 != reg278))) ?
                  (wire273[4'b10111000:3'b011101] >> ((^reg280) ?
                      $unsigned(wire4) : (reg282 < reg277))) : ((8'haa) ?
                      $signed($unsigned((8'h9c))) : $unsigned({reg277}))));
            end
          else
            begin
              reg287 <= $signed((wire271 >>> ({wire275[3'b100111:3'b11101]} <<< reg283[4'b01011110:1'b01])));
              reg288 <= $signed(((8'hb3) ?
                  $unsigned(wire4[4'b01101110:2'b1011]) : ((^~$signed(reg287)) == reg285[2'b1010:1'b11])));
              reg289 <= ((8'hbb) >>> reg286);
              reg290 <= $signed((reg281[4'b11011110:4'b10011011] ?
                  $unsigned($signed((reg280 && wire4))) : (^~wire1)));
            end
          if ({(~{reg278[3'b000100:1'b10],
                  ({wire1, reg276} ? $signed(reg288) : reg282)}),
              {(reg281 > ((reg286 ? wire275 : reg290) >> (reg289 ?
                      wire3 : wire4)))}})
            begin
              reg291 <= ((reg286 ?
                      (~|(wire3[2'b0111:2'b1011] & reg285[3'b111101:3'b010101])) : reg286[3'b100:2'b0110]) ?
                  $unsigned($unsigned(((reg289 <<< reg276) || (+reg286)))) : {wire271});
              reg292 <= {{($signed(wire0) | {{reg289}}),
                      ((+$unsigned(reg290)) ?
                          ($signed(wire74) ^ (|wire273)) : ((reg283 ?
                              wire0 : wire0) ~^ (reg283 ? wire273 : reg287)))}};
              reg293 <= $unsigned($signed((8'h9d)));
            end
          else
            begin
              reg291 <= reg282[2'b1110:2'b0110];
              reg292 <= reg281;
            end
          reg294 <= ($signed((^reg276)) <= {{$unsigned(reg277)}, reg289});
          reg295 <= ($signed(reg289[4'b00111100:1'b10]) != (|wire273[2'b1010:1'b11]));
        end
    end
  always
    @(posedge clk) begin
      if (reg276[2'b1110:2'b0110])
        begin
          reg296 <= $signed({reg284[2'b0111:2'b10], reg295});
          reg297 <= $signed(reg285);
          reg298 <= ((reg295 ? reg281 : $unsigned(reg286[5'b0000010000:1'b11])) ?
              {(!reg278)} : $signed((8'h9d)));
          reg299 <= (!(^(wire4 ?
              $signed({reg278, reg292}) : $unsigned(reg294))));
          reg300 <= reg285;
        end
      else
        begin
          reg296 <= ((reg281[4'b00111011:3'b110110] && $unsigned($unsigned($unsigned(wire2)))) && ((~$unsigned((reg292 ?
              reg279 : reg288))) > (+(reg288 ?
              $signed(wire273) : ((8'hb6) ? wire2 : reg299)))));
          reg297 <= {({($signed(reg293) ?
                          (wire1 ? reg287 : wire74) : $signed(wire271)),
                      (~&$signed(reg297))} ?
                  ($signed((reg295 <= wire4)) | (~$signed(wire0))) : (($signed(reg279) & (reg286 ?
                          reg282 : (8'had))) ?
                      ((wire273 ? reg296 : reg297) ?
                          (reg285 ^ reg299) : (-(8'hb9))) : $unsigned(reg283))),
              $unsigned((-$unsigned($signed(reg287))))};
          reg298 <= ($signed($unsigned((reg297[1'b01:1'b11] + reg297))) ?
              {reg292[4'b1110:4'b10101001],
                  (|(|(reg299 ?
                      reg291 : wire1)))} : ($signed(reg294[5'b0001110011:3'b100100]) >>> ((&wire74[4'b11001001:2'b0110]) ?
                  reg280 : (7'h40))));
          reg299 <= wire0;
        end
      reg301 <= (&reg279);
      reg302 <= wire271;
      reg303 <= {($signed(reg284[2'b010:1'b10]) - ($unsigned($signed(reg276)) + ((wire271 ?
                  reg279 : reg295) ?
              (-(8'h9c)) : $unsigned(reg301)))),
          reg291[5'b0000110011:2'b0011]};
      if (reg283[3'b000100:1'b01])
        begin
          reg304 <= (-(8'hb3));
          if ({reg300})
            begin
              reg305 <= reg289[3'b000110:1'b00];
              reg306 <= reg294[4'b01011001:4'b00111001];
              reg307 <= wire273;
            end
          else
            begin
              reg305 <= {reg293};
            end
        end
      else
        begin
          reg304 <= reg307[1'b10:1'b10];
          reg305 <= reg290[3'b111111:2'b0111];
          if ($unsigned({reg301[3'b001100:3'b001100]}))
            begin
              reg306 <= {({($unsigned(reg284) * {reg299})} & $unsigned((reg283 << $signed(reg290)))),
                  (wire271 < $unsigned(((reg306 ?
                      reg300 : wire3) || $unsigned(reg305))))};
              reg307 <= (~^{$signed($unsigned(((8'hb4) | reg287)))});
            end
          else
            begin
              reg306 <= (($signed(reg281[2'b0111:2'b10]) ~^ $signed({wire1[2'b0111:2'b10]})) ?
                  (~^wire2[1'b10:1'b10]) : {$signed((8'haf)),
                      reg290[3'b000101:1'b00]});
              reg307 <= ((~|reg286) & $signed(reg290));
              reg308 <= (8'hb5);
              reg309 <= $signed(($signed($unsigned(reg292)) >>> (|$signed($signed(wire273)))));
            end
          reg310 <= $signed((&(reg288[3'b000101:1'b00] ?
              ($unsigned(reg303) ?
                  wire0[4'b11111100:3'b101111] : (reg289 ?
                      (8'hb3) : wire4)) : $signed((8'hb1)))));
        end
    end
  assign wire311 = ({reg282} >= reg280[4'b10111001:2'b1111]);
  assign wire312 = ($signed((($signed(reg297) ?
                       $signed(wire2) : reg303[3'b001110:1'b01]) ^ reg303)) != $unsigned(($unsigned((reg310 ^~ reg306)) || {reg305})));
  assign wire313 = {$unsigned((!((reg283 ? wire275 : reg289) * (~^wire0)))),
                       reg303[3'b111101:3'b010101]};
  assign wire314 = (wire275 ^ $unsigned((|(reg283 != reg286))));
  assign wire315 = $unsigned($unsigned(reg297));
  assign wire316 = reg287;
  assign wire317 = $unsigned($unsigned(reg281[4'b00101011:3'b100101]));
  module131 modinst319 (wire318, clk, wire311, reg310, reg282, wire1, reg301);
  always
    @(posedge clk) begin
      if ((reg296 > reg276[4'b1110:4'b10101001]))
        begin
          reg320 <= (~^($unsigned($unsigned($signed(reg291))) ?
              reg299[3'b100:2'b0110] : (!reg306)));
        end
      else
        begin
          reg320 <= wire271[4'b1010:1'b10];
          reg321 <= $signed($signed((|$unsigned((reg308 ? wire0 : (8'h9f))))));
          reg322 <= ({((-{reg277, reg294}) ?
                      reg289[3'b110110:3'b101101] : ((reg277 | (8'h9c)) ?
                          ((8'hbd) && reg284) : wire318[1'b01:1'b11])),
                  (reg281 << ((|reg309) ?
                      wire271[3'b110110:3'b101101] : wire315[4'b10111000:3'b001100]))} ?
              ({(wire275 ~^ (8'ha9)),
                  ((wire271 != wire2) ^~ (reg288 ?
                      reg296 : wire313))} ^ ($signed($unsigned((8'haf))) << ($signed((8'hb9)) ?
                  reg300[3'b000100:1'b10] : $unsigned(reg299)))) : $signed((~$unsigned((reg294 == reg287)))));
          reg323 <= {({((wire4 << reg276) ~^ reg290)} ?
                  wire273 : ((reg279 + wire4[1'b11:1'b00]) << reg289))};
        end
      reg324 <= ((8'hb6) & reg280[5'b0010110011:4'b11001111]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module76
#( parameter param269 = ((&{(((8'h9c) ? (8'ha4) : (8'hbb)) ? (|(8'hac)) : (+(8'hab)))}) >>> (+((((7'h41) * (7'h42)) ? ((8'hbd) ? (8'hb2) : (8'hae)) : ((7'h43) ? (7'h43) : (8'haf))) ~^ {((7'h42) > (8'hb3))})))
, parameter param270 = ((|((!(param269 | (8'h9e))) ? param269 : {(param269 ? param269 : param269), {(8'ha7)}})) * ((param269 - param269) << (~((param269 ? param269 : (8'hb2)) ? ((7'h41) ? param269 : param269) : (param269 ? param269 : param269))))) )
(y, clk, wire81, wire80, wire79, wire78, wire77);
  output wire [32'b00000000000000000000000100100000:32'b00000000000000000000000000000000] y;
  input wire [1'b10:1'b10] clk;
  input wire signed [3'b001111:1'b00] wire81;
  input wire [4'b10101110:1'b10] wire80;
  input wire [5'b0001110101:1'b00] wire79;
  input wire signed [4'b10101110:1'b10] wire78;
  input wire signed [3'b001111:1'b00] wire77;
  wire [5'b0101010011:1'b10] wire267;
  wire signed [3'b000100:1'b10] wire250;
  wire signed [2'b1011:1'b00] wire249;
  reg [5'b0001010010:1'b10] reg248 = (1'h0);
  reg signed [4'b10101110:1'b10] reg247 = (1'h0);
  reg signed [4'b01001111:1'b10] reg246 = (1'h0);
  reg [5'b0101010011:1'b10] reg245 = (1'h0);
  reg signed [5'b1111010100:1'b00] reg244 = (1'h0);
  reg [2'b010:1'b10] reg243 = (1'h0);
  wire signed [4'b00101011:1'b00] wire242;
  wire [2'b010:1'b10] wire126;
  wire signed [4'b10101110:1'b10] wire89;
  wire signed [5'b0101010011:1'b10] wire88;
  wire [4'b10001101:1'b10] wire87;
  reg [5'b1000110000:1'b0] reg86 = (1'h0);
  reg [5'b1000110000:1'b0] reg85 = (1'h0);
  reg [4'b00111100:1'b10] reg84 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg83 = (1'h0);
  reg signed [4'b11011001:1'b10] reg82 = (1'h0);
  wire signed [3'b001111:1'b00] wire128;
  wire [4'b00111100:1'b10] wire129;
  wire signed [4'b1010:1'b10] wire130;
  wire signed [5'b1000110000:1'b0] wire240;
  assign y = {wire267,
                 wire250,
                 wire249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 wire242,
                 wire126,
                 wire89,
                 wire88,
                 wire87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 wire128,
                 wire129,
                 wire130,
                 wire240,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg82 <= wire78[1'b10:1'b10];
      if (wire78)
        begin
          reg83 <= ((|($unsigned((+(8'hb2))) - wire78[1'b11:1'b00])) != (~^(~|$unsigned(wire78))));
          reg84 <= $unsigned($signed(((~&$signed(wire77)) >= ((wire77 ?
              reg82 : (8'haa)) && (wire78 ? reg83 : wire78)))));
        end
      else
        begin
          reg83 <= {reg82[3'b100:2'b0110],
              ($signed(($unsigned((8'h9e)) ?
                  {reg82} : wire81)) | (&wire79[4'b01011000:4'b01001000]))};
          reg84 <= ($signed((~$signed((|wire79)))) * {(wire79[3'b000100:1'b10] && (reg82[2'b0111:2'b10] ?
                  (reg82 ? wire79 : reg84) : reg84[3'b000110:1'b00]))});
          reg85 <= $unsigned($unsigned(reg83[3'b011110:2'b1011]));
        end
      reg86 <= {($unsigned($unsigned($signed(reg83))) - (reg83 >= ($unsigned((7'h41)) || (wire77 ?
              wire80 : (8'ha2)))))};
    end
  assign wire87 = wire77;
  assign wire88 = (!($unsigned((+$signed(reg86))) ^ ($unsigned((reg85 ?
                          reg82 : wire79)) ?
                      (~&$signed(reg85)) : reg86[3'b100:2'b0110])));
  assign wire89 = $unsigned($unsigned((($signed((8'hb9)) ?
                      wire79 : (wire78 ^~ reg84)) * (wire87[4'b11101011:2'b1110] == reg83))));
  module90 modinst127 (wire126, clk, wire80, wire88, reg86, reg85, wire79);
  assign wire128 = ((reg85 && $signed((~(wire87 || (8'h9c))))) ?
                       (reg84[2'b0111:2'b10] * wire87[4'b01101001:3'b110110]) : wire77[3'b010110:2'b1010]);
  assign wire129 = $unsigned($signed({(~|$unsigned((8'ha3))),
                       ((-wire88) > (wire88 * reg84))}));
  assign wire130 = (((8'hb9) ? wire78 : wire77) ?
                       $signed(reg86[1'b10:1'b10]) : $unsigned($unsigned(((wire81 < wire129) != $unsigned(wire126)))));
  module131 modinst241 (.wire136(reg84), .wire132(wire87), .clk(clk), .wire134(wire128), .wire133(wire79), .wire135(wire129), .y(wire240));
  assign wire242 = $signed(({{(wire81 ? (8'haa) : reg86),
                               (wire240 ? reg83 : reg84)}} ?
                       (|wire129) : ((8'hb9) ?
                           {(wire87 ? reg82 : wire126),
                               wire88[2'b1110:2'b0110]} : {wire80[2'b1010:1'b11],
                               $signed(wire87)})));
  always
    @(posedge clk) begin
      reg243 <= $unsigned((&$unsigned($unsigned({wire81, wire129}))));
      if ({$unsigned($signed(wire89[1'b10:1'b10])), wire126})
        begin
          reg244 <= (((reg83[1'b10:1'b10] ?
                      $signed((reg243 ?
                          wire130 : wire89)) : (((8'ha6) & wire242) ^ wire89)) ?
                  wire78[4'b10011110:3'b101110] : ($signed($unsigned(wire77)) >= (wire81[3'b101101:2'b0110] ?
                      (reg243 ? wire240 : wire128) : (wire88 ?
                          reg82 : (8'hac))))) ?
              (reg86 ?
                  (^wire128[3'b000100:1'b01]) : ($unsigned($unsigned(wire128)) ?
                      $unsigned(wire77[3'b100:2'b0110]) : $unsigned({wire240,
                          reg84}))) : $unsigned($unsigned($unsigned({wire126}))));
          if (($signed((((|wire128) ?
                  ((8'had) ? wire242 : wire88) : $unsigned(wire129)) ?
              (wire89 ?
                  $unsigned((8'hbd)) : reg244[3'b010111:3'b100100]) : reg243)) & (~^wire77)))
            begin
              reg245 <= {wire89,
                  (~^(reg82[2'b1110:2'b0110] ?
                      $signed(wire129[4'b01111011:1'b01]) : (reg82 ?
                          reg244[3'b111111:1'b01] : ((8'hba) <= reg244))))};
              reg246 <= ((-wire89) ^~ wire126);
            end
          else
            begin
              reg245 <= wire130[1'b10:1'b10];
              reg246 <= (($signed(((reg83 ^ (8'hab)) ~^ (+(8'ha8)))) <= ($signed((reg86 ?
                  reg245 : reg244)) >> $signed(wire81[1'b11:1'b00]))) == wire129[4'b01011010:4'b10101000]);
            end
          reg247 <= (~^$signed(reg246[4'b00111011:3'b110110]));
        end
      else
        begin
          if ((reg82[3'b000100:2'b1011] ?
              ((-((wire126 ? wire80 : wire79) ? (8'ha7) : {wire80})) ?
                  wire126 : wire81) : wire81[3'b100111:3'b010110]))
            begin
              reg244 <= {$signed({reg83, reg245[2'b0111:2'b1011]}),
                  $signed(reg246[4'b01011000:4'b01001000])};
            end
          else
            begin
              reg244 <= $unsigned($unsigned($unsigned(reg83[2'b0111:2'b1011])));
              reg245 <= (($signed(((reg83 << reg83) >>> (wire78 * (8'ha4)))) || (reg244[4'b11011011:4'b01011000] ?
                  $signed(reg243) : ({reg82, reg83} ?
                      wire240[4'b00101010:4'b01111010] : {wire129}))) + $signed((8'h9f)));
              reg246 <= (-{$unsigned(($signed(reg245) ?
                      $signed(wire80) : ((8'hb0) + wire87))),
                  ($unsigned((wire129 ? wire81 : reg245)) ?
                      $unsigned((wire128 ? wire130 : wire78)) : reg86)});
              reg247 <= (wire80[4'b11111010:3'b100110] >> (&$signed(reg84)));
              reg248 <= wire77[2'b0111:2'b1011];
            end
        end
    end
  assign wire249 = ((8'ha0) ?
                       $signed(reg243) : {($unsigned((wire89 ?
                               (8'ha0) : reg84)) > ((7'h44) ? reg84 : reg82))});
  assign wire250 = reg84[2'b1010:1'b11];
  module251 modinst268 (.wire253(wire87), .clk(clk), .y(wire267), .wire255(wire79), .wire252(reg248), .wire254(wire89));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5
#( parameter param73 = {(((|((8'h9e) ? (8'hae) : (8'h9d))) ? {{(8'hbb)}, (~(8'ha3))} : ({(8'hb4)} ? ((8'had) && (8'hbd)) : (~^(8'ha1)))) >>> ({((8'hb7) ? (8'ha8) : (8'haa))} ? (~&((8'hb9) ? (7'h44) : (7'h43))) : (|((8'ha0) ? (7'h40) : (8'ha8)))))} )
(y, clk, wire6, wire7, wire8, wire9);
  output wire [32'b00000000000000000000000011011010:32'b00000000000000000000000000000000] y;
  input wire [1'b10:1'b10] clk;
  input wire signed [5'b1000110000:1'b0] wire6;
  input wire signed [5'b1111010100:1'b00] wire7;
  input wire signed [4'b10101110:1'b10] wire8;
  input wire signed [4'b00111100:1'b10] wire9;
  wire [2'b1011:1'b00] wire72;
  wire signed [4'b11011001:1'b10] wire71;
  wire [4'b00111100:1'b10] wire10;
  wire signed [3'b000110:1'b00] wire11;
  wire signed [5'b0101010011:1'b10] wire12;
  reg [4'b11111000:1'b00] reg13 = (1'h0);
  reg signed [4'b10001101:1'b10] reg14 = (1'h0);
  reg signed [4'b10001101:1'b10] reg15 = (1'h0);
  reg signed [4'b00111100:1'b10] reg16 = (1'h0);
  reg [4'b11011001:1'b10] reg17 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg18 = (1'h0);
  reg [2'b010:1'b10] reg19 = (1'h0);
  reg signed [2'b010:1'b10] reg20 = (1'h0);
  reg [5'b0101010011:1'b10] reg21 = (1'h0);
  reg signed [4'b10001101:1'b10] reg22 = (1'h0);
  wire [5'b1110001:1'b10] wire23;
  wire [4'b00111100:1'b10] wire24;
  wire signed [4'b01001111:1'b10] wire25;
  wire [5'b1110001:1'b10] wire69;
  assign y = {wire72,
                 wire71,
                 wire10,
                 wire11,
                 wire12,
                 reg13,
                 reg14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 wire23,
                 wire24,
                 wire25,
                 wire69,
                 (1'h0)};
  assign wire10 = $signed(wire9[3'b011111:3'b110111]);
  assign wire11 = wire9[3'b101110:3'b011110];
  assign wire12 = ($signed((~&{(|(8'ha5)),
                      (wire7 ? wire9 : (7'h44))})) >>> (({((8'had) ?
                                  wire8 : wire11)} ?
                          ((|wire8) ?
                              ((8'hb4) ?
                                  wire9 : wire9) : ((8'had) < wire7)) : $unsigned(wire11[2'b0111:2'b10])) ?
                      wire7 : wire11[2'b1110:2'b0110]));
  always
    @(posedge clk) begin
      reg13 <= wire7[1'b10:1'b10];
      if (wire9[3'b111101:3'b010101])
        begin
          if ({(wire10[4'b00111010:2'b0011] >>> wire7[3'b100111:2'b0010]),
              $signed($signed(((^wire8) << $signed((8'had)))))})
            begin
              reg14 <= $unsigned((~|{(-(^wire8)), $signed((&reg13))}));
              reg15 <= reg13[1'b11:1'b00];
            end
          else
            begin
              reg14 <= ($unsigned((8'h9e)) >>> $unsigned(($signed(wire6[3'b101110:3'b011110]) & wire11[1'b10:1'b10])));
              reg15 <= ({(+(-(wire8 ^ reg13)))} | ({(reg14 < (!wire12)),
                      ({wire12, wire8} ? wire10 : (reg13 | reg13))} ?
                  reg13 : ($unsigned($unsigned(wire10)) | ($unsigned(wire12) ?
                      (wire7 < (7'h41)) : $signed(wire11)))));
              reg16 <= ((({$unsigned(wire9),
                          $signed((8'hb5))} + $signed((+reg15))) ?
                      wire12[5'b1000110001:4'b10111001] : (reg13 ?
                          {{wire7},
                              wire8[4'b01101001:3'b110110]} : (~|$unsigned(reg15)))) ?
                  ($unsigned(((~^(8'hb0)) >>> (wire11 ? wire7 : wire6))) ?
                      ((+wire8) + wire7[4'b00101000:1'b11]) : wire6) : {($unsigned(wire10[2'b010:1'b10]) == ((wire9 != wire6) ?
                          (!reg15) : $unsigned(reg13))),
                      {(+(wire8 <<< wire11))}});
              reg17 <= (~$signed({reg13, wire8[3'b100111:2'b0010]}));
            end
          reg18 <= ((wire7[4'b01101001:3'b000111] ? (8'hae) : (8'ha2)) ?
              wire12 : (~^wire6[5'b1011110000:4'b10101000]));
          reg19 <= $unsigned((&$signed((wire12[3'b000101:1'b00] ?
              (reg16 ? reg15 : reg16) : (reg18 ? wire7 : wire8)))));
        end
      else
        begin
          if ((((|{$signed(reg18)}) ?
              $signed((~|$signed(reg19))) : $unsigned((wire9 ~^ wire8))) >= $signed(($signed(wire12[1'b11:1'b00]) ?
              {$unsigned(wire7)} : reg18[2'b1111:1'b11]))))
            begin
              reg14 <= (reg17[1'b10:1'b10] ?
                  $unsigned($unsigned((wire10 <= $unsigned(reg16)))) : $unsigned(($signed(wire6) ?
                      wire6 : (wire11 ? wire6[4'b01110:2'b1110] : reg16))));
              reg15 <= {wire8[4'b11111000:1'b00]};
            end
          else
            begin
              reg14 <= ((^$unsigned((~^$unsigned(reg17)))) ^~ (-$signed(wire6[4'b01101110:2'b1011])));
              reg15 <= wire9;
              reg16 <= reg13[3'b000100:2'b1011];
              reg17 <= (!wire11[3'b000101:2'b0111]);
            end
          reg18 <= $unsigned((reg16[4'b10111000:3'b011101] ?
              wire7[1'b11:1'b00] : wire10[3'b001111:1'b00]));
          reg19 <= {(~^$unsigned($signed({reg19, reg18})))};
          reg20 <= wire8[2'b0111:2'b10];
          reg21 <= (~&$unsigned(($signed(wire9) + reg13)));
        end
      reg22 <= $unsigned(reg17[2'b1010:1'b11]);
    end
  assign wire23 = $signed($signed((^~(wire11 + reg20[2'b1110:2'b0110]))));
  assign wire24 = reg19;
  assign wire25 = (^(8'hb9));
  module26 modinst70 (wire69, clk, wire7, reg18, reg16, wire23, wire8);
  assign wire71 = ($unsigned(reg14) ^~ ($signed($signed($unsigned(reg21))) ?
                      (&$unsigned(wire9)) : (^(^wire9[3'b110101:1'b11]))));
  assign wire72 = ($signed(wire12) >> wire23);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module26  (y, clk, wire31, wire30, wire29, wire28, wire27);
  output wire [32'b00000000000000000000000110101111:32'b00000000000000000000000000000000] y;
  input wire [1'b10:1'b10] clk;
  input wire signed [5'b1111010100:1'b00] wire31;
  input wire [4'b10101110:1'b10] wire30;
  input wire signed [4'b00111100:1'b10] wire29;
  input wire [5'b1110001:1'b10] wire28;
  input wire [3'b000100:1'b10] wire27;
  wire signed [3'b000101:1'b00] wire68;
  wire [3'b000101:1'b00] wire67;
  wire signed [4'b01001111:1'b10] wire66;
  wire [5'b1110001:1'b10] wire65;
  wire [4'b11011001:1'b10] wire64;
  wire [3'b000100:1'b10] wire63;
  wire [5'b1111010100:1'b00] wire62;
  wire signed [5'b0001110101:1'b00] wire61;
  wire signed [4'b01001111:1'b10] wire60;
  reg signed [4'b1010:1'b10] reg59 = (1'h0);
  wire signed [4'b00111100:1'b10] wire58;
  wire [5'b0001010010:1'b10] wire57;
  wire [5'b0101010011:1'b10] wire56;
  wire signed [3'b000101:1'b00] wire55;
  wire [2'b1011:1'b00] wire54;
  reg signed [3'b000100:1'b10] reg53 = (1'h0);
  reg [3'b001111:1'b00] reg52 = (1'h0);
  wire [4'b11011001:1'b10] wire51;
  wire [2'b1011:1'b00] wire50;
  reg signed [5'b0001110101:1'b00] reg49 = (1'h0);
  reg signed [4'b11111000:1'b00] reg48 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg47 = (1'h0);
  reg [5'b0001110101:1'b00] reg46 = (1'h0);
  reg [4'b00101011:1'b00] reg45 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg44 = (1'h0);
  reg signed [4'b01001111:1'b10] reg43 = (1'h0);
  reg [4'b00111100:1'b10] reg42 = (1'h0);
  reg [4'b00101011:1'b00] reg41 = (1'h0);
  reg signed [3'b000110:1'b00] reg40 = (1'h0);
  reg signed [4'b1010:1'b10] reg39 = (1'h0);
  reg signed [4'b00101011:1'b00] reg38 = (1'h0);
  reg signed [3'b000101:1'b00] reg37 = (1'h0);
  reg signed [4'b11111000:1'b00] reg36 = (1'h0);
  wire [4'b11011001:1'b10] wire35;
  wire signed [5'b0001010010:1'b10] wire34;
  wire [4'b11011001:1'b10] wire33;
  wire [5'b0101010011:1'b10] wire32;
  assign y = {wire68,
                 wire67,
                 wire66,
                 wire65,
                 wire64,
                 wire63,
                 wire62,
                 wire61,
                 wire60,
                 reg59,
                 wire58,
                 wire57,
                 wire56,
                 wire55,
                 wire54,
                 reg53,
                 reg52,
                 wire51,
                 wire50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 (1'h0)};
  assign wire32 = (($signed($unsigned($signed(wire28))) ?
                      (-$signed(wire28)) : {$unsigned(wire27[3'b001100:3'b001100]),
                          (8'h9c)}) - {((~|wire29[4'b01111100:3'b011101]) ?
                          $signed((wire31 ? wire31 : wire27)) : wire31),
                      {((wire29 ? wire30 : (8'hb7)) ?
                              wire31 : $unsigned(wire27))}});
  assign wire33 = (~|$signed(wire27));
  assign wire34 = (~^(~&wire33[4'b00101000:1'b11]));
  assign wire35 = ($signed(wire33) || $signed({($unsigned(wire30) ?
                          (wire28 ? wire28 : wire28) : (wire32 < (8'ha9)))}));
  always
    @(posedge clk) begin
      reg36 <= $signed(({(8'h9d),
              ($unsigned(wire27) ? wire29[3'b001111:1'b00] : {wire34})} ?
          $signed(wire32) : (wire30[4'b11101011:2'b1110] ?
              wire35[2'b1111:1'b11] : ((^wire33) ?
                  ((8'hbe) ? wire29 : wire31) : wire27[1'b10:1'b10]))));
      reg37 <= (~|$signed(($signed((|wire35)) ^~ wire33[2'b1010:1'b11])));
      if ($signed(((reg37 ? wire28[1'b01:1'b11] : (^~(wire34 << wire33))) ?
          wire28 : reg36[3'b011110:2'b1011])))
        begin
          if ((8'hbe))
            begin
              reg38 <= (wire32 <= {$signed((~(-wire30)))});
              reg39 <= (wire35[2'b1111:1'b11] ?
                  ((~|wire29[1'b10:1'b10]) + wire32[5'b0001110010:3'b101110]) : (~wire32[4'b01011110:4'b001110]));
              reg40 <= $signed((wire27[3'b001100:3'b001100] ?
                  $unsigned($signed(wire34[1'b01:1'b11])) : (($signed((8'hb5)) >= $signed(wire34)) || $signed($signed(wire31)))));
              reg41 <= {reg36[2'b1110:2'b0110], (^wire35)};
              reg42 <= reg39;
            end
          else
            begin
              reg38 <= (!$signed(wire32));
              reg39 <= (8'ha8);
            end
        end
      else
        begin
          reg38 <= reg36;
          reg39 <= ((!$signed(reg38[2'b1010:1'b11])) * $signed($unsigned(reg40)));
          if (wire29[4'b0111100:4'b00011001])
            begin
              reg40 <= ((reg38 & $unsigned((~|(!wire33)))) >>> wire34[2'b1011:1'b00]);
            end
          else
            begin
              reg40 <= (wire28[4'b00101110:3'b110100] ?
                  ({$unsigned($unsigned(reg40)),
                      $unsigned($unsigned(wire29))} && $signed((8'hb4))) : ($signed($signed($signed(wire29))) - (((|wire28) ?
                      $signed(wire28) : {wire33}) & (8'hb8))));
              reg41 <= (~|(~|reg38[3'b000100:1'b01]));
              reg42 <= ($signed($signed((wire31 <= {(8'haa), wire32}))) ?
                  $unsigned(reg42) : (~|$unsigned((reg38[4'b11001011:4'b10101011] ?
                      (reg38 != wire31) : (reg40 ? reg36 : (8'ha3))))));
              reg43 <= (8'hbf);
            end
          reg44 <= $signed((&reg43[4'b01111100:3'b011101]));
          if (reg42[3'b101110:3'b011110])
            begin
              reg45 <= $unsigned(({(reg39 ?
                      wire28 : (wire29 || wire31))} || $unsigned((~^$signed((8'hb3))))));
              reg46 <= $unsigned(reg45[3'b000100:1'b10]);
              reg47 <= $unsigned(reg38);
              reg48 <= $unsigned({((^~(^(8'ha2))) ?
                      $signed($unsigned(wire30)) : ((&wire34) != reg42[1'b01:1'b11])),
                  {wire28, $signed($signed(reg38))}});
              reg49 <= ({(~^$unsigned((wire32 > reg37))),
                  (8'hb6)} & wire33[3'b011110:2'b1011]);
            end
          else
            begin
              reg45 <= (^~$signed(($signed((wire27 ? wire28 : reg41)) ?
                  ($signed(reg38) + {reg41}) : ((wire33 == wire30) ?
                      (^reg41) : (reg43 ^~ (8'ha7))))));
            end
        end
    end
  assign wire50 = {$signed((&reg48[3'b011111:3'b110111])),
                      {(wire29[3'b111111:1'b01] ?
                              reg43 : $signed((reg39 ? wire32 : wire32))),
                          (8'hbe)}};
  assign wire51 = (!wire34);
  always
    @(posedge clk) begin
      reg52 <= reg49[3'b000101:1'b00];
      reg53 <= reg42[1'b11:1'b00];
    end
  assign wire54 = reg46[5'b1011110011:4'b10111011];
  assign wire55 = $unsigned($unsigned($unsigned(reg47)));
  assign wire56 = ($signed((&{(|reg46)})) | (~$signed($signed((reg40 ?
                      wire54 : reg44)))));
  assign wire57 = (~(reg45 ?
                      ((!$signed(reg45)) ?
                          (~(+reg39)) : (|$unsigned(wire56))) : reg37));
  assign wire58 = (-(wire32 ?
                      (wire35 ^~ reg43[4'b10011101:4'b01000]) : (($signed(reg36) | $unsigned(reg41)) ?
                          ({wire30} ~^ $unsigned(wire50)) : reg41[3'b100111:3'b010110])));
  always
    @(posedge clk) begin
      reg59 <= $signed((((~|(|reg46)) >> (~|$unsigned((8'hb7)))) ?
          (reg47 >= reg36) : (~^$unsigned($unsigned(reg52)))));
    end
  assign wire60 = (wire35 == (-wire34[3'b000100:1'b10]));
  assign wire61 = {((+$signed(((8'hac) + reg48))) || ($signed(reg48[3'b110110:3'b101101]) ?
                          reg49 : (reg43[1'b01:1'b11] >> (reg42 >> reg41)))),
                      {($unsigned((wire60 ? reg46 : reg45)) ?
                              {reg47} : (wire57 ?
                                  (reg38 <<< (8'hb3)) : $unsigned(reg37)))}};
  assign wire62 = $unsigned(reg47[4'b11011001:1'b10]);
  assign wire63 = ($signed((((!wire30) ?
                              wire62[4'b11101011:2'b1110] : $unsigned(wire28)) ?
                          wire29[4'b01101001:3'b000111] : {(reg37 | wire50),
                              $signed(wire34)})) ?
                      (-(wire29[3'b001111:1'b00] ?
                          reg41[2'b1110:2'b0110] : reg48[3'b011110:2'b1011])) : (reg42 ?
                          (~|(|$unsigned(wire30))) : (&$signed((wire60 ?
                              wire60 : wire55)))));
  assign wire64 = {reg38[1'b01:1'b11]};
  assign wire65 = {reg42, (&{(&((8'hb5) == wire28))})};
  assign wire66 = $unsigned(($signed((~&((8'h9e) ^~ (8'hb8)))) > reg46[4'b10011110:3'b111111]));
  assign wire67 = (wire60[4'b1110:4'b10101001] >= reg42[4'b10111001:2'b1111]);
  assign wire68 = ({(($signed(reg42) | {wire32}) ?
                          {(reg48 ? wire33 : reg45),
                              $unsigned(wire33)} : wire65[3'b100111:3'b11101])} >= (reg48 || ($signed($unsigned(wire65)) ?
                      ($unsigned(wire60) ?
                          (wire63 ?
                              wire57 : wire62) : (reg49 | wire30)) : ($unsigned(reg53) <<< $signed(wire33)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module251  (y, clk, wire255, wire254, wire253, wire252);
  output wire [32'b00000000000000000000000001100001:32'b00000000000000000000000000000000] y;
  input wire [1'b10:1'b10] clk;
  input wire signed [3'b000101:1'b00] wire255;
  input wire signed [4'b10101110:1'b10] wire254;
  input wire signed [3'b001111:1'b00] wire253;
  input wire [5'b0001010010:1'b10] wire252;
  wire [5'b0101010011:1'b10] wire266;
  wire [5'b0001010010:1'b10] wire265;
  wire signed [4'b1010:1'b10] wire264;
  wire [2'b010:1'b10] wire263;
  wire signed [4'b00111100:1'b10] wire262;
  reg [3'b000110:1'b00] reg261 = (1'h0);
  wire signed [4'b00111100:1'b10] wire260;
  wire [3'b001111:1'b00] wire259;
  wire signed [2'b1011:1'b00] wire258;
  wire signed [2'b010:1'b10] wire257;
  wire [3'b000101:1'b00] wire256;
  assign y = {wire266,
                 wire265,
                 wire264,
                 wire263,
                 wire262,
                 reg261,
                 wire260,
                 wire259,
                 wire258,
                 wire257,
                 wire256,
                 (1'h0)};
  assign wire256 = wire252;
  assign wire257 = {{wire255[2'b1111:1'b11],
                           (wire253[1'b01:1'b11] ?
                               ((~^wire253) ?
                                   wire253[1'b01:1'b11] : (~|wire254)) : $signed((wire254 >>> wire252)))},
                       (~$signed((wire252 ?
                           $unsigned(wire253) : wire256[3'b100:2'b0110])))};
  assign wire258 = ((8'hbd) <= $signed(wire256[3'b000100:1'b01]));
  assign wire259 = wire253[3'b100:2'b0110];
  assign wire260 = $signed(($signed($signed(wire255[2'b0111:2'b1011])) ~^ (wire252 == $signed($unsigned(wire254)))));
  always
    @(posedge clk) begin
      reg261 <= (wire253 <<< $signed($signed($signed((wire257 ?
          wire257 : wire255)))));
    end
  assign wire262 = ((reg261 ^ {$signed((~|wire258)),
                           ((~wire252) >= {wire260, (8'ha4)})}) ?
                       ($signed((wire252 ~^ $signed(wire260))) || ($unsigned($unsigned(wire255)) != reg261[2'b010:1'b10])) : ($unsigned((reg261[3'b000100:1'b01] ?
                               (8'hb1) : ((8'hb6) ? wire259 : wire255))) ?
                           wire259[2'b0111:2'b1011] : ($signed(wire255) ?
                               (~|wire253) : ((|reg261) - reg261))));
  assign wire263 = (wire254 || $unsigned(wire258[2'b1010:1'b11]));
  assign wire264 = (^~{((wire256 <= reg261[1'b11:1'b00]) ?
                           wire258[1'b10:1'b10] : ((8'hb5) >>> wire262[3'b111111:2'b0111]))});
  assign wire265 = (8'hb5);
  assign wire266 = $signed(wire260[2'b1111:1'b11]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module131
#( parameter param238 = (((^(((8'ha7) ? (7'h43) : (8'hba)) ? (8'h9e) : ((8'hb3) ? (8'h9c) : (8'hac)))) ~^ (!(|((8'hbb) ? (8'ha9) : (8'hbd))))) >> (~(((+(7'h43)) >>> (|(8'hbf))) & (~|(~&(8'hb0))))))
, parameter param239 = param238 )
(y, clk, wire136, wire135, wire134, wire133, wire132);
  output wire [32'b00000000000000000000010010010110:32'b00000000000000000000000000000000] y;
  input wire [1'b10:1'b10] clk;
  input wire signed [4'b00111100:1'b10] wire136;
  input wire [4'b00111100:1'b10] wire135;
  input wire [3'b001111:1'b00] wire134;
  input wire [5'b0001110101:1'b00] wire133;
  input wire [2'b010:1'b10] wire132;
  wire signed [4'b10001101:1'b10] wire237;
  reg [4'b11111000:1'b00] reg236 = (1'h0);
  reg [3'b000101:1'b00] reg235 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg234 = (1'h0);
  reg [5'b1110001:1'b10] reg233 = (1'h0);
  reg signed [4'b1010:1'b10] reg232 = (1'h0);
  reg [3'b000110:1'b00] reg231 = (1'h0);
  reg signed [4'b11011001:1'b10] reg230 = (1'h0);
  reg [5'b0001010010:1'b10] reg229 = (1'h0);
  reg [4'b10101110:1'b10] reg228 = (1'h0);
  reg signed [3'b000100:1'b10] reg227 = (1'h0);
  reg signed [2'b1011:1'b00] reg226 = (1'h0);
  reg signed [4'b01001111:1'b10] reg225 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg224 = (1'h0);
  reg signed [3'b000110:1'b00] reg223 = (1'h0);
  reg [4'b1010:1'b10] reg222 = (1'h0);
  reg [4'b10001101:1'b10] reg221 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg220 = (1'h0);
  reg signed [5'b1111010100:1'b00] reg219 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg218 = (1'h0);
  reg signed [2'b010:1'b10] reg217 = (1'h0);
  wire signed [3'b000100:1'b10] wire216;
  wire signed [2'b1011:1'b00] wire215;
  reg signed [5'b1110001:1'b10] reg214 = (1'h0);
  reg signed [4'b10001101:1'b10] reg213 = (1'h0);
  reg signed [5'b0001010010:1'b10] reg212 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg211 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg210 = (1'h0);
  reg [3'b001111:1'b00] reg209 = (1'h0);
  reg signed [2'b1011:1'b00] reg208 = (1'h0);
  reg [5'b1111010100:1'b00] reg207 = (1'h0);
  reg signed [5'b1111010100:1'b00] reg206 = (1'h0);
  wire [3'b000100:1'b10] wire205;
  reg signed [3'b000110:1'b00] reg204 = (1'h0);
  reg [5'b1000110000:1'b0] reg203 = (1'h0);
  reg [3'b000110:1'b00] reg202 = (1'h0);
  reg signed [4'b00101011:1'b00] reg201 = (1'h0);
  reg [4'b00101011:1'b00] reg200 = (1'h0);
  reg [5'b1111010100:1'b00] reg199 = (1'h0);
  wire signed [4'b00101011:1'b00] wire198;
  reg signed [3'b000101:1'b00] reg197 = (1'h0);
  wire [3'b001111:1'b00] wire196;
  reg signed [5'b0001010010:1'b10] reg195 = (1'h0);
  reg [5'b1111010100:1'b00] reg194 = (1'h0);
  reg signed [4'b10101110:1'b10] reg193 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg192 = (1'h0);
  reg [3'b000110:1'b00] reg191 = (1'h0);
  reg signed [4'b11111000:1'b00] reg190 = (1'h0);
  reg signed [3'b001111:1'b00] reg189 = (1'h0);
  reg signed [3'b000100:1'b10] reg188 = (1'h0);
  reg signed [4'b00111100:1'b10] reg187 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg186 = (1'h0);
  reg signed [4'b1010:1'b10] reg185 = (1'h0);
  wire [2'b010:1'b10] wire184;
  wire signed [3'b000110:1'b00] wire183;
  reg signed [4'b11111000:1'b00] reg182 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg181 = (1'h0);
  reg signed [4'b1010:1'b10] reg180 = (1'h0);
  reg [5'b1110001:1'b10] reg179 = (1'h0);
  reg signed [5'b0001110101:1'b00] reg178 = (1'h0);
  reg signed [5'b0001010010:1'b10] reg177 = (1'h0);
  reg [3'b000100:1'b10] reg176 = (1'h0);
  reg [4'b11111000:1'b00] reg175 = (1'h0);
  reg [2'b1011:1'b00] reg174 = (1'h0);
  reg [4'b10101110:1'b10] reg173 = (1'h0);
  reg signed [4'b00101011:1'b00] reg172 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg171 = (1'h0);
  reg [5'b0001010010:1'b10] reg170 = (1'h0);
  reg [3'b000100:1'b10] reg169 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg168 = (1'h0);
  reg signed [3'b000110:1'b00] reg167 = (1'h0);
  reg signed [5'b0001110101:1'b00] reg166 = (1'h0);
  reg [3'b000100:1'b10] reg165 = (1'h0);
  reg signed [4'b10001101:1'b10] reg164 = (1'h0);
  reg [4'b00101011:1'b00] reg163 = (1'h0);
  reg [4'b11111000:1'b00] reg162 = (1'h0);
  reg [5'b0001010010:1'b10] reg161 = (1'h0);
  reg [4'b11111000:1'b00] reg160 = (1'h0);
  reg signed [3'b000100:1'b10] reg159 = (1'h0);
  reg [5'b1000110000:1'b0] reg158 = (1'h0);
  reg signed [3'b000110:1'b00] reg157 = (1'h0);
  reg signed [4'b00111100:1'b10] reg156 = (1'h0);
  reg signed [4'b10101110:1'b10] reg155 = (1'h0);
  reg [5'b1000110000:1'b0] reg154 = (1'h0);
  reg [5'b1000110000:1'b0] reg153 = (1'h0);
  reg signed [3'b001111:1'b00] reg152 = (1'h0);
  reg [3'b001111:1'b00] reg151 = (1'h0);
  reg signed [4'b11111000:1'b00] reg150 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg149 = (1'h0);
  reg signed [5'b1000110000:1'b0] reg148 = (1'h0);
  reg [5'b1111010100:1'b00] reg147 = (1'h0);
  reg signed [5'b1110001:1'b10] reg146 = (1'h0);
  reg signed [5'b1111010100:1'b00] reg145 = (1'h0);
  reg signed [4'b10101110:1'b10] reg144 = (1'h0);
  reg signed [5'b1110001:1'b10] reg143 = (1'h0);
  wire signed [4'b1010:1'b10] wire142;
  wire signed [2'b1011:1'b00] wire141;
  reg [5'b1111010100:1'b00] reg140 = (1'h0);
  reg [3'b001111:1'b00] reg139 = (1'h0);
  reg signed [2'b010:1'b10] reg138 = (1'h0);
  wire [3'b000100:1'b10] wire137;
  assign y = {wire237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg217,
                 wire216,
                 wire215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 wire205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 wire198,
                 reg197,
                 wire196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 wire184,
                 wire183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 wire142,
                 wire141,
                 reg140,
                 reg139,
                 reg138,
                 wire137,
                 (1'h0)};
  assign wire137 = $signed(wire136[4'b01111011:1'b01]);
  always
    @(posedge clk) begin
      reg138 <= wire133[4'b11111010:3'b100110];
      reg139 <= (~^(~&$signed(((reg138 <= wire137) && (wire136 ?
          (8'hb4) : (8'hb1))))));
      reg140 <= $signed(($unsigned(reg138[2'b1110:2'b0110]) != $unsigned(wire137)));
    end
  assign wire141 = $signed(({$unsigned($unsigned(wire133)),
                       wire135[1'b01:1'b11]} >> ($signed((8'hb8)) >= ($signed(wire135) || (wire137 > reg138)))));
  assign wire142 = $signed(wire136[3'b100:2'b0110]);
  always
    @(posedge clk) begin
      reg143 <= wire136;
      reg144 <= {(!(|wire142[3'b111101:3'b010101]))};
      if (wire141[2'b010:1'b10])
        begin
          reg145 <= ((({wire135[2'b1111:1'b11]} ?
                      (!(^wire135)) : $signed((wire136 != wire136))) ?
                  (^$unsigned($unsigned(reg144))) : ($unsigned($unsigned((8'h9e))) | {(wire142 | wire135)})) ?
              $signed(wire141[2'b010:1'b10]) : wire137);
          if (wire133[4'b01111000:3'b100111])
            begin
              reg146 <= reg139[3'b111111:2'b0111];
            end
          else
            begin
              reg146 <= (reg146[3'b100:2'b0110] > ((($signed(wire141) ?
                      $unsigned((8'hae)) : wire136) ?
                  (wire136[4'b10001100:2'b1111] ?
                      $unsigned((8'hb9)) : (wire142 & wire142)) : ((8'hb4) ?
                      {reg144} : {reg143, wire137})) ^~ reg138[1'b01:1'b11]));
              reg147 <= $unsigned(wire135);
            end
          if (reg138[1'b11:1'b00])
            begin
              reg148 <= {wire141[2'b010:1'b10],
                  $signed((reg145[4'b1100:1'b11] & $signed((^~wire136))))};
            end
          else
            begin
              reg148 <= (^(~&(({wire135, (8'hb0)} ?
                  (^~reg147) : reg139) >>> (!wire134[3'b001110:1'b01]))));
              reg149 <= ($signed($signed({(wire142 && (8'hbb))})) < reg145);
              reg150 <= (reg147 ?
                  $unsigned($signed((wire135 >> $signed((8'ha9))))) : (reg145 ?
                      (wire135[4'b11111100:4'b10111100] + {{wire136}}) : ((wire136 ?
                              {(8'h9d)} : reg148) ?
                          (reg139 ? (^(8'hb8)) : $signed((7'h40))) : {(reg144 ?
                                  reg147 : wire137)})));
              reg151 <= (reg150[2'b1011:1'b00] && (~^$signed($unsigned(reg148))));
              reg152 <= wire136;
            end
          if ((~$signed(({wire135[3'b110101:1'b11]} | $unsigned((wire137 == reg145))))))
            begin
              reg153 <= ({$unsigned($unsigned($unsigned(reg152)))} ?
                  reg139 : $unsigned((&reg138)));
              reg154 <= reg146[4'b1011100:3'b101110];
              reg155 <= ({{(|{reg149, (8'hb4)})}} ?
                  (~&wire141) : {(((reg139 <= (8'hb9)) == $unsigned(reg138)) <<< reg148[3'b110101:1'b11])});
            end
          else
            begin
              reg153 <= $signed($unsigned((reg149 >> ($signed(reg153) ?
                  reg148 : (~&reg147)))));
              reg154 <= $signed(((wire141[2'b0111:2'b10] == reg139) ?
                  $unsigned(reg152) : (reg139[2'b1111:1'b11] ?
                      $unsigned((reg140 * reg145)) : $unsigned($signed(reg143)))));
              reg155 <= ((!$signed(reg152[1'b10:1'b10])) ?
                  $unsigned(($unsigned($signed(wire132)) >>> $unsigned(reg155))) : $unsigned((-$unsigned((reg139 ?
                      reg145 : reg153)))));
            end
        end
      else
        begin
          reg145 <= ((+reg147[4'b01011001:4'b00111001]) ?
              $unsigned(reg152) : (reg150[1'b11:1'b00] >> ((8'hbc) ?
                  {$unsigned(reg153),
                      $unsigned(reg148)} : reg153[4'b10111110:4'b10101000])));
        end
      if (reg152[3'b000110:1'b00])
        begin
          reg156 <= ({$signed((8'h9d)),
                  {((reg144 <= wire142) <<< $unsigned((7'h43)))}} ?
              $signed((&((~^(8'ha0)) & {reg154,
                  reg146}))) : $signed($unsigned($signed(wire133))));
          if ((reg155[4'b01011000:4'b01001000] ?
              (wire135[4'b00101000:1'b11] ?
                  (8'haf) : (~^($signed((8'haf)) | (wire141 ?
                      wire132 : reg145)))) : (((!wire132) ?
                      $signed((reg140 <<< (8'hb5))) : $signed((-reg144))) ?
                  ($unsigned((wire141 ^ reg154)) ^~ ((8'ha0) == reg155)) : reg140)))
            begin
              reg157 <= reg150[1'b11:1'b00];
              reg158 <= $signed(((reg154 || wire132[2'b1110:2'b0110]) >= reg156[1'b10:1'b10]));
              reg159 <= (|(($unsigned($signed(reg143)) ?
                  reg155 : wire133[4'b11111011:3'b110111]) | reg138[1'b11:1'b00]));
              reg160 <= {(^~reg140)};
            end
          else
            begin
              reg157 <= ($signed((reg144[4'b01011001:4'b00111001] ?
                      {(reg138 ? wire136 : wire132),
                          $unsigned(reg138)} : ($unsigned(reg153) > (reg154 ?
                          reg154 : reg138)))) ?
                  (^~(reg149[4'b00101010:4'b01111010] ?
                      (^~reg143) : (reg158[4'b1010:1'b10] - $signed(reg154)))) : wire142);
            end
          reg161 <= reg154[4'b11011111:3'b100101];
          reg162 <= reg145;
          reg163 <= (7'h43);
        end
      else
        begin
          reg156 <= $unsigned(((($signed((8'hb7)) ?
              $signed(reg163) : (reg146 ?
                  reg158 : wire136)) <<< $signed($unsigned((8'had)))) > (($signed(reg157) - (&reg144)) ?
              (-((8'hb3) ^ reg154)) : $unsigned((wire135 ?
                  reg139 : wire133)))));
          reg157 <= (reg160 != $signed($unsigned({(~&reg154)})));
          reg158 <= $unsigned(wire135[2'b010:1'b10]);
          reg159 <= ((-(reg158[3'b000100:1'b10] < (^~(reg147 ?
              (8'ha5) : reg143)))) == (+(reg148[4'b00111111:4'b10101111] ?
              (reg155 ?
                  (reg152 ?
                      reg143 : (8'ha7)) : $signed(reg145)) : $unsigned((wire134 ?
                  reg161 : wire134)))));
          reg160 <= $signed((reg158 ? wire132[2'b1110:2'b0110] : (~^(7'h42))));
        end
      reg164 <= {(-reg140[4'b01011111:4'b11111110])};
    end
  always
    @(posedge clk) begin
      if ($unsigned((~|$unsigned(reg157))))
        begin
          reg165 <= $signed((8'ha2));
          if ($signed(($unsigned(reg139) ?
              ({(reg157 ^ reg145)} != {(!wire142),
                  $unsigned((8'ha4))}) : $unsigned({(+wire135),
                  (wire133 ? reg143 : reg154)}))))
            begin
              reg166 <= (~reg165[2'b0111:2'b1011]);
              reg167 <= {($unsigned(($unsigned(reg161) ?
                      reg165 : (8'hbf))) ^~ reg151),
                  reg149};
              reg168 <= wire134[3'b100:2'b0110];
            end
          else
            begin
              reg166 <= (reg155[1'b10:1'b10] << reg168);
              reg167 <= $unsigned($signed(({reg153} ?
                  ({reg152} ? $signed(reg158) : $signed(reg167)) : (reg152 ?
                      (~^(8'hb6)) : (reg167 && reg145)))));
            end
          reg169 <= $signed(reg154);
        end
      else
        begin
          reg165 <= ({(!((wire141 ~^ (8'hab)) * $signed(reg168)))} ?
              wire132[1'b10:1'b10] : (($unsigned(reg152) ?
                      (reg140[3'b010110:2'b1010] == (~&wire141)) : (reg163 ?
                          reg156[1'b01:1'b11] : reg151)) ?
                  (reg147[3'b010101:3'b110100] & $signed({reg151})) : {($unsigned(reg156) < reg161[4'b01011001:4'b00111001])}));
        end
    end
  always
    @(posedge clk) begin
      if (reg139)
        begin
          reg170 <= ({(~&$unsigned(reg150)), $unsigned($signed(reg167))} ?
              (wire137[1'b10:1'b10] ?
                  reg148[4'b00011101:4'b01101] : (8'ha8)) : ($signed($unsigned({reg147,
                  (8'hb9)})) - $signed(reg143)));
        end
      else
        begin
          if (reg154[2'b1111:1'b11])
            begin
              reg170 <= reg155;
              reg171 <= ((8'hbb) ~^ (($signed($signed(reg165)) ?
                      $signed((~&wire132)) : reg153) ?
                  (^reg156[4'b00101010:1'b11]) : reg151[3'b000100:1'b01]));
            end
          else
            begin
              reg170 <= (wire142 == reg154);
            end
          reg172 <= {reg168[4'b11111000:1'b00]};
        end
      if (reg150)
        begin
          reg173 <= reg144[4'b00101101:3'b000100];
          if (wire133[4'b00011101:4'b11111010])
            begin
              reg174 <= wire132;
              reg175 <= (~^({$signed($unsigned(reg148)),
                  (reg158[4'b11011110:4'b10011011] <= (~reg170))} ^ $unsigned({(!wire134)})));
              reg176 <= ($unsigned(({(reg145 ?
                      reg172 : reg145)} - $signed($unsigned((8'haa))))) != (~reg168));
              reg177 <= (~&reg166);
            end
          else
            begin
              reg174 <= $unsigned((~&(wire133 ?
                  (((8'h9d) >> reg153) ?
                      reg174[1'b01:1'b11] : {reg152}) : (^~wire133))));
              reg175 <= (8'hb3);
              reg176 <= ((~|reg174) ^~ (($signed(reg158[4'b00101010:1'b11]) ^~ $unsigned((reg165 ?
                      wire142 : reg165))) ?
                  reg171[4'b1100:1'b11] : (reg138 < wire141)));
              reg177 <= {(reg172[1'b10:1'b10] >= $unsigned(reg144[3'b011111:3'b110111])),
                  reg148};
            end
          reg178 <= $signed(reg173);
          reg179 <= $unsigned((+((~&wire137) ?
              (^~((7'h42) <<< reg178)) : (~|(reg155 << (8'hb3))))));
        end
      else
        begin
          reg173 <= (reg165[3'b000100:2'b1011] <<< ($signed($signed(((8'ha5) | reg167))) ?
              $signed(wire142[1'b10:1'b10]) : $unsigned(reg173[4'b00001101:2'b1010])));
        end
      reg180 <= ($signed(((reg151 ?
                  reg161[5'b010010:5'b110110000] : $unsigned(wire134)) ?
              {((8'hba) ? wire142 : wire134), $unsigned(reg151)} : {reg172})) ?
          ((^~$unsigned({(8'h9f), reg165})) ?
              reg140[1'b10:1'b10] : ($signed($signed(wire137)) - (8'hbd))) : ((8'ha2) && ($signed($unsigned(wire136)) < (~(+reg150)))));
      reg181 <= $unsigned(($unsigned(((reg162 >>> reg140) ?
              (reg155 > (8'ha4)) : (8'hae))) ?
          (&($signed(reg146) ? reg158 : $unsigned(reg160))) : ((reg162 ?
              {reg146} : (reg162 ?
                  reg165 : reg178)) && $unsigned($signed(reg152)))));
      reg182 <= $signed($unsigned((reg139 != ($unsigned(reg154) ^ reg180))));
    end
  assign wire183 = reg169;
  assign wire184 = ((reg150 ?
                       (((+(8'hb5)) ?
                           $signed(reg157) : $signed(wire137)) * reg166) : reg169) ~^ $unsigned($signed($unsigned((reg160 < reg181)))));
  always
    @(posedge clk) begin
      reg185 <= {$signed($unsigned(((reg167 ? reg138 : reg169) * (~reg164))))};
      reg186 <= (((~&(&reg152)) ?
              (reg156[3'b010101:3'b110100] ?
                  $signed($signed((8'ha0))) : (|(reg171 ?
                      reg173 : wire141))) : reg160) ?
          reg175[4'b00101000:1'b11] : (((((8'hb3) ? reg162 : (8'ha9)) <<< (8'haf)) ?
              $signed((~&reg177)) : ((wire142 ?
                  reg175 : (8'hb2)) * $unsigned(reg148))) < reg143));
      if ((8'ha5))
        begin
          reg187 <= reg158[5'b0000010000:1'b11];
          reg188 <= reg163[4'b1010:3'b100101];
          reg189 <= $signed(($unsigned({$signed(reg147),
              (8'hb6)}) && $signed((^~(wire137 ? reg162 : wire136)))));
          if ($unsigned(($signed($unsigned((reg172 ?
              reg150 : (8'ha3)))) << $unsigned(reg181))))
            begin
              reg190 <= $unsigned({reg178[5'b0110110100:4'b01011], reg178});
              reg191 <= ((reg138[1'b10:1'b10] >>> $signed(((reg173 ?
                  reg172 : (8'h9c)) ~^ $unsigned((8'h9d))))) ^~ (|$signed($signed((wire133 ~^ (8'ha1))))));
              reg192 <= ({reg154} ?
                  reg178[2'b1110:2'b0110] : (~^reg171[3'b000100:1'b10]));
              reg193 <= wire133[4'b00111011:4'b00011001];
              reg194 <= reg154[3'b010110:2'b1010];
            end
          else
            begin
              reg190 <= reg179;
              reg191 <= reg166[5'b0011010000:4'b10101010];
              reg192 <= (8'hba);
              reg193 <= (&(|reg160[3'b101101:2'b0110]));
              reg194 <= reg172[4'b00011001:3'b010101];
            end
          reg195 <= ((~reg150) == $unsigned(reg165[1'b01:1'b11]));
        end
      else
        begin
          if (($signed({reg160,
              $signed((^reg194))}) << ({(reg188 < (reg192 >>> reg158)),
                  ((reg187 ? reg171 : wire132) >> (&wire136))} ?
              (((!reg169) & $signed((8'ha0))) ?
                  $unsigned((reg146 ? wire142 : (7'h42))) : ($unsigned(reg147) ?
                      (^(8'hb9)) : $signed(reg154))) : (reg140[2'b0111:2'b1011] <= reg189))))
            begin
              reg187 <= (reg180 && reg182);
              reg188 <= {$signed(reg164)};
            end
          else
            begin
              reg187 <= $signed((reg172[3'b001111:1'b00] ?
                  $unsigned((8'ha0)) : {$signed((reg176 ? reg171 : reg149))}));
            end
          reg189 <= {$unsigned($signed((reg138 ?
                  $signed(wire141) : (~|reg167))))};
          reg190 <= {$signed(reg150), (^reg186[4'b01101011:4'b11010])};
        end
    end
  assign wire196 = (~&$unsigned((reg178[4'b10011101:4'b01000] ^~ (~|$signed((8'hbd))))));
  always
    @(posedge clk) begin
      reg197 <= (~($unsigned(reg164[3'b000101:1'b00]) ?
          ((reg191[1'b01:1'b11] <<< ((8'hbb) | (8'hb5))) ?
              reg192 : $unsigned($unsigned(wire141))) : (~(reg157[3'b010110:2'b1010] ?
              $signed(reg155) : $unsigned((8'hba))))));
    end
  assign wire198 = (+((^~reg163[2'b0111:2'b1011]) ^ (((!reg178) * reg170) ?
                       {{reg166}} : reg182)));
  always
    @(posedge clk) begin
      reg199 <= ((reg147[4'b10001111:4'b01101100] ?
          {reg188[2'b1011:1'b00]} : wire141[1'b01:1'b11]) >> reg187[4'b01011010:4'b10101000]);
      reg200 <= reg158[3'b000100:2'b1011];
      if (($unsigned((^$unsigned((reg169 ?
          wire134 : (8'hae))))) & $signed((reg188[2'b1010:1'b11] ?
          (8'hb3) : (^(|(8'ha2)))))))
        begin
          reg201 <= (-{$unsigned((^~$signed(reg151)))});
          if ($unsigned($unsigned($signed($unsigned(reg188)))))
            begin
              reg202 <= ($unsigned($unsigned(reg177)) > $signed((8'ha0)));
            end
          else
            begin
              reg202 <= ($unsigned($unsigned((wire136[4'b01101001:3'b110110] <<< $signed(reg138)))) && {wire136[2'b1110:2'b0110]});
            end
          reg203 <= (reg193[1'b10:1'b10] ?
              reg150[3'b001111:1'b00] : reg164[3'b010101:3'b110100]);
          reg204 <= $signed(reg177);
        end
      else
        begin
          if ({($unsigned((8'hb1)) >> reg169[3'b100:2'b0110])})
            begin
              reg201 <= wire183[3'b101101:2'b0110];
              reg202 <= $signed(wire136[3'b000101:2'b0111]);
              reg203 <= reg202;
            end
          else
            begin
              reg201 <= (reg168[2'b0111:2'b10] & $signed($unsigned(reg174)));
            end
          reg204 <= reg155;
        end
    end
  assign wire205 = reg163[1'b01:1'b11];
  always
    @(posedge clk) begin
      reg206 <= (reg177 ?
          $signed($signed(($unsigned(reg190) ?
              wire205[1'b10:1'b10] : (~&(7'h40))))) : reg153[4'b01110:3'b101101]);
      if (($unsigned(reg145) + $signed(reg206)))
        begin
          if ($unsigned($signed(reg177)))
            begin
              reg207 <= ($signed({reg149, reg180[3'b011111:3'b110111]}) ?
                  ({((reg169 ? wire141 : reg147) <= (reg147 ?
                          reg197 : reg172))} < reg148) : reg153);
              reg208 <= ((&{$signed((!wire142)), {(wire205 == reg202)}}) ?
                  reg204[3'b010110:2'b1010] : reg161[4'b11011001:1'b10]);
              reg209 <= $unsigned(wire205[2'b1111:1'b11]);
            end
          else
            begin
              reg207 <= $signed(reg195);
            end
          reg210 <= $unsigned(reg152[3'b001110:1'b01]);
          reg211 <= $signed((^~((~|$signed((8'ha4))) && $unsigned((-reg171)))));
        end
      else
        begin
          if (wire196)
            begin
              reg207 <= {(!(reg163[2'b1011:1'b00] >= reg206[3'b111101:3'b010101]))};
            end
          else
            begin
              reg207 <= (^wire137);
              reg208 <= ($unsigned($unsigned((~&reg210))) ~^ ((((8'hbe) ?
                          $signed((8'hb5)) : $signed(reg194)) ?
                      reg185 : ({reg147} <= (reg201 < reg140))) ?
                  {reg204[1'b10:1'b10],
                      (~|reg143[2'b0111:2'b10])} : ($unsigned((reg147 ?
                      reg171 : wire184)) < (8'ha8))));
              reg209 <= $unsigned(({((reg139 >= reg202) ?
                          reg168 : $signed(reg197))} ?
                  (8'hb3) : (reg191[3'b000100:2'b1011] ?
                      reg206[5'b1011110100:3'b101110] : $signed($unsigned(reg160)))));
              reg210 <= ((reg147 < {$unsigned(wire184),
                      reg172[2'b0111:2'b10]}) ?
                  $signed($signed($unsigned(wire136))) : reg204);
              reg211 <= $signed(reg201);
            end
          reg212 <= reg178;
          reg213 <= ($signed($signed($signed(reg192[3'b100111:3'b11101]))) > {reg179,
              (reg208[2'b010:1'b10] ?
                  (reg161 ?
                      (reg178 ? reg144 : (8'hb8)) : (-reg201)) : (8'hb6))});
        end
      if ((reg177[4'b11101110:4'b10001010] ^~ (reg208 ?
          (reg186[3'b111111:2'b0111] <<< $signed({(8'hbb)})) : reg149)))
        begin
          reg214 <= $unsigned($unsigned($signed($unsigned(wire141))));
        end
      else
        begin
          reg214 <= {{$signed(reg157)}};
        end
    end
  assign wire215 = $unsigned(reg213);
  assign wire216 = $unsigned((!{$unsigned({reg181, reg155})}));
  always
    @(posedge clk) begin
      if (reg138[1'b11:1'b00])
        begin
          reg217 <= reg168;
          reg218 <= ({(reg180 > ($unsigned(wire142) ?
                      $signed(reg153) : (reg146 ^ reg176)))} ?
              (reg176 ? reg207[3'b110110:3'b101101] : reg144) : ($unsigned({(+reg140),
                      (reg178 >>> reg177)}) ?
                  reg139 : (!($signed((8'ha0)) ?
                      (reg139 * (8'hb9)) : (^~(8'had))))));
          if (((+reg217) ?
              $signed((&$unsigned($unsigned(reg157)))) : wire184[2'b1110:2'b0110]))
            begin
              reg219 <= $unsigned(wire142[1'b10:1'b10]);
              reg220 <= (reg180 ?
                  $unsigned($unsigned((+(reg174 ? reg201 : reg162)))) : reg194);
            end
          else
            begin
              reg219 <= (~&((reg160[1'b10:1'b10] ?
                      ((!reg188) ^ (~&(7'h40))) : $unsigned({reg208, reg180})) ?
                  wire133 : ($signed({reg160,
                      (8'hb9)}) >> $signed($signed(wire216)))));
              reg220 <= reg148;
              reg221 <= ((wire205[1'b01:1'b11] != $unsigned($signed((|wire135)))) ?
                  $unsigned((wire137 >= reg155[1'b11:1'b00])) : ({{(~&wire215),
                              wire216[2'b0111:2'b1011]},
                          $unsigned(reg154[4'b01011001:4'b00111001])} ?
                      (8'hb1) : wire136));
            end
        end
      else
        begin
          reg217 <= wire135;
          reg218 <= (-$signed((^(reg185[3'b101110:3'b011110] << reg164))));
        end
      reg222 <= reg217;
      if ((($signed($unsigned(reg197)) == (($unsigned(wire132) ?
              (reg180 <= reg163) : (reg193 ? reg154 : reg164)) ?
          $unsigned(reg138[2'b1110:2'b0110]) : (-(wire133 ?
              wire216 : reg164)))) >> reg176[1'b01:1'b11]))
        begin
          reg223 <= wire216;
          if ({(&{(reg155 && {reg189, reg190}),
                  (reg201[4'b01011010:4'b10101000] ? {reg175} : (reg146 >= reg171))}),
              (!{$signed({reg181})})})
            begin
              reg224 <= reg202[2'b010:1'b10];
              reg225 <= ((wire184[2'b010:1'b10] ?
                  reg151[3'b000100:1'b10] : $signed($unsigned((8'h9e)))) <<< $unsigned(reg154[4'b00111010:2'b0011]));
              reg226 <= $unsigned(reg164);
              reg227 <= reg166[4'b00011111:3'b001111];
            end
          else
            begin
              reg224 <= {(reg172[3'b000100:1'b01] >>> ($unsigned((^(8'hb0))) - ((wire134 ?
                      reg165 : reg222) <= $unsigned(reg224))))};
              reg225 <= reg224;
              reg226 <= $unsigned(wire183);
              reg227 <= (^{$signed($unsigned((reg178 ? (8'hab) : (7'h40)))),
                  reg143[4'b01011110:4'b001110]});
            end
          if (((reg221[4'b00111010:2'b0011] ?
              (reg172[3'b100111:3'b010110] ?
                  reg150 : reg208) : $unsigned(reg203[1'b01:1'b11])) >>> {wire132[1'b01:1'b11]}))
            begin
              reg228 <= $unsigned(($unsigned($unsigned((|reg176))) >> reg150[3'b100111:3'b010110]));
              reg229 <= $unsigned((^$signed((^~wire196))));
            end
          else
            begin
              reg228 <= $unsigned(($signed(reg210) ?
                  (|$signed((reg203 ?
                      (8'haa) : reg204))) : (((reg226 * reg168) + (~(8'h9c))) ?
                      reg195[4'b00101101:3'b000100] : $unsigned((reg154 == wire216)))));
            end
          if ($unsigned($unsigned(reg138[1'b11:1'b00])))
            begin
              reg230 <= (8'hb6);
              reg231 <= ($signed($signed($unsigned(reg153))) > {reg162[1'b01:1'b11]});
              reg232 <= reg156;
              reg233 <= wire216[2'b1010:1'b11];
              reg234 <= reg210[3'b010101:3'b110100];
            end
          else
            begin
              reg230 <= reg223[1'b10:1'b10];
            end
        end
      else
        begin
          reg223 <= (&{reg202, reg146});
        end
      reg235 <= $signed({(!reg143[4'b00111001:1'b01])});
      reg236 <= $signed((reg146[4'b11001011:4'b10101011] & reg153[3'b100111:2'b0010]));
    end
  assign wire237 = $unsigned(({reg189,
                       ((~|reg166) <= $signed(reg150))} >>> $unsigned($signed($unsigned(reg194)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module90
#( parameter param124 = (-((&((+(8'ha9)) ~^ ((7'h43) ~^ (8'haa)))) ? (+((~&(8'hb3)) > {(8'ha6)})) : {(-((8'hae) ? (8'hb1) : (8'hb1))), (~&((8'hbe) & (8'hbb)))}))
, parameter param125 = (({(param124 ? (param124 * param124) : param124), param124} < param124) > ({(|(^~param124))} == (~|((+(8'hb3)) ? (param124 ? param124 : param124) : param124)))) )
(y, clk, wire95, wire94, wire93, wire92, wire91);
  output wire [32'b00000000000000000000000101100000:32'b00000000000000000000000000000000] y;
  input wire [1'b10:1'b10] clk;
  input wire [4'b10101110:1'b10] wire95;
  input wire [5'b0101010011:1'b10] wire94;
  input wire [5'b1000110000:1'b0] wire93;
  input wire signed [3'b000100:1'b10] wire92;
  input wire signed [3'b000110:1'b00] wire91;
  wire [3'b000100:1'b10] wire123;
  wire signed [4'b10101110:1'b10] wire122;
  wire [3'b000101:1'b00] wire121;
  reg [3'b000101:1'b00] reg120 = (1'h0);
  reg [4'b10001101:1'b10] reg119 = (1'h0);
  reg signed [5'b0101010011:1'b10] reg118 = (1'h0);
  reg [3'b001111:1'b00] reg117 = (1'h0);
  reg signed [4'b01001111:1'b10] reg116 = (1'h0);
  reg [4'b10101110:1'b10] reg115 = (1'h0);
  reg [4'b00111100:1'b10] reg114 = (1'h0);
  reg [5'b1000110000:1'b0] reg113 = (1'h0);
  reg [5'b0101010011:1'b10] reg112 = (1'h0);
  reg [3'b000101:1'b00] reg111 = (1'h0);
  reg [5'b0001010010:1'b10] reg110 = (1'h0);
  reg [4'b01001111:1'b10] reg109 = (1'h0);
  reg [2'b1011:1'b00] reg108 = (1'h0);
  reg signed [4'b01001111:1'b10] reg107 = (1'h0);
  wire [5'b1110001:1'b10] wire106;
  reg signed [4'b11111000:1'b00] reg105 = (1'h0);
  reg [5'b1111010100:1'b00] reg104 = (1'h0);
  reg signed [5'b0001110101:1'b00] reg103 = (1'h0);
  reg signed [5'b0001010010:1'b10] reg102 = (1'h0);
  wire [2'b1011:1'b00] wire101;
  wire signed [4'b11111000:1'b00] wire100;
  wire [4'b00111100:1'b10] wire99;
  wire signed [5'b1000110000:1'b0] wire98;
  reg signed [5'b1000110000:1'b0] reg97 = (1'h0);
  reg signed [4'b10001101:1'b10] reg96 = (1'h0);
  assign y = {wire123,
                 wire122,
                 wire121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 wire106,
                 reg105,
                 reg104,
                 reg103,
                 reg102,
                 wire101,
                 wire100,
                 wire99,
                 wire98,
                 reg97,
                 reg96,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg96 <= ($unsigned(wire94) ^~ wire93[4'b11101000:3'b010110]);
      reg97 <= {$signed({reg96[3'b000100:2'b1011], wire92[2'b1111:1'b11]}), wire95};
    end
  assign wire98 = $unsigned((wire95 & ($unsigned(reg97) < wire92)));
  assign wire99 = ((8'ha0) ? (7'h44) : wire94);
  assign wire100 = (($signed(wire95[1'b10:1'b10]) ?
                       ($unsigned({wire91,
                           reg97}) <<< $unsigned($signed(wire94))) : wire98) ~^ wire98[4'b01011111:4'b11111110]);
  assign wire101 = wire98[1'b10:1'b10];
  always
    @(posedge clk) begin
      if (wire99)
        begin
          reg102 <= $signed($signed(wire99));
        end
      else
        begin
          if ({(~^reg102)})
            begin
              reg102 <= ({wire100} <= wire93[1'b10:1'b10]);
              reg103 <= $unsigned($unsigned(wire94[3'b000100:2'b1011]));
            end
          else
            begin
              reg102 <= ($signed({$signed((wire94 > wire99)),
                      $signed($unsigned(wire100))}) ?
                  {$unsigned(wire101)} : ((~|$unsigned((wire95 << wire95))) ?
                      wire100[3'b100111:3'b11101] : (wire101[1'b01:1'b11] >>> $signed((wire101 ?
                          wire100 : wire98)))));
            end
          reg104 <= ($signed($unsigned((wire91[3'b010101:3'b110100] == (wire94 ?
              wire101 : wire94)))) != $signed((wire100[2'b1111:1'b11] ?
              ((wire92 ^~ reg103) >>> (reg96 ^~ reg103)) : wire91[3'b110101:1'b11])));
          reg105 <= wire93;
        end
    end
  assign wire106 = (8'h9d);
  always
    @(posedge clk) begin
      if ($unsigned(wire106[4'b00001101:2'b1010]))
        begin
          reg107 <= (~^(+($signed(wire100[3'b001100:3'b001100]) ?
              (~$unsigned(reg103)) : wire95)));
        end
      else
        begin
          if ($unsigned({$signed((!(-(8'hbf))))}))
            begin
              reg107 <= wire98[4'b11101000:3'b010110];
              reg108 <= (~^$unsigned(wire100[3'b100:2'b0110]));
              reg109 <= (&wire101[1'b01:1'b11]);
              reg110 <= $unsigned(({(+wire100[4'b01111000:3'b100111])} + (~(wire91 ?
                  (8'hbc) : $unsigned(reg109)))));
            end
          else
            begin
              reg107 <= (((|(8'h9f)) ?
                      wire94[4'b11111000:1'b00] : (~|(reg105[3'b101110:3'b011110] + (wire106 ?
                          reg110 : (7'h43))))) ?
                  (~(!((wire106 ~^ wire91) ^~ wire95[4'b11011011:4'b01011000]))) : $unsigned($signed($unsigned($unsigned(wire95)))));
              reg108 <= (|((+($unsigned(reg96) ?
                  (wire99 ?
                      reg105 : (8'hae)) : $unsigned(reg109))) >= $signed((|{wire98,
                  reg97}))));
            end
        end
      reg111 <= $signed((&(((wire106 ^~ wire106) == (8'hbd)) ?
          $signed(reg104[4'b01101000:2'b0110]) : ($unsigned(reg102) <<< {(8'hac),
              wire91}))));
      reg112 <= $unsigned(wire101[1'b01:1'b11]);
      if ((7'h44))
        begin
          if ($signed(((~|reg107[4'b01101000:2'b0011]) ^ ((~^(wire93 >> reg109)) ?
              (reg104[5'b0001110001:2'b1011] || (wire93 ?
                  reg111 : wire106)) : ((|(8'ha1)) ?
                  wire93[4'b01011010:3'b100] : (~^reg103))))))
            begin
              reg113 <= $signed(wire95[1'b11:1'b00]);
              reg114 <= $unsigned(wire106);
              reg115 <= wire91;
              reg116 <= reg114[3'b001110:1'b01];
              reg117 <= reg97[4'b01111000:3'b100111];
            end
          else
            begin
              reg113 <= (wire101 ?
                  reg107[4'b11111100:4'b10111100] : ((~&$signed({reg113,
                      wire95})) ^ ($signed((reg110 + reg116)) ?
                      (~&(wire92 ? reg109 : reg107)) : (8'ha6))));
            end
          reg118 <= (&$signed((^$signed({wire93}))));
          reg119 <= reg107[4'b11111011:3'b110111];
          reg120 <= (8'hbf);
        end
      else
        begin
          reg113 <= reg113[4'b00101011:3'b100101];
          reg114 <= (|(reg104[3'b000101:1'b00] ^~ $signed({{wire106, wire98}})));
          reg115 <= reg116;
          if (reg97)
            begin
              reg116 <= reg108[2'b0111:2'b10];
              reg117 <= wire99[4'b00101010:1'b11];
              reg118 <= $unsigned($signed(($signed((8'hac)) ?
                  wire101 : ((wire94 * reg114) || (!wire93)))));
              reg119 <= reg107[4'b01101011:4'b11010];
            end
          else
            begin
              reg116 <= wire95;
              reg117 <= {({{reg102[2'b1010:1'b11], (^reg103)},
                      {(^wire99), reg107[4'b11101000:3'b010110]}} & {(7'h40)}),
                  ($signed(((reg118 * reg110) & $signed((8'had)))) ?
                      (^{(reg120 || reg108),
                          reg118}) : ($signed(wire92[1'b01:1'b11]) ~^ ((8'h9e) >= {reg116})))};
              reg118 <= (reg117[1'b10:1'b10] ?
                  {({$signed(wire91)} - $signed({wire100,
                          wire94}))} : $unsigned(reg105[1'b10:1'b10]));
              reg119 <= (reg104[5'b1001010010:4'b01001010] << wire99[2'b0111:2'b10]);
              reg120 <= ($unsigned($unsigned($signed($signed(wire95)))) ?
                  $signed((($signed(reg109) >> (reg119 ?
                      reg102 : (8'hb6))) || reg116[3'b100111:3'b010110])) : $signed($unsigned((reg96 < {reg112}))));
            end
        end
    end
  assign wire121 = {wire99[3'b000100:1'b10]};
  assign wire122 = ($signed($unsigned((~wire121))) ?
                       {(8'hb1),
                           reg105[2'b0111:2'b10]} : (((+reg103) ^~ (+$unsigned(wire101))) * wire94));
  assign wire123 = ((^~($signed((reg113 << reg113)) ?
                       ($signed(wire94) ?
                           wire93[4'b10101110:1'b10] : (&wire98)) : $signed(reg107))) ^~ $signed(reg103));
endmodule