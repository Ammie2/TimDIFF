(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param4556 = {((^~(|(8'hab))) ? ({(8'haa)} ? ((8'hae) ? (8'haa) : (8'ha7)) : (~|(8'hb6))) : (((8'hb2) ^ (8'ha3)) ^~ (^~(8'hb1))))} )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h7ea):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire3;
  input wire [(4'h9):(1'h0)] wire2;
  input wire signed [(4'hf):(1'h0)] wire1;
  input wire signed [(3'h5):(1'h0)] wire0;
  wire signed [(4'h8):(1'h0)] wire4555;
  wire signed [(4'h9):(1'h0)] wire4554;
  wire signed [(3'h6):(1'h0)] wire4553;
  reg signed [(4'h8):(1'h0)] reg4552 = (1'h0);
  reg [(5'h10):(1'h0)] reg4551 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4550 = (1'h0);
  reg [(4'hc):(1'h0)] reg4549 = (1'h0);
  reg [(2'h3):(1'h0)] reg4548 = (1'h0);
  reg [(2'h3):(1'h0)] reg4547 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4546 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4545 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4543 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4545 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4544 = (1'h0);
  reg [(3'h7):(1'h0)] reg4543 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4542 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4541 = (1'h0);
  reg [(4'h9):(1'h0)] reg4540 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4539 = (1'h0);
  reg [(4'h8):(1'h0)] reg4538 = (1'h0);
  reg [(4'h8):(1'h0)] reg4537 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4536 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4535 = (1'h0);
  reg [(4'hf):(1'h0)] reg4534 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4533 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4532 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4531 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4530 = (1'h0);
  reg [(4'h8):(1'h0)] reg4526 = (1'h0);
  reg [(4'h9):(1'h0)] reg4522 = (1'h0);
  reg [(4'he):(1'h0)] forvar4521 = (1'h0);
  reg [(4'he):(1'h0)] reg4529 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4528 = (1'h0);
  reg [(4'h9):(1'h0)] reg4527 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4526 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4525 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4524 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4523 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4522 = (1'h0);
  reg [(4'ha):(1'h0)] reg4521 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4520 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4519 = (1'h0);
  reg [(4'ha):(1'h0)] reg4518 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4517 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4516 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4515 = (1'h0);
  reg [(2'h2):(1'h0)] reg4514 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4513 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4511 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4510 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4512 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4511 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4510 = (1'h0);
  reg [(3'h5):(1'h0)] reg4509 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4508 = (1'h0);
  reg [(3'h5):(1'h0)] reg4507 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4506 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4505 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4504 = (1'h0);
  reg [(4'hb):(1'h0)] reg4494 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4493 = (1'h0);
  reg [(3'h5):(1'h0)] reg4503 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4502 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4501 = (1'h0);
  reg [(4'hb):(1'h0)] reg4500 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4499 = (1'h0);
  reg [(4'h8):(1'h0)] reg4498 = (1'h0);
  reg [(4'hd):(1'h0)] reg4497 = (1'h0);
  reg [(2'h3):(1'h0)] reg4496 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4495 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4494 = (1'h0);
  reg [(4'ha):(1'h0)] reg4493 = (1'h0);
  reg [(3'h6):(1'h0)] reg4492 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4491 = (1'h0);
  reg [(2'h2):(1'h0)] reg4490 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4489 = (1'h0);
  reg [(4'hf):(1'h0)] reg4488 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4487 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4486 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4485 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4484 = (1'h0);
  reg [(4'he):(1'h0)] reg4483 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4482 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4481 = (1'h0);
  reg [(3'h4):(1'h0)] reg4480 = (1'h0);
  reg [(4'he):(1'h0)] reg4479 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4478 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4477 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4475 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4472 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4476 = (1'h0);
  reg [(4'hc):(1'h0)] reg4475 = (1'h0);
  reg [(4'h9):(1'h0)] reg4474 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4473 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4472 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4471 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4470 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4469 = (1'h0);
  reg [(5'h10):(1'h0)] reg4468 = (1'h0);
  reg [(3'h7):(1'h0)] reg4467 = (1'h0);
  reg [(3'h7):(1'h0)] reg4466 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4465 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4464 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4462 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4457 = (1'h0);
  reg [(4'ha):(1'h0)] reg4464 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4463 = (1'h0);
  reg [(4'ha):(1'h0)] reg4462 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4458 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4455 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4454 = (1'h0);
  reg [(3'h5):(1'h0)] reg4453 = (1'h0);
  reg [(4'he):(1'h0)] reg4451 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4443 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4441 = (1'h0);
  reg [(3'h7):(1'h0)] reg4440 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4432 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4461 = (1'h0);
  reg [(4'hb):(1'h0)] reg4460 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4459 = (1'h0);
  reg [(4'ha):(1'h0)] reg4458 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4457 = (1'h0);
  reg [(4'hc):(1'h0)] reg4456 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4455 = (1'h0);
  reg [(4'hf):(1'h0)] reg4454 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4453 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4452 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4451 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4450 = (1'h0);
  reg [(3'h6):(1'h0)] reg4449 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4448 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4447 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4446 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4445 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4444 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4443 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4442 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4441 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4440 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4439 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4438 = (1'h0);
  reg [(4'hc):(1'h0)] reg4437 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4436 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4435 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4431 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4429 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4427 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4434 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4433 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4432 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4431 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4430 = (1'h0);
  reg [(4'hb):(1'h0)] reg4429 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4428 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4427 = (1'h0);
  reg [(2'h3):(1'h0)] reg4421 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4414 = (1'h0);
  reg [(4'h8):(1'h0)] reg4413 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4409 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4405 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4402 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4400 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4426 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4425 = (1'h0);
  reg [(5'h10):(1'h0)] reg4424 = (1'h0);
  reg [(4'ha):(1'h0)] reg4423 = (1'h0);
  reg [(3'h4):(1'h0)] reg4422 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4421 = (1'h0);
  reg [(3'h5):(1'h0)] reg4420 = (1'h0);
  reg [(4'h8):(1'h0)] reg4419 = (1'h0);
  reg [(4'he):(1'h0)] reg4418 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4417 = (1'h0);
  reg [(2'h3):(1'h0)] reg4416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4415 = (1'h0);
  reg [(4'h9):(1'h0)] reg4414 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4413 = (1'h0);
  reg [(5'h10):(1'h0)] reg4412 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4407 = (1'h0);
  reg [(5'h10):(1'h0)] reg4411 = (1'h0);
  reg [(4'he):(1'h0)] reg4410 = (1'h0);
  reg [(4'ha):(1'h0)] reg4409 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4408 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4407 = (1'h0);
  reg [(3'h6):(1'h0)] reg4406 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4405 = (1'h0);
  reg [(3'h4):(1'h0)] reg4404 = (1'h0);
  reg [(4'hb):(1'h0)] reg4403 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4402 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4401 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4400 = (1'h0);
  reg [(2'h2):(1'h0)] reg4399 = (1'h0);
  reg [(4'h8):(1'h0)] reg4398 = (1'h0);
  reg [(2'h3):(1'h0)] reg4397 = (1'h0);
  reg [(3'h5):(1'h0)] reg4396 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4395 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4394 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4393 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4392 = (1'h0);
  reg [(3'h5):(1'h0)] reg4391 = (1'h0);
  reg [(4'he):(1'h0)] forvar4390 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4389 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4388 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire4386;
  wire [(4'h8):(1'h0)] wire629;
  wire signed [(4'hf):(1'h0)] wire628;
  wire [(4'hc):(1'h0)] wire627;
  wire signed [(3'h5):(1'h0)] wire626;
  wire signed [(4'hb):(1'h0)] wire625;
  wire signed [(4'h8):(1'h0)] wire624;
  wire signed [(2'h3):(1'h0)] wire623;
  wire [(4'hb):(1'h0)] wire621;
  wire signed [(5'h10):(1'h0)] wire8;
  wire [(4'hb):(1'h0)] wire7;
  wire signed [(5'h10):(1'h0)] wire6;
  wire signed [(4'hf):(1'h0)] wire5;
  wire [(3'h6):(1'h0)] wire4;
  assign y = {wire4555,
                 wire4554,
                 wire4553,
                 reg4552,
                 reg4551,
                 reg4550,
                 reg4549,
                 reg4548,
                 reg4547,
                 reg4546,
                 forvar4545,
                 forvar4543,
                 reg4545,
                 reg4544,
                 reg4543,
                 reg4542,
                 forvar4541,
                 reg4540,
                 forvar4539,
                 reg4538,
                 reg4537,
                 reg4536,
                 reg4535,
                 reg4534,
                 reg4533,
                 forvar4532,
                 reg4531,
                 reg4530,
                 reg4526,
                 reg4522,
                 forvar4521,
                 reg4529,
                 reg4528,
                 reg4527,
                 forvar4526,
                 reg4525,
                 reg4524,
                 reg4523,
                 forvar4522,
                 reg4521,
                 forvar4520,
                 reg4519,
                 reg4518,
                 forvar4517,
                 reg4516,
                 reg4515,
                 reg4514,
                 reg4513,
                 forvar4511,
                 reg4510,
                 reg4512,
                 reg4511,
                 forvar4510,
                 reg4509,
                 reg4508,
                 reg4507,
                 reg4506,
                 forvar4505,
                 forvar4504,
                 reg4494,
                 forvar4493,
                 reg4503,
                 reg4502,
                 reg4501,
                 reg4500,
                 forvar4499,
                 reg4498,
                 reg4497,
                 reg4496,
                 reg4495,
                 forvar4494,
                 reg4493,
                 reg4492,
                 reg4491,
                 reg4490,
                 forvar4489,
                 reg4488,
                 reg4487,
                 reg4486,
                 reg4485,
                 reg4484,
                 reg4483,
                 reg4482,
                 reg4481,
                 reg4480,
                 reg4479,
                 forvar4478,
                 forvar4477,
                 forvar4475,
                 reg4472,
                 reg4476,
                 reg4475,
                 reg4474,
                 reg4473,
                 forvar4472,
                 reg4471,
                 forvar4470,
                 forvar4469,
                 reg4468,
                 reg4467,
                 reg4466,
                 reg4465,
                 forvar4464,
                 forvar4462,
                 forvar4457,
                 reg4464,
                 reg4463,
                 reg4462,
                 forvar4458,
                 forvar4455,
                 forvar4454,
                 reg4453,
                 reg4451,
                 forvar4443,
                 reg4441,
                 reg4440,
                 forvar4432,
                 reg4461,
                 reg4460,
                 reg4459,
                 reg4458,
                 reg4457,
                 reg4456,
                 reg4455,
                 reg4454,
                 forvar4453,
                 reg4452,
                 forvar4451,
                 reg4450,
                 reg4449,
                 reg4448,
                 reg4447,
                 reg4446,
                 reg4445,
                 forvar4444,
                 reg4443,
                 reg4442,
                 forvar4441,
                 forvar4440,
                 reg4439,
                 reg4438,
                 reg4437,
                 reg4436,
                 reg4435,
                 forvar4431,
                 forvar4429,
                 forvar4427,
                 reg4434,
                 reg4433,
                 reg4432,
                 reg4431,
                 reg4430,
                 reg4429,
                 reg4428,
                 reg4427,
                 reg4421,
                 forvar4414,
                 reg4413,
                 forvar4409,
                 forvar4405,
                 reg4402,
                 reg4400,
                 reg4426,
                 reg4425,
                 reg4424,
                 reg4423,
                 reg4422,
                 forvar4421,
                 reg4420,
                 reg4419,
                 reg4418,
                 forvar4417,
                 reg4416,
                 reg4415,
                 reg4414,
                 forvar4413,
                 reg4412,
                 forvar4407,
                 reg4411,
                 reg4410,
                 reg4409,
                 reg4408,
                 reg4407,
                 reg4406,
                 reg4405,
                 reg4404,
                 reg4403,
                 forvar4402,
                 reg4401,
                 forvar4400,
                 reg4399,
                 reg4398,
                 reg4397,
                 reg4396,
                 forvar4395,
                 reg4394,
                 reg4393,
                 reg4392,
                 reg4391,
                 forvar4390,
                 forvar4389,
                 forvar4388,
                 wire4386,
                 wire629,
                 wire628,
                 wire627,
                 wire626,
                 wire625,
                 wire624,
                 wire623,
                 wire621,
                 wire8,
                 wire7,
                 wire6,
                 wire5,
                 wire4,
                 (1'h0)};
  assign wire4 = $unsigned($signed($unsigned((wire0 ? wire2 : wire3))));
  assign wire5 = wire4[(2'h2):(1'h0)];
  assign wire6 = ($signed($signed((~|wire3))) <= wire3[(3'h4):(2'h2)]);
  assign wire7 = ($unsigned(wire3) ^~ (wire3[(4'he):(4'ha)] >> $signed((|(8'hb2)))));
  assign wire8 = $unsigned((wire5[(4'he):(3'h6)] ?
                     $unsigned(wire6) : wire0[(1'h0):(1'h0)]));
  module9 modinst622 (wire621, clk, wire4, wire0, wire8, wire2);
  assign wire623 = ((&wire8) ?
                       wire1 : ($signed($signed(wire621)) <= wire0[(3'h5):(2'h2)]));
  assign wire624 = $signed(wire3[(2'h2):(1'h1)]);
  assign wire625 = $signed({((-wire624) ?
                           $unsigned(wire624) : (wire7 ? wire7 : (8'hae)))});
  assign wire626 = $unsigned((~$unsigned($signed(wire1))));
  assign wire627 = ((((wire4 ? wire0 : wire7) ?
                           (~&(8'ha8)) : wire3[(4'hf):(2'h3)]) ?
                       (wire623[(2'h3):(2'h2)] >> (&wire623)) : $unsigned((!wire621))) && wire0[(1'h1):(1'h1)]);
  assign wire628 = wire624[(1'h0):(1'h0)];
  assign wire629 = {({(&wire4)} ?
                           (wire627 >>> $unsigned(wire6)) : $unsigned((wire624 == wire628)))};
  module630 modinst4387 (wire4386, clk, wire7, wire5, wire8, wire629);
  always
    @(posedge clk) begin
      for (forvar4388 = (1'h0); (forvar4388 < (2'h3)); forvar4388 = (forvar4388 + (1'h1)))
        begin
          if ({($unsigned(wire5[(2'h2):(1'h1)]) ?
                  wire0[(1'h0):(1'h0)] : wire621[(4'hb):(2'h3)])})
            begin
              for (forvar4389 = (1'h0); (forvar4389 < (1'h0)); forvar4389 = (forvar4389 + (1'h1)))
                begin
                  for (forvar4390 = (1'h0); (forvar4390 < (2'h2)); forvar4390 = (forvar4390 + (1'h1)))
                    begin
                      reg4391 <= $signed(wire627);
                      reg4392 <= wire625;
                      reg4393 <= (|(~^forvar4388));
                      reg4394 <= $signed($unsigned($signed($signed((8'hab)))));
                    end
                  for (forvar4395 = (1'h0); (forvar4395 < (1'h0)); forvar4395 = (forvar4395 + (1'h1)))
                    begin
                      reg4396 <= $signed($unsigned((^wire629[(4'h8):(3'h6)])));
                      reg4397 <= $signed((($signed(forvar4388) != forvar4390) ?
                          (^~(^~(8'h9f))) : $signed($signed(wire628))));
                      reg4398 <= (^~wire629[(2'h3):(2'h3)]);
                      reg4399 <= (~|$signed($unsigned($signed(wire623))));
                    end
                  for (forvar4400 = (1'h0); (forvar4400 < (1'h1)); forvar4400 = (forvar4400 + (1'h1)))
                    begin
                      reg4401 <= (wire4386 >>> ($unsigned((wire621 || forvar4389)) ?
                          $unsigned(wire624) : $unsigned({wire623})));
                    end
                  for (forvar4402 = (1'h0); (forvar4402 < (1'h1)); forvar4402 = (forvar4402 + (1'h1)))
                    begin
                      reg4403 <= forvar4390[(4'hb):(3'h4)];
                      reg4404 <= ($signed(((reg4399 + wire2) ?
                              $signed((8'hae)) : forvar4400[(3'h4):(1'h0)])) ?
                          $signed((+(forvar4390 ?
                              wire625 : wire7))) : (~|$signed(wire6)));
                      reg4405 <= (^$signed((~^(~&reg4403))));
                    end
                end
              if (((({(8'hae)} == wire624) ? reg4394 : wire3[(4'h8):(3'h4)]) ?
                  forvar4402[(2'h2):(1'h0)] : $unsigned($unsigned(reg4392))))
                begin
                  reg4406 <= wire621;
                  if ((wire0 ?
                      (reg4394 <<< $unsigned($signed(reg4403))) : ($unsigned((~|reg4403)) >>> (wire627[(1'h0):(1'h0)] ?
                          (wire625 - wire0) : (forvar4400 ~^ reg4394)))))
                    begin
                      reg4407 <= {$signed(forvar4400)};
                      reg4408 <= (^reg4391);
                      reg4409 <= $signed(wire624[(4'h8):(1'h1)]);
                    end
                  else
                    begin
                      reg4407 <= $unsigned($signed(((8'hb6) >= reg4392)));
                      reg4408 <= (+reg4404);
                      reg4409 <= reg4401[(1'h1):(1'h1)];
                      reg4410 <= {(8'hb8)};
                    end
                  reg4411 <= ($signed($unsigned((-(8'ha0)))) ?
                      (wire626[(2'h3):(1'h1)] ?
                          wire0[(1'h0):(1'h0)] : wire2) : $signed(wire3));
                end
              else
                begin
                  reg4406 <= (8'had);
                  for (forvar4407 = (1'h0); (forvar4407 < (2'h2)); forvar4407 = (forvar4407 + (1'h1)))
                    begin
                      reg4408 <= ((8'ha8) ?
                          (^~$signed((~wire8))) : (^(reg4410[(1'h0):(1'h0)] ?
                              (+forvar4390) : forvar4395)));
                    end
                end
              if ((forvar4400 ~^ ((wire624 ? (forvar4400 ~^ wire0) : reg4398) ?
                  forvar4400 : $signed(forvar4400[(3'h6):(3'h4)]))))
                begin
                  reg4412 <= $signed(forvar4388);
                end
              else
                begin
                  reg4412 <= (^{($unsigned(forvar4407) ?
                          (|wire627) : reg4409[(4'h8):(4'h8)])});
                  for (forvar4413 = (1'h0); (forvar4413 < (2'h3)); forvar4413 = (forvar4413 + (1'h1)))
                    begin
                      reg4414 <= (8'ha8);
                      reg4415 <= wire624[(1'h1):(1'h0)];
                      reg4416 <= (|$signed(reg4398));
                    end
                  for (forvar4417 = (1'h0); (forvar4417 < (2'h3)); forvar4417 = (forvar4417 + (1'h1)))
                    begin
                      reg4418 <= wire629[(4'h8):(3'h5)];
                      reg4419 <= ($signed($signed((reg4393 ?
                              reg4393 : reg4406))) ?
                          ((reg4397 >= {forvar4390}) & wire6) : forvar4390[(4'hd):(3'h5)]);
                      reg4420 <= ((wire4 << $signed($unsigned(forvar4417))) ?
                          $unsigned((+$unsigned(wire6))) : (^~($signed(forvar4402) ?
                              wire628[(3'h4):(3'h4)] : {wire629})));
                    end
                  for (forvar4421 = (1'h0); (forvar4421 < (1'h0)); forvar4421 = (forvar4421 + (1'h1)))
                    begin
                      reg4422 <= wire5;
                      reg4423 <= reg4409;
                      reg4424 <= reg4410;
                      reg4425 <= wire623[(1'h1):(1'h0)];
                    end
                end
              reg4426 <= wire7[(3'h4):(1'h1)];
            end
          else
            begin
              for (forvar4389 = (1'h0); (forvar4389 < (1'h1)); forvar4389 = (forvar4389 + (1'h1)))
                begin
                  for (forvar4390 = (1'h0); (forvar4390 < (2'h3)); forvar4390 = (forvar4390 + (1'h1)))
                    begin
                      reg4391 <= $signed(wire6[(3'h4):(3'h4)]);
                      reg4392 <= wire626;
                      reg4393 <= $signed((!(~reg4425)));
                      reg4394 <= reg4420[(2'h3):(1'h1)];
                    end
                  for (forvar4395 = (1'h0); (forvar4395 < (2'h2)); forvar4395 = (forvar4395 + (1'h1)))
                    begin
                      reg4396 <= $unsigned((reg4391 * $signed(reg4425)));
                      reg4397 <= reg4420;
                      reg4398 <= reg4401;
                      reg4399 <= (!(~|(+(reg4396 || (8'ha6)))));
                    end
                  if (wire628)
                    begin
                      reg4400 <= reg4398[(3'h7):(3'h5)];
                    end
                  else
                    begin
                      reg4400 <= $signed((((reg4425 ? reg4424 : forvar4417) ?
                              (wire3 == forvar4388) : forvar4388) ?
                          (wire628 ?
                              forvar4402[(2'h2):(1'h1)] : $unsigned(wire7)) : ((forvar4407 >= wire623) ?
                              wire8[(4'ha):(3'h4)] : (forvar4388 <<< reg4391))));
                      reg4401 <= ((~|forvar4417[(3'h6):(3'h5)]) ?
                          ($signed($unsigned(forvar4402)) ^ wire621) : forvar4390);
                      reg4402 <= $signed(($unsigned($unsigned(reg4416)) ?
                          $signed((reg4408 ?
                              forvar4417 : forvar4400)) : reg4396[(3'h4):(1'h0)]));
                    end
                  reg4403 <= reg4414;
                end
              reg4404 <= reg4424[(5'h10):(1'h1)];
              for (forvar4405 = (1'h0); (forvar4405 < (2'h3)); forvar4405 = (forvar4405 + (1'h1)))
                begin
                  if ((^reg4409))
                    begin
                      reg4406 <= (^{{{reg4403}}});
                    end
                  else
                    begin
                      reg4406 <= $signed(wire628[(2'h3):(2'h3)]);
                      reg4407 <= (|{wire1[(4'ha):(1'h1)]});
                      reg4408 <= wire3;
                    end
                  for (forvar4409 = (1'h0); (forvar4409 < (2'h2)); forvar4409 = (forvar4409 + (1'h1)))
                    begin
                      reg4410 <= wire1;
                      reg4411 <= ((((~&reg4397) || ((8'h9f) << reg4398)) ?
                          $signed($signed((8'hb5))) : wire625) + (8'h9f));
                      reg4412 <= $unsigned($signed($unsigned($signed(reg4415))));
                      reg4413 <= ((!(+(reg4412 ?
                          (8'h9d) : reg4397))) * (wire0[(3'h4):(1'h1)] ?
                          reg4398 : ($signed(reg4398) >> (!wire626))));
                    end
                  for (forvar4414 = (1'h0); (forvar4414 < (1'h0)); forvar4414 = (forvar4414 + (1'h1)))
                    begin
                      reg4415 <= (~^{(((8'hb8) ?
                              reg4424 : reg4399) ^ $signed(reg4397))});
                      reg4416 <= reg4404[(1'h0):(1'h0)];
                    end
                  for (forvar4417 = (1'h0); (forvar4417 < (2'h3)); forvar4417 = (forvar4417 + (1'h1)))
                    begin
                      reg4418 <= (8'hb6);
                      reg4419 <= wire0;
                      reg4420 <= $signed($signed((~&(reg4410 + forvar4407))));
                      reg4421 <= {$unsigned(forvar4395[(3'h5):(1'h0)])};
                    end
                end
            end
          if (($signed((8'ha8)) >>> $signed({(~^(8'hb0))})))
            begin
              if ({(~|reg4408)})
                begin
                  if ((reg4404[(2'h3):(1'h0)] ? reg4426[(4'h8):(4'h8)] : wire0))
                    begin
                      reg4427 <= (8'had);
                      reg4428 <= wire623[(1'h0):(1'h0)];
                      reg4429 <= $signed(wire624);
                    end
                  else
                    begin
                      reg4427 <= $signed(reg4400[(4'h8):(4'h8)]);
                    end
                  if (reg4423)
                    begin
                      reg4430 <= (({reg4415} <= wire4386) ?
                          forvar4407 : reg4424);
                    end
                  else
                    begin
                      reg4430 <= $unsigned(reg4429[(3'h6):(1'h1)]);
                      reg4431 <= ((&((wire625 ? reg4420 : reg4408) ?
                              wire5[(3'h5):(1'h1)] : (forvar4389 ~^ reg4400))) ?
                          $unsigned(($signed(reg4421) || $signed(reg4427))) : forvar4409[(4'hc):(2'h3)]);
                    end
                  reg4432 <= $unsigned(wire4386);
                  if ((|(-reg4420)))
                    begin
                      reg4433 <= reg4399[(1'h1):(1'h1)];
                      reg4434 <= $signed($unsigned($signed(reg4415[(3'h4):(2'h2)])));
                    end
                  else
                    begin
                      reg4433 <= {(!{$signed(forvar4407)})};
                    end
                end
              else
                begin
                  for (forvar4427 = (1'h0); (forvar4427 < (1'h0)); forvar4427 = (forvar4427 + (1'h1)))
                    begin
                      reg4428 <= reg4404;
                    end
                  for (forvar4429 = (1'h0); (forvar4429 < (2'h2)); forvar4429 = (forvar4429 + (1'h1)))
                    begin
                      reg4430 <= reg4431[(4'hb):(3'h6)];
                    end
                  for (forvar4431 = (1'h0); (forvar4431 < (1'h0)); forvar4431 = (forvar4431 + (1'h1)))
                    begin
                      reg4432 <= forvar4395[(3'h5):(1'h1)];
                      reg4433 <= $unsigned((forvar4390 ?
                          $unsigned($signed(reg4408)) : reg4399));
                      reg4434 <= wire0[(3'h5):(3'h4)];
                      reg4435 <= ((8'haf) ?
                          $unsigned(reg4405) : (~^($unsigned(reg4421) ?
                              (wire5 ?
                                  reg4427 : reg4392) : $unsigned(reg4422))));
                    end
                  if ((+reg4391[(3'h5):(1'h1)]))
                    begin
                      reg4436 <= ({(^reg4414)} ~^ reg4404[(3'h4):(1'h0)]);
                      reg4437 <= ((reg4403[(3'h6):(1'h1)] >>> forvar4417) ?
                          $signed($signed(reg4424)) : (reg4432[(4'h8):(3'h6)] > ($signed((8'had)) >> $unsigned(reg4391))));
                      reg4438 <= (|(~{$signed((8'ha7))}));
                    end
                  else
                    begin
                      reg4436 <= (^~($signed($unsigned(reg4410)) ?
                          (^(forvar4409 ^ wire0)) : (reg4430 * $unsigned((8'ha2)))));
                      reg4437 <= $unsigned((~|reg4432));
                      reg4438 <= ((((wire623 ^ forvar4409) & reg4428[(4'h9):(3'h6)]) ?
                          (!wire8[(4'ha):(2'h2)]) : (~&wire4386)) ^~ reg4412[(4'he):(3'h5)]);
                    end
                end
              reg4439 <= reg4428;
              for (forvar4440 = (1'h0); (forvar4440 < (2'h3)); forvar4440 = (forvar4440 + (1'h1)))
                begin
                  for (forvar4441 = (1'h0); (forvar4441 < (1'h1)); forvar4441 = (forvar4441 + (1'h1)))
                    begin
                      reg4442 <= (|{(8'haf)});
                      reg4443 <= forvar4395;
                    end
                  for (forvar4444 = (1'h0); (forvar4444 < (2'h3)); forvar4444 = (forvar4444 + (1'h1)))
                    begin
                      reg4445 <= ((($signed((8'hb6)) ? reg4391 : (^reg4400)) ?
                          (!$signed((8'hb5))) : {{reg4431}}) ~^ (!$unsigned((!(8'hb8)))));
                      reg4446 <= (wire629 ?
                          (^~{$unsigned(reg4400)}) : (^reg4419));
                      reg4447 <= $signed(reg4406[(1'h1):(1'h1)]);
                    end
                  if (($signed(reg4437) * $signed((8'ha9))))
                    begin
                      reg4448 <= wire6;
                      reg4449 <= {reg4419};
                    end
                  else
                    begin
                      reg4448 <= ($unsigned(((wire621 <<< wire629) ?
                              (reg4448 ?
                                  wire623 : forvar4388) : (forvar4402 - wire0))) ?
                          ((~^((8'hb4) != forvar4444)) == (8'h9e)) : $unsigned(reg4449));
                      reg4449 <= $signed($signed(((8'hae) ?
                          (reg4400 ?
                              wire6 : reg4402) : reg4424[(3'h6):(2'h2)])));
                      reg4450 <= (((reg4391 >> $unsigned((8'hb7))) ?
                          ({forvar4414} ?
                              $unsigned(reg4447) : (forvar4429 * reg4421)) : {$unsigned(wire627)}) >= forvar4405);
                    end
                end
              for (forvar4451 = (1'h0); (forvar4451 < (2'h2)); forvar4451 = (forvar4451 + (1'h1)))
                begin
                  reg4452 <= (!reg4414[(4'h9):(2'h2)]);
                  for (forvar4453 = (1'h0); (forvar4453 < (2'h2)); forvar4453 = (forvar4453 + (1'h1)))
                    begin
                      reg4454 <= reg4433;
                      reg4455 <= (~|reg4397[(1'h0):(1'h0)]);
                      reg4456 <= wire628[(3'h6):(3'h6)];
                      reg4457 <= $signed((~&$signed((forvar4451 <= reg4442))));
                    end
                  if (((($unsigned((8'ha8)) ^ reg4407[(3'h6):(2'h2)]) || {$signed(reg4455)}) ?
                      (reg4442[(4'h9):(1'h1)] ~^ $signed((wire3 ?
                          reg4402 : wire6))) : reg4433))
                    begin
                      reg4458 <= $signed((((^reg4439) + wire5[(4'hd):(3'h7)]) ?
                          (~^((8'hab) ~^ reg4411)) : $unsigned((8'h9d))));
                      reg4459 <= {$signed(forvar4427[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg4458 <= reg4434[(3'h6):(3'h4)];
                      reg4459 <= {$unsigned({$signed(reg4455)})};
                    end
                  if (forvar4427[(4'hb):(3'h7)])
                    begin
                      reg4460 <= $unsigned((reg4443 ?
                          ((|reg4429) ?
                              {wire6} : reg4458) : (|$signed(forvar4444))));
                      reg4461 <= reg4394;
                    end
                  else
                    begin
                      reg4460 <= {((^~(^~reg4433)) || $signed(((8'hb9) ?
                              forvar4421 : wire628)))};
                    end
                end
            end
          else
            begin
              for (forvar4427 = (1'h0); (forvar4427 < (1'h1)); forvar4427 = (forvar4427 + (1'h1)))
                begin
                  if ((&$unsigned($signed(wire625))))
                    begin
                      reg4428 <= {reg4404[(1'h0):(1'h0)]};
                      reg4429 <= wire8[(4'h8):(4'h8)];
                      reg4430 <= reg4415;
                      reg4431 <= reg4458[(3'h7):(3'h6)];
                    end
                  else
                    begin
                      reg4428 <= (^((~|$signed(forvar4413)) ?
                          ($signed(reg4391) == (|reg4393)) : $signed($signed(reg4397))));
                    end
                  for (forvar4432 = (1'h0); (forvar4432 < (2'h3)); forvar4432 = (forvar4432 + (1'h1)))
                    begin
                      reg4433 <= ((forvar4421 ~^ forvar4407) | $unsigned(reg4429[(4'h9):(4'h9)]));
                      reg4434 <= (forvar4429[(3'h5):(1'h0)] ?
                          (((reg4392 || reg4399) && {forvar4453}) || wire8) : $unsigned((reg4454 && $unsigned((8'hb5)))));
                      reg4435 <= $signed(((!(wire0 ~^ reg4447)) ?
                          wire624 : forvar4388[(1'h1):(1'h1)]));
                      reg4436 <= {($unsigned((|(8'had))) ?
                              (&wire625) : (reg4407[(3'h6):(3'h5)] ?
                                  {wire625} : $signed(reg4446)))};
                    end
                  if ((|(forvar4389 <= forvar4407[(2'h2):(1'h0)])))
                    begin
                      reg4437 <= (^forvar4388[(3'h4):(2'h3)]);
                      reg4438 <= forvar4440;
                      reg4439 <= {reg4415};
                    end
                  else
                    begin
                      reg4437 <= (8'h9c);
                    end
                  if ((8'hb0))
                    begin
                      reg4440 <= ((forvar4421[(3'h5):(2'h2)] ?
                              reg4413[(2'h2):(2'h2)] : $signed((~^wire621))) ?
                          reg4436 : $unsigned(forvar4451[(4'ha):(3'h7)]));
                      reg4441 <= {(8'ha2)};
                      reg4442 <= ((~((^~(8'ha4)) ?
                          {forvar4407} : $unsigned(reg4393))) <= wire4386);
                    end
                  else
                    begin
                      reg4440 <= ((~&forvar4402[(2'h2):(1'h1)]) ?
                          $signed($unsigned((&forvar4453))) : (!(!{reg4431})));
                      reg4441 <= $unsigned((reg4447[(1'h0):(1'h0)] ?
                          ($unsigned(forvar4441) <= wire3[(4'h8):(3'h6)]) : $signed({reg4433})));
                    end
                end
              for (forvar4443 = (1'h0); (forvar4443 < (2'h2)); forvar4443 = (forvar4443 + (1'h1)))
                begin
                  for (forvar4444 = (1'h0); (forvar4444 < (1'h1)); forvar4444 = (forvar4444 + (1'h1)))
                    begin
                      reg4445 <= ($signed($signed($unsigned(reg4436))) ?
                          $unsigned($unsigned($unsigned(reg4402))) : $unsigned($signed((reg4448 ^~ forvar4440))));
                      reg4446 <= $unsigned(reg4393[(3'h5):(2'h2)]);
                      reg4447 <= reg4455[(2'h3):(1'h1)];
                    end
                  reg4448 <= $unsigned(((!$unsigned(wire4)) != $unsigned((reg4402 ?
                      reg4409 : reg4460))));
                  reg4449 <= reg4427;
                  if ({reg4396[(1'h1):(1'h1)]})
                    begin
                      reg4450 <= (~|{reg4421[(1'h0):(1'h0)]});
                      reg4451 <= (($unsigned(reg4413[(3'h7):(1'h0)]) ^ {(reg4407 >= (8'hab))}) ?
                          (8'hb8) : ($signed($signed(reg4455)) ?
                              reg4410 : ($signed(reg4441) ?
                                  $unsigned(reg4450) : (~|reg4419))));
                      reg4452 <= $unsigned($unsigned({$unsigned(forvar4407)}));
                      reg4453 <= {wire629};
                    end
                  else
                    begin
                      reg4450 <= $signed($unsigned($signed(wire627[(1'h0):(1'h0)])));
                      reg4451 <= ((wire621[(3'h7):(2'h3)] ^~ $signed(reg4428)) ?
                          {$unsigned((^~reg4418))} : $unsigned(forvar4441[(4'ha):(1'h1)]));
                    end
                end
              for (forvar4454 = (1'h0); (forvar4454 < (2'h2)); forvar4454 = (forvar4454 + (1'h1)))
                begin
                  for (forvar4455 = (1'h0); (forvar4455 < (1'h1)); forvar4455 = (forvar4455 + (1'h1)))
                    begin
                      reg4456 <= $signed(wire0);
                    end
                end
              if ({(((!reg4410) ? $unsigned((8'ha2)) : {reg4425}) && reg4404)})
                begin
                  reg4457 <= ((8'hb1) - (^~forvar4388));
                  for (forvar4458 = (1'h0); (forvar4458 < (2'h3)); forvar4458 = (forvar4458 + (1'h1)))
                    begin
                      reg4459 <= reg4447;
                      reg4460 <= (^~($signed((+reg4423)) <<< ((reg4451 * reg4404) ?
                          reg4409[(3'h6):(2'h3)] : (^reg4452))));
                    end
                  if ((+(reg4435[(2'h3):(2'h2)] <= ($unsigned(forvar4431) ^~ (forvar4427 ?
                      wire625 : wire8)))))
                    begin
                      reg4461 <= ({$unsigned(wire7[(4'hb):(4'ha)])} * $signed(((reg4425 < reg4436) != $unsigned((8'had)))));
                      reg4462 <= $unsigned(reg4438);
                      reg4463 <= reg4455[(1'h1):(1'h1)];
                      reg4464 <= reg4430;
                    end
                  else
                    begin
                      reg4461 <= (-(^($signed(reg4421) >> reg4461[(4'he):(3'h7)])));
                      reg4462 <= $unsigned($unsigned(reg4452[(2'h2):(1'h0)]));
                      reg4463 <= $signed($signed(($signed(reg4448) ?
                          (+reg4397) : $unsigned((8'hb7)))));
                    end
                end
              else
                begin
                  for (forvar4457 = (1'h0); (forvar4457 < (2'h3)); forvar4457 = (forvar4457 + (1'h1)))
                    begin
                      reg4458 <= $signed(((~|reg4453) ?
                          (reg4448[(2'h3):(1'h0)] || (&forvar4431)) : (+$unsigned(reg4428))));
                      reg4459 <= $unsigned((^(reg4438 ?
                          {reg4456} : (~^(8'hac)))));
                      reg4460 <= reg4436[(3'h7):(2'h3)];
                      reg4461 <= reg4405[(3'h7):(2'h2)];
                    end
                  for (forvar4462 = (1'h0); (forvar4462 < (2'h2)); forvar4462 = (forvar4462 + (1'h1)))
                    begin
                      reg4463 <= reg4414;
                    end
                  for (forvar4464 = (1'h0); (forvar4464 < (2'h2)); forvar4464 = (forvar4464 + (1'h1)))
                    begin
                      reg4465 <= $unsigned((8'h9c));
                      reg4466 <= ((~|((reg4453 ? reg4411 : reg4392) ?
                          reg4433[(3'h4):(2'h3)] : (forvar4414 ?
                              wire629 : forvar4388))) + ((~^(!reg4418)) == $unsigned(reg4436[(1'h0):(1'h0)])));
                      reg4467 <= (reg4410[(4'hc):(1'h0)] ?
                          forvar4402 : (~(~&$signed((8'hb1)))));
                      reg4468 <= ((({forvar4417} ?
                                  (~&reg4449) : $signed(reg4451)) ?
                              (reg4423[(4'h8):(2'h2)] ^ {forvar4440}) : reg4425) ?
                          $unsigned({reg4398}) : $signed({forvar4441}));
                    end
                end
            end
        end
      for (forvar4469 = (1'h0); (forvar4469 < (2'h2)); forvar4469 = (forvar4469 + (1'h1)))
        begin
          for (forvar4470 = (1'h0); (forvar4470 < (2'h3)); forvar4470 = (forvar4470 + (1'h1)))
            begin
              if ($signed($unsigned(((reg4396 ? (8'haa) : forvar4429) ?
                  $signed((8'hb1)) : forvar4431))))
                begin
                  reg4471 <= (((reg4440 ^ $unsigned(reg4462)) | (~^wire0)) ?
                      {(8'hb0)} : $signed(((|forvar4414) <= (reg4425 ?
                          forvar4427 : wire4))));
                  for (forvar4472 = (1'h0); (forvar4472 < (2'h2)); forvar4472 = (forvar4472 + (1'h1)))
                    begin
                      reg4473 <= $unsigned((($signed(reg4411) && reg4466[(3'h6):(3'h4)]) ?
                          ($unsigned(forvar4395) ?
                              reg4453[(1'h1):(1'h0)] : $signed(reg4393)) : reg4471));
                    end
                  if (((($signed((8'had)) && (forvar4469 << (8'hac))) & ((~|forvar4400) << (forvar4453 >>> reg4416))) | $unsigned({((8'h9e) ?
                          reg4405 : forvar4443)})))
                    begin
                      reg4474 <= $signed((~(wire6[(4'hf):(4'he)] ?
                          $unsigned(wire627) : {reg4455})));
                      reg4475 <= $signed((reg4397 && $signed((+reg4397))));
                      reg4476 <= {(~^(~$signed(reg4452)))};
                    end
                  else
                    begin
                      reg4474 <= wire621;
                    end
                end
              else
                begin
                  if (wire625[(3'h5):(1'h1)])
                    begin
                      reg4471 <= (~^(((forvar4390 >= reg4468) ?
                              forvar4443[(1'h1):(1'h1)] : reg4468) ?
                          forvar4389[(3'h5):(2'h2)] : ($signed((8'hb8)) ?
                              reg4415[(2'h2):(2'h2)] : (wire623 && reg4434))));
                      reg4472 <= (8'hba);
                      reg4473 <= reg4410;
                    end
                  else
                    begin
                      reg4471 <= $unsigned(reg4422[(2'h2):(1'h0)]);
                      reg4472 <= reg4465[(1'h0):(1'h0)];
                      reg4473 <= forvar4413;
                      reg4474 <= (~&(&$signed((|reg4441))));
                    end
                  for (forvar4475 = (1'h0); (forvar4475 < (2'h2)); forvar4475 = (forvar4475 + (1'h1)))
                    begin
                      reg4476 <= wire7[(3'h4):(2'h3)];
                    end
                end
              for (forvar4477 = (1'h0); (forvar4477 < (1'h1)); forvar4477 = (forvar4477 + (1'h1)))
                begin
                  for (forvar4478 = (1'h0); (forvar4478 < (2'h3)); forvar4478 = (forvar4478 + (1'h1)))
                    begin
                      reg4479 <= (~&forvar4470);
                      reg4480 <= $unsigned((((forvar4454 ?
                              forvar4454 : reg4471) ?
                          (!reg4430) : (~|reg4432)) >> ($signed(reg4465) && $unsigned(reg4473))));
                      reg4481 <= $unsigned((($unsigned(reg4472) <<< (forvar4390 ?
                              reg4456 : reg4460)) ?
                          $signed($signed((8'hb4))) : $unsigned((~^forvar4395))));
                      reg4482 <= (^forvar4440[(3'h7):(1'h0)]);
                    end
                  if ($signed(reg4393[(3'h6):(2'h2)]))
                    begin
                      reg4483 <= (~$unsigned(reg4437[(4'hc):(1'h1)]));
                    end
                  else
                    begin
                      reg4483 <= $unsigned(wire6[(3'h7):(2'h2)]);
                      reg4484 <= forvar4431[(1'h1):(1'h0)];
                      reg4485 <= {forvar4441};
                      reg4486 <= {reg4450[(2'h2):(1'h1)]};
                    end
                  if ($signed($unsigned(forvar4431[(1'h1):(1'h1)])))
                    begin
                      reg4487 <= ($unsigned($unsigned((8'h9e))) >= $signed(reg4416[(1'h0):(1'h0)]));
                      reg4488 <= (wire3[(4'he):(4'he)] || (-$signed(reg4391[(3'h5):(2'h3)])));
                    end
                  else
                    begin
                      reg4487 <= $unsigned($signed((~|$signed(reg4475))));
                    end
                  for (forvar4489 = (1'h0); (forvar4489 < (2'h3)); forvar4489 = (forvar4489 + (1'h1)))
                    begin
                      reg4490 <= (((8'ha7) >>> (reg4432 ?
                              (!reg4453) : reg4459)) ?
                          $unsigned($signed((reg4432 ?
                              reg4468 : reg4394))) : reg4418[(2'h2):(1'h0)]);
                      reg4491 <= reg4474[(2'h3):(2'h2)];
                      reg4492 <= (((8'hae) < (reg4428[(3'h7):(3'h4)] != {(8'had)})) >> $signed($unsigned($signed((8'hb1)))));
                    end
                end
              if (({$unsigned((reg4425 << reg4462))} < ((^~{reg4415}) ?
                  wire5 : $unsigned(reg4423))))
                begin
                  if ($signed(((^reg4414) ? $unsigned({(8'haf)}) : reg4396)))
                    begin
                      reg4493 <= ((((reg4401 != (8'h9f)) ?
                              $unsigned(forvar4455) : (-forvar4429)) >> (+wire1[(4'hc):(4'h8)])) ?
                          reg4416 : ((+(reg4464 ?
                              (8'hb8) : forvar4427)) <= reg4404));
                    end
                  else
                    begin
                      reg4493 <= ($signed((reg4468 ^ ((8'h9d) ?
                          forvar4407 : reg4462))) == ((~&reg4402) ?
                          (~(forvar4405 <<< reg4466)) : (-reg4488[(3'h5):(3'h5)])));
                    end
                  for (forvar4494 = (1'h0); (forvar4494 < (1'h1)); forvar4494 = (forvar4494 + (1'h1)))
                    begin
                      reg4495 <= {$unsigned(((~|wire4) ?
                              reg4474[(4'h9):(4'h9)] : (+forvar4462)))};
                      reg4496 <= (~&$signed(reg4463));
                      reg4497 <= (forvar4432 == $unsigned($signed($unsigned(reg4393))));
                      reg4498 <= (8'h9e);
                    end
                  for (forvar4499 = (1'h0); (forvar4499 < (1'h0)); forvar4499 = (forvar4499 + (1'h1)))
                    begin
                      reg4500 <= wire0[(1'h0):(1'h0)];
                      reg4501 <= forvar4413[(2'h2):(1'h1)];
                      reg4502 <= ((reg4393[(2'h3):(1'h1)] ?
                              (8'h9d) : reg4427[(2'h3):(2'h2)]) ?
                          (reg4433 ?
                              reg4402[(3'h5):(3'h5)] : (reg4447 ?
                                  reg4398 : $unsigned(wire623))) : $unsigned(wire4[(3'h6):(2'h2)]));
                      reg4503 <= {(^((wire4386 & (8'ha2)) >= (~|reg4474)))};
                    end
                end
              else
                begin
                  for (forvar4493 = (1'h0); (forvar4493 < (2'h3)); forvar4493 = (forvar4493 + (1'h1)))
                    begin
                      reg4494 <= forvar4455[(2'h2):(1'h1)];
                    end
                end
            end
          for (forvar4504 = (1'h0); (forvar4504 < (1'h1)); forvar4504 = (forvar4504 + (1'h1)))
            begin
              if (forvar4405)
                begin
                  for (forvar4505 = (1'h0); (forvar4505 < (2'h2)); forvar4505 = (forvar4505 + (1'h1)))
                    begin
                      reg4506 <= $unsigned((!reg4399));
                      reg4507 <= reg4474;
                      reg4508 <= wire4386[(1'h0):(1'h0)];
                      reg4509 <= (((&reg4462) ?
                              $unsigned((reg4502 ?
                                  (8'hba) : reg4419)) : (^~(forvar4388 == wire623))) ?
                          $unsigned($unsigned($signed(reg4438))) : reg4399);
                    end
                  for (forvar4510 = (1'h0); (forvar4510 < (1'h0)); forvar4510 = (forvar4510 + (1'h1)))
                    begin
                      reg4511 <= ({(^(forvar4489 | reg4412))} ?
                          $signed((reg4474 << $signed(wire624))) : {$signed(reg4403[(4'ha):(2'h3)])});
                      reg4512 <= (!$signed(((^~forvar4407) ?
                          $unsigned(reg4485) : reg4443[(2'h2):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar4505 = (1'h0); (forvar4505 < (1'h0)); forvar4505 = (forvar4505 + (1'h1)))
                    begin
                      reg4506 <= $signed({(|wire1[(1'h1):(1'h1)])});
                      reg4507 <= wire623;
                      reg4508 <= ($unsigned(((wire7 | reg4441) ?
                              (wire627 ?
                                  forvar4432 : reg4493) : {forvar4455})) ?
                          reg4496[(2'h2):(1'h0)] : ((forvar4477 ?
                              (8'hac) : $unsigned((8'ha3))) > ((forvar4494 ?
                                  reg4450 : reg4447) ?
                              (reg4428 ?
                                  reg4468 : reg4468) : reg4413[(4'h8):(4'h8)])));
                      reg4509 <= ((((reg4484 ^ (8'hb5)) ?
                                  $signed((8'h9c)) : wire627[(3'h6):(1'h0)]) ?
                              $signed((reg4439 * forvar4475)) : (reg4460[(4'h9):(3'h4)] | reg4453[(3'h5):(2'h3)])) ?
                          $signed(reg4488) : (8'haf));
                    end
                  reg4510 <= $signed($unsigned($unsigned(((8'ha8) ?
                      reg4453 : reg4485))));
                  for (forvar4511 = (1'h0); (forvar4511 < (1'h1)); forvar4511 = (forvar4511 + (1'h1)))
                    begin
                      reg4512 <= {(8'ha5)};
                      reg4513 <= reg4453[(2'h3):(2'h2)];
                      reg4514 <= (reg4451[(4'he):(4'ha)] ?
                          (8'ha1) : (^~reg4475[(1'h0):(1'h0)]));
                      reg4515 <= $unsigned(reg4420[(2'h3):(1'h1)]);
                    end
                  reg4516 <= $unsigned($unsigned((~(+reg4495))));
                end
            end
          for (forvar4517 = (1'h0); (forvar4517 < (2'h3)); forvar4517 = (forvar4517 + (1'h1)))
            begin
              if (($unsigned(forvar4429[(4'h8):(1'h1)]) ?
                  ((~|(reg4408 ? reg4514 : reg4472)) ?
                      reg4460[(4'h9):(3'h6)] : ((forvar4427 && reg4416) + (reg4484 ?
                          (8'hb2) : forvar4414))) : $signed(($signed(wire621) ?
                      $signed(reg4391) : (+forvar4499)))))
                begin
                  if ((&$signed($signed({(8'hac)}))))
                    begin
                      reg4518 <= reg4438;
                      reg4519 <= (reg4442 ?
                          reg4501[(2'h3):(2'h3)] : reg4423[(3'h6):(1'h1)]);
                    end
                  else
                    begin
                      reg4518 <= {{reg4509[(3'h4):(2'h3)]}};
                    end
                end
              else
                begin
                  reg4518 <= reg4443;
                  reg4519 <= $unsigned(forvar4470);
                end
            end
          for (forvar4520 = (1'h0); (forvar4520 < (1'h1)); forvar4520 = (forvar4520 + (1'h1)))
            begin
              if (reg4406)
                begin
                  reg4521 <= reg4408;
                  for (forvar4522 = (1'h0); (forvar4522 < (2'h2)); forvar4522 = (forvar4522 + (1'h1)))
                    begin
                      reg4523 <= $unsigned((^reg4501));
                      reg4524 <= ($unsigned($signed(forvar4413[(2'h2):(1'h0)])) && {$unsigned({forvar4510})});
                    end
                  reg4525 <= (8'ha1);
                  for (forvar4526 = (1'h0); (forvar4526 < (2'h2)); forvar4526 = (forvar4526 + (1'h1)))
                    begin
                      reg4527 <= ((^~reg4411[(3'h6):(3'h4)]) > $unsigned((+$signed(forvar4402))));
                      reg4528 <= $signed((~|{wire621}));
                      reg4529 <= (!(8'ha1));
                    end
                end
              else
                begin
                  for (forvar4521 = (1'h0); (forvar4521 < (1'h0)); forvar4521 = (forvar4521 + (1'h1)))
                    begin
                      reg4522 <= reg4434;
                      reg4523 <= reg4414;
                    end
                  if (forvar4432[(4'hc):(2'h3)])
                    begin
                      reg4524 <= ($unsigned(($signed((8'hae)) >>> $signed(reg4472))) ?
                          reg4414[(4'h8):(2'h2)] : $unsigned($unsigned($signed((8'hac)))));
                      reg4525 <= {$signed({(reg4497 ? forvar4413 : reg4391)})};
                      reg4526 <= forvar4520[(3'h7):(3'h5)];
                      reg4527 <= (^~$signed(reg4396));
                    end
                  else
                    begin
                      reg4524 <= (&(($unsigned((8'ha8)) ^~ (reg4456 > (8'hae))) ?
                          $signed(forvar4478[(1'h0):(1'h0)]) : $unsigned({reg4448})));
                    end
                  if ($unsigned(forvar4499))
                    begin
                      reg4528 <= reg4481;
                      reg4529 <= reg4494[(4'hb):(1'h1)];
                      reg4530 <= {(((&forvar4388) ?
                              (^reg4456) : (~reg4495)) || ((reg4467 ?
                                  forvar4395 : forvar4389) ?
                              {forvar4443} : reg4432))};
                      reg4531 <= {$signed((forvar4427 ?
                              forvar4414[(3'h7):(1'h0)] : (forvar4405 ?
                                  (8'hb3) : reg4445)))};
                    end
                  else
                    begin
                      reg4528 <= $signed($signed(((reg4429 ?
                          reg4450 : reg4493) < (reg4531 ? (8'ha0) : reg4524))));
                    end
                end
              for (forvar4532 = (1'h0); (forvar4532 < (2'h2)); forvar4532 = (forvar4532 + (1'h1)))
                begin
                  if ($signed((($unsigned(forvar4505) ?
                          reg4454 : (reg4392 ? reg4523 : reg4514)) ?
                      ((reg4429 << reg4450) | $unsigned(forvar4489)) : (reg4495[(1'h0):(1'h0)] >= (!reg4460)))))
                    begin
                      reg4533 <= (^$unsigned($signed((^~reg4432))));
                      reg4534 <= {{((reg4516 ?
                                  reg4393 : reg4433) + (forvar4432 ~^ wire628))}};
                    end
                  else
                    begin
                      reg4533 <= $unsigned((forvar4429 != (^~(wire4386 >>> (8'hab)))));
                      reg4534 <= forvar4443;
                      reg4535 <= ($unsigned({reg4484}) == $signed(forvar4522[(3'h5):(3'h4)]));
                    end
                  if (reg4473[(3'h6):(2'h3)])
                    begin
                      reg4536 <= (reg4427 != reg4396[(1'h1):(1'h0)]);
                      reg4537 <= $signed(($signed($unsigned(forvar4470)) ?
                          ((reg4500 + reg4391) ?
                              ((8'h9e) & wire0) : $unsigned(reg4433)) : $unsigned(reg4519[(3'h6):(2'h2)])));
                      reg4538 <= (~(|$unsigned($signed((8'h9c)))));
                    end
                  else
                    begin
                      reg4536 <= reg4420[(2'h3):(2'h2)];
                      reg4537 <= (-({reg4454[(4'ha):(1'h0)]} >>> (reg4423 ?
                          (reg4506 ^ reg4466) : ((8'hb5) <= (8'hba)))));
                    end
                end
              for (forvar4539 = (1'h0); (forvar4539 < (1'h1)); forvar4539 = (forvar4539 + (1'h1)))
                begin
                  reg4540 <= $signed(($signed($unsigned(reg4446)) ?
                      reg4391[(1'h1):(1'h0)] : ({(8'haa)} + (wire6 ?
                          forvar4389 : (8'ha8)))));
                  for (forvar4541 = (1'h0); (forvar4541 < (1'h1)); forvar4541 = (forvar4541 + (1'h1)))
                    begin
                      reg4542 <= reg4436;
                    end
                end
              if (wire0[(2'h3):(2'h2)])
                begin
                  if ($unsigned(((reg4482[(3'h5):(2'h3)] >> (forvar4517 >>> forvar4431)) < reg4441)))
                    begin
                      reg4543 <= ($unsigned(wire1) ?
                          forvar4511 : $unsigned($signed({reg4530})));
                      reg4544 <= (reg4427 <<< reg4528[(2'h3):(2'h3)]);
                      reg4545 <= ($unsigned(reg4442) ?
                          $signed($signed($unsigned(reg4400))) : reg4506);
                    end
                  else
                    begin
                      reg4543 <= $unsigned(reg4393);
                    end
                end
              else
                begin
                  for (forvar4543 = (1'h0); (forvar4543 < (2'h2)); forvar4543 = (forvar4543 + (1'h1)))
                    begin
                      reg4544 <= $unsigned($unsigned(wire7));
                    end
                  for (forvar4545 = (1'h0); (forvar4545 < (2'h3)); forvar4545 = (forvar4545 + (1'h1)))
                    begin
                      reg4546 <= $unsigned($unsigned(((+reg4436) < forvar4520[(2'h3):(2'h3)])));
                      reg4547 <= $unsigned((8'ha4));
                    end
                  if ({(^$unsigned((&forvar4511)))})
                    begin
                      reg4548 <= {((&reg4411[(4'ha):(2'h2)]) < (^~reg4540[(3'h6):(3'h5)]))};
                      reg4549 <= $unsigned(((~^(reg4400 ?
                              reg4413 : forvar4405)) ?
                          ({wire625} ?
                              (reg4430 ?
                                  reg4528 : forvar4478) : (reg4392 ^ forvar4440)) : (reg4442 ?
                              (reg4500 ^ reg4514) : ((8'hb6) - reg4405))));
                      reg4550 <= reg4451;
                      reg4551 <= {(({reg4409} && (^reg4407)) * reg4461)};
                    end
                  else
                    begin
                      reg4548 <= (8'haf);
                      reg4549 <= (((forvar4493 > reg4548) ?
                          reg4420 : (~^wire623[(1'h0):(1'h0)])) * (~^{(forvar4545 == reg4446)}));
                    end
                end
            end
        end
      if ((reg4460[(1'h0):(1'h0)] ?
          $unsigned((8'hb5)) : ($signed($unsigned(reg4403)) ?
              reg4433[(2'h2):(1'h1)] : (+$signed(reg4459)))))
        begin
          reg4552 <= (forvar4494 != (^(+(8'hb0))));
        end
      else
        begin
          reg4552 <= $signed(reg4476);
        end
    end
  assign wire4553 = reg4430[(1'h1):(1'h0)];
  assign wire4554 = $unsigned((8'ha7));
  assign wire4555 = (((&{forvar4444}) ?
                        $unsigned((reg4513 ? reg4542 : reg4536)) : {((8'hb0) ?
                                reg4473 : forvar4444)}) != (!reg4472));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module630
#( parameter param4385 = ({(~((8'h9e) ? (8'hae) : (8'had)))} ? ((((8'ha8) ^~ (8'hb3)) ? (!(8'hb9)) : ((8'ha9) >>> (8'ha5))) + {{(8'haa)}}) : (-{(-(8'ha1))})) )
(y, clk, wire634, wire633, wire632, wire631);
  output wire [(32'h941):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire634;
  input wire signed [(4'hf):(1'h0)] wire633;
  input wire [(3'h4):(1'h0)] wire632;
  input wire [(3'h5):(1'h0)] wire631;
  wire [(3'h7):(1'h0)] wire4384;
  wire [(4'he):(1'h0)] wire4383;
  reg signed [(4'hb):(1'h0)] reg4382 = (1'h0);
  reg [(4'h8):(1'h0)] reg4381 = (1'h0);
  reg [(3'h5):(1'h0)] reg4380 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4379 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4378 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4377 = (1'h0);
  reg [(5'h10):(1'h0)] reg4376 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4375 = (1'h0);
  reg [(3'h7):(1'h0)] reg4373 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4368 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4365 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4375 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4374 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4373 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4372 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4371 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4370 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4369 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4368 = (1'h0);
  reg [(4'hf):(1'h0)] reg4367 = (1'h0);
  reg [(4'ha):(1'h0)] reg4366 = (1'h0);
  reg [(4'hf):(1'h0)] reg4365 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4356 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4364 = (1'h0);
  reg [(3'h7):(1'h0)] reg4363 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4362 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4361 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4360 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4359 = (1'h0);
  reg [(2'h3):(1'h0)] reg4358 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4357 = (1'h0);
  reg [(4'hf):(1'h0)] reg4356 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4355 = (1'h0);
  reg [(3'h6):(1'h0)] reg4354 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4353 = (1'h0);
  reg [(3'h7):(1'h0)] reg4352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4351 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4350 = (1'h0);
  reg [(3'h5):(1'h0)] reg4349 = (1'h0);
  reg [(4'hd):(1'h0)] reg4348 = (1'h0);
  reg [(4'hb):(1'h0)] reg4347 = (1'h0);
  reg [(4'hc):(1'h0)] reg4346 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4345 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4344 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4343 = (1'h0);
  reg [(4'ha):(1'h0)] reg4342 = (1'h0);
  reg [(4'hc):(1'h0)] reg4341 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4340 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4339 = (1'h0);
  reg [(4'h8):(1'h0)] reg4338 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4337 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4336 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4335 = (1'h0);
  reg [(4'hb):(1'h0)] reg4334 = (1'h0);
  reg [(4'h9):(1'h0)] reg4333 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4331 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4332 = (1'h0);
  reg [(4'h8):(1'h0)] reg4331 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4330 = (1'h0);
  reg [(4'he):(1'h0)] forvar4329 = (1'h0);
  reg [(4'ha):(1'h0)] reg4328 = (1'h0);
  reg [(4'ha):(1'h0)] reg4327 = (1'h0);
  reg [(4'h8):(1'h0)] reg4326 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4325 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4324 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4323 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4322 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4300 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4306 = (1'h0);
  reg [(4'hc):(1'h0)] reg4321 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4320 = (1'h0);
  reg [(2'h2):(1'h0)] reg4319 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4318 = (1'h0);
  reg [(4'hb):(1'h0)] reg4317 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4316 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4315 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4314 = (1'h0);
  reg [(4'he):(1'h0)] reg4313 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4312 = (1'h0);
  reg [(4'h9):(1'h0)] reg4311 = (1'h0);
  reg [(4'hc):(1'h0)] reg4310 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4309 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4308 = (1'h0);
  reg [(4'h9):(1'h0)] reg4307 = (1'h0);
  reg [(3'h5):(1'h0)] reg4306 = (1'h0);
  reg [(3'h5):(1'h0)] reg4305 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4304 = (1'h0);
  reg [(4'hb):(1'h0)] reg4303 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4302 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4301 = (1'h0);
  reg [(5'h10):(1'h0)] reg4300 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4299 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4298 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4297 = (1'h0);
  reg [(4'hf):(1'h0)] reg4290 = (1'h0);
  reg [(3'h7):(1'h0)] reg4296 = (1'h0);
  reg [(4'h9):(1'h0)] reg4295 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4294 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4293 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4292 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4291 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4290 = (1'h0);
  reg [(3'h6):(1'h0)] reg4289 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4288 = (1'h0);
  reg [(4'h9):(1'h0)] reg4287 = (1'h0);
  reg [(4'h9):(1'h0)] reg4286 = (1'h0);
  reg [(2'h2):(1'h0)] reg4285 = (1'h0);
  reg [(4'he):(1'h0)] forvar4284 = (1'h0);
  reg [(2'h3):(1'h0)] reg4283 = (1'h0);
  reg [(4'h9):(1'h0)] reg4282 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4281 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4280 = (1'h0);
  reg [(3'h4):(1'h0)] reg4279 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4278 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4277 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4276 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4275 = (1'h0);
  reg [(4'hb):(1'h0)] reg4274 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4273 = (1'h0);
  reg [(4'h9):(1'h0)] reg4272 = (1'h0);
  reg [(2'h2):(1'h0)] reg4271 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4270 = (1'h0);
  reg [(4'h9):(1'h0)] reg4269 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4268 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4267 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4266 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4265 = (1'h0);
  reg [(4'hf):(1'h0)] reg4264 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4263 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4247 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4262 = (1'h0);
  reg [(4'ha):(1'h0)] reg4261 = (1'h0);
  reg [(3'h5):(1'h0)] reg4260 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4259 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4258 = (1'h0);
  reg [(4'ha):(1'h0)] reg4257 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4256 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4255 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4254 = (1'h0);
  reg [(4'hb):(1'h0)] reg4253 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4252 = (1'h0);
  reg [(4'h8):(1'h0)] reg4251 = (1'h0);
  reg [(4'hd):(1'h0)] reg4250 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4249 = (1'h0);
  reg [(3'h5):(1'h0)] reg4248 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4247 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4246 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4245 = (1'h0);
  reg [(3'h6):(1'h0)] reg4244 = (1'h0);
  reg [(4'hc):(1'h0)] reg4243 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4242 = (1'h0);
  reg [(4'hb):(1'h0)] reg4241 = (1'h0);
  reg [(3'h5):(1'h0)] reg4240 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4239 = (1'h0);
  reg [(4'he):(1'h0)] reg4238 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4237 = (1'h0);
  reg [(4'hb):(1'h0)] reg4236 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4235 = (1'h0);
  reg [(4'he):(1'h0)] reg4234 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4233 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4232 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4231 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4230 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4229 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4228 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4227 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4226 = (1'h0);
  reg [(3'h4):(1'h0)] reg4225 = (1'h0);
  reg [(4'hb):(1'h0)] reg4224 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4223 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4222 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4221 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4220 = (1'h0);
  reg [(4'h8):(1'h0)] reg4219 = (1'h0);
  reg [(3'h6):(1'h0)] reg4218 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4217 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4216 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4215 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4214 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4213 = (1'h0);
  reg [(5'h10):(1'h0)] reg4212 = (1'h0);
  reg [(2'h2):(1'h0)] reg4211 = (1'h0);
  reg [(2'h3):(1'h0)] reg4210 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4209 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4208 = (1'h0);
  reg [(2'h2):(1'h0)] reg4207 = (1'h0);
  reg [(4'hf):(1'h0)] reg4206 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4205 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4204 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4203 = (1'h0);
  reg [(3'h4):(1'h0)] reg4202 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4201 = (1'h0);
  reg [(4'hb):(1'h0)] reg4200 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4199 = (1'h0);
  reg [(4'h8):(1'h0)] reg4198 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4197 = (1'h0);
  reg [(4'he):(1'h0)] reg4196 = (1'h0);
  reg [(4'hb):(1'h0)] reg4195 = (1'h0);
  reg [(3'h5):(1'h0)] reg4194 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4193 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4192 = (1'h0);
  reg [(5'h10):(1'h0)] reg4191 = (1'h0);
  reg [(5'h10):(1'h0)] reg4190 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4189 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4188 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4187 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4186 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4185 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4184 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4183 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4182 = (1'h0);
  reg [(3'h7):(1'h0)] reg4181 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4180 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4179 = (1'h0);
  reg [(2'h2):(1'h0)] reg4178 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4177 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4176 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4175 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4174 = (1'h0);
  reg [(4'hd):(1'h0)] reg4173 = (1'h0);
  reg [(4'hb):(1'h0)] reg4172 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4171 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4170 = (1'h0);
  reg [(3'h5):(1'h0)] reg4169 = (1'h0);
  reg [(2'h2):(1'h0)] reg4168 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4167 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4165 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4161 = (1'h0);
  reg [(4'he):(1'h0)] reg4157 = (1'h0);
  reg [(2'h2):(1'h0)] reg4155 = (1'h0);
  reg [(4'h9):(1'h0)] reg4153 = (1'h0);
  reg [(4'hc):(1'h0)] reg4167 = (1'h0);
  reg [(5'h10):(1'h0)] reg4166 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4165 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4164 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4163 = (1'h0);
  reg [(3'h6):(1'h0)] reg4162 = (1'h0);
  reg [(4'h9):(1'h0)] reg4161 = (1'h0);
  reg [(4'hc):(1'h0)] reg4160 = (1'h0);
  reg [(4'he):(1'h0)] reg4159 = (1'h0);
  reg [(3'h7):(1'h0)] reg4158 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4157 = (1'h0);
  reg [(2'h2):(1'h0)] reg4156 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4155 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4154 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4153 = (1'h0);
  wire [(4'ha):(1'h0)] wire4152;
  wire [(4'h9):(1'h0)] wire4151;
  wire [(4'h8):(1'h0)] wire4150;
  wire signed [(5'h10):(1'h0)] wire4149;
  wire signed [(2'h2):(1'h0)] wire4148;
  wire signed [(4'ha):(1'h0)] wire4146;
  wire signed [(3'h4):(1'h0)] wire640;
  wire signed [(4'h8):(1'h0)] wire639;
  wire signed [(4'h9):(1'h0)] wire638;
  wire signed [(4'h8):(1'h0)] wire637;
  wire [(4'ha):(1'h0)] wire636;
  wire [(4'hf):(1'h0)] wire635;
  assign y = {wire4384,
                 wire4383,
                 reg4382,
                 reg4381,
                 reg4380,
                 forvar4379,
                 forvar4378,
                 forvar4377,
                 reg4376,
                 forvar4375,
                 reg4373,
                 reg4368,
                 forvar4365,
                 reg4375,
                 reg4374,
                 forvar4373,
                 reg4372,
                 reg4371,
                 reg4370,
                 reg4369,
                 forvar4368,
                 reg4367,
                 reg4366,
                 reg4365,
                 forvar4356,
                 reg4364,
                 reg4363,
                 reg4362,
                 reg4361,
                 reg4360,
                 reg4359,
                 reg4358,
                 reg4357,
                 reg4356,
                 reg4355,
                 reg4354,
                 forvar4353,
                 reg4352,
                 reg4351,
                 reg4350,
                 reg4349,
                 reg4348,
                 reg4347,
                 reg4346,
                 forvar4345,
                 reg4344,
                 reg4343,
                 reg4342,
                 reg4341,
                 forvar4340,
                 reg4339,
                 reg4338,
                 reg4337,
                 forvar4336,
                 reg4335,
                 reg4334,
                 reg4333,
                 forvar4331,
                 reg4332,
                 reg4331,
                 reg4330,
                 forvar4329,
                 reg4328,
                 reg4327,
                 reg4326,
                 reg4325,
                 forvar4324,
                 forvar4323,
                 forvar4322,
                 forvar4300,
                 forvar4306,
                 reg4321,
                 reg4320,
                 reg4319,
                 reg4318,
                 reg4317,
                 reg4316,
                 reg4315,
                 reg4314,
                 reg4313,
                 forvar4312,
                 reg4311,
                 reg4310,
                 reg4309,
                 forvar4308,
                 reg4307,
                 reg4306,
                 reg4305,
                 reg4304,
                 reg4303,
                 reg4302,
                 reg4301,
                 reg4300,
                 reg4299,
                 forvar4298,
                 reg4297,
                 reg4290,
                 reg4296,
                 reg4295,
                 reg4294,
                 reg4293,
                 reg4292,
                 reg4291,
                 forvar4290,
                 reg4289,
                 reg4288,
                 reg4287,
                 reg4286,
                 reg4285,
                 forvar4284,
                 reg4283,
                 reg4282,
                 reg4281,
                 reg4280,
                 reg4279,
                 forvar4278,
                 forvar4277,
                 forvar4276,
                 reg4275,
                 reg4274,
                 reg4273,
                 reg4272,
                 reg4271,
                 reg4270,
                 reg4269,
                 forvar4268,
                 reg4267,
                 reg4266,
                 forvar4265,
                 reg4264,
                 forvar4263,
                 forvar4247,
                 reg4262,
                 reg4261,
                 reg4260,
                 forvar4259,
                 reg4258,
                 reg4257,
                 reg4256,
                 reg4255,
                 forvar4254,
                 reg4253,
                 reg4252,
                 reg4251,
                 reg4250,
                 reg4249,
                 reg4248,
                 reg4247,
                 forvar4246,
                 forvar4245,
                 reg4244,
                 reg4243,
                 reg4242,
                 reg4241,
                 reg4240,
                 forvar4239,
                 reg4238,
                 reg4237,
                 reg4236,
                 forvar4235,
                 reg4234,
                 forvar4233,
                 reg4232,
                 reg4231,
                 reg4230,
                 forvar4229,
                 forvar4228,
                 forvar4227,
                 reg4226,
                 reg4225,
                 reg4224,
                 reg4223,
                 reg4222,
                 reg4221,
                 forvar4220,
                 reg4219,
                 reg4218,
                 reg4217,
                 forvar4216,
                 reg4215,
                 forvar4214,
                 forvar4213,
                 reg4212,
                 reg4211,
                 reg4210,
                 reg4209,
                 forvar4208,
                 reg4207,
                 reg4206,
                 reg4205,
                 forvar4204,
                 reg4203,
                 reg4202,
                 reg4201,
                 reg4200,
                 forvar4199,
                 reg4198,
                 forvar4197,
                 reg4196,
                 reg4195,
                 reg4194,
                 forvar4193,
                 forvar4192,
                 reg4191,
                 reg4190,
                 reg4189,
                 reg4188,
                 reg4187,
                 reg4186,
                 reg4185,
                 forvar4184,
                 reg4183,
                 reg4182,
                 reg4181,
                 reg4180,
                 forvar4179,
                 reg4178,
                 reg4177,
                 forvar4176,
                 forvar4175,
                 forvar4174,
                 reg4173,
                 reg4172,
                 reg4171,
                 reg4170,
                 reg4169,
                 reg4168,
                 forvar4167,
                 reg4165,
                 forvar4161,
                 reg4157,
                 reg4155,
                 reg4153,
                 reg4167,
                 reg4166,
                 forvar4165,
                 reg4164,
                 reg4163,
                 reg4162,
                 reg4161,
                 reg4160,
                 reg4159,
                 reg4158,
                 forvar4157,
                 reg4156,
                 forvar4155,
                 reg4154,
                 forvar4153,
                 wire4152,
                 wire4151,
                 wire4150,
                 wire4149,
                 wire4148,
                 wire4146,
                 wire640,
                 wire639,
                 wire638,
                 wire637,
                 wire636,
                 wire635,
                 (1'h0)};
  assign wire635 = (wire632 | $unsigned({$signed(wire631)}));
  assign wire636 = wire635[(2'h2):(1'h1)];
  assign wire637 = wire632[(3'h4):(3'h4)];
  assign wire638 = (((~|wire634[(3'h4):(1'h0)]) ?
                           ((wire631 ? wire636 : wire631) ?
                               (wire635 ?
                                   wire631 : (8'hae)) : wire632) : ($signed(wire634) ?
                               {wire633} : (wire632 * wire633))) ?
                       $signed(wire637) : (~&(&{wire635})));
  assign wire639 = ($signed($unsigned(wire631)) ^~ (+($unsigned(wire635) ?
                       ((8'hb8) ?
                           wire638 : wire633) : wire636[(3'h7):(3'h5)])));
  assign wire640 = (~^($signed((~&wire635)) >>> ((wire631 + wire632) ?
                       (wire631 ? wire634 : wire634) : {wire639})));
  module641 modinst4147 (wire4146, clk, wire638, wire637, wire635, wire639);
  assign wire4148 = $unsigned(wire638[(4'h8):(1'h1)]);
  assign wire4149 = (wire635[(4'hc):(3'h7)] ?
                        (~((~|wire634) ?
                            (wire639 <= wire637) : $signed(wire638))) : $signed(wire637));
  assign wire4150 = $signed((^wire634[(2'h2):(1'h1)]));
  assign wire4151 = wire634[(3'h4):(3'h4)];
  assign wire4152 = wire4148[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      if ((wire637 & wire4151))
        begin
          for (forvar4153 = (1'h0); (forvar4153 < (2'h3)); forvar4153 = (forvar4153 + (1'h1)))
            begin
              reg4154 <= $unsigned((((&(8'h9f)) < $unsigned(wire4151)) > (~|{wire635})));
            end
          for (forvar4155 = (1'h0); (forvar4155 < (2'h3)); forvar4155 = (forvar4155 + (1'h1)))
            begin
              reg4156 <= (wire635 ? {wire4150} : forvar4153);
              for (forvar4157 = (1'h0); (forvar4157 < (1'h0)); forvar4157 = (forvar4157 + (1'h1)))
                begin
                  reg4158 <= {$unsigned(reg4154[(2'h2):(1'h0)])};
                  if (($unsigned($signed(reg4158[(3'h7):(3'h4)])) ?
                      $signed(($unsigned((8'ha2)) >= (wire632 * wire4148))) : (wire4150[(2'h2):(1'h1)] <<< $unsigned($unsigned(reg4156)))))
                    begin
                      reg4159 <= $signed({wire631[(1'h1):(1'h1)]});
                      reg4160 <= ((8'ha8) ? wire4150 : {(^$unsigned((8'hae)))});
                      reg4161 <= {(((reg4154 ^~ forvar4155) ?
                              (wire633 ? wire639 : reg4160) : (wire4148 ?
                                  wire640 : wire639)) << ({reg4159} == wire4149[(3'h7):(1'h1)]))};
                    end
                  else
                    begin
                      reg4159 <= (reg4160 >> reg4154);
                      reg4160 <= ($unsigned(wire631[(1'h0):(1'h0)]) ?
                          {wire634} : $signed($unsigned((wire4152 ?
                              (8'ha2) : reg4156))));
                    end
                  if ({wire634[(3'h5):(2'h3)]})
                    begin
                      reg4162 <= forvar4157;
                      reg4163 <= ($signed(($unsigned(wire4150) ?
                          (8'ha0) : (wire4146 << wire638))) >>> $unsigned($unsigned(reg4156)));
                    end
                  else
                    begin
                      reg4162 <= (((-((8'ha3) ?
                              wire4152 : wire637)) > ((8'ha8) ?
                              wire638[(1'h0):(1'h0)] : {(8'ha9)})) ?
                          wire640[(2'h2):(1'h0)] : wire634[(2'h2):(2'h2)]);
                      reg4163 <= wire4150;
                      reg4164 <= wire4152[(4'h8):(3'h6)];
                    end
                  for (forvar4165 = (1'h0); (forvar4165 < (2'h3)); forvar4165 = (forvar4165 + (1'h1)))
                    begin
                      reg4166 <= reg4159[(4'hb):(3'h5)];
                    end
                end
            end
          reg4167 <= (~|(-({forvar4155} ^~ wire4148)));
        end
      else
        begin
          if (wire4152)
            begin
              if ((wire633 ^ $unsigned(wire635)))
                begin
                  if (({($signed(forvar4157) + (wire4149 >>> (8'ha4)))} ?
                      $unsigned(wire631[(3'h5):(3'h5)]) : ((wire631[(3'h5):(2'h3)] ?
                          wire636 : (wire631 * wire4146)) >>> ($unsigned(reg4156) ?
                          forvar4157 : ((8'hb1) ? forvar4157 : wire637)))))
                    begin
                      reg4153 <= $unsigned($unsigned($signed($unsigned(forvar4157))));
                    end
                  else
                    begin
                      reg4153 <= (((~^reg4154) > (((8'ha3) ?
                                  wire637 : wire638) ?
                              wire631 : {wire637})) ?
                          (8'had) : $signed(($signed(wire4149) ?
                              (+reg4154) : (reg4159 ? (8'hb5) : (8'haa)))));
                      reg4154 <= reg4162;
                      reg4155 <= reg4159;
                      reg4156 <= $unsigned(($unsigned($unsigned((8'ha6))) << (^~(reg4164 ?
                          wire638 : reg4166))));
                    end
                  if ($unsigned(wire632[(2'h2):(1'h0)]))
                    begin
                      reg4157 <= (reg4160[(2'h2):(1'h1)] - $unsigned((~^forvar4157)));
                    end
                  else
                    begin
                      reg4157 <= (reg4161 << wire634);
                      reg4158 <= $unsigned((|{{(8'hb6)}}));
                      reg4159 <= wire4148[(2'h2):(1'h0)];
                      reg4160 <= $unsigned(($signed((forvar4157 ?
                          wire4151 : reg4159)) && (reg4164 & wire633[(4'he):(3'h4)])));
                    end
                  for (forvar4161 = (1'h0); (forvar4161 < (2'h2)); forvar4161 = (forvar4161 + (1'h1)))
                    begin
                      reg4162 <= (({wire4148[(1'h0):(1'h0)]} && ($signed(forvar4155) ?
                          $unsigned(wire638) : (~&wire640))) == (~^$signed(reg4160)));
                      reg4163 <= $unsigned($signed(wire635[(1'h0):(1'h0)]));
                      reg4164 <= wire633;
                      reg4165 <= ({$signed($signed(reg4166))} ?
                          $signed(wire639[(3'h6):(2'h2)]) : reg4166[(3'h7):(3'h5)]);
                    end
                end
              else
                begin
                  for (forvar4153 = (1'h0); (forvar4153 < (2'h2)); forvar4153 = (forvar4153 + (1'h1)))
                    begin
                      reg4154 <= reg4164;
                      reg4155 <= wire639[(3'h6):(1'h1)];
                    end
                end
              reg4166 <= {($signed((+(8'h9f))) >= forvar4161[(1'h1):(1'h1)])};
              if ($signed(wire631))
                begin
                  for (forvar4167 = (1'h0); (forvar4167 < (1'h1)); forvar4167 = (forvar4167 + (1'h1)))
                    begin
                      reg4168 <= (8'ha1);
                      reg4169 <= ((8'hac) ? reg4160 : wire4146[(2'h3):(2'h2)]);
                      reg4170 <= (reg4164[(2'h2):(1'h1)] ^ wire634);
                    end
                end
              else
                begin
                  reg4167 <= ($unsigned(forvar4155[(3'h4):(2'h3)]) ?
                      $unsigned($unsigned($signed(reg4170))) : $signed(reg4159[(3'h4):(1'h1)]));
                  reg4168 <= $unsigned(reg4157);
                  if ((reg4155[(2'h2):(1'h0)] + ((~(wire4148 ?
                          reg4169 : forvar4153)) ?
                      $unsigned($signed(reg4165)) : ((wire636 ?
                              wire4146 : reg4156) ?
                          (reg4168 >> wire632) : forvar4155[(3'h7):(2'h2)]))))
                    begin
                      reg4169 <= {$signed($signed(forvar4153))};
                    end
                  else
                    begin
                      reg4169 <= $signed($unsigned($unsigned($signed(reg4169))));
                      reg4170 <= {$unsigned(($signed(reg4157) | {wire4146}))};
                      reg4171 <= wire4146;
                    end
                end
              reg4172 <= (^(wire4148[(1'h0):(1'h0)] ?
                  ($signed(wire632) << wire632[(2'h2):(1'h1)]) : $unsigned((8'hb6))));
            end
          else
            begin
              reg4153 <= (({forvar4167} ?
                      (((8'ha3) ^~ wire639) > (reg4153 ?
                          reg4169 : (8'had))) : {(forvar4153 ~^ wire634)}) ?
                  ($unsigned((-forvar4157)) ?
                      (-{wire639}) : {wire4149[(3'h6):(3'h4)]}) : (|((&(8'hb3)) ^ wire639)));
            end
          reg4173 <= $signed($unsigned(((8'ha7) ^~ {(8'ha4)})));
          for (forvar4174 = (1'h0); (forvar4174 < (1'h0)); forvar4174 = (forvar4174 + (1'h1)))
            begin
              for (forvar4175 = (1'h0); (forvar4175 < (1'h0)); forvar4175 = (forvar4175 + (1'h1)))
                begin
                  for (forvar4176 = (1'h0); (forvar4176 < (1'h0)); forvar4176 = (forvar4176 + (1'h1)))
                    begin
                      reg4177 <= (!forvar4155);
                      reg4178 <= reg4172;
                    end
                  for (forvar4179 = (1'h0); (forvar4179 < (2'h3)); forvar4179 = (forvar4179 + (1'h1)))
                    begin
                      reg4180 <= reg4171[(1'h0):(1'h0)];
                      reg4181 <= ((8'hb2) < reg4160);
                      reg4182 <= reg4157[(4'hc):(1'h1)];
                      reg4183 <= $unsigned((8'hba));
                    end
                  for (forvar4184 = (1'h0); (forvar4184 < (1'h1)); forvar4184 = (forvar4184 + (1'h1)))
                    begin
                      reg4185 <= forvar4161[(2'h2):(2'h2)];
                      reg4186 <= reg4168[(2'h2):(1'h0)];
                      reg4187 <= (^$unsigned($signed(reg4164[(1'h1):(1'h0)])));
                    end
                  if ($unsigned(wire632[(2'h3):(2'h3)]))
                    begin
                      reg4188 <= wire4150[(3'h7):(3'h5)];
                      reg4189 <= ($signed((|$unsigned(forvar4184))) << (wire4146 ~^ $signed(reg4181)));
                      reg4190 <= $signed((8'hba));
                      reg4191 <= {(|forvar4167)};
                    end
                  else
                    begin
                      reg4188 <= $unsigned((((reg4189 ? (8'hb6) : wire639) ?
                              (reg4168 ? forvar4161 : wire4148) : wire640) ?
                          reg4173[(3'h5):(2'h2)] : reg4163[(1'h1):(1'h1)]));
                    end
                end
              for (forvar4192 = (1'h0); (forvar4192 < (1'h0)); forvar4192 = (forvar4192 + (1'h1)))
                begin
                  for (forvar4193 = (1'h0); (forvar4193 < (1'h0)); forvar4193 = (forvar4193 + (1'h1)))
                    begin
                      reg4194 <= $unsigned(((+(|(8'hb8))) ^ ((~^reg4186) ?
                          $signed(reg4172) : (wire4150 >= wire631))));
                      reg4195 <= wire4152;
                      reg4196 <= (8'hb9);
                    end
                end
              for (forvar4197 = (1'h0); (forvar4197 < (2'h2)); forvar4197 = (forvar4197 + (1'h1)))
                begin
                  reg4198 <= ((+((+reg4191) ?
                      {wire4149} : $signed(wire640))) >>> ($signed((&forvar4175)) ?
                      ((!(8'ha0)) && $signed((8'ha8))) : {$signed(reg4161)}));
                  for (forvar4199 = (1'h0); (forvar4199 < (1'h0)); forvar4199 = (forvar4199 + (1'h1)))
                    begin
                      reg4200 <= (+reg4154[(1'h0):(1'h0)]);
                      reg4201 <= $signed(reg4194);
                      reg4202 <= {$signed((8'ha6))};
                      reg4203 <= $signed($unsigned($signed((forvar4197 - reg4202))));
                    end
                  for (forvar4204 = (1'h0); (forvar4204 < (2'h3)); forvar4204 = (forvar4204 + (1'h1)))
                    begin
                      reg4205 <= {reg4172};
                      reg4206 <= reg4177;
                      reg4207 <= $unsigned((!$unsigned((8'hb9))));
                    end
                  for (forvar4208 = (1'h0); (forvar4208 < (2'h3)); forvar4208 = (forvar4208 + (1'h1)))
                    begin
                      reg4209 <= reg4160[(1'h0):(1'h0)];
                      reg4210 <= $unsigned({$unsigned((^~wire632))});
                      reg4211 <= ((((reg4195 <= reg4162) ?
                          $unsigned(reg4160) : (wire4146 & forvar4179)) ^~ reg4186) <<< forvar4199);
                      reg4212 <= forvar4204;
                    end
                end
              for (forvar4213 = (1'h0); (forvar4213 < (1'h1)); forvar4213 = (forvar4213 + (1'h1)))
                begin
                  for (forvar4214 = (1'h0); (forvar4214 < (2'h2)); forvar4214 = (forvar4214 + (1'h1)))
                    begin
                      reg4215 <= {wire632};
                    end
                  for (forvar4216 = (1'h0); (forvar4216 < (2'h3)); forvar4216 = (forvar4216 + (1'h1)))
                    begin
                      reg4217 <= forvar4184[(4'h8):(3'h6)];
                      reg4218 <= (8'h9c);
                      reg4219 <= (((~&(forvar4216 | wire4150)) ?
                              reg4194 : $signed(wire4148)) ?
                          ($unsigned(reg4206) >= reg4155) : (((reg4189 ?
                                  forvar4174 : reg4170) ?
                              (reg4189 ^ forvar4153) : (wire4151 & reg4202)) <= (8'hba)));
                    end
                  for (forvar4220 = (1'h0); (forvar4220 < (2'h2)); forvar4220 = (forvar4220 + (1'h1)))
                    begin
                      reg4221 <= (+(8'hae));
                      reg4222 <= (^~reg4183);
                      reg4223 <= wire631;
                      reg4224 <= (($unsigned((reg4190 ? reg4191 : reg4205)) ?
                          (^wire4150[(2'h3):(1'h0)]) : ($signed((8'ha2)) ?
                              {forvar4153} : ((8'h9e) ?
                                  (8'hb3) : forvar4216))) == (^($signed(reg4170) >>> {reg4156})));
                    end
                  reg4225 <= (-(wire631[(1'h0):(1'h0)] ?
                      $unsigned((reg4221 ? wire632 : wire4149)) : (wire635 ?
                          (!forvar4216) : ((8'haa) * reg4188))));
                end
            end
          reg4226 <= ((-((^~reg4212) != $signed(reg4186))) ?
              (($unsigned(reg4177) ?
                  $signed(forvar4192) : reg4172) ^~ $signed((reg4161 ?
                  forvar4197 : forvar4204))) : (|($unsigned(reg4162) ~^ reg4202)));
        end
      for (forvar4227 = (1'h0); (forvar4227 < (1'h0)); forvar4227 = (forvar4227 + (1'h1)))
        begin
          for (forvar4228 = (1'h0); (forvar4228 < (1'h1)); forvar4228 = (forvar4228 + (1'h1)))
            begin
              if (reg4158)
                begin
                  for (forvar4229 = (1'h0); (forvar4229 < (2'h2)); forvar4229 = (forvar4229 + (1'h1)))
                    begin
                      reg4230 <= $signed($unsigned($unsigned((forvar4228 ?
                          (8'hb3) : wire634))));
                      reg4231 <= reg4163;
                      reg4232 <= {$unsigned(reg4188)};
                    end
                end
              else
                begin
                  for (forvar4229 = (1'h0); (forvar4229 < (1'h0)); forvar4229 = (forvar4229 + (1'h1)))
                    begin
                      reg4230 <= (~|($signed(wire4151[(1'h0):(1'h0)]) ?
                          (8'hac) : $unsigned(reg4157)));
                      reg4231 <= ((forvar4213 ?
                              ($unsigned(forvar4155) ?
                                  $unsigned(wire4151) : (&reg4158)) : (^{forvar4176})) ?
                          (forvar4229[(4'hd):(4'hb)] ^ (^~(reg4207 ?
                              forvar4204 : reg4156))) : reg4230[(2'h2):(2'h2)]);
                    end
                end
              for (forvar4233 = (1'h0); (forvar4233 < (2'h2)); forvar4233 = (forvar4233 + (1'h1)))
                begin
                  reg4234 <= (reg4177[(3'h5):(2'h2)] ?
                      {({reg4156} + reg4164[(1'h0):(1'h0)])} : $signed(((~&wire633) >> (reg4230 < reg4153))));
                end
              for (forvar4235 = (1'h0); (forvar4235 < (2'h3)); forvar4235 = (forvar4235 + (1'h1)))
                begin
                  if ($signed($unsigned(((reg4188 ^~ forvar4227) ?
                      $signed(reg4201) : (&reg4159)))))
                    begin
                      reg4236 <= wire636[(4'ha):(3'h5)];
                      reg4237 <= $unsigned($signed($unsigned((forvar4184 && wire640))));
                      reg4238 <= (((forvar4214 ?
                              reg4191 : (|(8'h9e))) - $unsigned((forvar4208 ?
                              reg4219 : reg4218))) ?
                          {(8'ha2)} : $unsigned({(!reg4232)}));
                    end
                  else
                    begin
                      reg4236 <= $signed($signed(((reg4234 ?
                          wire4148 : wire640) << (wire4146 ?
                          reg4154 : forvar4208))));
                      reg4237 <= $signed(((reg4207 & reg4230) ?
                          reg4172[(3'h6):(1'h0)] : $unsigned((wire637 ?
                              (8'hac) : forvar4204))));
                    end
                  for (forvar4239 = (1'h0); (forvar4239 < (1'h1)); forvar4239 = (forvar4239 + (1'h1)))
                    begin
                      reg4240 <= (reg4191[(5'h10):(4'he)] ?
                          reg4210[(2'h3):(1'h0)] : ($signed($signed((8'hb9))) + (~|(~(8'hb1)))));
                      reg4241 <= $signed((-$signed(wire4149[(4'he):(3'h6)])));
                      reg4242 <= ($signed($signed((~wire634))) ?
                          reg4226[(4'hc):(4'ha)] : reg4167[(1'h1):(1'h1)]);
                      reg4243 <= $signed(forvar4197[(2'h2):(1'h0)]);
                    end
                end
              reg4244 <= {forvar4167[(3'h6):(3'h5)]};
            end
        end
      for (forvar4245 = (1'h0); (forvar4245 < (1'h1)); forvar4245 = (forvar4245 + (1'h1)))
        begin
          for (forvar4246 = (1'h0); (forvar4246 < (2'h3)); forvar4246 = (forvar4246 + (1'h1)))
            begin
              if (reg4170)
                begin
                  if ({$signed(($unsigned(reg4238) ?
                          wire636[(3'h7):(3'h5)] : reg4170))})
                    begin
                      reg4247 <= {{$unsigned($signed((8'h9c)))}};
                      reg4248 <= {$unsigned($signed((^~reg4165)))};
                    end
                  else
                    begin
                      reg4247 <= (((^reg4222[(1'h0):(1'h0)]) | {$signed(wire4149)}) ?
                          (reg4218 ?
                              reg4181[(2'h2):(2'h2)] : $signed($signed(reg4203))) : ((reg4221 < $unsigned(reg4224)) + {(|(8'hb9))}));
                      reg4248 <= ($unsigned(reg4205) || ($unsigned((reg4191 ?
                          reg4155 : wire638)) == $unsigned($signed((8'ha4)))));
                      reg4249 <= $signed($signed(reg4153[(3'h7):(2'h3)]));
                    end
                  if (($unsigned($unsigned($unsigned(reg4169))) ?
                      (~^reg4249) : $unsigned((!wire4151))))
                    begin
                      reg4250 <= ((8'ha8) > $unsigned(((forvar4246 || (8'ha6)) != (wire4152 - wire636))));
                      reg4251 <= ($unsigned((reg4238 | (reg4250 ?
                          reg4190 : forvar4175))) <<< (^~{((8'hb1) ?
                              reg4181 : (8'hb7))}));
                      reg4252 <= wire4151;
                    end
                  else
                    begin
                      reg4250 <= forvar4165;
                      reg4251 <= (reg4172 << reg4247[(2'h2):(1'h1)]);
                      reg4252 <= forvar4179;
                      reg4253 <= $signed(reg4212);
                    end
                  for (forvar4254 = (1'h0); (forvar4254 < (2'h2)); forvar4254 = (forvar4254 + (1'h1)))
                    begin
                      reg4255 <= (~^$unsigned((|forvar4167[(1'h0):(1'h0)])));
                      reg4256 <= (reg4207[(1'h0):(1'h0)] ?
                          (+(+$unsigned(reg4249))) : (forvar4228[(3'h4):(1'h1)] ?
                              $signed(reg4212) : {(&(8'haa))}));
                      reg4257 <= reg4166;
                      reg4258 <= reg4219;
                    end
                  for (forvar4259 = (1'h0); (forvar4259 < (1'h1)); forvar4259 = (forvar4259 + (1'h1)))
                    begin
                      reg4260 <= (-({(8'ha5)} ?
                          {reg4183} : wire636[(3'h7):(2'h2)]));
                      reg4261 <= $unsigned((8'hae));
                      reg4262 <= $signed((!(8'hac)));
                    end
                end
              else
                begin
                  for (forvar4247 = (1'h0); (forvar4247 < (1'h1)); forvar4247 = (forvar4247 + (1'h1)))
                    begin
                      reg4248 <= forvar4235;
                      reg4249 <= (8'had);
                      reg4250 <= $signed(wire640);
                      reg4251 <= reg4217[(1'h1):(1'h0)];
                    end
                end
            end
          for (forvar4263 = (1'h0); (forvar4263 < (1'h1)); forvar4263 = (forvar4263 + (1'h1)))
            begin
              reg4264 <= reg4180[(1'h0):(1'h0)];
              for (forvar4265 = (1'h0); (forvar4265 < (1'h0)); forvar4265 = (forvar4265 + (1'h1)))
                begin
                  reg4266 <= reg4183;
                end
              reg4267 <= forvar4214;
              for (forvar4268 = (1'h0); (forvar4268 < (2'h3)); forvar4268 = (forvar4268 + (1'h1)))
                begin
                  reg4269 <= ((forvar4192 ?
                      (|((8'ha3) + reg4264)) : (^~reg4161[(3'h4):(2'h3)])) > forvar4254[(1'h1):(1'h0)]);
                  if ((reg4247 ^~ (+$unsigned($unsigned(reg4262)))))
                    begin
                      reg4270 <= (forvar4161 ?
                          (-((reg4167 ? reg4210 : wire638) ?
                              {reg4219} : (forvar4157 && reg4261))) : reg4264);
                      reg4271 <= reg4219[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg4270 <= forvar4245[(2'h3):(1'h1)];
                      reg4271 <= (~^$signed(($unsigned(reg4201) >>> (reg4182 ?
                          forvar4233 : reg4253))));
                      reg4272 <= ($signed((&(+wire634))) == (!((^~wire632) ?
                          $unsigned(reg4164) : $signed(reg4237))));
                    end
                  if (((reg4219 ?
                      (!$signed(reg4225)) : forvar4227[(4'hc):(2'h3)]) >>> (-(^~reg4169[(1'h1):(1'h0)]))))
                    begin
                      reg4273 <= reg4262[(2'h3):(1'h0)];
                      reg4274 <= {$signed(forvar4220)};
                    end
                  else
                    begin
                      reg4273 <= $unsigned(((reg4154[(1'h1):(1'h0)] != {reg4269}) ?
                          ((^reg4231) ?
                              $unsigned((8'hb0)) : forvar4246) : ((reg4154 ?
                                  reg4187 : reg4177) ?
                              (^(8'hb4)) : (wire637 ? reg4172 : (8'ha2)))));
                      reg4274 <= ((forvar4246 || (~&reg4168)) ~^ (~|$signed($unsigned(reg4224))));
                    end
                  reg4275 <= forvar4246[(1'h0):(1'h0)];
                end
            end
          for (forvar4276 = (1'h0); (forvar4276 < (1'h1)); forvar4276 = (forvar4276 + (1'h1)))
            begin
              for (forvar4277 = (1'h0); (forvar4277 < (1'h0)); forvar4277 = (forvar4277 + (1'h1)))
                begin
                  for (forvar4278 = (1'h0); (forvar4278 < (2'h3)); forvar4278 = (forvar4278 + (1'h1)))
                    begin
                      reg4279 <= forvar4175[(4'h8):(1'h1)];
                      reg4280 <= (+reg4230);
                    end
                  if (({$signed((reg4275 ? reg4275 : reg4232))} <<< forvar4259))
                    begin
                      reg4281 <= (reg4244 - $signed($signed(reg4243[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg4281 <= reg4166[(1'h1):(1'h0)];
                      reg4282 <= (~&reg4178);
                    end
                  reg4283 <= reg4162[(1'h1):(1'h1)];
                  for (forvar4284 = (1'h0); (forvar4284 < (1'h1)); forvar4284 = (forvar4284 + (1'h1)))
                    begin
                      reg4285 <= $signed((!$signed(forvar4193[(4'h8):(2'h3)])));
                      reg4286 <= $signed($unsigned({reg4177[(4'h8):(4'h8)]}));
                      reg4287 <= ($signed((8'haf)) >>> (reg4269 ?
                          wire635[(3'h7):(3'h5)] : forvar4278));
                      reg4288 <= (!$signed((reg4209 ?
                          (reg4187 << reg4244) : reg4252)));
                    end
                end
              reg4289 <= reg4218[(3'h5):(3'h5)];
              if (reg4161[(1'h1):(1'h0)])
                begin
                  for (forvar4290 = (1'h0); (forvar4290 < (1'h0)); forvar4290 = (forvar4290 + (1'h1)))
                    begin
                      reg4291 <= wire4150[(4'h8):(4'h8)];
                    end
                  reg4292 <= ((($signed(reg4234) ? reg4260 : {reg4177}) ?
                          ((forvar4247 ?
                              reg4282 : reg4215) > {(8'h9f)}) : $unsigned((&reg4241))) ?
                      reg4171 : (+(forvar4214 ? reg4159 : $signed((8'ha6)))));
                  if ($signed(reg4289[(1'h1):(1'h1)]))
                    begin
                      reg4293 <= (reg4198 > reg4248);
                      reg4294 <= (reg4250[(4'hb):(3'h6)] <= ($signed($unsigned(reg4252)) ?
                          ((~&reg4178) <<< (~&reg4191)) : $unsigned(reg4219[(3'h7):(2'h3)])));
                      reg4295 <= $unsigned(reg4158[(3'h6):(2'h2)]);
                      reg4296 <= (&reg4215);
                    end
                  else
                    begin
                      reg4293 <= $unsigned(({reg4251} && {(+forvar4247)}));
                      reg4294 <= ($unsigned((8'ha7)) | (reg4240 | reg4286));
                      reg4295 <= $unsigned(reg4257[(4'h9):(1'h0)]);
                      reg4296 <= ($signed((&forvar4247)) || ((wire4151[(3'h7):(1'h0)] ?
                          (^~forvar4214) : $unsigned((8'ha0))) <= $signed($signed(forvar4184))));
                    end
                end
              else
                begin
                  reg4290 <= (-forvar4247);
                  if ((+(~^reg4159[(3'h6):(2'h2)])))
                    begin
                      reg4291 <= forvar4153;
                      reg4292 <= forvar4254;
                      reg4293 <= (({{(8'hb8)}} >>> forvar4277) ?
                          (|$unsigned(forvar4235[(1'h0):(1'h0)])) : reg4255);
                    end
                  else
                    begin
                      reg4291 <= reg4156;
                      reg4292 <= forvar4278;
                    end
                end
              reg4297 <= reg4287[(1'h1):(1'h0)];
            end
        end
      for (forvar4298 = (1'h0); (forvar4298 < (2'h3)); forvar4298 = (forvar4298 + (1'h1)))
        begin
          if (reg4274[(1'h1):(1'h0)])
            begin
              reg4299 <= reg4279;
              if (reg4279[(1'h0):(1'h0)])
                begin
                  if ($signed(reg4271))
                    begin
                      reg4300 <= $unsigned(($unsigned(reg4171[(2'h3):(1'h0)]) ?
                          ({reg4171} || reg4281) : (|reg4258)));
                      reg4301 <= $signed($unsigned(($unsigned((8'ha8)) ?
                          (reg4210 && (8'hb2)) : (wire4149 ?
                              forvar4174 : forvar4184))));
                      reg4302 <= ($signed(((-wire4148) != {forvar4284})) == {($unsigned(reg4244) ?
                              (reg4224 ?
                                  wire636 : wire640) : $signed(reg4182))});
                    end
                  else
                    begin
                      reg4300 <= (-$unsigned($unsigned({(8'hb6)})));
                      reg4301 <= ($signed((!$unsigned(reg4302))) | (reg4173[(3'h4):(2'h3)] <<< ({reg4211} ?
                          reg4224 : forvar4204)));
                    end
                end
              else
                begin
                  if ({(reg4262 ?
                          (~(forvar4179 ?
                              forvar4155 : forvar4254)) : $unsigned(reg4266[(4'h8):(3'h6)]))})
                    begin
                      reg4300 <= (forvar4213 <= (!$unsigned((&(8'ha0)))));
                      reg4301 <= $signed((~&($unsigned(forvar4213) ^ (^~reg4258))));
                      reg4302 <= (($signed(forvar4284) ?
                              (^(~&reg4157)) : (8'hb1)) ?
                          ($unsigned((reg4285 ? wire638 : (8'haf))) ?
                              (|(reg4264 ?
                                  wire4151 : reg4299)) : reg4222[(4'h8):(2'h3)]) : $unsigned($unsigned($signed(reg4158))));
                      reg4303 <= (&((8'hb5) <<< (~&(^(8'ha0)))));
                    end
                  else
                    begin
                      reg4300 <= $unsigned(forvar4265);
                      reg4301 <= (+{wire4150});
                    end
                  if ({(reg4288 & reg4194[(3'h4):(1'h0)])})
                    begin
                      reg4304 <= (~(~^$unsigned($signed(reg4299))));
                      reg4305 <= ((($unsigned((8'ha6)) * (wire4150 ?
                              reg4172 : reg4165)) && forvar4298[(2'h3):(1'h0)]) ?
                          ((|(forvar4208 ? reg4262 : reg4211)) ?
                              reg4244[(2'h2):(2'h2)] : (~^forvar4176[(2'h2):(1'h1)])) : (8'ha1));
                    end
                  else
                    begin
                      reg4304 <= ({((reg4231 ?
                              reg4251 : reg4256) * forvar4290[(1'h0):(1'h0)])} - (($unsigned(forvar4197) ?
                              (^reg4247) : (reg4264 ? reg4221 : reg4269)) ?
                          $unsigned(forvar4197) : $signed((~forvar4239))));
                      reg4305 <= ({($signed((8'h9e)) ?
                                  reg4240[(3'h4):(1'h1)] : {forvar4276})} ?
                          (+reg4238[(2'h2):(1'h0)]) : $unsigned((reg4181 ?
                              reg4282[(2'h2):(1'h0)] : forvar4214)));
                      reg4306 <= (-$unsigned({$signed(reg4223)}));
                      reg4307 <= $unsigned((&$signed($unsigned(forvar4228))));
                    end
                  for (forvar4308 = (1'h0); (forvar4308 < (1'h0)); forvar4308 = (forvar4308 + (1'h1)))
                    begin
                      reg4309 <= $unsigned($unsigned(((reg4292 ?
                              (8'haf) : forvar4155) ?
                          {reg4266} : {forvar4308})));
                      reg4310 <= reg4238;
                      reg4311 <= reg4297[(1'h1):(1'h0)];
                    end
                  for (forvar4312 = (1'h0); (forvar4312 < (1'h0)); forvar4312 = (forvar4312 + (1'h1)))
                    begin
                      reg4313 <= reg4291;
                      reg4314 <= reg4244[(2'h2):(2'h2)];
                      reg4315 <= reg4200[(3'h4):(3'h4)];
                    end
                end
              if (reg4181)
                begin
                  reg4316 <= reg4182[(3'h6):(3'h4)];
                end
              else
                begin
                  if (forvar4167)
                    begin
                      reg4316 <= $signed($unsigned(((reg4188 ?
                          reg4205 : reg4159) == $signed((8'hb1)))));
                    end
                  else
                    begin
                      reg4316 <= {reg4316};
                      reg4317 <= {forvar4228};
                      reg4318 <= $unsigned((($unsigned((8'hb5)) == reg4164) ?
                          (~|{forvar4290}) : wire640[(2'h2):(1'h0)]));
                    end
                  if (forvar4220)
                    begin
                      reg4319 <= ((+(|(reg4290 | reg4170))) ?
                          $unsigned((^(forvar4167 ?
                              reg4236 : reg4264))) : reg4162);
                      reg4320 <= $unsigned(forvar4246[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg4319 <= $unsigned(forvar4229[(2'h3):(2'h3)]);
                    end
                  reg4321 <= ((~(forvar4263 >>> (wire638 ^ forvar4184))) ?
                      reg4313[(4'ha):(4'h8)] : reg4217);
                end
            end
          else
            begin
              if (($unsigned((forvar4284[(4'hd):(2'h3)] ^~ ((8'hba) ?
                  (8'h9c) : (8'h9d)))) > (~&reg4269[(2'h2):(1'h0)])))
                begin
                  if (reg4256)
                    begin
                      reg4299 <= ($signed(forvar4246) ?
                          {((reg4190 - reg4293) ?
                                  (reg4223 ?
                                      reg4188 : forvar4165) : (forvar4155 ?
                                      reg4311 : reg4283))} : (~({wire4151} ~^ $signed(forvar4161))));
                      reg4300 <= $unsigned($signed(($unsigned(reg4296) ^ wire631)));
                      reg4301 <= (&reg4164[(3'h7):(3'h6)]);
                    end
                  else
                    begin
                      reg4299 <= (&forvar4213);
                      reg4300 <= (~&$signed(((forvar4153 >= wire4148) <= (+(8'hb6)))));
                      reg4301 <= $unsigned($unsigned(((reg4161 ?
                              reg4258 : reg4159) ?
                          $unsigned(reg4301) : (8'h9f))));
                    end
                  if ($unsigned(forvar4199))
                    begin
                      reg4302 <= $signed($signed(((~&reg4243) ?
                          $signed((8'ha0)) : (8'ha3))));
                    end
                  else
                    begin
                      reg4302 <= reg4296[(3'h5):(1'h0)];
                      reg4303 <= $unsigned($signed((~^$signed(reg4169))));
                      reg4304 <= reg4305;
                      reg4305 <= (8'hae);
                    end
                  for (forvar4306 = (1'h0); (forvar4306 < (1'h1)); forvar4306 = (forvar4306 + (1'h1)))
                    begin
                      reg4307 <= (8'ha9);
                    end
                end
              else
                begin
                  reg4299 <= ((~&reg4185[(1'h0):(1'h0)]) ?
                      (forvar4245[(4'h8):(3'h4)] & $signed(reg4292[(1'h1):(1'h0)])) : reg4232);
                  for (forvar4300 = (1'h0); (forvar4300 < (1'h1)); forvar4300 = (forvar4300 + (1'h1)))
                    begin
                      reg4301 <= {$unsigned(($unsigned(reg4318) ?
                              (reg4171 ?
                                  reg4261 : reg4195) : reg4222[(4'hb):(1'h0)]))};
                    end
                end
            end
          for (forvar4322 = (1'h0); (forvar4322 < (1'h1)); forvar4322 = (forvar4322 + (1'h1)))
            begin
              for (forvar4323 = (1'h0); (forvar4323 < (2'h3)); forvar4323 = (forvar4323 + (1'h1)))
                begin
                  for (forvar4324 = (1'h0); (forvar4324 < (1'h0)); forvar4324 = (forvar4324 + (1'h1)))
                    begin
                      reg4325 <= forvar4214[(3'h7):(2'h3)];
                      reg4326 <= reg4160;
                    end
                end
              reg4327 <= ($signed(reg4238) <= $unsigned(reg4300[(4'hb):(4'hb)]));
              reg4328 <= (reg4286[(4'h8):(3'h4)] <<< forvar4259);
            end
          if (reg4261[(3'h7):(3'h5)])
            begin
              for (forvar4329 = (1'h0); (forvar4329 < (1'h0)); forvar4329 = (forvar4329 + (1'h1)))
                begin
                  if (((&((wire4150 ? reg4251 : reg4215) << $signed(wire631))) ?
                      (~|reg4258[(2'h2):(2'h2)]) : (reg4285[(2'h2):(2'h2)] ?
                          $signed(reg4252) : forvar4306)))
                    begin
                      reg4330 <= (~$signed($unsigned($unsigned(reg4158))));
                      reg4331 <= ($unsigned({((8'ha7) >= (8'h9d))}) ^~ ($unsigned($unsigned(reg4212)) ~^ reg4159[(3'h6):(3'h5)]));
                      reg4332 <= $signed((({reg4301} ?
                              $unsigned(forvar4268) : (forvar4214 >= reg4273)) ?
                          {forvar4157[(1'h1):(1'h0)]} : $signed((reg4196 ?
                              (8'hba) : reg4326))));
                    end
                  else
                    begin
                      reg4330 <= $signed(reg4302[(3'h6):(3'h4)]);
                      reg4331 <= {(~^$unsigned($signed(reg4330)))};
                      reg4332 <= reg4230[(1'h0):(1'h0)];
                    end
                end
            end
          else
            begin
              if ((reg4200[(1'h1):(1'h0)] << $signed(($signed(reg4321) ?
                  reg4171[(4'h9):(2'h3)] : (8'hb8)))))
                begin
                  for (forvar4329 = (1'h0); (forvar4329 < (2'h3)); forvar4329 = (forvar4329 + (1'h1)))
                    begin
                      reg4330 <= $unsigned(forvar4298[(4'ha):(1'h0)]);
                    end
                  for (forvar4331 = (1'h0); (forvar4331 < (2'h2)); forvar4331 = (forvar4331 + (1'h1)))
                    begin
                      reg4332 <= wire635;
                      reg4333 <= (8'ha8);
                      reg4334 <= (~&reg4163);
                      reg4335 <= reg4221;
                    end
                  for (forvar4336 = (1'h0); (forvar4336 < (2'h3)); forvar4336 = (forvar4336 + (1'h1)))
                    begin
                      reg4337 <= forvar4308[(4'hd):(1'h1)];
                      reg4338 <= reg4337[(4'hf):(4'hf)];
                    end
                  reg4339 <= $unsigned((^~$signed($unsigned(forvar4278))));
                end
              else
                begin
                  for (forvar4329 = (1'h0); (forvar4329 < (2'h3)); forvar4329 = (forvar4329 + (1'h1)))
                    begin
                      reg4330 <= reg4234;
                      reg4331 <= {(~&reg4189[(3'h5):(1'h0)])};
                      reg4332 <= (|(|reg4232[(3'h4):(2'h2)]));
                      reg4333 <= (~$signed((forvar4235[(1'h0):(1'h0)] || reg4186[(4'hb):(2'h3)])));
                    end
                  reg4334 <= reg4231[(1'h0):(1'h0)];
                end
              for (forvar4340 = (1'h0); (forvar4340 < (2'h3)); forvar4340 = (forvar4340 + (1'h1)))
                begin
                  if ($signed((^reg4225[(1'h0):(1'h0)])))
                    begin
                      reg4341 <= forvar4239;
                      reg4342 <= ((+(|$signed(forvar4197))) ?
                          (((~|reg4306) ?
                              (~^wire637) : (&reg4273)) << $unsigned(reg4301)) : (8'h9e));
                      reg4343 <= $signed(reg4207);
                    end
                  else
                    begin
                      reg4341 <= (~($signed((reg4241 || forvar4174)) ?
                          {{reg4251}} : reg4291));
                      reg4342 <= $signed((&{(~|reg4262)}));
                      reg4343 <= $unsigned((reg4293 | ($unsigned((8'h9f)) ?
                          forvar4245 : (reg4275 ? reg4170 : reg4157))));
                      reg4344 <= (!forvar4213);
                    end
                  for (forvar4345 = (1'h0); (forvar4345 < (1'h0)); forvar4345 = (forvar4345 + (1'h1)))
                    begin
                      reg4346 <= {({(reg4331 ? reg4285 : (8'hb1))} ?
                              $unsigned((reg4159 ?
                                  reg4331 : forvar4175)) : (-(reg4222 << (8'ha3))))};
                      reg4347 <= (^~$unsigned($signed(reg4173)));
                      reg4348 <= {reg4167};
                      reg4349 <= reg4320;
                    end
                  if (reg4157)
                    begin
                      reg4350 <= (|$signed(((reg4347 == reg4343) + (&reg4185))));
                      reg4351 <= (reg4195[(3'h5):(3'h4)] ?
                          reg4327 : $signed(reg4251));
                      reg4352 <= ($unsigned(reg4244[(3'h5):(3'h4)]) ?
                          ({(8'ha5)} ?
                              reg4270 : ($signed(reg4290) ?
                                  reg4264[(4'ha):(2'h2)] : (reg4162 ?
                                      reg4273 : forvar4300))) : reg4225[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg4350 <= (~|forvar4323);
                    end
                end
              if (forvar4308[(3'h4):(2'h3)])
                begin
                  for (forvar4353 = (1'h0); (forvar4353 < (1'h1)); forvar4353 = (forvar4353 + (1'h1)))
                    begin
                      reg4354 <= $unsigned((~(reg4185 ?
                          reg4163[(3'h7):(1'h1)] : reg4279[(3'h4):(3'h4)])));
                      reg4355 <= $unsigned((+$signed(((8'haf) ?
                          reg4155 : (8'hb7)))));
                      reg4356 <= reg4279;
                    end
                  if (reg4351)
                    begin
                      reg4357 <= (($signed($signed(reg4296)) && $signed(reg4183)) >>> $signed($signed((&reg4200))));
                      reg4358 <= reg4330;
                      reg4359 <= (((^reg4261) <= reg4183) ?
                          (&(!(^forvar4174))) : {(~|$unsigned(forvar4353))});
                      reg4360 <= ((!reg4219) <<< forvar4184);
                    end
                  else
                    begin
                      reg4357 <= $unsigned(forvar4312);
                      reg4358 <= reg4357[(3'h4):(3'h4)];
                      reg4359 <= (|$unsigned(($unsigned(reg4237) ^~ $signed(reg4196))));
                    end
                  if (forvar4193)
                    begin
                      reg4361 <= {(reg4186[(4'h8):(3'h4)] ?
                              {(~&(8'hb6))} : reg4332)};
                      reg4362 <= reg4191[(2'h3):(2'h2)];
                      reg4363 <= $signed((reg4162[(2'h3):(1'h1)] <<< (reg4330[(4'h9):(2'h2)] && ((8'hb2) ^ forvar4197))));
                    end
                  else
                    begin
                      reg4361 <= ({($signed(forvar4308) ?
                              (|forvar4323) : (reg4288 && reg4275))} >> {(~&(reg4301 > reg4211))});
                      reg4362 <= forvar4247[(2'h3):(2'h3)];
                      reg4363 <= (reg4240 ?
                          ({{(8'ha6)}} || ((forvar4153 ?
                              forvar4331 : reg4348) * {reg4181})) : $signed($signed((^reg4260))));
                    end
                  reg4364 <= $unsigned(($unsigned($unsigned(forvar4254)) ?
                      {$signed((8'h9c))} : reg4181[(1'h1):(1'h0)]));
                end
              else
                begin
                  for (forvar4353 = (1'h0); (forvar4353 < (1'h0)); forvar4353 = (forvar4353 + (1'h1)))
                    begin
                      reg4354 <= (~|((&forvar4176) ? reg4223 : forvar4336));
                    end
                  reg4355 <= $signed((reg4360 ?
                      reg4304[(3'h4):(2'h2)] : {(+reg4244)}));
                  for (forvar4356 = (1'h0); (forvar4356 < (2'h2)); forvar4356 = (forvar4356 + (1'h1)))
                    begin
                      reg4357 <= (-$unsigned($signed(reg4250)));
                    end
                  reg4358 <= (((reg4166 ?
                          $unsigned(reg4354) : $unsigned((8'h9e))) || forvar4254) ?
                      (forvar4184 ?
                          (reg4364 ?
                              $unsigned((8'hb7)) : $unsigned((8'haa))) : (+{reg4188})) : (((!forvar4208) && {reg4202}) <= ((reg4352 << (8'hba)) && (8'hb3))));
                end
              if (((-reg4349[(2'h3):(2'h3)]) ?
                  $signed({(~reg4346)}) : {reg4339}))
                begin
                  if ($unsigned($signed(reg4360[(1'h1):(1'h1)])))
                    begin
                      reg4365 <= (+(reg4343[(1'h0):(1'h0)] >> $signed((8'hb0))));
                      reg4366 <= ((((reg4166 >> (8'ha1)) ?
                              (~|forvar4161) : (reg4236 ? reg4359 : (8'haf))) ?
                          $unsigned($signed(reg4264)) : $signed($signed(reg4273))) >> $unsigned((8'h9e)));
                      reg4367 <= reg4234[(4'hd):(4'h8)];
                    end
                  else
                    begin
                      reg4365 <= ($unsigned((!(wire632 ?
                              (8'ha3) : forvar4239))) ?
                          ((^forvar4153) ~^ $unsigned((forvar4356 > (8'h9c)))) : wire638[(4'h8):(4'h8)]);
                      reg4366 <= (-(((reg4156 == reg4333) >>> (8'hae)) || reg4315));
                    end
                  for (forvar4368 = (1'h0); (forvar4368 < (2'h3)); forvar4368 = (forvar4368 + (1'h1)))
                    begin
                      reg4369 <= (|(~^forvar4199[(3'h7):(2'h2)]));
                      reg4370 <= $unsigned((!forvar4199));
                      reg4371 <= reg4173;
                    end
                  reg4372 <= $signed($signed((((8'hb4) ?
                      (8'hb9) : reg4186) == $signed(reg4297))));
                  for (forvar4373 = (1'h0); (forvar4373 < (2'h3)); forvar4373 = (forvar4373 + (1'h1)))
                    begin
                      reg4374 <= (^(forvar4276[(3'h6):(2'h3)] << {reg4160}));
                      reg4375 <= {(~|(!((8'haf) ? reg4302 : (8'h9c))))};
                    end
                end
              else
                begin
                  for (forvar4365 = (1'h0); (forvar4365 < (1'h0)); forvar4365 = (forvar4365 + (1'h1)))
                    begin
                      reg4366 <= (reg4168 * forvar4312[(4'ha):(4'h9)]);
                      reg4367 <= forvar4373[(2'h2):(1'h1)];
                    end
                  if ((^$signed((-reg4356[(4'hb):(2'h2)]))))
                    begin
                      reg4368 <= ((&((reg4230 | reg4198) ?
                              $unsigned(reg4361) : reg4264)) ?
                          $signed(forvar4155[(4'h8):(2'h3)]) : ($unsigned(reg4355) ?
                              reg4350 : (-(reg4201 ? reg4158 : forvar4199))));
                      reg4369 <= reg4319[(2'h2):(1'h1)];
                      reg4370 <= reg4280;
                    end
                  else
                    begin
                      reg4368 <= forvar4278[(3'h6):(3'h4)];
                      reg4369 <= {(8'ha6)};
                      reg4370 <= $unsigned($unsigned(reg4300[(1'h0):(1'h0)]));
                      reg4371 <= forvar4277;
                    end
                  if ((!reg4250))
                    begin
                      reg4372 <= $unsigned((reg4170 <<< (8'ha2)));
                      reg4373 <= (~|{{((8'hab) ~^ forvar4246)}});
                      reg4374 <= forvar4277[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg4372 <= forvar4268[(3'h4):(1'h0)];
                      reg4373 <= {{({(8'hb2)} <= (reg4286 ?
                                  reg4309 : (8'hb0)))}};
                      reg4374 <= (8'hab);
                    end
                  for (forvar4375 = (1'h0); (forvar4375 < (2'h2)); forvar4375 = (forvar4375 + (1'h1)))
                    begin
                      reg4376 <= ({(+((8'ha4) ?
                              forvar4153 : forvar4247))} * reg4317[(4'h9):(3'h6)]);
                    end
                end
            end
          for (forvar4377 = (1'h0); (forvar4377 < (2'h3)); forvar4377 = (forvar4377 + (1'h1)))
            begin
              for (forvar4378 = (1'h0); (forvar4378 < (1'h1)); forvar4378 = (forvar4378 + (1'h1)))
                begin
                  for (forvar4379 = (1'h0); (forvar4379 < (2'h3)); forvar4379 = (forvar4379 + (1'h1)))
                    begin
                      reg4380 <= ({forvar4208} ?
                          $unsigned({reg4299}) : $signed(reg4206));
                      reg4381 <= reg4370[(2'h2):(1'h1)];
                    end
                  reg4382 <= {$signed(reg4182)};
                end
            end
        end
    end
  assign wire4383 = $unsigned(reg4300);
  assign wire4384 = $signed($signed($signed($signed((8'hb1)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module9  (y, clk, wire13, wire12, wire11, wire10);
  output wire [(32'h99f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire13;
  input wire [(3'h5):(1'h0)] wire12;
  input wire [(4'h9):(1'h0)] wire11;
  input wire [(3'h5):(1'h0)] wire10;
  wire [(3'h6):(1'h0)] wire620;
  wire [(4'he):(1'h0)] wire618;
  wire signed [(3'h6):(1'h0)] wire205;
  wire signed [(4'he):(1'h0)] wire204;
  wire [(4'ha):(1'h0)] wire203;
  wire [(3'h6):(1'h0)] wire202;
  wire signed [(4'hf):(1'h0)] wire201;
  wire signed [(4'h9):(1'h0)] wire200;
  wire signed [(3'h7):(1'h0)] wire199;
  wire [(4'hd):(1'h0)] wire198;
  wire signed [(4'hc):(1'h0)] wire197;
  wire signed [(3'h4):(1'h0)] wire196;
  wire [(4'hf):(1'h0)] wire195;
  reg signed [(4'hc):(1'h0)] reg194 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar185 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg184 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg179 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar176 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg174 = (1'h0);
  reg [(2'h2):(1'h0)] reg173 = (1'h0);
  reg [(3'h6):(1'h0)] reg170 = (1'h0);
  reg [(4'hf):(1'h0)] reg193 = (1'h0);
  reg signed [(4'he):(1'h0)] reg192 = (1'h0);
  reg [(4'hf):(1'h0)] reg191 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg190 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg189 = (1'h0);
  reg [(4'hd):(1'h0)] forvar188 = (1'h0);
  reg [(4'hb):(1'h0)] reg187 = (1'h0);
  reg [(4'hc):(1'h0)] forvar186 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg185 = (1'h0);
  reg [(4'hc):(1'h0)] forvar184 = (1'h0);
  reg [(2'h3):(1'h0)] reg183 = (1'h0);
  reg signed [(4'he):(1'h0)] reg182 = (1'h0);
  reg [(5'h10):(1'h0)] reg181 = (1'h0);
  reg [(3'h6):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar179 = (1'h0);
  reg [(3'h5):(1'h0)] reg178 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg177 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg175 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar174 = (1'h0);
  reg [(4'hc):(1'h0)] forvar173 = (1'h0);
  reg [(3'h6):(1'h0)] reg172 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar171 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar170 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar132 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar133 = (1'h0);
  reg [(2'h3):(1'h0)] forvar131 = (1'h0);
  reg [(4'hc):(1'h0)] forvar126 = (1'h0);
  reg [(2'h2):(1'h0)] reg125 = (1'h0);
  reg [(3'h6):(1'h0)] reg129 = (1'h0);
  reg [(4'he):(1'h0)] reg128 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg168 = (1'h0);
  reg [(4'hd):(1'h0)] reg167 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar166 = (1'h0);
  reg [(5'h10):(1'h0)] reg165 = (1'h0);
  reg [(4'he):(1'h0)] reg164 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar163 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar162 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg161 = (1'h0);
  reg [(4'h9):(1'h0)] reg160 = (1'h0);
  reg [(4'h8):(1'h0)] forvar159 = (1'h0);
  reg [(2'h2):(1'h0)] reg158 = (1'h0);
  reg [(5'h10):(1'h0)] reg157 = (1'h0);
  reg [(3'h6):(1'h0)] reg156 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg155 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg153 = (1'h0);
  reg [(4'hc):(1'h0)] reg152 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar151 = (1'h0);
  reg [(4'hc):(1'h0)] reg150 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar149 = (1'h0);
  reg [(4'h9):(1'h0)] reg148 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar147 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar146 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg145 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg143 = (1'h0);
  reg [(5'h10):(1'h0)] forvar142 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg141 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg140 = (1'h0);
  reg [(3'h6):(1'h0)] reg139 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar138 = (1'h0);
  reg [(4'he):(1'h0)] reg137 = (1'h0);
  reg [(4'hd):(1'h0)] reg136 = (1'h0);
  reg [(3'h5):(1'h0)] reg135 = (1'h0);
  reg [(4'h9):(1'h0)] reg134 = (1'h0);
  reg [(4'ha):(1'h0)] reg133 = (1'h0);
  reg [(5'h10):(1'h0)] reg132 = (1'h0);
  reg [(3'h5):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg130 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar129 = (1'h0);
  reg [(4'h8):(1'h0)] forvar128 = (1'h0);
  reg signed [(4'he):(1'h0)] reg127 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg126 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar125 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg123 = (1'h0);
  reg [(2'h3):(1'h0)] reg122 = (1'h0);
  reg [(3'h6):(1'h0)] reg121 = (1'h0);
  reg signed [(4'he):(1'h0)] reg120 = (1'h0);
  reg [(4'h9):(1'h0)] reg119 = (1'h0);
  reg [(4'hd):(1'h0)] reg118 = (1'h0);
  reg [(4'hf):(1'h0)] reg117 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar116 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar115 = (1'h0);
  reg [(4'ha):(1'h0)] reg114 = (1'h0);
  reg [(4'hd):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar112 = (1'h0);
  reg [(4'hc):(1'h0)] reg111 = (1'h0);
  reg signed [(4'he):(1'h0)] reg110 = (1'h0);
  reg [(4'h8):(1'h0)] forvar102 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg96 = (1'h0);
  reg signed [(4'he):(1'h0)] reg109 = (1'h0);
  reg [(4'hb):(1'h0)] reg108 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar107 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg106 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg105 = (1'h0);
  reg signed [(4'he):(1'h0)] reg104 = (1'h0);
  reg signed [(4'he):(1'h0)] reg103 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg98 = (1'h0);
  reg [(4'h8):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg101 = (1'h0);
  reg [(5'h10):(1'h0)] reg100 = (1'h0);
  reg [(5'h10):(1'h0)] reg99 = (1'h0);
  reg [(4'ha):(1'h0)] forvar98 = (1'h0);
  reg [(5'h10):(1'h0)] reg97 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar96 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar95 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg94 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg93 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar90 = (1'h0);
  reg [(4'hf):(1'h0)] forvar85 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg81 = (1'h0);
  reg [(4'h8):(1'h0)] forvar80 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg77 = (1'h0);
  reg [(2'h2):(1'h0)] forvar76 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar75 = (1'h0);
  reg [(3'h7):(1'h0)] reg72 = (1'h0);
  reg [(4'h9):(1'h0)] reg71 = (1'h0);
  reg [(3'h6):(1'h0)] forvar69 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg60 = (1'h0);
  reg [(4'ha):(1'h0)] forvar55 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg91 = (1'h0);
  reg [(2'h2):(1'h0)] reg90 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg89 = (1'h0);
  reg [(4'he):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg87 = (1'h0);
  reg [(4'hb):(1'h0)] reg86 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg85 = (1'h0);
  reg [(4'h9):(1'h0)] reg84 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg83 = (1'h0);
  reg signed [(4'he):(1'h0)] reg82 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar81 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg80 = (1'h0);
  reg [(4'hf):(1'h0)] reg79 = (1'h0);
  reg [(4'hc):(1'h0)] reg78 = (1'h0);
  reg [(2'h2):(1'h0)] forvar77 = (1'h0);
  reg [(3'h7):(1'h0)] reg76 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg75 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg74 = (1'h0);
  reg signed [(4'he):(1'h0)] reg73 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar72 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar71 = (1'h0);
  reg [(3'h5):(1'h0)] reg70 = (1'h0);
  reg signed [(4'he):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg68 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar66 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg64 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar63 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg61 = (1'h0);
  reg [(4'hd):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg53 = (1'h0);
  reg [(5'h10):(1'h0)] forvar52 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar51 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg50 = (1'h0);
  reg [(2'h3):(1'h0)] reg49 = (1'h0);
  reg signed [(4'he):(1'h0)] reg48 = (1'h0);
  reg [(4'ha):(1'h0)] forvar42 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar36 = (1'h0);
  reg [(4'hb):(1'h0)] forvar34 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar28 = (1'h0);
  reg [(4'hb):(1'h0)] reg40 = (1'h0);
  reg [(4'h9):(1'h0)] reg39 = (1'h0);
  reg [(4'hc):(1'h0)] forvar38 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar35 = (1'h0);
  reg [(4'h8):(1'h0)] forvar30 = (1'h0);
  reg signed [(4'he):(1'h0)] reg29 = (1'h0);
  reg [(4'hc):(1'h0)] forvar27 = (1'h0);
  reg signed [(4'he):(1'h0)] reg25 = (1'h0);
  reg [(2'h3):(1'h0)] forvar22 = (1'h0);
  reg [(4'hb):(1'h0)] reg20 = (1'h0);
  reg [(4'hf):(1'h0)] reg19 = (1'h0);
  reg [(4'hf):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg66 = (1'h0);
  reg [(4'hc):(1'h0)] reg65 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar64 = (1'h0);
  reg [(3'h7):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg62 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar61 = (1'h0);
  reg [(4'hf):(1'h0)] forvar60 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg58 = (1'h0);
  reg [(4'hf):(1'h0)] forvar57 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg56 = (1'h0);
  reg [(3'h5):(1'h0)] reg55 = (1'h0);
  reg [(5'h10):(1'h0)] reg54 = (1'h0);
  reg [(2'h3):(1'h0)] forvar53 = (1'h0);
  reg [(3'h4):(1'h0)] reg52 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg51 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar50 = (1'h0);
  reg [(3'h5):(1'h0)] forvar49 = (1'h0);
  reg [(3'h6):(1'h0)] forvar48 = (1'h0);
  reg [(4'hd):(1'h0)] reg47 = (1'h0);
  reg [(5'h10):(1'h0)] reg46 = (1'h0);
  reg [(2'h3):(1'h0)] reg45 = (1'h0);
  reg [(3'h5):(1'h0)] reg44 = (1'h0);
  reg [(4'he):(1'h0)] reg43 = (1'h0);
  reg [(3'h7):(1'h0)] reg42 = (1'h0);
  reg [(4'ha):(1'h0)] reg41 = (1'h0);
  reg [(4'hd):(1'h0)] forvar40 = (1'h0);
  reg [(2'h2):(1'h0)] forvar39 = (1'h0);
  reg [(5'h10):(1'h0)] reg38 = (1'h0);
  reg [(5'h10):(1'h0)] reg37 = (1'h0);
  reg [(4'hd):(1'h0)] reg36 = (1'h0);
  reg [(4'h8):(1'h0)] reg35 = (1'h0);
  reg [(3'h4):(1'h0)] reg34 = (1'h0);
  reg [(5'h10):(1'h0)] reg33 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg32 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg31 = (1'h0);
  reg [(4'hb):(1'h0)] reg30 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar29 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg28 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg27 = (1'h0);
  reg [(3'h6):(1'h0)] reg26 = (1'h0);
  reg [(4'h8):(1'h0)] forvar25 = (1'h0);
  reg [(4'ha):(1'h0)] reg24 = (1'h0);
  reg [(2'h3):(1'h0)] reg23 = (1'h0);
  reg [(4'hd):(1'h0)] reg22 = (1'h0);
  reg signed [(4'he):(1'h0)] reg21 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar20 = (1'h0);
  reg [(4'hb):(1'h0)] forvar19 = (1'h0);
  reg [(4'hd):(1'h0)] forvar18 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire17;
  wire signed [(4'hf):(1'h0)] wire16;
  wire signed [(3'h6):(1'h0)] wire15;
  wire [(4'hc):(1'h0)] wire14;
  assign y = {wire620,
                 wire618,
                 wire205,
                 wire204,
                 wire203,
                 wire202,
                 wire201,
                 wire200,
                 wire199,
                 wire198,
                 wire197,
                 wire196,
                 wire195,
                 reg194,
                 forvar185,
                 reg184,
                 reg179,
                 forvar176,
                 reg174,
                 reg173,
                 reg170,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 forvar188,
                 reg187,
                 forvar186,
                 reg185,
                 forvar184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 forvar179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 forvar174,
                 forvar173,
                 reg172,
                 forvar171,
                 forvar170,
                 forvar132,
                 forvar133,
                 forvar131,
                 forvar126,
                 reg125,
                 reg129,
                 reg128,
                 reg169,
                 reg168,
                 reg167,
                 forvar166,
                 reg165,
                 reg164,
                 forvar163,
                 forvar162,
                 reg161,
                 reg160,
                 forvar159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 forvar151,
                 reg150,
                 forvar149,
                 reg148,
                 forvar147,
                 forvar146,
                 reg145,
                 reg144,
                 reg143,
                 forvar142,
                 reg141,
                 reg140,
                 reg139,
                 forvar138,
                 reg137,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 forvar129,
                 forvar128,
                 reg127,
                 reg126,
                 forvar125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 forvar116,
                 forvar115,
                 reg114,
                 reg113,
                 forvar112,
                 reg111,
                 reg110,
                 forvar102,
                 reg96,
                 reg109,
                 reg108,
                 forvar107,
                 reg106,
                 reg105,
                 reg104,
                 reg103,
                 reg98,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 forvar98,
                 reg97,
                 forvar96,
                 forvar95,
                 reg94,
                 reg93,
                 forvar90,
                 forvar85,
                 reg81,
                 forvar80,
                 reg77,
                 forvar76,
                 forvar75,
                 reg72,
                 reg71,
                 forvar69,
                 reg60,
                 forvar55,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 forvar81,
                 reg80,
                 reg79,
                 reg78,
                 forvar77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 forvar72,
                 forvar71,
                 reg70,
                 reg69,
                 reg68,
                 forvar66,
                 reg64,
                 forvar63,
                 reg61,
                 reg57,
                 reg53,
                 forvar52,
                 forvar51,
                 reg50,
                 reg49,
                 reg48,
                 forvar42,
                 forvar36,
                 forvar34,
                 forvar28,
                 reg40,
                 reg39,
                 forvar38,
                 forvar35,
                 forvar30,
                 reg29,
                 forvar27,
                 reg25,
                 forvar22,
                 reg20,
                 reg19,
                 reg67,
                 reg66,
                 reg65,
                 forvar64,
                 reg63,
                 reg62,
                 forvar61,
                 forvar60,
                 reg59,
                 reg58,
                 forvar57,
                 reg56,
                 reg55,
                 reg54,
                 forvar53,
                 reg52,
                 reg51,
                 forvar50,
                 forvar49,
                 forvar48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 forvar40,
                 forvar39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 forvar29,
                 reg28,
                 reg27,
                 reg26,
                 forvar25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 forvar20,
                 forvar19,
                 forvar18,
                 wire17,
                 wire16,
                 wire15,
                 wire14,
                 (1'h0)};
  assign wire14 = wire11[(3'h6):(3'h6)];
  assign wire15 = (^~wire13);
  assign wire16 = wire12[(1'h1):(1'h0)];
  assign wire17 = wire15[(2'h3):(1'h1)];
  always
    @(posedge clk) begin
      if (($signed($unsigned(((8'ha2) ? wire17 : (8'ha6)))) ?
          $signed(($signed(wire11) == (wire17 <<< (8'hb2)))) : ((wire11[(4'h9):(2'h3)] << ((8'hb2) ?
              wire14 : wire14)) & $signed((wire11 <= wire15)))))
        begin
          for (forvar18 = (1'h0); (forvar18 < (1'h0)); forvar18 = (forvar18 + (1'h1)))
            begin
              for (forvar19 = (1'h0); (forvar19 < (2'h2)); forvar19 = (forvar19 + (1'h1)))
                begin
                  for (forvar20 = (1'h0); (forvar20 < (2'h3)); forvar20 = (forvar20 + (1'h1)))
                    begin
                      reg21 <= forvar18;
                      reg22 <= wire14;
                      reg23 <= wire14[(4'ha):(1'h1)];
                      reg24 <= {(forvar20[(2'h2):(1'h1)] ?
                              wire15[(3'h4):(2'h3)] : (+(reg21 & wire11)))};
                    end
                  for (forvar25 = (1'h0); (forvar25 < (1'h0)); forvar25 = (forvar25 + (1'h1)))
                    begin
                      reg26 <= (!forvar25);
                      reg27 <= forvar19[(4'h8):(1'h1)];
                      reg28 <= wire13[(1'h1):(1'h0)];
                    end
                  for (forvar29 = (1'h0); (forvar29 < (2'h2)); forvar29 = (forvar29 + (1'h1)))
                    begin
                      reg30 <= ($signed(((^~wire17) ?
                          (forvar29 ?
                              wire16 : wire10) : (forvar18 >>> wire15))) >>> (&$signed((forvar18 >> reg23))));
                      reg31 <= wire16;
                    end
                  if ($unsigned((forvar18 ?
                      reg23[(1'h1):(1'h1)] : (forvar19[(4'hb):(4'h8)] ?
                          (wire13 ? reg24 : reg31) : (wire17 & reg28)))))
                    begin
                      reg32 <= ((-$signed((reg26 - reg26))) * {reg30[(3'h5):(2'h3)]});
                      reg33 <= reg26[(2'h2):(1'h0)];
                      reg34 <= reg23;
                    end
                  else
                    begin
                      reg32 <= $signed($signed((^~$signed((8'hb1)))));
                      reg33 <= (^~$signed((|(8'ha1))));
                    end
                end
              if (((reg21 ?
                  (|((8'ha5) ? reg23 : wire17)) : ((|wire12) ?
                      (reg22 ? forvar25 : (8'hb0)) : (reg34 ?
                          (8'ha0) : reg26))) ^~ (reg34[(2'h2):(1'h0)] ?
                  (reg23 ?
                      ((8'h9e) ?
                          reg27 : reg21) : $unsigned(wire13)) : forvar20[(1'h1):(1'h0)])))
                begin
                  if (wire14[(4'hb):(4'h8)])
                    begin
                      reg35 <= (-$signed(reg22));
                    end
                  else
                    begin
                      reg35 <= $signed(reg28[(4'h8):(2'h3)]);
                      reg36 <= (^~{wire15[(3'h5):(3'h5)]});
                      reg37 <= ({($unsigned(reg31) <= (~&wire11))} >> $unsigned($signed($signed(reg31))));
                    end
                  if (((^~reg21) ?
                      reg23[(1'h0):(1'h0)] : wire14[(3'h6):(2'h3)]))
                    begin
                      reg38 <= (^(-wire15[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg38 <= {(((-reg37) ?
                              $signed((8'had)) : (reg32 != wire10)) + (forvar19[(2'h3):(2'h2)] ?
                              (forvar19 >>> reg28) : {reg32}))};
                    end
                end
              else
                begin
                  if ((8'ha3))
                    begin
                      reg35 <= reg35[(2'h2):(1'h1)];
                      reg36 <= reg35[(3'h7):(2'h2)];
                    end
                  else
                    begin
                      reg35 <= (((&(forvar29 ?
                          forvar18 : wire15)) >> $unsigned(wire13[(2'h3):(2'h3)])) || $signed(reg38));
                    end
                end
              for (forvar39 = (1'h0); (forvar39 < (2'h3)); forvar39 = (forvar39 + (1'h1)))
                begin
                  for (forvar40 = (1'h0); (forvar40 < (2'h2)); forvar40 = (forvar40 + (1'h1)))
                    begin
                      reg41 <= $signed($unsigned(wire13[(1'h1):(1'h1)]));
                      reg42 <= (~&forvar19);
                      reg43 <= reg21[(4'h8):(3'h5)];
                    end
                  if (((reg37 ? $unsigned({wire13}) : forvar20) ?
                      ({(~^(8'hb2))} ?
                          reg41 : (forvar19 >>> $signed(reg41))) : (^{$signed(wire16)})))
                    begin
                      reg44 <= ($signed(reg27) ^ $unsigned(((~&reg24) << reg38[(4'ha):(3'h7)])));
                      reg45 <= wire14;
                      reg46 <= reg27[(4'h9):(2'h3)];
                      reg47 <= $unsigned(reg30);
                    end
                  else
                    begin
                      reg44 <= ({reg32} ?
                          $unsigned(((~^reg28) ?
                              $signed(reg33) : $unsigned((8'hb3)))) : ({((8'hb2) != reg23)} >> $unsigned((wire13 <<< reg47))));
                      reg45 <= (~&{forvar40});
                      reg46 <= ($unsigned((~&reg43)) & (reg46[(4'hd):(3'h4)] > $signed((reg44 > (8'hb3)))));
                      reg47 <= ($signed(($unsigned(forvar20) >= $signed(forvar18))) | ((~^$unsigned(reg36)) ?
                          reg23 : {forvar39}));
                    end
                end
            end
          for (forvar48 = (1'h0); (forvar48 < (2'h2)); forvar48 = (forvar48 + (1'h1)))
            begin
              for (forvar49 = (1'h0); (forvar49 < (1'h1)); forvar49 = (forvar49 + (1'h1)))
                begin
                  for (forvar50 = (1'h0); (forvar50 < (1'h1)); forvar50 = (forvar50 + (1'h1)))
                    begin
                      reg51 <= $signed(({reg28} ?
                          (~&reg34[(1'h1):(1'h1)]) : (((8'h9f) ?
                                  reg35 : reg30) ?
                              $unsigned(wire11) : wire17)));
                      reg52 <= $signed({(!(8'hb1))});
                    end
                  for (forvar53 = (1'h0); (forvar53 < (1'h1)); forvar53 = (forvar53 + (1'h1)))
                    begin
                      reg54 <= $unsigned(forvar49);
                      reg55 <= reg54;
                      reg56 <= $unsigned(reg21);
                    end
                end
              for (forvar57 = (1'h0); (forvar57 < (1'h1)); forvar57 = (forvar57 + (1'h1)))
                begin
                  if (forvar48[(3'h6):(3'h5)])
                    begin
                      reg58 <= $signed($signed($signed(((8'h9c) ?
                          reg45 : reg31))));
                    end
                  else
                    begin
                      reg58 <= (8'hb2);
                      reg59 <= $unsigned((8'ha4));
                    end
                end
              for (forvar60 = (1'h0); (forvar60 < (1'h1)); forvar60 = (forvar60 + (1'h1)))
                begin
                  for (forvar61 = (1'h0); (forvar61 < (2'h3)); forvar61 = (forvar61 + (1'h1)))
                    begin
                      reg62 <= (~^((-reg51[(1'h0):(1'h0)]) <<< ((forvar48 || (8'hae)) > $unsigned(reg37))));
                      reg63 <= (($unsigned($signed(forvar25)) <<< $unsigned(wire16[(4'hc):(4'hb)])) ?
                          wire16[(1'h1):(1'h0)] : $signed({(&wire15)}));
                    end
                  for (forvar64 = (1'h0); (forvar64 < (1'h0)); forvar64 = (forvar64 + (1'h1)))
                    begin
                      reg65 <= ($unsigned((reg22[(3'h6):(1'h1)] & wire11)) ?
                          (reg24 | (-reg52[(1'h1):(1'h1)])) : (~$unsigned($signed(wire17))));
                    end
                end
            end
          reg66 <= (8'ha8);
          reg67 <= {(^$signed($signed(reg65)))};
        end
      else
        begin
          for (forvar18 = (1'h0); (forvar18 < (1'h1)); forvar18 = (forvar18 + (1'h1)))
            begin
              if (({(reg63[(3'h4):(2'h3)] != $signed(reg38))} || (+(wire12 ?
                  reg21 : (!forvar19)))))
                begin
                  if (reg31[(3'h6):(1'h0)])
                    begin
                      reg19 <= ((+reg44) ?
                          (&(reg47[(3'h6):(2'h2)] ?
                              $unsigned(forvar25) : forvar64[(1'h0):(1'h0)])) : (forvar18[(2'h3):(2'h2)] ?
                              ((^forvar48) ?
                                  $unsigned(forvar39) : ((8'hae) ?
                                      reg27 : reg32)) : forvar64));
                      reg20 <= ((~|({wire15} ?
                              (~&reg43) : (reg41 ^~ (8'ha3)))) ?
                          $unsigned($unsigned((reg36 ?
                              wire17 : reg26))) : $signed($unsigned(wire12)));
                    end
                  else
                    begin
                      reg19 <= (+$signed($unsigned($signed(forvar20))));
                      reg20 <= {reg47[(3'h5):(3'h5)]};
                    end
                end
              else
                begin
                  reg19 <= (&$unsigned($unsigned(forvar50[(4'h9):(1'h0)])));
                  if (reg55)
                    begin
                      reg20 <= (reg59 < $signed(forvar49[(2'h2):(1'h1)]));
                      reg21 <= $unsigned($signed(reg67));
                    end
                  else
                    begin
                      reg20 <= $unsigned(reg54[(3'h4):(1'h1)]);
                    end
                  for (forvar22 = (1'h0); (forvar22 < (1'h1)); forvar22 = (forvar22 + (1'h1)))
                    begin
                      reg23 <= {reg43};
                      reg24 <= (~^($unsigned((reg58 - reg42)) ?
                          $unsigned(reg23) : reg23[(1'h1):(1'h1)]));
                      reg25 <= ((-(~&(&forvar53))) >= (-$unsigned((forvar48 ?
                          reg36 : (8'had)))));
                    end
                end
              reg26 <= $unsigned(reg23);
            end
          if ($unsigned(($signed($signed((8'ha2))) ? reg23 : $signed(reg46))))
            begin
              if ((~($unsigned((reg21 ?
                  reg25 : reg30)) == $unsigned((reg41 <<< wire11)))))
                begin
                  for (forvar27 = (1'h0); (forvar27 < (1'h0)); forvar27 = (forvar27 + (1'h1)))
                    begin
                      reg28 <= (($unsigned(reg31[(3'h7):(3'h5)]) ?
                              $signed(forvar25) : ({wire14} <<< reg20[(2'h3):(1'h0)])) ?
                          (|$unsigned((forvar19 && reg32))) : (|wire14));
                      reg29 <= ({$unsigned($signed(reg62))} ?
                          (8'ha4) : wire13[(1'h1):(1'h0)]);
                      reg30 <= forvar22;
                    end
                end
              else
                begin
                  if ((^(^~((reg54 ? (8'hac) : reg59) & (wire15 ?
                      reg54 : forvar57)))))
                    begin
                      reg27 <= $signed({reg58});
                      reg28 <= $unsigned(wire15[(1'h1):(1'h1)]);
                      reg29 <= reg37;
                    end
                  else
                    begin
                      reg27 <= $unsigned(reg27[(4'hf):(4'he)]);
                      reg28 <= reg23[(2'h3):(2'h3)];
                    end
                  for (forvar30 = (1'h0); (forvar30 < (2'h3)); forvar30 = (forvar30 + (1'h1)))
                    begin
                      reg31 <= (|($unsigned($signed(reg22)) ?
                          forvar29[(3'h6):(3'h6)] : (8'ha3)));
                      reg32 <= (&(&forvar20));
                      reg33 <= (~|(reg32 >>> $signed(reg23[(1'h1):(1'h1)])));
                      reg34 <= {wire13[(2'h2):(2'h2)]};
                    end
                  for (forvar35 = (1'h0); (forvar35 < (2'h3)); forvar35 = (forvar35 + (1'h1)))
                    begin
                      reg36 <= $unsigned($unsigned({reg31[(3'h5):(1'h1)]}));
                      reg37 <= reg42;
                    end
                  for (forvar38 = (1'h0); (forvar38 < (1'h1)); forvar38 = (forvar38 + (1'h1)))
                    begin
                      reg39 <= reg38;
                      reg40 <= reg26;
                      reg41 <= ((-$signed((^~reg34))) * $unsigned(wire10[(3'h4):(2'h2)]));
                      reg42 <= (&(!$unsigned($signed(reg58))));
                    end
                end
            end
          else
            begin
              for (forvar27 = (1'h0); (forvar27 < (1'h1)); forvar27 = (forvar27 + (1'h1)))
                begin
                  for (forvar28 = (1'h0); (forvar28 < (1'h0)); forvar28 = (forvar28 + (1'h1)))
                    begin
                      reg29 <= reg20[(4'h8):(3'h7)];
                    end
                end
              if ((!reg52[(2'h2):(2'h2)]))
                begin
                  for (forvar30 = (1'h0); (forvar30 < (1'h0)); forvar30 = (forvar30 + (1'h1)))
                    begin
                      reg31 <= (((+$unsigned(reg24)) ?
                              reg32 : $signed((wire15 ? wire14 : reg29))) ?
                          $signed(($signed(reg31) ^ (&reg56))) : $unsigned($unsigned((-reg46))));
                      reg32 <= $unsigned($signed(forvar38));
                      reg33 <= $unsigned($unsigned((-$unsigned((8'hb3)))));
                    end
                  if (reg38[(5'h10):(3'h6)])
                    begin
                      reg34 <= $signed((~&reg30[(3'h7):(2'h3)]));
                      reg35 <= $signed($signed((8'hb2)));
                      reg36 <= (-(reg47 ?
                          forvar39 : ($signed((8'hb8)) ~^ (forvar53 - forvar61))));
                    end
                  else
                    begin
                      reg34 <= reg67;
                    end
                  if ((forvar18[(1'h1):(1'h1)] < (-(forvar22[(2'h2):(1'h1)] ?
                      $signed(forvar38) : $unsigned(wire17)))))
                    begin
                      reg37 <= (((forvar28[(3'h4):(1'h0)] <= $unsigned(reg21)) ?
                              ($signed((8'hac)) ?
                                  {reg39} : forvar30) : $signed((+reg58))) ?
                          reg35[(3'h5):(2'h3)] : $unsigned(reg20[(4'ha):(2'h2)]));
                    end
                  else
                    begin
                      reg37 <= (&{($unsigned(reg34) != (~^wire10))});
                      reg38 <= $unsigned($signed(($unsigned(reg19) | $unsigned((8'hb1)))));
                      reg39 <= ({$unsigned((8'hb3))} < $signed($unsigned(reg26[(3'h5):(1'h1)])));
                    end
                end
              else
                begin
                  if ($signed(reg47[(4'h9):(4'h9)]))
                    begin
                      reg30 <= forvar64[(3'h6):(1'h1)];
                      reg31 <= forvar35;
                    end
                  else
                    begin
                      reg30 <= ($signed(reg54[(3'h4):(3'h4)]) ?
                          $signed((-(+wire10))) : $unsigned(wire17));
                      reg31 <= {reg42[(1'h0):(1'h0)]};
                      reg32 <= $signed(reg27);
                      reg33 <= {{$unsigned((+forvar53))}};
                    end
                  for (forvar34 = (1'h0); (forvar34 < (2'h3)); forvar34 = (forvar34 + (1'h1)))
                    begin
                      reg35 <= reg56;
                    end
                  for (forvar36 = (1'h0); (forvar36 < (2'h3)); forvar36 = (forvar36 + (1'h1)))
                    begin
                      reg37 <= ((forvar40[(3'h7):(1'h1)] ?
                              $signed((reg66 ? reg47 : reg22)) : (wire11 ?
                                  (forvar20 * wire13) : (forvar22 & (8'hb4)))) ?
                          (!reg28[(4'h8):(2'h2)]) : reg27[(4'he):(4'h8)]);
                      reg38 <= (($signed($signed(wire17)) ?
                              ((forvar50 ?
                                  reg51 : wire12) & (!reg44)) : (~$unsigned(reg30))) ?
                          ($unsigned($signed(wire13)) - ((forvar35 <<< forvar40) ?
                              $unsigned(reg31) : {(8'ha3)})) : (+(~&(reg40 > reg45))));
                      reg39 <= (8'hb6);
                    end
                  for (forvar40 = (1'h0); (forvar40 < (1'h1)); forvar40 = (forvar40 + (1'h1)))
                    begin
                      reg41 <= (^~{($unsigned(reg62) ? wire16 : (~|forvar30))});
                    end
                end
              for (forvar42 = (1'h0); (forvar42 < (1'h1)); forvar42 = (forvar42 + (1'h1)))
                begin
                  if ((~|reg22[(4'hd):(4'h8)]))
                    begin
                      reg43 <= (-(^(((8'hb6) ? (8'ha0) : forvar25) ?
                          ((8'hb5) ? reg28 : wire13) : (|forvar22))));
                      reg44 <= (reg52 || forvar35);
                      reg45 <= ($signed((~&reg38)) ?
                          (forvar27 ?
                              (&forvar20) : ($unsigned(forvar50) ^ (|wire11))) : {($signed(reg46) ?
                                  (reg27 ?
                                      reg37 : reg36) : (forvar29 ~^ (8'hb2)))});
                    end
                  else
                    begin
                      reg43 <= forvar29[(4'h9):(3'h6)];
                      reg44 <= $signed($unsigned(reg46[(2'h3):(2'h3)]));
                      reg45 <= ($signed($unsigned($unsigned(forvar53))) ?
                          (((reg43 | (8'hb7)) ~^ ((8'haa) >> wire17)) ?
                              $signed((^forvar39)) : reg46[(4'h9):(2'h2)]) : ((~&(8'hb9)) ?
                              $signed(reg56) : (~&{(8'haa)})));
                      reg46 <= ((((8'ha3) ?
                              (+(8'ha5)) : (reg33 >>> reg67)) == $signed({reg31})) ?
                          forvar50[(4'ha):(3'h5)] : (^~reg30));
                    end
                  if ({{(~|(reg45 ? reg31 : (8'h9d)))}})
                    begin
                      reg47 <= ((((~reg65) ?
                                  ((8'had) ? reg67 : forvar30) : forvar30) ?
                              ($unsigned((8'hb2)) ?
                                  (~^reg66) : (~&reg58)) : (^~wire14)) ?
                          (forvar64 == $unsigned($unsigned(reg56))) : reg63);
                      reg48 <= reg34;
                      reg49 <= $unsigned(reg66[(1'h0):(1'h0)]);
                      reg50 <= {reg59};
                    end
                  else
                    begin
                      reg47 <= ($signed($unsigned($signed((8'hb4)))) ~^ reg28[(1'h0):(1'h0)]);
                      reg48 <= (reg25[(3'h5):(1'h1)] < $signed($unsigned((reg23 ^ forvar57))));
                      reg49 <= (~^reg34[(3'h4):(1'h1)]);
                      reg50 <= reg28[(2'h2):(2'h2)];
                    end
                end
            end
          if ((-((~reg43[(2'h2):(1'h0)]) ?
              $unsigned(forvar49) : (-((8'had) ? forvar19 : forvar27)))))
            begin
              for (forvar51 = (1'h0); (forvar51 < (1'h0)); forvar51 = (forvar51 + (1'h1)))
                begin
                  for (forvar52 = (1'h0); (forvar52 < (1'h1)); forvar52 = (forvar52 + (1'h1)))
                    begin
                      reg53 <= (-$unsigned((&$unsigned(forvar25))));
                      reg54 <= (reg58[(3'h4):(2'h3)] ?
                          $unsigned(reg32) : ((reg28 - $signed(forvar48)) == forvar64[(2'h3):(1'h1)]));
                      reg55 <= {wire16[(4'h9):(4'h8)]};
                    end
                  if ({{reg52}})
                    begin
                      reg56 <= $signed(forvar25[(2'h2):(1'h0)]);
                      reg57 <= forvar38;
                      reg58 <= $unsigned(wire17[(1'h1):(1'h1)]);
                      reg59 <= (((~^(wire12 << forvar29)) ?
                          ($unsigned(reg51) ?
                              reg65[(2'h3):(1'h1)] : $unsigned(forvar40)) : ((~&(8'hb2)) ?
                              ((8'hba) ?
                                  forvar20 : wire10) : reg45[(2'h2):(2'h2)])) == (((reg25 > (8'had)) && $signed(forvar39)) & (reg36[(1'h0):(1'h0)] ?
                          (reg48 ? reg30 : forvar20) : ((8'hb7) << reg53))));
                    end
                  else
                    begin
                      reg56 <= (-(reg20 == $signed(wire16)));
                      reg57 <= $unsigned($unsigned($unsigned($signed(reg58))));
                      reg58 <= ((~&wire13[(2'h2):(1'h1)]) ?
                          (&($signed(forvar39) ^~ $signed(reg45))) : $unsigned({(forvar42 && reg62)}));
                      reg59 <= (8'ha3);
                    end
                end
              for (forvar60 = (1'h0); (forvar60 < (2'h3)); forvar60 = (forvar60 + (1'h1)))
                begin
                  reg61 <= (~|(reg39[(4'h9):(2'h3)] ^~ $unsigned($unsigned(reg63))));
                  reg62 <= ((~&(^~$unsigned(forvar36))) ?
                      $signed($unsigned((~&(8'h9f)))) : {(reg32 ?
                              reg66[(3'h7):(3'h7)] : wire15)});
                  for (forvar63 = (1'h0); (forvar63 < (2'h2)); forvar63 = (forvar63 + (1'h1)))
                    begin
                      reg64 <= reg33;
                      reg65 <= reg58;
                    end
                  for (forvar66 = (1'h0); (forvar66 < (2'h2)); forvar66 = (forvar66 + (1'h1)))
                    begin
                      reg67 <= (&forvar53);
                      reg68 <= (reg62 ?
                          (~&$signed((~reg45))) : wire15[(3'h4):(3'h4)]);
                      reg69 <= ($signed(((reg30 + (8'hba)) ?
                              ((8'hb6) ?
                                  reg40 : wire16) : reg54[(4'h8):(3'h6)])) ?
                          $unsigned(wire10) : (~(8'h9e)));
                      reg70 <= $unsigned($signed($signed((&forvar60))));
                    end
                end
              for (forvar71 = (1'h0); (forvar71 < (2'h3)); forvar71 = (forvar71 + (1'h1)))
                begin
                  for (forvar72 = (1'h0); (forvar72 < (1'h0)); forvar72 = (forvar72 + (1'h1)))
                    begin
                      reg73 <= $signed(forvar61);
                      reg74 <= reg52;
                      reg75 <= ($unsigned(forvar18[(4'hb):(2'h3)]) && ((((8'h9e) ?
                              reg73 : (8'h9c)) || $unsigned(forvar49)) ?
                          {$unsigned(reg24)} : (((8'h9d) ?
                              forvar57 : forvar49) > (reg70 >> wire12))));
                    end
                  reg76 <= $signed(forvar36);
                  for (forvar77 = (1'h0); (forvar77 < (2'h2)); forvar77 = (forvar77 + (1'h1)))
                    begin
                      reg78 <= $signed(reg61[(4'ha):(2'h2)]);
                      reg79 <= (reg61 ? reg46 : (-reg26));
                      reg80 <= $signed($unsigned((+$unsigned(forvar40))));
                    end
                end
              for (forvar81 = (1'h0); (forvar81 < (1'h0)); forvar81 = (forvar81 + (1'h1)))
                begin
                  if (((8'ha5) < reg51))
                    begin
                      reg82 <= {(reg52 ^~ reg54[(3'h6):(3'h5)])};
                      reg83 <= $unsigned($signed((+$signed(reg28))));
                      reg84 <= forvar71;
                    end
                  else
                    begin
                      reg82 <= forvar34[(3'h4):(2'h3)];
                    end
                  if (reg50[(4'h9):(2'h2)])
                    begin
                      reg85 <= reg57;
                      reg86 <= {$signed(forvar20)};
                    end
                  else
                    begin
                      reg85 <= reg54[(1'h0):(1'h0)];
                    end
                  if ($unsigned((~&$unsigned((|reg24)))))
                    begin
                      reg87 <= $unsigned($unsigned((forvar29[(4'h8):(4'h8)] ?
                          $signed(reg66) : forvar20[(4'ha):(4'ha)])));
                    end
                  else
                    begin
                      reg87 <= ({$unsigned($signed(forvar77))} ^~ (((forvar22 >= reg31) ?
                          reg61 : (forvar25 | reg56)) >= $signed($signed(reg74))));
                      reg88 <= ($unsigned(reg39[(3'h6):(1'h1)]) ?
                          reg75[(2'h2):(1'h0)] : (reg39 ? reg40 : (~^{reg87})));
                    end
                  if (({reg33} >>> $unsigned({$unsigned(reg34)})))
                    begin
                      reg89 <= $signed((^(8'ha5)));
                      reg90 <= $unsigned({reg69[(3'h7):(3'h6)]});
                      reg91 <= ((reg39 ?
                              $unsigned($signed(reg51)) : ((^(8'h9f)) >= (forvar63 > reg40))) ?
                          {forvar64[(3'h6):(3'h5)]} : reg34[(1'h1):(1'h1)]);
                      reg92 <= (|$signed(wire14));
                    end
                  else
                    begin
                      reg89 <= $signed((~(&$signed(reg35))));
                      reg90 <= (8'hb1);
                      reg91 <= ((reg24[(4'ha):(3'h4)] || (forvar48 ?
                          reg52 : $signed(forvar18))) < (^(wire14 ^ reg48[(3'h5):(2'h3)])));
                      reg92 <= $unsigned({((~|reg78) == (reg63 ?
                              reg87 : forvar19))});
                    end
                end
            end
          else
            begin
              if ({reg42[(3'h7):(3'h4)]})
                begin
                  for (forvar51 = (1'h0); (forvar51 < (2'h2)); forvar51 = (forvar51 + (1'h1)))
                    begin
                      reg52 <= $unsigned({($unsigned(forvar52) ?
                              $signed((8'hb6)) : $signed(reg42))});
                      reg53 <= $signed(((forvar48[(3'h5):(2'h3)] ?
                          $unsigned(forvar20) : reg49) ^ $signed((~reg88))));
                      reg54 <= $signed((|((~&(8'hb8)) + ((8'hb4) ^~ reg40))));
                    end
                  for (forvar55 = (1'h0); (forvar55 < (2'h3)); forvar55 = (forvar55 + (1'h1)))
                    begin
                      reg56 <= $unsigned(reg50[(3'h7):(2'h2)]);
                      reg57 <= $unsigned((+$signed(reg50[(2'h2):(1'h0)])));
                      reg58 <= (($signed(reg37) >> ((reg42 + reg52) && $unsigned(reg25))) >>> $unsigned(reg31));
                    end
                  if ($signed(forvar27[(3'h5):(1'h0)]))
                    begin
                      reg59 <= ((!{(reg56 ?
                              forvar39 : reg20)}) == reg80[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg59 <= ((reg49 < forvar71) ?
                          (reg92 ?
                              $signed((^reg52)) : {{reg19}}) : $unsigned($signed(reg57)));
                      reg60 <= (&$signed({$unsigned(reg58)}));
                      reg61 <= $signed($signed((^(8'hac))));
                    end
                  if (forvar39[(1'h0):(1'h0)])
                    begin
                      reg62 <= (~$unsigned($unsigned((+(8'h9c)))));
                      reg63 <= $signed(forvar81[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg62 <= $signed(reg39);
                      reg63 <= $signed((~({forvar63} ^~ reg35)));
                      reg64 <= (~&(^(!(reg33 ^ reg37))));
                      reg65 <= reg82;
                    end
                end
              else
                begin
                  if ($unsigned(($unsigned($unsigned(reg64)) << forvar60[(4'hf):(1'h1)])))
                    begin
                      reg51 <= $unsigned(forvar61);
                      reg52 <= (^reg24[(4'ha):(4'ha)]);
                      reg53 <= (($unsigned($unsigned((8'ha8))) == ({reg87} * $signed(reg60))) && ((8'hb7) ?
                          $signed(reg21) : forvar72));
                      reg54 <= $unsigned($signed(((reg25 ? (8'hb0) : (8'hb6)) ?
                          {reg19} : $unsigned((8'h9c)))));
                    end
                  else
                    begin
                      reg51 <= $unsigned($unsigned((reg26[(3'h6):(2'h3)] <= $signed(reg40))));
                    end
                end
              if ($unsigned(reg32))
                begin
                  reg66 <= (~|$signed(reg79));
                  reg67 <= $signed((({reg39} ?
                          (reg30 > forvar77) : {forvar51}) ?
                      reg24[(3'h7):(2'h3)] : (^~$unsigned(reg73))));
                  if (((($signed(reg24) >> $unsigned(forvar25)) ?
                      reg62[(2'h2):(1'h1)] : reg78[(2'h2):(1'h0)]) ^~ ({$signed(forvar20)} ?
                      (~(reg89 ? (8'hab) : reg32)) : reg45[(2'h3):(2'h3)])))
                    begin
                      reg68 <= forvar18[(3'h6):(2'h2)];
                      reg69 <= reg64[(4'h9):(3'h6)];
                      reg70 <= forvar49[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg68 <= $signed(reg53);
                    end
                end
              else
                begin
                  if (($signed(($unsigned(reg26) ? (!(8'had)) : (8'hb9))) ?
                      (&$signed((+reg19))) : $signed(reg87)))
                    begin
                      reg66 <= $unsigned((((&forvar35) ?
                              ((8'h9c) * forvar48) : reg19[(1'h1):(1'h0)]) ?
                          {$signed(forvar20)} : $unsigned($unsigned(reg37))));
                    end
                  else
                    begin
                      reg66 <= $signed($unsigned(reg19[(4'hc):(4'ha)]));
                      reg67 <= reg78[(4'hb):(1'h1)];
                      reg68 <= reg29[(4'he):(2'h3)];
                    end
                  for (forvar69 = (1'h0); (forvar69 < (1'h0)); forvar69 = (forvar69 + (1'h1)))
                    begin
                      reg70 <= (-(-$unsigned($signed(reg76))));
                    end
                  reg71 <= (&((reg78 && forvar50) & {forvar19[(3'h7):(1'h0)]}));
                  if (reg75[(1'h0):(1'h0)])
                    begin
                      reg72 <= $signed($unsigned((reg65[(1'h0):(1'h0)] ?
                          (+(8'hb7)) : reg87[(3'h7):(1'h0)])));
                    end
                  else
                    begin
                      reg72 <= reg27[(1'h0):(1'h0)];
                      reg73 <= (reg91 ? (~(~|(^reg21))) : {(8'hb5)});
                      reg74 <= $signed(($signed((~|reg44)) != reg71));
                    end
                end
              for (forvar75 = (1'h0); (forvar75 < (1'h1)); forvar75 = (forvar75 + (1'h1)))
                begin
                  for (forvar76 = (1'h0); (forvar76 < (1'h0)); forvar76 = (forvar76 + (1'h1)))
                    begin
                      reg77 <= ((8'hb7) ?
                          $unsigned(forvar50) : $unsigned(reg90));
                      reg78 <= ($unsigned((-$signed(reg85))) ?
                          (-($signed(wire11) ?
                              (reg59 < reg87) : {(8'ha8)})) : (wire14 ?
                              (forvar63 <= {wire14}) : reg38));
                      reg79 <= $unsigned($signed(reg65[(2'h2):(1'h1)]));
                    end
                  for (forvar80 = (1'h0); (forvar80 < (2'h2)); forvar80 = (forvar80 + (1'h1)))
                    begin
                      reg81 <= reg62[(3'h5):(3'h5)];
                      reg82 <= (reg65 << reg64[(4'hd):(4'h8)]);
                      reg83 <= (~$unsigned($signed($unsigned(reg55))));
                      reg84 <= $signed({$signed(reg63[(1'h0):(1'h0)])});
                    end
                end
              for (forvar85 = (1'h0); (forvar85 < (2'h3)); forvar85 = (forvar85 + (1'h1)))
                begin
                  reg86 <= $unsigned(reg61);
                  if ({$unsigned($signed(wire11[(3'h7):(3'h6)]))})
                    begin
                      reg87 <= (~|$unsigned(reg90));
                    end
                  else
                    begin
                      reg87 <= ($signed(((reg40 & forvar35) ?
                          reg47 : (8'ha7))) ^~ reg76);
                      reg88 <= $unsigned(((-{reg79}) ?
                          forvar66[(4'hb):(2'h3)] : $unsigned((forvar80 ?
                              (8'haf) : forvar81))));
                      reg89 <= ({forvar57} >>> ($signed($signed(forvar20)) ?
                          $signed(reg23) : $signed((~|wire13))));
                    end
                  for (forvar90 = (1'h0); (forvar90 < (2'h2)); forvar90 = (forvar90 + (1'h1)))
                    begin
                      reg91 <= (^~(8'hb5));
                      reg92 <= reg62;
                      reg93 <= ((^reg28[(3'h7):(3'h6)]) | $signed(forvar85));
                      reg94 <= ((forvar49[(3'h5):(1'h1)] & {$signed(reg24)}) ?
                          (-(forvar35[(2'h3):(2'h3)] ?
                              (reg74 ?
                                  wire14 : (8'hb6)) : $unsigned((8'ha8)))) : (~|$unsigned((reg31 ?
                              (8'hb2) : forvar19))));
                    end
                end
            end
          if (wire17[(1'h1):(1'h0)])
            begin
              for (forvar95 = (1'h0); (forvar95 < (2'h3)); forvar95 = (forvar95 + (1'h1)))
                begin
                  for (forvar96 = (1'h0); (forvar96 < (1'h0)); forvar96 = (forvar96 + (1'h1)))
                    begin
                      reg97 <= $signed((8'ha9));
                    end
                end
              if ((8'h9d))
                begin
                  for (forvar98 = (1'h0); (forvar98 < (1'h0)); forvar98 = (forvar98 + (1'h1)))
                    begin
                      reg99 <= (forvar35[(2'h3):(1'h0)] != (reg48 <<< reg27));
                      reg100 <= (($unsigned((reg72 ? reg44 : forvar95)) ?
                              (+reg26) : $signed((reg82 <= reg40))) ?
                          (~&forvar64) : ($unsigned($signed(forvar64)) << (|$unsigned(reg84))));
                      reg101 <= ($signed({$signed((8'hba))}) ~^ {$signed(forvar40)});
                      reg102 <= (~&$signed(($unsigned(reg74) ?
                          $signed(forvar50) : $signed(reg35))));
                    end
                end
              else
                begin
                  reg98 <= (($unsigned(reg45) != (~forvar61[(1'h0):(1'h0)])) * forvar42[(4'ha):(4'h8)]);
                  if ((^~((~reg62) == forvar85)))
                    begin
                      reg99 <= {(~&((~|wire15) ?
                              (forvar20 ? reg87 : reg47) : (forvar90 ?
                                  reg28 : reg31)))};
                      reg100 <= reg82;
                      reg101 <= {(((reg24 < reg81) ~^ {reg43}) ?
                              reg48[(4'h8):(4'h8)] : ($signed(wire16) ?
                                  $unsigned(reg46) : (reg55 && reg21)))};
                      reg102 <= (reg79[(3'h6):(3'h6)] >= reg46[(4'hf):(3'h5)]);
                    end
                  else
                    begin
                      reg99 <= ($unsigned(($unsigned(forvar22) ?
                          (8'hba) : $unsigned((8'hb0)))) || reg59[(3'h7):(1'h1)]);
                      reg100 <= $unsigned((-forvar80[(1'h0):(1'h0)]));
                    end
                  if ((~^reg88))
                    begin
                      reg103 <= (wire15[(1'h1):(1'h0)] ?
                          reg68[(1'h1):(1'h1)] : reg21[(1'h0):(1'h0)]);
                      reg104 <= $unsigned({forvar52[(2'h3):(2'h3)]});
                      reg105 <= $unsigned($unsigned(($signed(reg91) ~^ {forvar69})));
                      reg106 <= $signed($signed((+$unsigned(reg77))));
                    end
                  else
                    begin
                      reg103 <= $signed(reg40);
                      reg104 <= ({reg71} ?
                          (|$unsigned(reg59[(2'h3):(1'h0)])) : $unsigned((-((8'ha8) ?
                              forvar22 : forvar38))));
                      reg105 <= ($signed(((reg99 <= forvar39) ?
                              {forvar27} : {reg103})) ?
                          (reg20 ?
                              {((8'hae) < forvar57)} : wire17[(3'h7):(3'h7)]) : $signed($signed((reg50 * forvar19))));
                      reg106 <= (8'hb2);
                    end
                end
              if ($signed(((reg41 * $unsigned(forvar60)) ?
                  {forvar52} : forvar53)))
                begin
                  for (forvar107 = (1'h0); (forvar107 < (2'h3)); forvar107 = (forvar107 + (1'h1)))
                    begin
                      reg108 <= $signed((($signed(forvar52) ?
                              forvar48[(3'h6):(2'h3)] : (~reg67)) ?
                          (8'haf) : ($unsigned(reg56) ?
                              (reg104 != reg40) : {(8'haa)})));
                      reg109 <= ($unsigned($signed((8'had))) - $signed(($signed(reg25) ?
                          (~reg45) : $unsigned(reg57))));
                    end
                end
              else
                begin
                  for (forvar107 = (1'h0); (forvar107 < (2'h3)); forvar107 = (forvar107 + (1'h1)))
                    begin
                      reg108 <= forvar72;
                      reg109 <= (~|((forvar28[(4'h8):(2'h3)] || $unsigned(forvar69)) ^~ (&{reg20})));
                    end
                end
            end
          else
            begin
              for (forvar95 = (1'h0); (forvar95 < (2'h2)); forvar95 = (forvar95 + (1'h1)))
                begin
                  if (forvar27[(4'ha):(1'h0)])
                    begin
                      reg96 <= forvar20[(4'h8):(3'h6)];
                      reg97 <= $signed($unsigned((^$unsigned(forvar30))));
                      reg98 <= reg31;
                      reg99 <= ($unsigned((forvar60 & reg42[(3'h5):(1'h0)])) ?
                          reg91 : $unsigned((8'h9e)));
                    end
                  else
                    begin
                      reg96 <= ((^$signed($signed(reg53))) ?
                          reg84[(3'h7):(1'h0)] : $unsigned($signed({reg58})));
                      reg97 <= {(~(reg98 ? wire17 : ((8'hb2) | reg77)))};
                    end
                  reg100 <= ($unsigned(forvar22) > reg99);
                  reg101 <= $unsigned(reg90);
                end
              for (forvar102 = (1'h0); (forvar102 < (2'h2)); forvar102 = (forvar102 + (1'h1)))
                begin
                  if (((((+reg74) > $unsigned(forvar75)) ?
                          (reg74 ?
                              (forvar63 && (8'ha2)) : $unsigned(wire13)) : reg58[(2'h2):(1'h1)]) ?
                      (&($signed(forvar69) ?
                          (reg101 ?
                              wire12 : reg46) : $unsigned((8'hb1)))) : forvar107[(3'h4):(3'h4)]))
                    begin
                      reg103 <= ((reg52[(1'h0):(1'h0)] ?
                              ({reg60} != ((8'hb3) ?
                                  (8'ha6) : (8'h9d))) : reg34[(1'h1):(1'h1)]) ?
                          forvar51 : ((!(reg33 ? wire14 : reg37)) <= forvar22));
                    end
                  else
                    begin
                      reg103 <= forvar40;
                      reg104 <= reg92;
                      reg105 <= reg100[(2'h3):(2'h2)];
                      reg106 <= reg71;
                    end
                  for (forvar107 = (1'h0); (forvar107 < (2'h2)); forvar107 = (forvar107 + (1'h1)))
                    begin
                      reg108 <= {$signed(((+forvar64) ?
                              (^reg40) : forvar27[(4'h9):(4'h9)]))};
                      reg109 <= $unsigned($unsigned(((reg90 ?
                          forvar50 : forvar19) >= wire12)));
                    end
                  if (reg45)
                    begin
                      reg110 <= ((({reg56} ? (-wire16) : {(8'ha4)}) ?
                              (reg35 ?
                                  (wire13 ?
                                      reg34 : forvar48) : (reg48 < reg80)) : ((8'h9f) >> (!(8'hb0)))) ?
                          $unsigned((8'hac)) : reg47);
                      reg111 <= $unsigned((~&$unsigned(reg86)));
                    end
                  else
                    begin
                      reg110 <= $unsigned($unsigned({{reg41}}));
                    end
                  for (forvar112 = (1'h0); (forvar112 < (2'h2)); forvar112 = (forvar112 + (1'h1)))
                    begin
                      reg113 <= forvar66[(4'h9):(4'h9)];
                      reg114 <= (~|$unsigned({(~|forvar102)}));
                    end
                end
            end
        end
      for (forvar115 = (1'h0); (forvar115 < (2'h3)); forvar115 = (forvar115 + (1'h1)))
        begin
          for (forvar116 = (1'h0); (forvar116 < (1'h1)); forvar116 = (forvar116 + (1'h1)))
            begin
              reg117 <= ((~reg34) ^ wire16[(4'h9):(3'h7)]);
              if ($signed((+($unsigned((8'ha2)) ?
                  {(8'had)} : (forvar29 + reg25)))))
                begin
                  if ({({{forvar64}} == reg35)})
                    begin
                      reg118 <= ($unsigned((8'ha2)) ?
                          {$signed(reg26[(3'h6):(3'h4)])} : $unsigned((forvar76[(2'h2):(1'h0)] ?
                              reg89[(3'h7):(2'h2)] : forvar42[(3'h4):(1'h1)])));
                    end
                  else
                    begin
                      reg118 <= (reg20 + $signed(((reg98 ? (8'hb1) : reg40) ?
                          (~|reg101) : $unsigned(reg70))));
                      reg119 <= ($unsigned($signed((^~reg39))) ?
                          $signed(reg80) : reg79);
                      reg120 <= $signed(reg63[(3'h4):(2'h2)]);
                      reg121 <= $unsigned({(^~(forvar55 ? reg49 : reg109))});
                    end
                end
              else
                begin
                  reg118 <= ($signed((^~forvar25[(3'h7):(3'h7)])) ?
                      ((!(reg88 <<< forvar116)) ?
                          (&$signed(forvar51)) : (^~(reg25 ?
                              reg89 : forvar55))) : $signed((~^(forvar29 ?
                          (8'ha1) : (8'hb9)))));
                  reg119 <= (|wire16[(4'hc):(2'h2)]);
                  if ((reg109[(3'h5):(1'h0)] ?
                      ($signed(reg77) <= (forvar81[(1'h0):(1'h0)] | {reg29})) : (|forvar71[(2'h3):(2'h2)])))
                    begin
                      reg120 <= (~^(^~forvar63));
                    end
                  else
                    begin
                      reg120 <= forvar98;
                      reg121 <= forvar25[(3'h6):(1'h1)];
                      reg122 <= (|$unsigned((reg32 ?
                          reg97 : reg89[(3'h6):(1'h0)])));
                    end
                  reg123 <= ($signed(forvar42[(4'ha):(2'h2)]) ?
                      forvar34 : wire13);
                end
              reg124 <= reg104;
            end
        end
      if ($unsigned({reg59[(4'hc):(4'ha)]}))
        begin
          for (forvar125 = (1'h0); (forvar125 < (1'h0)); forvar125 = (forvar125 + (1'h1)))
            begin
              reg126 <= (&{({wire11} | reg46)});
            end
          reg127 <= $unsigned(($unsigned(((8'ha8) - reg79)) ?
              ((8'ha6) << $signed(reg67)) : (reg21[(4'h9):(2'h3)] ?
                  ((8'ha8) * reg51) : reg39[(4'h8):(2'h2)])));
          for (forvar128 = (1'h0); (forvar128 < (1'h1)); forvar128 = (forvar128 + (1'h1)))
            begin
              for (forvar129 = (1'h0); (forvar129 < (2'h3)); forvar129 = (forvar129 + (1'h1)))
                begin
                  if ((8'hb3))
                    begin
                      reg130 <= (reg23[(1'h0):(1'h0)] ?
                          (|reg57) : (((~|wire13) - forvar53) >= (forvar76 * (reg113 == forvar115))));
                      reg131 <= (^$unsigned({(reg37 >> reg34)}));
                      reg132 <= $signed((!($unsigned(reg126) ?
                          wire16[(4'h8):(3'h4)] : ((8'hb5) ? reg49 : reg43))));
                      reg133 <= reg91;
                    end
                  else
                    begin
                      reg130 <= reg23;
                      reg131 <= (&$unsigned($signed((8'hb3))));
                    end
                  if ((reg106[(4'h9):(3'h6)] && forvar76[(2'h2):(1'h0)]))
                    begin
                      reg134 <= {reg133[(4'h8):(1'h0)]};
                    end
                  else
                    begin
                      reg134 <= ((((forvar52 >> reg46) ?
                                  (reg80 >> reg97) : $unsigned(forvar19)) ?
                              ((!reg114) * forvar29[(2'h3):(1'h1)]) : $signed(((8'hac) >> (8'hab)))) ?
                          $unsigned((8'hae)) : reg79);
                      reg135 <= reg120[(3'h7):(1'h1)];
                      reg136 <= ($unsigned((~|$signed(reg100))) ?
                          $unsigned({(|reg89)}) : (reg110[(4'h8):(4'h8)] & (8'hae)));
                      reg137 <= $signed((|$signed((~reg29))));
                    end
                  for (forvar138 = (1'h0); (forvar138 < (2'h3)); forvar138 = (forvar138 + (1'h1)))
                    begin
                      reg139 <= {{forvar55}};
                      reg140 <= (^forvar61[(1'h0):(1'h0)]);
                      reg141 <= ($signed(reg118[(1'h1):(1'h1)]) ?
                          reg127[(3'h5):(3'h5)] : (~(!(reg29 && reg63))));
                    end
                  for (forvar142 = (1'h0); (forvar142 < (2'h2)); forvar142 = (forvar142 + (1'h1)))
                    begin
                      reg143 <= ($unsigned(((8'hae) ?
                              (~&reg22) : (reg86 ? reg127 : (8'hb4)))) ?
                          (&((8'hb9) ? $unsigned(reg80) : (|wire15))) : reg71);
                      reg144 <= (-{reg90[(2'h2):(2'h2)]});
                    end
                end
              reg145 <= ((reg63[(2'h2):(1'h1)] ?
                  ((reg45 || reg43) ?
                      (reg84 > reg63) : wire12) : $signed((!(8'h9f)))) + reg86[(2'h3):(2'h2)]);
              for (forvar146 = (1'h0); (forvar146 < (2'h3)); forvar146 = (forvar146 + (1'h1)))
                begin
                  for (forvar147 = (1'h0); (forvar147 < (2'h3)); forvar147 = (forvar147 + (1'h1)))
                    begin
                      reg148 <= $unsigned($unsigned($unsigned({(8'ha5)})));
                    end
                  for (forvar149 = (1'h0); (forvar149 < (1'h0)); forvar149 = (forvar149 + (1'h1)))
                    begin
                      reg150 <= $signed(((reg94 ?
                              (reg148 | (8'ha9)) : $unsigned(reg66)) ?
                          ($signed((8'hab)) ?
                              {reg25} : (forvar85 ?
                                  reg94 : forvar149)) : $unsigned(reg76)));
                    end
                end
              for (forvar151 = (1'h0); (forvar151 < (2'h2)); forvar151 = (forvar151 + (1'h1)))
                begin
                  if (((8'hba) ?
                      ({(+forvar76)} <<< forvar115[(1'h1):(1'h1)]) : $unsigned((reg98 ?
                          reg120 : (8'ha0)))))
                    begin
                      reg152 <= $unsigned(({wire17[(2'h2):(1'h0)]} ~^ (forvar38[(4'hb):(1'h1)] ?
                          reg27 : (^reg23))));
                      reg153 <= ($unsigned($signed($unsigned((8'hba)))) ?
                          forvar72[(1'h0):(1'h0)] : forvar95[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg152 <= (((8'haf) * reg91) ?
                          $signed($signed($signed((8'had)))) : (8'hb4));
                      reg153 <= ($signed($unsigned(forvar20[(1'h1):(1'h0)])) ?
                          reg32[(1'h0):(1'h0)] : {($unsigned(reg143) ?
                                  ((8'hae) ?
                                      (8'hb7) : (8'hb5)) : forvar20[(3'h5):(3'h5)])});
                      reg154 <= $unsigned((-$unsigned(forvar142)));
                    end
                  reg155 <= {reg70};
                  if ((~&reg121))
                    begin
                      reg156 <= (wire11 ?
                          (~^((reg123 ? forvar49 : reg93) ?
                              (reg137 < reg153) : $signed(reg30))) : ((reg106[(4'ha):(4'h9)] ?
                              (reg100 ? reg72 : reg43) : (forvar49 ?
                                  reg28 : reg36)) >>> {{(8'hb4)}}));
                    end
                  else
                    begin
                      reg156 <= $unsigned(wire17[(1'h1):(1'h0)]);
                      reg157 <= (~^reg57[(3'h4):(2'h3)]);
                      reg158 <= (8'hb2);
                    end
                end
            end
          for (forvar159 = (1'h0); (forvar159 < (1'h1)); forvar159 = (forvar159 + (1'h1)))
            begin
              reg160 <= $signed({(~&(reg45 * (8'hb6)))});
              reg161 <= (~&$unsigned(({reg66} ?
                  $unsigned(forvar19) : {forvar29})));
              for (forvar162 = (1'h0); (forvar162 < (1'h0)); forvar162 = (forvar162 + (1'h1)))
                begin
                  for (forvar163 = (1'h0); (forvar163 < (2'h3)); forvar163 = (forvar163 + (1'h1)))
                    begin
                      reg164 <= (+(&$signed((reg100 ? (8'hb7) : forvar125))));
                      reg165 <= reg65[(3'h5):(2'h2)];
                    end
                  for (forvar166 = (1'h0); (forvar166 < (1'h0)); forvar166 = (forvar166 + (1'h1)))
                    begin
                      reg167 <= ({reg73} ?
                          $unsigned((forvar129[(3'h7):(1'h1)] ?
                              forvar166[(2'h2):(2'h2)] : $signed(forvar166))) : reg119[(4'h9):(3'h5)]);
                      reg168 <= (^wire11);
                      reg169 <= reg67[(4'h9):(3'h7)];
                    end
                end
            end
        end
      else
        begin
          if ($signed(forvar63[(3'h4):(2'h2)]))
            begin
              for (forvar125 = (1'h0); (forvar125 < (2'h2)); forvar125 = (forvar125 + (1'h1)))
                begin
                  if (((|reg122[(1'h1):(1'h1)]) ^ {($signed(forvar63) & (forvar142 - (8'ha1)))}))
                    begin
                      reg126 <= {{$unsigned(reg102[(1'h1):(1'h0)])}};
                    end
                  else
                    begin
                      reg126 <= $signed((forvar163 ^~ $unsigned((reg91 << reg157))));
                      reg127 <= reg74[(3'h5):(2'h3)];
                      reg128 <= ((forvar75 != $unsigned($unsigned((8'ha2)))) + $unsigned($unsigned({reg39})));
                    end
                  if ($unsigned({$unsigned((reg108 >> (8'h9d)))}))
                    begin
                      reg129 <= ((forvar69 ^~ $unsigned((reg47 ?
                          forvar72 : reg132))) * $signed(({reg111} == (reg43 >>> forvar51))));
                    end
                  else
                    begin
                      reg129 <= $signed(forvar85);
                    end
                end
              reg130 <= reg64;
            end
          else
            begin
              reg125 <= reg51[(1'h0):(1'h0)];
              if ($signed($unsigned(((forvar63 <= reg136) ?
                  $unsigned(reg51) : (wire17 ~^ forvar36)))))
                begin
                  for (forvar126 = (1'h0); (forvar126 < (2'h2)); forvar126 = (forvar126 + (1'h1)))
                    begin
                      reg127 <= (&(reg41 || $signed($signed(reg114))));
                      reg128 <= $unsigned($unsigned({{reg58}}));
                      reg129 <= {(&($signed(reg44) ~^ (^~reg84)))};
                      reg130 <= (forvar116 < ((!(reg156 && (8'hb9))) << (reg91[(4'h9):(2'h2)] ?
                          {(8'ha3)} : (|(8'ha8)))));
                    end
                  for (forvar131 = (1'h0); (forvar131 < (2'h2)); forvar131 = (forvar131 + (1'h1)))
                    begin
                      reg132 <= reg140[(1'h1):(1'h1)];
                    end
                  for (forvar133 = (1'h0); (forvar133 < (2'h3)); forvar133 = (forvar133 + (1'h1)))
                    begin
                      reg134 <= ({forvar66} && (forvar96[(3'h7):(3'h5)] ?
                          (~|(reg93 ? reg47 : reg52)) : $signed((~|forvar66))));
                      reg135 <= ($signed(($unsigned(forvar128) ^~ {(8'hb7)})) & forvar48);
                      reg136 <= {$unsigned(reg26)};
                      reg137 <= forvar95[(1'h0):(1'h0)];
                    end
                  for (forvar138 = (1'h0); (forvar138 < (1'h0)); forvar138 = (forvar138 + (1'h1)))
                    begin
                      reg139 <= $unsigned(forvar163[(3'h4):(1'h1)]);
                      reg140 <= ($signed($signed($signed(forvar151))) ?
                          $signed($unsigned($signed(reg78))) : (|(((8'hb0) * reg60) ?
                              (forvar166 ?
                                  reg169 : reg72) : (reg42 || wire13))));
                    end
                end
              else
                begin
                  if (((&(^~$signed(reg137))) - (reg42 ?
                      $signed(reg167) : reg158)))
                    begin
                      reg126 <= wire15[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg126 <= {$unsigned($signed($signed(forvar159)))};
                      reg127 <= ($signed(((reg133 ?
                          (8'haf) : forvar39) == $unsigned(forvar125))) >> $signed((~&(8'hb5))));
                    end
                  for (forvar128 = (1'h0); (forvar128 < (2'h3)); forvar128 = (forvar128 + (1'h1)))
                    begin
                      reg129 <= (!(reg57[(4'hb):(3'h6)] >>> (reg32[(1'h0):(1'h0)] ?
                          {reg55} : (reg124 == (8'ha2)))));
                    end
                  if ((reg56 ~^ $unsigned(reg71[(2'h2):(1'h1)])))
                    begin
                      reg130 <= forvar115;
                      reg131 <= {((+(reg150 ? wire17 : (8'hb5))) ?
                              reg23[(1'h0):(1'h0)] : {forvar128[(3'h6):(1'h1)]})};
                    end
                  else
                    begin
                      reg130 <= reg97[(1'h1):(1'h1)];
                      reg131 <= ((((reg125 ? forvar128 : (8'h9f)) ?
                                  $signed(reg23) : $unsigned((8'ha3))) ?
                              (reg32[(2'h2):(1'h0)] | (reg127 ~^ reg100)) : reg156) ?
                          reg119 : (~reg30));
                    end
                  for (forvar132 = (1'h0); (forvar132 < (2'h3)); forvar132 = (forvar132 + (1'h1)))
                    begin
                      reg133 <= reg128;
                      reg134 <= reg153;
                      reg135 <= $signed((((~reg93) | (8'ha5)) + reg70[(3'h5):(3'h5)]));
                    end
                end
              reg141 <= (forvar71 == $signed($unsigned(forvar112[(1'h0):(1'h0)])));
            end
        end
      if (((8'haf) ? $unsigned((8'hb8)) : (&{forvar49[(2'h3):(1'h1)]})))
        begin
          for (forvar170 = (1'h0); (forvar170 < (1'h1)); forvar170 = (forvar170 + (1'h1)))
            begin
              for (forvar171 = (1'h0); (forvar171 < (1'h0)); forvar171 = (forvar171 + (1'h1)))
                begin
                  reg172 <= forvar126;
                end
              for (forvar173 = (1'h0); (forvar173 < (2'h2)); forvar173 = (forvar173 + (1'h1)))
                begin
                  for (forvar174 = (1'h0); (forvar174 < (1'h1)); forvar174 = (forvar174 + (1'h1)))
                    begin
                      reg175 <= (^reg145[(2'h2):(2'h2)]);
                      reg176 <= {{({reg148} ? {reg84} : (^forvar18))}};
                      reg177 <= reg38[(4'hd):(3'h4)];
                      reg178 <= $signed((&$signed((-forvar60))));
                    end
                  for (forvar179 = (1'h0); (forvar179 < (1'h1)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= reg108;
                      reg181 <= $signed((reg25[(4'he):(3'h4)] || forvar50[(2'h3):(2'h3)]));
                      reg182 <= $signed($unsigned((-(~|(8'ha8)))));
                      reg183 <= {(~^$unsigned({(8'ha6)}))};
                    end
                end
              for (forvar184 = (1'h0); (forvar184 < (2'h3)); forvar184 = (forvar184 + (1'h1)))
                begin
                  reg185 <= reg73[(4'ha):(3'h4)];
                  for (forvar186 = (1'h0); (forvar186 < (2'h3)); forvar186 = (forvar186 + (1'h1)))
                    begin
                      reg187 <= reg114;
                    end
                  for (forvar188 = (1'h0); (forvar188 < (2'h2)); forvar188 = (forvar188 + (1'h1)))
                    begin
                      reg189 <= ((reg35 <<< ((reg183 ?
                              forvar96 : reg102) > reg101[(5'h10):(4'h8)])) ?
                          ((reg156 ? {reg127} : (-(8'ha7))) ?
                              {(reg81 ?
                                      reg100 : reg46)} : ((reg29 << forvar63) >> $signed((8'ha7)))) : {$signed(reg177)});
                      reg190 <= $signed(reg76);
                      reg191 <= reg82;
                    end
                end
              reg192 <= $signed(reg81);
            end
          reg193 <= $signed({($unsigned((8'hb1)) ?
                  (forvar149 ? forvar29 : reg169) : (reg47 ?
                      forvar20 : forvar96))});
        end
      else
        begin
          reg170 <= forvar81;
          for (forvar171 = (1'h0); (forvar171 < (1'h0)); forvar171 = (forvar171 + (1'h1)))
            begin
              if ((+$unsigned(reg28[(3'h6):(3'h5)])))
                begin
                  if ((|({$signed((8'ha8))} ?
                      ((reg99 != wire10) ?
                          (8'ha6) : reg65[(3'h6):(3'h4)]) : forvar163[(2'h2):(1'h1)])))
                    begin
                      reg172 <= reg27;
                      reg173 <= $unsigned($unsigned($unsigned((reg123 >= reg124))));
                      reg174 <= reg167;
                      reg175 <= reg54[(4'hb):(2'h2)];
                    end
                  else
                    begin
                      reg172 <= reg156[(3'h6):(1'h0)];
                      reg173 <= forvar112[(1'h0):(1'h0)];
                      reg174 <= (reg37 ^ (^~reg128));
                    end
                  for (forvar176 = (1'h0); (forvar176 < (1'h0)); forvar176 = (forvar176 + (1'h1)))
                    begin
                      reg177 <= $unsigned((forvar76[(1'h0):(1'h0)] ?
                          $unsigned((reg85 < reg169)) : forvar30));
                      reg178 <= ($signed((+reg124[(4'h9):(3'h7)])) ?
                          forvar64[(1'h1):(1'h1)] : forvar39);
                      reg179 <= (forvar138[(2'h3):(1'h1)] <<< reg137[(1'h1):(1'h1)]);
                      reg180 <= {forvar18};
                    end
                  if ($unsigned(forvar35[(1'h0):(1'h0)]))
                    begin
                      reg181 <= ((reg39 | (|{reg59})) < reg133[(4'h8):(2'h2)]);
                      reg182 <= ($signed((!(+forvar133))) && $signed(forvar146[(1'h1):(1'h1)]));
                      reg183 <= reg85[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg181 <= (^~reg148[(3'h6):(3'h6)]);
                    end
                  reg184 <= $unsigned(((-forvar112) ~^ forvar163));
                end
              else
                begin
                  if ((forvar29[(4'h9):(3'h5)] ?
                      forvar63[(3'h6):(1'h1)] : ((forvar48 < reg37[(3'h6):(2'h2)]) ?
                          $signed(forvar176) : reg189[(1'h0):(1'h0)])))
                    begin
                      reg172 <= forvar102[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg172 <= reg114[(2'h2):(1'h1)];
                    end
                  reg173 <= (~&($signed($signed(reg117)) <= $unsigned(forvar18)));
                  if ($unsigned($unsigned((forvar159 ?
                      reg102[(2'h2):(2'h2)] : forvar57))))
                    begin
                      reg174 <= (!{($signed(reg45) - $unsigned(forvar20))});
                      reg175 <= ($unsigned(reg184) ^ $unsigned(((~forvar176) ?
                          (reg127 ? reg92 : reg79) : reg104)));
                      reg176 <= (forvar128[(3'h5):(1'h0)] ?
                          ((-forvar90) + $signed((8'hae))) : (({(8'hb4)} ?
                              (~&forvar77) : (forvar81 ^~ forvar63)) != $unsigned(forvar49)));
                      reg177 <= $unsigned(($unsigned({reg59}) ?
                          reg169 : $unsigned((reg179 ? reg60 : reg83))));
                    end
                  else
                    begin
                      reg174 <= $signed((&(+(~|reg124))));
                    end
                end
              for (forvar185 = (1'h0); (forvar185 < (1'h0)); forvar185 = (forvar185 + (1'h1)))
                begin
                  for (forvar186 = (1'h0); (forvar186 < (2'h3)); forvar186 = (forvar186 + (1'h1)))
                    begin
                      reg187 <= $signed((-(~|(reg64 ^ reg136))));
                    end
                  for (forvar188 = (1'h0); (forvar188 < (1'h1)); forvar188 = (forvar188 + (1'h1)))
                    begin
                      reg189 <= (reg172[(2'h2):(1'h0)] ?
                          reg158 : {reg44[(3'h4):(1'h1)]});
                      reg190 <= (((~^(forvar174 && (8'hba))) ?
                              {(~reg64)} : (^reg98[(4'hc):(1'h0)])) ?
                          (reg23 ?
                              ({forvar77} ?
                                  (forvar29 ?
                                      forvar81 : forvar25) : reg136[(2'h2):(2'h2)]) : forvar149) : (-(-{reg192})));
                      reg191 <= (reg165[(1'h1):(1'h0)] ?
                          ((&$unsigned(reg20)) ~^ reg76[(1'h0):(1'h0)]) : (((~|(8'ha0)) + {reg160}) & (&reg20)));
                      reg192 <= forvar55;
                    end
                  if (reg177[(3'h7):(3'h6)])
                    begin
                      reg193 <= reg123[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg193 <= reg185[(4'h9):(3'h7)];
                      reg194 <= reg192;
                    end
                end
            end
        end
    end
  assign wire195 = ($signed($unsigned((forvar147 >= reg117))) | forvar179[(2'h2):(2'h2)]);
  assign wire196 = ((~&(8'hb9)) + ($signed($unsigned(reg91)) <<< $unsigned(reg96[(2'h2):(2'h2)])));
  assign wire197 = (!reg109);
  assign wire198 = (+(-{$unsigned(reg140)}));
  assign wire199 = ((!$signed(forvar48)) ?
                       (reg42[(3'h5):(1'h1)] ^ reg181) : reg58[(2'h3):(1'h0)]);
  assign wire200 = $unsigned($signed((reg178[(3'h5):(2'h2)] ^~ ((8'hb5) ?
                       (8'hb9) : reg140))));
  assign wire201 = $signed((reg80 || reg81[(2'h3):(1'h0)]));
  assign wire202 = $signed(forvar90);
  assign wire203 = (reg50 ?
                       {{(!reg40)}} : ($unsigned(forvar116[(5'h10):(3'h5)]) ?
                           forvar131 : ((reg144 ? forvar53 : (8'ha4)) ?
                               (8'ha5) : (~^reg90))));
  assign wire204 = ($unsigned((reg132 ? reg31[(3'h6):(3'h6)] : {forvar85})) ?
                       $unsigned((^~$signed(reg50))) : ((~&reg117) ?
                           $signed({(8'hba)}) : (+reg135[(2'h2):(1'h0)])));
  assign wire205 = $signed(reg94);
  module206 modinst619 (wire618, clk, forvar51, reg150, wire204, forvar25);
  assign wire620 = $signed({reg77[(3'h6):(3'h6)]});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module206
#( parameter param617 = ((~(((8'hac) ? (8'haf) : (8'hab)) != {(8'hb8)})) ? (((~(8'ha7)) ? (^(8'hb1)) : ((8'hb2) <<< (8'ha2))) ? (((8'ha5) | (8'hae)) >> ((8'h9f) | (8'ha1))) : ({(8'ha3)} ? {(8'haf)} : ((8'hb8) >= (8'ha6)))) : ((!((8'ha4) ? (8'hab) : (8'hac))) ? (((8'haa) <= (8'hb3)) ? ((8'ha3) ^ (8'haa)) : ((8'had) ? (8'hb1) : (8'had))) : ((~&(8'ha2)) ? ((8'hb5) ? (8'had) : (8'hac)) : (^~(8'hab))))) )
(y, clk, wire210, wire209, wire208, wire207);
  output wire [(32'h1d9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire210;
  input wire [(4'hc):(1'h0)] wire209;
  input wire [(4'he):(1'h0)] wire208;
  input wire signed [(4'h8):(1'h0)] wire207;
  wire signed [(4'hc):(1'h0)] wire616;
  wire signed [(4'he):(1'h0)] wire615;
  wire [(4'h9):(1'h0)] wire614;
  wire signed [(3'h7):(1'h0)] wire613;
  wire [(5'h10):(1'h0)] wire612;
  reg signed [(2'h2):(1'h0)] reg611 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg610 = (1'h0);
  reg [(4'h9):(1'h0)] reg580 = (1'h0);
  reg [(4'hb):(1'h0)] forvar578 = (1'h0);
  reg [(2'h2):(1'h0)] reg577 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar576 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg575 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar574 = (1'h0);
  reg [(4'h9):(1'h0)] reg572 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg609 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg608 = (1'h0);
  reg [(3'h6):(1'h0)] reg607 = (1'h0);
  reg [(3'h5):(1'h0)] reg606 = (1'h0);
  reg [(4'hc):(1'h0)] reg605 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar604 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg603 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg602 = (1'h0);
  reg [(4'hf):(1'h0)] reg601 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar600 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar599 = (1'h0);
  reg [(3'h4):(1'h0)] reg598 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar597 = (1'h0);
  reg [(4'hd):(1'h0)] reg596 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg595 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar594 = (1'h0);
  reg [(4'ha):(1'h0)] reg593 = (1'h0);
  reg [(4'hd):(1'h0)] reg592 = (1'h0);
  reg [(5'h10):(1'h0)] reg591 = (1'h0);
  reg [(4'h8):(1'h0)] reg590 = (1'h0);
  reg [(2'h2):(1'h0)] forvar589 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar588 = (1'h0);
  reg [(4'hc):(1'h0)] forvar587 = (1'h0);
  reg [(3'h6):(1'h0)] reg586 = (1'h0);
  reg [(3'h5):(1'h0)] reg585 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg584 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar583 = (1'h0);
  reg [(3'h5):(1'h0)] reg582 = (1'h0);
  reg [(4'hc):(1'h0)] reg581 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar580 = (1'h0);
  reg [(4'h8):(1'h0)] reg579 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg578 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar577 = (1'h0);
  reg [(4'hc):(1'h0)] reg576 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar575 = (1'h0);
  reg [(3'h4):(1'h0)] reg574 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar573 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar572 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire570;
  assign y = {wire616,
                 wire615,
                 wire614,
                 wire613,
                 wire612,
                 reg611,
                 reg610,
                 reg580,
                 forvar578,
                 reg577,
                 forvar576,
                 reg575,
                 forvar574,
                 reg572,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 forvar604,
                 reg603,
                 reg602,
                 reg601,
                 forvar600,
                 forvar599,
                 reg598,
                 forvar597,
                 reg596,
                 reg595,
                 forvar594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 forvar589,
                 forvar588,
                 forvar587,
                 reg586,
                 reg585,
                 reg584,
                 forvar583,
                 reg582,
                 reg581,
                 forvar580,
                 reg579,
                 reg578,
                 forvar577,
                 reg576,
                 forvar575,
                 reg574,
                 forvar573,
                 forvar572,
                 wire570,
                 (1'h0)};
  module211 modinst571 (.wire213(wire208), .clk(clk), .wire215(wire207), .wire212(wire210), .y(wire570), .wire214(wire209));
  always
    @(posedge clk) begin
      if (wire208[(4'ha):(2'h3)])
        begin
          for (forvar572 = (1'h0); (forvar572 < (2'h3)); forvar572 = (forvar572 + (1'h1)))
            begin
              for (forvar573 = (1'h0); (forvar573 < (1'h1)); forvar573 = (forvar573 + (1'h1)))
                begin
                  reg574 <= wire207;
                end
              for (forvar575 = (1'h0); (forvar575 < (2'h2)); forvar575 = (forvar575 + (1'h1)))
                begin
                  reg576 <= ({((|(8'ha4)) << wire207[(2'h3):(2'h3)])} ?
                      $unsigned(forvar575) : (~&forvar572[(1'h1):(1'h0)]));
                end
              for (forvar577 = (1'h0); (forvar577 < (1'h1)); forvar577 = (forvar577 + (1'h1)))
                begin
                  if (wire208)
                    begin
                      reg578 <= ($unsigned(wire208[(4'hd):(3'h5)]) ?
                          (8'h9f) : wire208);
                    end
                  else
                    begin
                      reg578 <= $signed((reg576 ?
                          wire570 : wire210[(4'ha):(3'h5)]));
                      reg579 <= $signed(wire208[(4'hd):(4'hc)]);
                    end
                  for (forvar580 = (1'h0); (forvar580 < (2'h2)); forvar580 = (forvar580 + (1'h1)))
                    begin
                      reg581 <= $unsigned(($signed((forvar577 && reg574)) ?
                          ($signed(wire210) >>> (8'ha1)) : $signed((8'hb5))));
                      reg582 <= forvar573[(2'h2):(1'h1)];
                    end
                  for (forvar583 = (1'h0); (forvar583 < (1'h0)); forvar583 = (forvar583 + (1'h1)))
                    begin
                      reg584 <= $unsigned((wire208[(3'h6):(1'h0)] ?
                          ((wire210 ?
                              reg576 : forvar577) >> $signed(reg576)) : reg581));
                    end
                  if (((&reg578[(3'h6):(3'h5)]) != $signed((!(~&reg578)))))
                    begin
                      reg585 <= ($signed((~{wire570})) ?
                          wire207 : $signed($signed((~^forvar577))));
                    end
                  else
                    begin
                      reg585 <= $signed((!forvar572[(1'h1):(1'h1)]));
                      reg586 <= ((((wire209 <<< forvar575) ^ $signed(forvar580)) <= ({forvar575} ?
                          $signed(reg574) : $unsigned(forvar580))) << (reg574[(1'h0):(1'h0)] ?
                          (-(wire570 ^~ (8'ha5))) : ((-reg585) ?
                              (-reg579) : $signed((8'hac)))));
                    end
                end
            end
          for (forvar587 = (1'h0); (forvar587 < (2'h2)); forvar587 = (forvar587 + (1'h1)))
            begin
              for (forvar588 = (1'h0); (forvar588 < (2'h3)); forvar588 = (forvar588 + (1'h1)))
                begin
                  for (forvar589 = (1'h0); (forvar589 < (1'h1)); forvar589 = (forvar589 + (1'h1)))
                    begin
                      reg590 <= $unsigned(((~&(forvar588 ?
                              forvar588 : reg582)) ?
                          reg576 : {(reg582 ? reg586 : wire570)}));
                      reg591 <= {{(~reg578[(4'h8):(3'h7)])}};
                      reg592 <= reg586;
                      reg593 <= $unsigned((($unsigned(reg582) ?
                              $unsigned(reg574) : {wire208}) ?
                          reg581 : ($signed(forvar580) ?
                              forvar580[(4'hf):(2'h3)] : forvar587)));
                    end
                  for (forvar594 = (1'h0); (forvar594 < (2'h3)); forvar594 = (forvar594 + (1'h1)))
                    begin
                      reg595 <= ((~^{(|wire210)}) ?
                          forvar587[(1'h0):(1'h0)] : (~|$unsigned((reg582 ?
                              (8'hb8) : forvar594))));
                      reg596 <= (8'h9f);
                    end
                  for (forvar597 = (1'h0); (forvar597 < (2'h2)); forvar597 = (forvar597 + (1'h1)))
                    begin
                      reg598 <= reg581;
                    end
                end
              for (forvar599 = (1'h0); (forvar599 < (1'h0)); forvar599 = (forvar599 + (1'h1)))
                begin
                  for (forvar600 = (1'h0); (forvar600 < (1'h1)); forvar600 = (forvar600 + (1'h1)))
                    begin
                      reg601 <= (($signed(wire207) ?
                              reg592[(4'h8):(2'h3)] : (^$signed((8'h9d)))) ?
                          reg579[(3'h7):(3'h4)] : $signed((8'hba)));
                      reg602 <= (((^~(forvar572 ~^ forvar573)) ?
                              (+{forvar587}) : forvar572[(1'h0):(1'h0)]) ?
                          $unsigned((forvar589 ?
                              {forvar600} : forvar575[(1'h1):(1'h0)])) : (reg590[(2'h3):(2'h2)] ?
                              (|(^(8'haa))) : reg598));
                    end
                  reg603 <= ($signed(reg579[(3'h4):(2'h3)]) | forvar589[(1'h1):(1'h1)]);
                  for (forvar604 = (1'h0); (forvar604 < (1'h1)); forvar604 = (forvar604 + (1'h1)))
                    begin
                      reg605 <= ($unsigned((|reg598)) - ((forvar573[(4'hb):(4'hb)] <= $signed(reg585)) ?
                          forvar587 : $unsigned($signed(forvar587))));
                      reg606 <= $unsigned(wire209);
                      reg607 <= reg593;
                      reg608 <= (8'had);
                    end
                  reg609 <= forvar573[(2'h3):(2'h3)];
                end
            end
        end
      else
        begin
          reg572 <= {{($signed(reg574) & $signed((8'hb3)))}};
          for (forvar573 = (1'h0); (forvar573 < (2'h3)); forvar573 = (forvar573 + (1'h1)))
            begin
              for (forvar574 = (1'h0); (forvar574 < (2'h2)); forvar574 = (forvar574 + (1'h1)))
                begin
                  reg575 <= reg593[(1'h1):(1'h0)];
                  for (forvar576 = (1'h0); (forvar576 < (2'h2)); forvar576 = (forvar576 + (1'h1)))
                    begin
                      reg577 <= (((&(forvar572 ? reg609 : reg606)) + ((reg572 ?
                              (8'hb7) : wire210) ?
                          reg593[(2'h3):(2'h3)] : $signed(reg598))) << $unsigned($unsigned((reg605 && reg602))));
                    end
                  for (forvar578 = (1'h0); (forvar578 < (1'h0)); forvar578 = (forvar578 + (1'h1)))
                    begin
                      reg579 <= $signed((($signed(reg574) < {reg603}) * forvar588[(1'h0):(1'h0)]));
                      reg580 <= $unsigned(($signed($signed(reg591)) ?
                          $signed((-(8'ha6))) : $unsigned((reg606 ?
                              (8'hb8) : reg601))));
                      reg581 <= reg598;
                      reg582 <= (8'had);
                    end
                  for (forvar583 = (1'h0); (forvar583 < (1'h1)); forvar583 = (forvar583 + (1'h1)))
                    begin
                      reg584 <= (({$unsigned((8'ha1))} ?
                              $signed((^~reg608)) : forvar574) ?
                          {reg591} : reg575[(4'hc):(4'hc)]);
                      reg585 <= $signed(((forvar604[(3'h6):(3'h6)] | forvar573) ?
                          reg582[(1'h1):(1'h0)] : reg593[(4'h8):(1'h1)]));
                    end
                end
            end
          reg586 <= reg592[(3'h7):(3'h5)];
        end
      reg610 <= reg592[(1'h1):(1'h0)];
      reg611 <= $signed({wire210});
    end
  assign wire612 = $unsigned($unsigned($unsigned(wire570)));
  assign wire613 = (8'h9f);
  assign wire614 = wire570;
  assign wire615 = (((~^(reg601 >> (8'hb8))) ?
                           {{reg579}} : ($unsigned(forvar589) ?
                               (reg610 ? reg582 : (8'hae)) : (~&forvar600))) ?
                       reg608[(1'h1):(1'h1)] : wire208);
  assign wire616 = (reg601 + (forvar577 ?
                       (-$signed(forvar600)) : $unsigned((8'ha3))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module211
#( parameter param569 = ((~&(((8'haa) ? (8'haa) : (8'hba)) >> (|(8'haf)))) >> (^(((8'hb5) ^~ (8'hae)) ? ((8'hab) ? (8'hb9) : (8'h9d)) : (~|(8'hb4))))) )
(y, clk, wire215, wire214, wire213, wire212);
  output wire [(32'hef4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire215;
  input wire [(4'hc):(1'h0)] wire214;
  input wire signed [(4'ha):(1'h0)] wire213;
  input wire [(4'hc):(1'h0)] wire212;
  wire signed [(3'h4):(1'h0)] wire568;
  wire [(4'h8):(1'h0)] wire567;
  wire signed [(3'h6):(1'h0)] wire566;
  wire [(4'hd):(1'h0)] wire565;
  wire signed [(3'h7):(1'h0)] wire564;
  reg signed [(2'h3):(1'h0)] forvar556 = (1'h0);
  reg [(4'hf):(1'h0)] forvar554 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg563 = (1'h0);
  reg [(5'h10):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar561 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg560 = (1'h0);
  reg [(3'h5):(1'h0)] reg559 = (1'h0);
  reg [(2'h2):(1'h0)] reg558 = (1'h0);
  reg [(3'h7):(1'h0)] reg557 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg556 = (1'h0);
  reg [(4'he):(1'h0)] reg555 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg554 = (1'h0);
  reg [(4'h8):(1'h0)] reg553 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg552 = (1'h0);
  reg [(4'hd):(1'h0)] forvar551 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar550 = (1'h0);
  reg [(4'hc):(1'h0)] forvar549 = (1'h0);
  reg [(3'h6):(1'h0)] reg548 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg547 = (1'h0);
  reg [(4'h8):(1'h0)] forvar546 = (1'h0);
  reg [(3'h5):(1'h0)] reg545 = (1'h0);
  reg [(5'h10):(1'h0)] reg544 = (1'h0);
  reg [(4'hb):(1'h0)] reg543 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar542 = (1'h0);
  reg [(3'h7):(1'h0)] reg541 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg540 = (1'h0);
  reg [(4'h9):(1'h0)] reg539 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar538 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg537 = (1'h0);
  reg [(2'h3):(1'h0)] reg536 = (1'h0);
  reg [(4'ha):(1'h0)] forvar535 = (1'h0);
  reg [(4'he):(1'h0)] reg529 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar527 = (1'h0);
  reg [(2'h2):(1'h0)] forvar525 = (1'h0);
  reg [(3'h4):(1'h0)] reg524 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar521 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg535 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg534 = (1'h0);
  reg [(3'h7):(1'h0)] reg533 = (1'h0);
  reg [(4'h9):(1'h0)] reg532 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar531 = (1'h0);
  reg [(5'h10):(1'h0)] reg530 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar529 = (1'h0);
  reg [(5'h10):(1'h0)] reg528 = (1'h0);
  reg [(2'h2):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg526 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg525 = (1'h0);
  reg [(3'h4):(1'h0)] forvar524 = (1'h0);
  reg [(3'h6):(1'h0)] reg523 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg522 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg521 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg520 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg519 = (1'h0);
  reg [(3'h4):(1'h0)] reg518 = (1'h0);
  reg [(5'h10):(1'h0)] reg514 = (1'h0);
  reg [(2'h2):(1'h0)] reg510 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar509 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar506 = (1'h0);
  reg [(4'hf):(1'h0)] reg517 = (1'h0);
  reg [(3'h5):(1'h0)] reg516 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg515 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar514 = (1'h0);
  reg [(3'h7):(1'h0)] reg513 = (1'h0);
  reg [(4'he):(1'h0)] reg512 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg511 = (1'h0);
  reg [(4'hb):(1'h0)] forvar510 = (1'h0);
  reg [(3'h4):(1'h0)] reg509 = (1'h0);
  reg [(4'hb):(1'h0)] reg508 = (1'h0);
  reg [(2'h3):(1'h0)] reg507 = (1'h0);
  reg [(3'h5):(1'h0)] reg506 = (1'h0);
  reg [(4'hc):(1'h0)] reg505 = (1'h0);
  reg [(4'ha):(1'h0)] reg504 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar503 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg502 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg501 = (1'h0);
  reg [(5'h10):(1'h0)] forvar500 = (1'h0);
  reg [(5'h10):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg498 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg497 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg496 = (1'h0);
  reg [(4'hf):(1'h0)] reg495 = (1'h0);
  reg [(3'h4):(1'h0)] forvar494 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg494 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar493 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg484 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar483 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar477 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar475 = (1'h0);
  reg [(4'hb):(1'h0)] forvar473 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar471 = (1'h0);
  reg [(4'hf):(1'h0)] reg492 = (1'h0);
  reg [(3'h5):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar486 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg490 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg489 = (1'h0);
  reg [(2'h3):(1'h0)] reg488 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg487 = (1'h0);
  reg [(4'h9):(1'h0)] reg486 = (1'h0);
  reg [(4'ha):(1'h0)] reg485 = (1'h0);
  reg [(4'ha):(1'h0)] forvar484 = (1'h0);
  reg [(3'h5):(1'h0)] reg483 = (1'h0);
  reg [(3'h4):(1'h0)] reg482 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg481 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg480 = (1'h0);
  reg [(4'hb):(1'h0)] reg479 = (1'h0);
  reg [(3'h4):(1'h0)] reg478 = (1'h0);
  reg [(2'h3):(1'h0)] reg477 = (1'h0);
  reg [(3'h6):(1'h0)] reg476 = (1'h0);
  reg [(3'h5):(1'h0)] reg475 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg474 = (1'h0);
  reg [(4'h9):(1'h0)] reg473 = (1'h0);
  reg [(4'ha):(1'h0)] reg472 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg471 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar470 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg469 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg468 = (1'h0);
  reg [(4'ha):(1'h0)] reg467 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg466 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg465 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg464 = (1'h0);
  reg signed [(4'he):(1'h0)] reg463 = (1'h0);
  reg [(4'hd):(1'h0)] forvar462 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg461 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg460 = (1'h0);
  reg [(4'he):(1'h0)] reg459 = (1'h0);
  reg [(4'he):(1'h0)] reg458 = (1'h0);
  reg [(2'h3):(1'h0)] forvar457 = (1'h0);
  reg [(2'h2):(1'h0)] reg457 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg456 = (1'h0);
  reg [(4'h9):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg454 = (1'h0);
  reg [(2'h2):(1'h0)] forvar453 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar451 = (1'h0);
  reg [(3'h6):(1'h0)] reg450 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg449 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg448 = (1'h0);
  reg [(4'hd):(1'h0)] reg447 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg446 = (1'h0);
  reg [(2'h3):(1'h0)] forvar445 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg444 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar443 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg442 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg441 = (1'h0);
  reg [(4'he):(1'h0)] forvar420 = (1'h0);
  reg [(2'h3):(1'h0)] forvar425 = (1'h0);
  reg [(2'h2):(1'h0)] reg440 = (1'h0);
  reg signed [(4'he):(1'h0)] reg439 = (1'h0);
  reg [(4'hf):(1'h0)] reg438 = (1'h0);
  reg [(4'hc):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar436 = (1'h0);
  reg [(3'h6):(1'h0)] forvar435 = (1'h0);
  reg [(3'h7):(1'h0)] reg434 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg433 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar430 = (1'h0);
  reg [(4'hc):(1'h0)] reg428 = (1'h0);
  reg [(4'hb):(1'h0)] forvar423 = (1'h0);
  reg [(2'h3):(1'h0)] reg432 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg430 = (1'h0);
  reg [(4'hd):(1'h0)] reg429 = (1'h0);
  reg [(4'he):(1'h0)] forvar428 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg427 = (1'h0);
  reg [(3'h7):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg425 = (1'h0);
  reg [(4'h8):(1'h0)] reg424 = (1'h0);
  reg [(3'h6):(1'h0)] reg423 = (1'h0);
  reg signed [(4'he):(1'h0)] reg422 = (1'h0);
  reg [(4'h8):(1'h0)] reg421 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg420 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg419 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg418 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg417 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg416 = (1'h0);
  reg [(4'hb):(1'h0)] reg415 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg414 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg413 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg412 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg411 = (1'h0);
  reg [(3'h5):(1'h0)] forvar410 = (1'h0);
  reg [(3'h7):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg408 = (1'h0);
  reg [(2'h3):(1'h0)] forvar407 = (1'h0);
  reg [(3'h5):(1'h0)] reg406 = (1'h0);
  reg [(3'h7):(1'h0)] forvar405 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg404 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar403 = (1'h0);
  reg [(2'h3):(1'h0)] reg402 = (1'h0);
  reg [(4'h9):(1'h0)] reg401 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg400 = (1'h0);
  reg [(5'h10):(1'h0)] forvar399 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg398 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg397 = (1'h0);
  reg [(3'h5):(1'h0)] reg396 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg395 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg389 = (1'h0);
  reg [(2'h3):(1'h0)] forvar388 = (1'h0);
  reg [(4'hb):(1'h0)] forvar387 = (1'h0);
  reg [(4'he):(1'h0)] forvar379 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg376 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg394 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg393 = (1'h0);
  reg [(4'hc):(1'h0)] reg392 = (1'h0);
  reg [(4'h8):(1'h0)] forvar391 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg390 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar389 = (1'h0);
  reg [(3'h5):(1'h0)] reg388 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar386 = (1'h0);
  reg [(4'he):(1'h0)] reg383 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar382 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg387 = (1'h0);
  reg [(3'h5):(1'h0)] reg386 = (1'h0);
  reg [(5'h10):(1'h0)] reg385 = (1'h0);
  reg [(4'ha):(1'h0)] reg384 = (1'h0);
  reg [(3'h7):(1'h0)] forvar383 = (1'h0);
  reg [(4'he):(1'h0)] reg382 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg381 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg380 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg379 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg378 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg377 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar376 = (1'h0);
  reg [(4'hb):(1'h0)] forvar375 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg374 = (1'h0);
  reg [(3'h7):(1'h0)] reg373 = (1'h0);
  reg [(5'h10):(1'h0)] reg372 = (1'h0);
  reg [(4'hf):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg370 = (1'h0);
  reg [(4'hb):(1'h0)] reg369 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar368 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg366 = (1'h0);
  reg [(4'ha):(1'h0)] forvar365 = (1'h0);
  reg [(4'ha):(1'h0)] forvar360 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg358 = (1'h0);
  reg [(4'hc):(1'h0)] reg355 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar351 = (1'h0);
  reg [(3'h7):(1'h0)] forvar346 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar345 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar344 = (1'h0);
  reg [(4'h8):(1'h0)] reg341 = (1'h0);
  reg [(5'h10):(1'h0)] forvar340 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg365 = (1'h0);
  reg [(4'ha):(1'h0)] reg364 = (1'h0);
  reg [(5'h10):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg362 = (1'h0);
  reg [(4'hb):(1'h0)] reg361 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg360 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar358 = (1'h0);
  reg signed [(4'he):(1'h0)] reg357 = (1'h0);
  reg [(4'hd):(1'h0)] reg356 = (1'h0);
  reg [(4'hf):(1'h0)] forvar355 = (1'h0);
  reg [(3'h6):(1'h0)] forvar354 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg350 = (1'h0);
  reg [(4'hf):(1'h0)] forvar348 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg347 = (1'h0);
  reg [(4'ha):(1'h0)] reg342 = (1'h0);
  reg [(4'h8):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg352 = (1'h0);
  reg [(2'h2):(1'h0)] reg351 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar350 = (1'h0);
  reg signed [(4'he):(1'h0)] reg349 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg348 = (1'h0);
  reg [(3'h6):(1'h0)] forvar347 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg346 = (1'h0);
  reg [(3'h5):(1'h0)] reg345 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg344 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg343 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar342 = (1'h0);
  reg [(3'h5):(1'h0)] forvar341 = (1'h0);
  reg [(4'hf):(1'h0)] reg340 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg339 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg338 = (1'h0);
  reg [(2'h2):(1'h0)] reg333 = (1'h0);
  reg [(4'hd):(1'h0)] forvar330 = (1'h0);
  reg [(4'hd):(1'h0)] forvar329 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar325 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg323 = (1'h0);
  reg [(3'h6):(1'h0)] forvar320 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg337 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg336 = (1'h0);
  reg [(4'hc):(1'h0)] reg335 = (1'h0);
  reg [(4'h8):(1'h0)] reg334 = (1'h0);
  reg [(4'he):(1'h0)] forvar333 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg332 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg331 = (1'h0);
  reg [(4'he):(1'h0)] reg330 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg329 = (1'h0);
  reg [(4'ha):(1'h0)] reg328 = (1'h0);
  reg [(4'hc):(1'h0)] reg327 = (1'h0);
  reg [(4'h9):(1'h0)] reg326 = (1'h0);
  reg [(4'hd):(1'h0)] reg325 = (1'h0);
  reg [(4'h8):(1'h0)] reg324 = (1'h0);
  reg [(4'he):(1'h0)] forvar323 = (1'h0);
  reg [(4'hd):(1'h0)] reg322 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg321 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg320 = (1'h0);
  reg [(4'h8):(1'h0)] reg319 = (1'h0);
  reg [(5'h10):(1'h0)] forvar318 = (1'h0);
  reg [(3'h5):(1'h0)] reg317 = (1'h0);
  wire [(4'hd):(1'h0)] wire316;
  wire [(3'h5):(1'h0)] wire315;
  wire signed [(4'h8):(1'h0)] wire314;
  reg [(3'h4):(1'h0)] reg285 = (1'h0);
  reg [(4'hc):(1'h0)] forvar283 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg279 = (1'h0);
  reg [(2'h2):(1'h0)] reg278 = (1'h0);
  reg [(4'hb):(1'h0)] forvar277 = (1'h0);
  reg [(4'he):(1'h0)] forvar272 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg274 = (1'h0);
  reg signed [(4'he):(1'h0)] reg273 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar264 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar261 = (1'h0);
  reg [(4'hb):(1'h0)] forvar260 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg258 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg313 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg312 = (1'h0);
  reg [(5'h10):(1'h0)] reg311 = (1'h0);
  reg [(4'h8):(1'h0)] forvar310 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg309 = (1'h0);
  reg [(2'h3):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar306 = (1'h0);
  reg [(3'h6):(1'h0)] reg305 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg304 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg303 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar302 = (1'h0);
  reg [(4'hb):(1'h0)] forvar301 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg297 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg300 = (1'h0);
  reg signed [(4'he):(1'h0)] reg299 = (1'h0);
  reg [(2'h2):(1'h0)] reg298 = (1'h0);
  reg [(2'h2):(1'h0)] forvar297 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar296 = (1'h0);
  reg [(4'h8):(1'h0)] reg276 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg295 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg293 = (1'h0);
  reg [(4'h8):(1'h0)] reg292 = (1'h0);
  reg [(4'h9):(1'h0)] forvar291 = (1'h0);
  reg [(3'h7):(1'h0)] reg290 = (1'h0);
  reg signed [(4'he):(1'h0)] reg289 = (1'h0);
  reg [(3'h5):(1'h0)] forvar288 = (1'h0);
  reg [(2'h2):(1'h0)] reg287 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg286 = (1'h0);
  reg [(4'hf):(1'h0)] forvar285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg284 = (1'h0);
  reg [(4'h9):(1'h0)] reg283 = (1'h0);
  reg [(3'h6):(1'h0)] reg282 = (1'h0);
  reg [(4'ha):(1'h0)] reg281 = (1'h0);
  reg signed [(4'he):(1'h0)] reg280 = (1'h0);
  reg [(4'h9):(1'h0)] forvar279 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg277 = (1'h0);
  reg [(3'h4):(1'h0)] forvar276 = (1'h0);
  reg [(4'hb):(1'h0)] reg259 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar274 = (1'h0);
  reg [(3'h4):(1'h0)] forvar273 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg272 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg271 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar270 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg269 = (1'h0);
  reg [(4'he):(1'h0)] reg268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg267 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg266 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar265 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg264 = (1'h0);
  reg [(4'ha):(1'h0)] reg263 = (1'h0);
  reg [(3'h5):(1'h0)] reg262 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg261 = (1'h0);
  reg [(4'h8):(1'h0)] reg260 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar259 = (1'h0);
  reg [(4'ha):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg238 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg257 = (1'h0);
  reg [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(4'h9):(1'h0)] forvar255 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar254 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg253 = (1'h0);
  reg [(4'h8):(1'h0)] forvar252 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg251 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg250 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar249 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar240 = (1'h0);
  reg [(4'hd):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg247 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg246 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg245 = (1'h0);
  reg [(5'h10):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg243 = (1'h0);
  reg [(4'hf):(1'h0)] reg242 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg241 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg240 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg239 = (1'h0);
  reg [(4'h9):(1'h0)] forvar238 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar237 = (1'h0);
  reg [(4'hf):(1'h0)] reg236 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg235 = (1'h0);
  reg [(2'h3):(1'h0)] reg234 = (1'h0);
  reg [(4'hf):(1'h0)] reg233 = (1'h0);
  reg [(3'h5):(1'h0)] reg232 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg231 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg229 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar228 = (1'h0);
  reg [(4'hd):(1'h0)] reg227 = (1'h0);
  reg [(3'h4):(1'h0)] reg226 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg225 = (1'h0);
  reg [(3'h7):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar222 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg221 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar220 = (1'h0);
  reg [(4'h9):(1'h0)] forvar219 = (1'h0);
  reg [(3'h4):(1'h0)] reg218 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire217;
  wire signed [(3'h5):(1'h0)] wire216;
  assign y = {wire568,
                 wire567,
                 wire566,
                 wire565,
                 wire564,
                 forvar556,
                 forvar554,
                 reg563,
                 reg562,
                 forvar561,
                 reg560,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 forvar551,
                 forvar550,
                 forvar549,
                 reg548,
                 reg547,
                 forvar546,
                 reg545,
                 reg544,
                 reg543,
                 forvar542,
                 reg541,
                 reg540,
                 reg539,
                 forvar538,
                 reg537,
                 reg536,
                 forvar535,
                 reg529,
                 forvar527,
                 forvar525,
                 reg524,
                 forvar521,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 forvar531,
                 reg530,
                 forvar529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 forvar524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg514,
                 reg510,
                 forvar509,
                 forvar506,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 reg513,
                 reg512,
                 reg511,
                 forvar510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 reg505,
                 reg504,
                 forvar503,
                 reg502,
                 reg501,
                 forvar500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 forvar494,
                 reg494,
                 forvar493,
                 reg484,
                 forvar483,
                 forvar477,
                 forvar475,
                 forvar473,
                 forvar471,
                 reg492,
                 reg491,
                 forvar486,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 forvar484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 forvar470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 forvar462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 forvar457,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 forvar453,
                 reg452,
                 forvar451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 forvar445,
                 reg444,
                 forvar443,
                 reg442,
                 reg441,
                 forvar420,
                 forvar425,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 forvar436,
                 forvar435,
                 reg434,
                 reg433,
                 forvar430,
                 reg428,
                 forvar423,
                 reg432,
                 reg431,
                 reg430,
                 reg429,
                 forvar428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg414,
                 reg413,
                 reg412,
                 reg411,
                 forvar410,
                 reg409,
                 reg408,
                 forvar407,
                 reg406,
                 forvar405,
                 reg404,
                 forvar403,
                 reg402,
                 reg401,
                 reg400,
                 forvar399,
                 reg398,
                 reg397,
                 reg396,
                 reg395,
                 reg389,
                 forvar388,
                 forvar387,
                 forvar379,
                 reg376,
                 reg394,
                 reg393,
                 reg392,
                 forvar391,
                 reg390,
                 forvar389,
                 reg388,
                 forvar386,
                 reg383,
                 forvar382,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 forvar383,
                 reg382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 forvar376,
                 forvar375,
                 reg368,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg369,
                 forvar368,
                 reg367,
                 reg366,
                 forvar365,
                 forvar360,
                 reg358,
                 reg355,
                 reg354,
                 forvar351,
                 forvar346,
                 forvar345,
                 forvar344,
                 reg341,
                 forvar340,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 forvar358,
                 reg357,
                 reg356,
                 forvar355,
                 forvar354,
                 reg350,
                 forvar348,
                 reg347,
                 reg342,
                 reg353,
                 reg352,
                 reg351,
                 forvar350,
                 reg349,
                 reg348,
                 forvar347,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 forvar342,
                 forvar341,
                 reg340,
                 reg339,
                 reg338,
                 reg333,
                 forvar330,
                 forvar329,
                 forvar325,
                 reg323,
                 forvar320,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 forvar333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 forvar323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 forvar318,
                 reg317,
                 wire316,
                 wire315,
                 wire314,
                 reg285,
                 forvar283,
                 reg279,
                 reg278,
                 forvar277,
                 forvar272,
                 reg274,
                 reg273,
                 reg270,
                 reg265,
                 forvar264,
                 forvar261,
                 forvar260,
                 reg258,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 reg309,
                 reg308,
                 reg307,
                 forvar306,
                 reg305,
                 reg304,
                 reg303,
                 forvar302,
                 forvar301,
                 reg297,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 forvar296,
                 reg276,
                 reg295,
                 reg294,
                 reg293,
                 reg292,
                 forvar291,
                 reg290,
                 reg289,
                 forvar288,
                 reg287,
                 reg286,
                 forvar285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 forvar279,
                 forvar278,
                 reg277,
                 forvar276,
                 reg259,
                 reg275,
                 forvar274,
                 forvar273,
                 reg272,
                 reg271,
                 forvar270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 forvar265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 forvar259,
                 forvar258,
                 reg238,
                 reg257,
                 reg256,
                 forvar255,
                 forvar254,
                 reg253,
                 forvar252,
                 reg251,
                 reg250,
                 forvar249,
                 forvar240,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 forvar238,
                 forvar237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 forvar228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 forvar222,
                 reg221,
                 forvar220,
                 forvar219,
                 reg218,
                 wire217,
                 wire216,
                 (1'h0)};
  assign wire216 = {$unsigned(($signed(wire212) ?
                           wire214[(4'ha):(3'h5)] : {wire212}))};
  assign wire217 = {$unsigned(wire213)};
  always
    @(posedge clk) begin
      reg218 <= ((wire213[(3'h5):(2'h3)] ?
              $signed($signed(wire217)) : ($signed(wire214) ?
                  (wire217 ? wire212 : wire213) : wire215[(1'h0):(1'h0)])) ?
          (((wire216 ? wire212 : wire215) ?
                  $unsigned((8'hb9)) : wire213[(2'h2):(1'h0)]) ?
              (8'hb1) : ((wire216 <<< wire213) > (wire216 != wire214))) : ((wire216[(1'h0):(1'h0)] & wire213) == (wire212[(4'ha):(3'h5)] ?
              wire212[(1'h1):(1'h1)] : wire212)));
      for (forvar219 = (1'h0); (forvar219 < (2'h3)); forvar219 = (forvar219 + (1'h1)))
        begin
          for (forvar220 = (1'h0); (forvar220 < (2'h2)); forvar220 = (forvar220 + (1'h1)))
            begin
              if ($unsigned(forvar219[(1'h0):(1'h0)]))
                begin
                  reg221 <= $unsigned($signed($unsigned((-(8'h9e)))));
                  for (forvar222 = (1'h0); (forvar222 < (2'h2)); forvar222 = (forvar222 + (1'h1)))
                    begin
                      reg223 <= $unsigned($signed((~(wire215 << wire215))));
                    end
                  if (forvar220)
                    begin
                      reg224 <= (^forvar220);
                    end
                  else
                    begin
                      reg224 <= ($unsigned(reg224[(3'h5):(3'h5)]) == (~forvar220[(3'h4):(1'h0)]));
                      reg225 <= wire215;
                      reg226 <= $unsigned((8'hb2));
                      reg227 <= ($unsigned($unsigned($signed(reg225))) ?
                          forvar219 : {({reg226} ? (~^wire217) : wire216)});
                    end
                  for (forvar228 = (1'h0); (forvar228 < (1'h0)); forvar228 = (forvar228 + (1'h1)))
                    begin
                      reg229 <= {((8'hab) ?
                              $signed(wire217) : ($unsigned((8'hb7)) ?
                                  $signed(reg225) : forvar222))};
                      reg230 <= ((wire213 + ((~&reg225) ?
                              (reg225 ? reg229 : forvar222) : (&(8'hab)))) ?
                          reg223 : reg227);
                      reg231 <= (wire216 ? wire213[(4'h8):(1'h0)] : reg225);
                      reg232 <= reg229[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  reg221 <= (^~wire217);
                end
              reg233 <= wire214;
              reg234 <= forvar222[(1'h0):(1'h0)];
            end
          reg235 <= ($unsigned((^~$signed(reg230))) ?
              $unsigned(($signed(reg224) == (^reg232))) : (|$unsigned(forvar220)));
          reg236 <= (wire216[(3'h5):(1'h1)] != $unsigned(forvar228));
        end
      for (forvar237 = (1'h0); (forvar237 < (1'h1)); forvar237 = (forvar237 + (1'h1)))
        begin
          if ($signed((8'ha4)))
            begin
              if (((^~(&(reg223 <<< (8'ha3)))) || {($signed((8'ha9)) ?
                      $unsigned(reg218) : wire216[(1'h1):(1'h0)])}))
                begin
                  for (forvar238 = (1'h0); (forvar238 < (1'h0)); forvar238 = (forvar238 + (1'h1)))
                    begin
                      reg239 <= $unsigned($unsigned((^~reg229[(2'h2):(1'h0)])));
                      reg240 <= ((wire216 ?
                          (-$unsigned(reg239)) : $signed(wire215)) + forvar238[(2'h2):(1'h1)]);
                      reg241 <= (~reg226);
                    end
                  if ($unsigned($unsigned(reg226)))
                    begin
                      reg242 <= (((8'hb9) ?
                          wire215 : {(reg235 ?
                                  forvar220 : (8'hab))}) | wire213[(3'h6):(3'h4)]);
                      reg243 <= (forvar222[(1'h0):(1'h0)] ?
                          $signed((reg235[(1'h1):(1'h0)] ?
                              (&reg241) : (reg241 ?
                                  wire214 : (8'hb6)))) : {(8'h9d)});
                      reg244 <= reg240[(4'hc):(4'hc)];
                      reg245 <= wire215;
                    end
                  else
                    begin
                      reg242 <= (((reg243 ?
                                  (-forvar228) : $unsigned(forvar228)) ?
                              (|(reg232 ?
                                  (8'hb6) : forvar219)) : reg233[(3'h4):(1'h1)]) ?
                          $signed((^~$unsigned(forvar237))) : $unsigned($signed(wire214[(4'ha):(1'h0)])));
                    end
                  if ($unsigned($signed(reg245)))
                    begin
                      reg246 <= ((~reg233) > (~&((reg234 * reg236) ?
                          $unsigned(wire212) : reg227[(4'h9):(2'h3)])));
                      reg247 <= reg234;
                    end
                  else
                    begin
                      reg246 <= (reg233 ?
                          $signed(reg225[(1'h0):(1'h0)]) : (^reg224));
                      reg247 <= $signed($signed($signed((reg239 + reg236))));
                      reg248 <= reg232;
                    end
                end
              else
                begin
                  for (forvar238 = (1'h0); (forvar238 < (1'h1)); forvar238 = (forvar238 + (1'h1)))
                    begin
                      reg239 <= $unsigned((reg245[(1'h0):(1'h0)] == (^((8'ha8) || reg244))));
                    end
                  for (forvar240 = (1'h0); (forvar240 < (1'h0)); forvar240 = (forvar240 + (1'h1)))
                    begin
                      reg241 <= ((($unsigned(reg242) || ((8'ha4) ?
                          (8'ha7) : reg247)) + $signed(reg242[(4'ha):(4'ha)])) << forvar228);
                      reg242 <= (reg229[(4'hb):(1'h0)] ?
                          ($signed($signed((8'hb5))) >= $unsigned((wire213 < reg227))) : ((^forvar228[(1'h1):(1'h0)]) ?
                              ($signed(reg242) ?
                                  ((8'hba) ?
                                      reg218 : forvar222) : {forvar237}) : (~((8'ha3) != forvar237))));
                      reg243 <= $signed((reg225[(3'h6):(3'h4)] == {$unsigned(forvar228)}));
                      reg244 <= (^(forvar237[(1'h1):(1'h1)] ?
                          ($signed(wire215) - $signed(reg241)) : $signed(reg235[(2'h2):(2'h2)])));
                    end
                  if (($signed((&forvar238)) <<< (|$unsigned($signed(wire216)))))
                    begin
                      reg245 <= (reg227[(2'h2):(1'h0)] ~^ ($unsigned((reg226 ?
                              (8'ha8) : reg218)) ?
                          (|$signed(forvar222)) : (~|(^~wire217))));
                      reg246 <= $signed($signed({(reg218 ^ reg247)}));
                      reg247 <= $unsigned((-(&forvar240)));
                    end
                  else
                    begin
                      reg245 <= ($signed(reg233[(4'h8):(3'h4)]) ?
                          reg242 : ({forvar238[(4'h8):(1'h0)]} ?
                              (-(wire214 ?
                                  reg223 : wire215)) : $unsigned(forvar238)));
                      reg246 <= (($signed({(8'ha3)}) < (forvar238 ?
                          (8'hab) : wire212[(4'hc):(3'h7)])) << reg223);
                      reg247 <= wire214[(3'h7):(3'h7)];
                    end
                end
              for (forvar249 = (1'h0); (forvar249 < (2'h2)); forvar249 = (forvar249 + (1'h1)))
                begin
                  if (reg241[(4'h9):(4'h9)])
                    begin
                      reg250 <= (wire213 ?
                          ($unsigned(forvar220) ^ reg230) : $signed(forvar249[(1'h0):(1'h0)]));
                      reg251 <= $unsigned({$unsigned((8'hb4))});
                    end
                  else
                    begin
                      reg250 <= $signed($unsigned(reg239));
                      reg251 <= ($unsigned(reg251[(4'h8):(3'h6)]) <= reg231);
                    end
                  for (forvar252 = (1'h0); (forvar252 < (2'h2)); forvar252 = (forvar252 + (1'h1)))
                    begin
                      reg253 <= reg233[(2'h3):(1'h1)];
                    end
                end
              for (forvar254 = (1'h0); (forvar254 < (2'h2)); forvar254 = (forvar254 + (1'h1)))
                begin
                  for (forvar255 = (1'h0); (forvar255 < (1'h0)); forvar255 = (forvar255 + (1'h1)))
                    begin
                      reg256 <= {reg226[(2'h3):(1'h0)]};
                      reg257 <= $unsigned((&$unsigned($signed(forvar238))));
                    end
                end
            end
          else
            begin
              reg238 <= (~^forvar255[(3'h7):(3'h4)]);
            end
        end
      if (($signed($unsigned((&reg230))) & $unsigned(forvar222)))
        begin
          if ((+{($unsigned(forvar255) ?
                  (reg229 ? reg223 : reg233) : ((8'hb8) ? reg218 : reg236))}))
            begin
              for (forvar258 = (1'h0); (forvar258 < (2'h3)); forvar258 = (forvar258 + (1'h1)))
                begin
                  for (forvar259 = (1'h0); (forvar259 < (1'h1)); forvar259 = (forvar259 + (1'h1)))
                    begin
                      reg260 <= ((+(8'hab)) << {wire216[(1'h1):(1'h0)]});
                      reg261 <= $unsigned($unsigned($unsigned((~^reg238))));
                      reg262 <= (((forvar258 + $unsigned((8'haa))) & $signed($unsigned(reg250))) || reg225[(4'h8):(2'h2)]);
                    end
                  if ($unsigned({forvar258}))
                    begin
                      reg263 <= $unsigned(reg243[(1'h0):(1'h0)]);
                      reg264 <= $signed($unsigned(reg223));
                    end
                  else
                    begin
                      reg263 <= forvar228[(3'h7):(3'h5)];
                      reg264 <= $signed(($signed($signed(reg261)) << (((8'ha6) || reg241) <<< forvar222[(1'h0):(1'h0)])));
                    end
                  for (forvar265 = (1'h0); (forvar265 < (2'h2)); forvar265 = (forvar265 + (1'h1)))
                    begin
                      reg266 <= $unsigned(reg243[(1'h0):(1'h0)]);
                      reg267 <= reg238;
                      reg268 <= (8'hb1);
                      reg269 <= forvar222;
                    end
                  for (forvar270 = (1'h0); (forvar270 < (2'h3)); forvar270 = (forvar270 + (1'h1)))
                    begin
                      reg271 <= $signed((!reg236[(1'h0):(1'h0)]));
                    end
                end
              reg272 <= forvar255[(3'h7):(1'h0)];
              for (forvar273 = (1'h0); (forvar273 < (1'h1)); forvar273 = (forvar273 + (1'h1)))
                begin
                  for (forvar274 = (1'h0); (forvar274 < (2'h2)); forvar274 = (forvar274 + (1'h1)))
                    begin
                      reg275 <= ((8'hab) & reg246[(2'h2):(1'h1)]);
                    end
                end
            end
          else
            begin
              if ($unsigned($signed($unsigned((~reg226)))))
                begin
                  for (forvar258 = (1'h0); (forvar258 < (1'h1)); forvar258 = (forvar258 + (1'h1)))
                    begin
                      reg259 <= reg247;
                      reg260 <= reg236;
                    end
                  reg261 <= forvar222[(1'h1):(1'h1)];
                end
              else
                begin
                  for (forvar258 = (1'h0); (forvar258 < (2'h3)); forvar258 = (forvar258 + (1'h1)))
                    begin
                      reg259 <= (((reg229 >> $signed(reg241)) == ((~^reg230) <<< {reg256})) ?
                          $signed(($unsigned(reg259) >> forvar219[(2'h2):(1'h0)])) : reg245);
                    end
                end
            end
          if (($signed($unsigned($unsigned(reg243))) >>> (wire216 << ((~^reg259) ?
              (+reg262) : $unsigned(wire217)))))
            begin
              for (forvar276 = (1'h0); (forvar276 < (1'h1)); forvar276 = (forvar276 + (1'h1)))
                begin
                  reg277 <= ($signed($signed($unsigned(wire212))) ?
                      reg246 : (({reg243} <= $unsigned(forvar228)) ?
                          (|{reg229}) : reg266));
                end
              for (forvar278 = (1'h0); (forvar278 < (1'h1)); forvar278 = (forvar278 + (1'h1)))
                begin
                  for (forvar279 = (1'h0); (forvar279 < (2'h3)); forvar279 = (forvar279 + (1'h1)))
                    begin
                      reg280 <= wire212;
                      reg281 <= reg261;
                      reg282 <= forvar238[(3'h7):(1'h1)];
                      reg283 <= (reg264[(2'h3):(2'h3)] && {$signed(((8'h9f) <= reg233))});
                    end
                  reg284 <= ((reg272[(2'h3):(1'h1)] == (((8'h9d) ?
                          reg236 : forvar279) ?
                      $unsigned(forvar276) : ((8'ha9) - reg242))) || $unsigned(forvar252));
                  for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
                    begin
                      reg286 <= reg283[(4'h8):(3'h6)];
                      reg287 <= $signed((|$signed({reg241})));
                    end
                  for (forvar288 = (1'h0); (forvar288 < (1'h0)); forvar288 = (forvar288 + (1'h1)))
                    begin
                      reg289 <= $signed(forvar273[(1'h0):(1'h0)]);
                      reg290 <= forvar240[(1'h0):(1'h0)];
                    end
                end
              for (forvar291 = (1'h0); (forvar291 < (2'h3)); forvar291 = (forvar291 + (1'h1)))
                begin
                  reg292 <= $unsigned({(8'ha3)});
                  if ($unsigned($unsigned(($signed(reg261) ?
                      $signed(reg231) : (reg280 < forvar258)))))
                    begin
                      reg293 <= $signed((reg233[(1'h1):(1'h0)] ?
                          reg229 : ($signed(reg275) >> (&(8'hb0)))));
                      reg294 <= reg242[(3'h6):(3'h5)];
                      reg295 <= (&wire216[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg293 <= forvar220;
                    end
                end
            end
          else
            begin
              reg276 <= $signed($unsigned((forvar274[(3'h5):(2'h2)] ?
                  $unsigned(forvar278) : (!(8'ha2)))));
            end
          for (forvar296 = (1'h0); (forvar296 < (2'h2)); forvar296 = (forvar296 + (1'h1)))
            begin
              if ((^$unsigned(((-(8'hb8)) <<< (forvar288 ? reg240 : (8'ha8))))))
                begin
                  for (forvar297 = (1'h0); (forvar297 < (1'h0)); forvar297 = (forvar297 + (1'h1)))
                    begin
                      reg298 <= reg284;
                      reg299 <= (~|$signed(($signed(forvar278) ?
                          $unsigned(reg289) : $unsigned(reg280))));
                      reg300 <= reg267;
                    end
                end
              else
                begin
                  if ({reg244})
                    begin
                      reg297 <= reg234;
                    end
                  else
                    begin
                      reg297 <= ($signed((reg225 << $unsigned(forvar219))) ?
                          reg227[(4'hc):(1'h1)] : (8'had));
                      reg298 <= (8'hb2);
                    end
                end
              for (forvar301 = (1'h0); (forvar301 < (1'h1)); forvar301 = (forvar301 + (1'h1)))
                begin
                  for (forvar302 = (1'h0); (forvar302 < (2'h3)); forvar302 = (forvar302 + (1'h1)))
                    begin
                      reg303 <= $signed({(^(8'hb6))});
                    end
                  if ((reg253 >>> forvar278[(2'h3):(1'h1)]))
                    begin
                      reg304 <= $unsigned($signed((8'haf)));
                      reg305 <= (reg269[(3'h7):(2'h2)] ?
                          ({$unsigned(reg244)} ?
                              ((wire212 | reg264) ?
                                  (-reg253) : forvar274[(3'h4):(2'h3)]) : ((~forvar279) << (reg295 >>> (8'h9d)))) : $signed(reg248));
                    end
                  else
                    begin
                      reg304 <= {(-$signed(forvar258))};
                      reg305 <= forvar276[(1'h1):(1'h0)];
                    end
                  for (forvar306 = (1'h0); (forvar306 < (1'h1)); forvar306 = (forvar306 + (1'h1)))
                    begin
                      reg307 <= $signed({$unsigned((!(8'h9f)))});
                      reg308 <= $signed(forvar265[(3'h6):(1'h0)]);
                      reg309 <= (reg226[(2'h3):(1'h0)] ~^ reg283[(3'h4):(2'h2)]);
                    end
                  for (forvar310 = (1'h0); (forvar310 < (1'h0)); forvar310 = (forvar310 + (1'h1)))
                    begin
                      reg311 <= (^~{((reg225 ? reg251 : (8'ha0)) ?
                              {(8'ha0)} : $unsigned((8'hb9)))});
                      reg312 <= (|(8'hb1));
                      reg313 <= forvar265[(4'hd):(1'h1)];
                    end
                end
            end
        end
      else
        begin
          reg258 <= $signed(((((8'ha0) ? forvar273 : reg247) ?
                  reg266[(4'hb):(3'h4)] : $unsigned(reg272)) ?
              (^reg240) : $signed((+reg242))));
          reg259 <= ((8'hb5) >= ($signed((wire217 * reg312)) ?
              ($unsigned(reg289) ?
                  $signed(forvar302) : reg232) : {forvar228[(1'h1):(1'h0)]}));
          if (reg311[(4'hc):(3'h4)])
            begin
              for (forvar260 = (1'h0); (forvar260 < (1'h1)); forvar260 = (forvar260 + (1'h1)))
                begin
                  for (forvar261 = (1'h0); (forvar261 < (1'h0)); forvar261 = (forvar261 + (1'h1)))
                    begin
                      reg262 <= (&($unsigned(((8'hb3) ?
                          (8'ha0) : reg245)) <= $signed(((8'hba) >>> reg266))));
                      reg263 <= ({{((8'haf) ?
                                  reg292 : (8'hb9))}} >>> wire213[(1'h1):(1'h0)]);
                    end
                end
              if ($unsigned($unsigned(reg269[(4'hf):(4'he)])))
                begin
                  for (forvar264 = (1'h0); (forvar264 < (1'h0)); forvar264 = (forvar264 + (1'h1)))
                    begin
                      reg265 <= reg272[(3'h4):(2'h3)];
                      reg266 <= $signed(reg313);
                      reg267 <= reg246[(1'h0):(1'h0)];
                      reg268 <= $signed(($unsigned((~forvar228)) || (^((8'hb1) - reg242))));
                    end
                  if ($signed($signed(($unsigned(forvar296) ^~ reg293))))
                    begin
                      reg269 <= $unsigned(forvar279);
                      reg270 <= reg218[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg269 <= ($unsigned(forvar259[(1'h0):(1'h0)]) ?
                          $unsigned($unsigned((8'ha8))) : ($signed((forvar259 ?
                                  reg309 : (8'h9e))) ?
                              {forvar285[(4'hd):(2'h3)]} : reg297[(2'h2):(2'h2)]));
                      reg270 <= {{forvar279}};
                      reg271 <= reg307;
                      reg272 <= reg304;
                    end
                  reg273 <= (reg245 ?
                      (8'ha2) : $unsigned(($signed(reg223) || $unsigned(reg234))));
                  reg274 <= $unsigned(reg264);
                end
              else
                begin
                  reg264 <= (&(+(~((8'ha7) ? reg264 : reg264))));
                  for (forvar265 = (1'h0); (forvar265 < (1'h1)); forvar265 = (forvar265 + (1'h1)))
                    begin
                      reg266 <= (reg244[(4'h8):(1'h0)] ?
                          {$unsigned($unsigned(forvar278))} : ((!reg309) + $unsigned((reg227 ?
                              reg256 : forvar270))));
                      reg267 <= (+reg271);
                      reg268 <= reg253[(2'h2):(1'h1)];
                      reg269 <= (reg294 ?
                          $signed(reg311) : (!$unsigned(((8'ha4) ?
                              forvar273 : reg276))));
                    end
                  if ({$signed({reg298[(2'h2):(2'h2)]})})
                    begin
                      reg270 <= (~|reg235[(2'h2):(2'h2)]);
                      reg271 <= ($signed((&$unsigned(reg241))) > ((reg235 <<< {(8'h9c)}) >> forvar296));
                    end
                  else
                    begin
                      reg270 <= reg246[(1'h0):(1'h0)];
                      reg271 <= $signed((forvar302 <= $signed(forvar264)));
                    end
                  for (forvar272 = (1'h0); (forvar272 < (2'h3)); forvar272 = (forvar272 + (1'h1)))
                    begin
                      reg273 <= forvar252;
                      reg274 <= reg298;
                      reg275 <= $signed(((((8'haa) ? reg272 : (8'hb1)) ?
                              $signed(reg274) : (^forvar220)) ?
                          ($unsigned((8'hac)) ?
                              reg287[(1'h0):(1'h0)] : ((8'ha2) ?
                                  reg312 : reg227)) : reg313));
                    end
                end
            end
          else
            begin
              for (forvar260 = (1'h0); (forvar260 < (2'h3)); forvar260 = (forvar260 + (1'h1)))
                begin
                  for (forvar261 = (1'h0); (forvar261 < (1'h0)); forvar261 = (forvar261 + (1'h1)))
                    begin
                      reg262 <= $unsigned($unsigned(reg294));
                      reg263 <= $signed(reg242[(2'h3):(2'h3)]);
                      reg264 <= (~|(8'h9f));
                    end
                end
              if (({$unsigned($unsigned(reg253))} ^ $signed(reg267)))
                begin
                  if (reg303[(1'h0):(1'h0)])
                    begin
                      reg265 <= (8'ha0);
                      reg266 <= reg289;
                    end
                  else
                    begin
                      reg265 <= {forvar276};
                    end
                end
              else
                begin
                  if (((^reg305[(3'h6):(2'h3)]) <<< $unsigned(reg313[(4'hc):(2'h3)])))
                    begin
                      reg265 <= (reg282 ?
                          $signed($unsigned(forvar252[(2'h2):(1'h1)])) : (reg239[(1'h0):(1'h0)] >= ((|forvar306) < $unsigned(reg230))));
                      reg266 <= $unsigned(((forvar240 ?
                              ((8'h9e) != reg268) : reg295) ?
                          {(&forvar219)} : ($unsigned(reg305) ?
                              (reg239 >= (8'hab)) : (wire217 ?
                                  reg225 : reg226))));
                      reg267 <= reg283;
                    end
                  else
                    begin
                      reg265 <= (((&{forvar302}) + {(^reg224)}) >> forvar264);
                    end
                  if (((~(^~(~&forvar265))) ^~ forvar260[(4'hb):(2'h3)]))
                    begin
                      reg268 <= $signed((^~$unsigned($signed(reg263))));
                      reg269 <= (^($signed($signed(reg242)) ?
                          $unsigned($signed(reg269)) : reg265));
                      reg270 <= {$signed((~^(~forvar219)))};
                    end
                  else
                    begin
                      reg268 <= $signed(reg224[(3'h7):(3'h7)]);
                    end
                  if ($signed($signed(($signed((8'hb1)) ?
                      (8'hb4) : (reg277 ? (8'hb5) : reg280)))))
                    begin
                      reg271 <= (^~$unsigned((forvar258[(4'h9):(3'h6)] != (reg261 ?
                          reg290 : (8'hb3)))));
                      reg272 <= ($signed($unsigned($signed(reg265))) ?
                          $signed(reg283[(1'h0):(1'h0)]) : (($unsigned(forvar254) * $signed(forvar255)) != (reg264[(3'h4):(2'h3)] >> $unsigned(forvar279))));
                    end
                  else
                    begin
                      reg271 <= reg308;
                      reg272 <= $signed(reg259[(2'h2):(1'h1)]);
                    end
                end
              for (forvar273 = (1'h0); (forvar273 < (1'h0)); forvar273 = (forvar273 + (1'h1)))
                begin
                  reg274 <= {(8'haa)};
                  if (((reg311[(3'h6):(1'h1)] ?
                          (&((8'hba) ? forvar297 : reg284)) : (-(reg261 ?
                              (8'haf) : reg224))) ?
                      $signed((8'haa)) : $signed(wire217)))
                    begin
                      reg275 <= $signed((((&(8'ha2)) ?
                              (reg276 ^~ forvar264) : (|forvar265)) ?
                          (!(-reg224)) : forvar302[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg275 <= reg308[(2'h3):(2'h2)];
                      reg276 <= ($signed((~&(~forvar288))) ?
                          $signed(((&(8'ha8)) ?
                              reg226[(2'h3):(1'h1)] : (~|(8'hb2)))) : {(~|$signed(reg275))});
                    end
                  for (forvar277 = (1'h0); (forvar277 < (1'h0)); forvar277 = (forvar277 + (1'h1)))
                    begin
                      reg278 <= {(+$signed($unsigned(reg262)))};
                    end
                  if (forvar249[(3'h7):(2'h2)])
                    begin
                      reg279 <= (($unsigned($signed(reg293)) ?
                          (forvar273 >>> $signed(reg256)) : $signed((-forvar237))) < {forvar237});
                      reg280 <= forvar297[(1'h1):(1'h0)];
                      reg281 <= reg304;
                    end
                  else
                    begin
                      reg279 <= {$unsigned((((8'h9c) ^~ reg272) ?
                              reg278[(1'h0):(1'h0)] : reg281[(1'h1):(1'h1)]))};
                      reg280 <= ((|(~|reg294[(1'h0):(1'h0)])) ?
                          forvar297 : {$signed({forvar219})});
                      reg281 <= $unsigned((+reg225[(4'h9):(2'h3)]));
                      reg282 <= wire217;
                    end
                end
              for (forvar283 = (1'h0); (forvar283 < (2'h2)); forvar283 = (forvar283 + (1'h1)))
                begin
                  if (reg312)
                    begin
                      reg284 <= reg223;
                      reg285 <= (reg281 > $signed(reg311[(3'h7):(2'h2)]));
                    end
                  else
                    begin
                      reg284 <= {$unsigned(reg309)};
                    end
                  if (reg244)
                    begin
                      reg286 <= reg307;
                    end
                  else
                    begin
                      reg286 <= forvar255[(2'h3):(2'h2)];
                      reg287 <= $signed((($signed(reg278) >>> forvar228[(1'h1):(1'h1)]) ^~ ($unsigned((8'had)) ?
                          {forvar259} : reg264[(2'h2):(1'h1)])));
                    end
                  for (forvar288 = (1'h0); (forvar288 < (2'h2)); forvar288 = (forvar288 + (1'h1)))
                    begin
                      reg289 <= $unsigned(forvar255[(1'h0):(1'h0)]);
                      reg290 <= ((($signed(forvar297) ?
                              (reg313 ?
                                  wire217 : reg286) : reg239[(4'h8):(2'h2)]) >> ($unsigned(reg271) ^~ (&reg232))) ?
                          $signed((~&$signed(reg290))) : $unsigned($unsigned($signed((8'ha2)))));
                    end
                  for (forvar291 = (1'h0); (forvar291 < (1'h1)); forvar291 = (forvar291 + (1'h1)))
                    begin
                      reg292 <= reg256[(4'hc):(4'ha)];
                      reg293 <= (~&(8'ha8));
                    end
                end
            end
          reg294 <= ($unsigned(forvar255[(1'h0):(1'h0)]) ?
              {(reg257[(3'h7):(1'h0)] ?
                      $unsigned(reg299) : $signed(reg236))} : (~reg305));
        end
    end
  assign wire314 = ({forvar297} ?
                       $unsigned($signed($unsigned(wire216))) : reg271[(3'h6):(1'h0)]);
  assign wire315 = {(8'ha2)};
  assign wire316 = reg313[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg317 <= reg272[(3'h6):(1'h1)];
      for (forvar318 = (1'h0); (forvar318 < (2'h2)); forvar318 = (forvar318 + (1'h1)))
        begin
          reg319 <= forvar277;
          if (($signed($unsigned((reg262 ^~ reg313))) ?
              forvar288[(1'h0):(1'h0)] : ({(reg294 ?
                      forvar254 : reg279)} - (^(forvar274 ?
                  reg226 : forvar219)))))
            begin
              if (($signed(reg258[(2'h2):(1'h1)]) << reg294[(3'h4):(1'h0)]))
                begin
                  if ({$unsigned((~^(forvar297 || reg304)))})
                    begin
                      reg320 <= reg305[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg320 <= reg262[(3'h5):(3'h5)];
                      reg321 <= ($unsigned({(reg270 > (8'hb7))}) ?
                          (&($unsigned(forvar249) ?
                              (~reg295) : wire212[(3'h5):(3'h5)])) : $signed(({forvar260} & {reg312})));
                      reg322 <= reg279[(1'h0):(1'h0)];
                    end
                  for (forvar323 = (1'h0); (forvar323 < (2'h3)); forvar323 = (forvar323 + (1'h1)))
                    begin
                      reg324 <= $unsigned((^reg232[(1'h1):(1'h0)]));
                      reg325 <= ($signed(reg221[(2'h2):(1'h0)]) == reg224[(3'h7):(1'h1)]);
                      reg326 <= {$signed(forvar291[(3'h4):(2'h2)])};
                      reg327 <= $signed((8'ha0));
                    end
                  reg328 <= forvar261[(3'h7):(3'h7)];
                end
              else
                begin
                  if ((-{reg311[(4'he):(1'h1)]}))
                    begin
                      reg320 <= reg270[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg320 <= $unsigned(reg289[(3'h7):(3'h4)]);
                      reg321 <= reg276[(1'h1):(1'h1)];
                      reg322 <= $signed((~|reg226[(2'h3):(1'h0)]));
                    end
                end
              if (reg230)
                begin
                  if ((forvar273[(1'h1):(1'h1)] == {(~^$unsigned(reg328))}))
                    begin
                      reg329 <= ($unsigned((reg275[(3'h7):(1'h0)] ?
                          reg243 : (reg232 ^ forvar219))) >= ((forvar222 >> forvar272[(4'h8):(3'h7)]) || ((reg227 ?
                              (8'haa) : reg243) ?
                          forvar306[(2'h3):(1'h0)] : forvar288[(2'h3):(2'h3)])));
                      reg330 <= reg259[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg329 <= ((^~reg272[(4'h8):(1'h1)]) ?
                          (reg311[(3'h5):(3'h4)] ?
                              {$signed(forvar255)} : (&(-(8'hb6)))) : reg235);
                      reg330 <= $unsigned(($unsigned((reg290 ?
                              reg284 : wire314)) ?
                          reg277[(2'h2):(2'h2)] : (|$signed(reg257))));
                    end
                end
              else
                begin
                  if ({({reg276[(3'h6):(1'h1)]} ?
                          reg266[(3'h6):(1'h0)] : $signed($signed(forvar240)))})
                    begin
                      reg329 <= $unsigned($unsigned(forvar265[(4'hb):(3'h6)]));
                      reg330 <= $unsigned((!reg250[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg329 <= $signed($signed((reg286[(3'h4):(1'h1)] ?
                          reg273 : $unsigned(forvar228))));
                      reg330 <= ((($unsigned(reg286) ?
                              forvar283[(4'hb):(4'hb)] : (reg268 ?
                                  reg273 : reg226)) - ($signed(reg238) ?
                              (reg269 != forvar291) : ((8'hb4) ?
                                  reg293 : reg268))) ?
                          $signed({(&reg270)}) : reg295[(3'h6):(3'h4)]);
                      reg331 <= $signed((forvar254[(4'h9):(2'h3)] ?
                          forvar297[(1'h1):(1'h1)] : $unsigned(forvar285)));
                      reg332 <= {$unsigned(forvar279)};
                    end
                  for (forvar333 = (1'h0); (forvar333 < (2'h3)); forvar333 = (forvar333 + (1'h1)))
                    begin
                      reg334 <= (8'hb6);
                      reg335 <= ((&($unsigned(reg218) << (reg290 >>> (8'ha7)))) ?
                          ($unsigned($signed(reg297)) ?
                              ((~^(8'ha3)) > (^~reg304)) : (-$signed(forvar277))) : (~forvar274));
                      reg336 <= reg239;
                      reg337 <= reg240;
                    end
                end
            end
          else
            begin
              for (forvar320 = (1'h0); (forvar320 < (1'h0)); forvar320 = (forvar320 + (1'h1)))
                begin
                  if ({(reg298 << (~&(forvar306 ? (8'h9f) : forvar291)))})
                    begin
                      reg321 <= (reg229 ?
                          ($signed(reg279[(4'hb):(4'h9)]) ?
                              reg224 : ((reg337 ~^ reg287) & $signed((8'haa)))) : reg335[(1'h1):(1'h0)]);
                      reg322 <= $signed($signed((reg308 ^ $signed(reg260))));
                      reg323 <= ((&((reg265 ?
                              forvar283 : reg292) && (^~reg265))) ?
                          ((reg337[(1'h0):(1'h0)] ?
                              (reg239 ? reg262 : reg232) : ((8'hb1) ?
                                  forvar265 : reg311)) & $unsigned({reg282})) : $unsigned(($signed(forvar261) * (~^wire217))));
                      reg324 <= (8'h9e);
                    end
                  else
                    begin
                      reg321 <= ({wire213[(3'h5):(2'h2)]} ^ $unsigned($signed(reg259)));
                    end
                  for (forvar325 = (1'h0); (forvar325 < (2'h2)); forvar325 = (forvar325 + (1'h1)))
                    begin
                      reg326 <= reg267;
                      reg327 <= $signed(($signed(forvar220[(2'h2):(1'h1)]) ?
                          (~(-forvar274)) : reg257[(4'ha):(2'h2)]));
                      reg328 <= (|$unsigned($signed($signed((8'ha1)))));
                    end
                end
              for (forvar329 = (1'h0); (forvar329 < (2'h3)); forvar329 = (forvar329 + (1'h1)))
                begin
                  for (forvar330 = (1'h0); (forvar330 < (1'h1)); forvar330 = (forvar330 + (1'h1)))
                    begin
                      reg331 <= reg234;
                      reg332 <= $signed(reg324[(3'h6):(3'h6)]);
                    end
                end
              reg333 <= reg230;
            end
          reg338 <= forvar306[(1'h0):(1'h0)];
          reg339 <= reg317;
        end
      if ($unsigned((forvar276 >= (|reg279[(4'hd):(2'h2)]))))
        begin
          reg340 <= forvar302;
          for (forvar341 = (1'h0); (forvar341 < (2'h3)); forvar341 = (forvar341 + (1'h1)))
            begin
              if (reg321)
                begin
                  for (forvar342 = (1'h0); (forvar342 < (2'h3)); forvar342 = (forvar342 + (1'h1)))
                    begin
                      reg343 <= reg311[(3'h4):(2'h3)];
                      reg344 <= ((^~reg290) ?
                          $signed({$signed(forvar252)}) : reg287[(1'h1):(1'h1)]);
                      reg345 <= $signed(reg243);
                      reg346 <= reg266;
                    end
                  for (forvar347 = (1'h0); (forvar347 < (2'h3)); forvar347 = (forvar347 + (1'h1)))
                    begin
                      reg348 <= (~&$unsigned((8'ha2)));
                      reg349 <= reg224;
                    end
                  for (forvar350 = (1'h0); (forvar350 < (2'h2)); forvar350 = (forvar350 + (1'h1)))
                    begin
                      reg351 <= $signed(((+(reg346 >= reg300)) - ((reg259 ?
                          forvar288 : reg227) << (+forvar220))));
                      reg352 <= (!{forvar265[(4'hb):(1'h0)]});
                      reg353 <= reg276;
                    end
                end
              else
                begin
                  if ($signed(($unsigned(reg261[(1'h0):(1'h0)]) ?
                      $unsigned(reg224[(3'h6):(1'h1)]) : {$unsigned(reg278)})))
                    begin
                      reg342 <= $signed((^~($signed(reg321) ?
                          reg294[(2'h3):(2'h3)] : $unsigned(reg297))));
                      reg343 <= $signed((&$unsigned(((8'ha3) << reg345))));
                    end
                  else
                    begin
                      reg342 <= $unsigned($unsigned(((forvar329 ?
                              reg238 : reg280) ?
                          forvar258[(3'h5):(2'h3)] : (+reg272))));
                      reg343 <= $unsigned($unsigned((-reg329)));
                    end
                  if ((forvar297[(2'h2):(2'h2)] ?
                      (~$signed((reg232 ?
                          reg344 : reg257))) : {(!$signed(reg293))}))
                    begin
                      reg344 <= {($signed({reg242}) ?
                              ($signed((8'ha2)) ?
                                  forvar272[(4'h9):(2'h2)] : ((8'hb7) ?
                                      reg337 : forvar310)) : {reg225})};
                      reg345 <= $unsigned(reg274);
                      reg346 <= wire212[(4'ha):(3'h6)];
                      reg347 <= (forvar254 >>> $unsigned($signed((reg279 < reg338))));
                    end
                  else
                    begin
                      reg344 <= ((~^reg331[(1'h1):(1'h0)]) ?
                          $signed($signed($signed(reg323))) : (($unsigned(reg282) <<< reg323[(1'h1):(1'h0)]) | reg331[(4'hb):(2'h3)]));
                      reg345 <= (reg352[(3'h7):(2'h2)] ?
                          $unsigned({reg236}) : $unsigned($signed((forvar270 ^~ reg309))));
                    end
                  for (forvar348 = (1'h0); (forvar348 < (2'h3)); forvar348 = (forvar348 + (1'h1)))
                    begin
                      reg349 <= $unsigned($unsigned(forvar260));
                      reg350 <= forvar318[(3'h7):(3'h4)];
                      reg351 <= $signed(($unsigned(reg309) ?
                          (((8'hb6) ? (8'hb2) : reg347) | ((8'ha4) ?
                              forvar341 : forvar254)) : (forvar288[(2'h2):(2'h2)] ?
                              forvar325 : (reg286 | (8'ha5)))));
                      reg352 <= ((-$unsigned($unsigned(reg244))) <<< reg339[(2'h2):(2'h2)]);
                    end
                end
              for (forvar354 = (1'h0); (forvar354 < (1'h0)); forvar354 = (forvar354 + (1'h1)))
                begin
                  for (forvar355 = (1'h0); (forvar355 < (1'h0)); forvar355 = (forvar355 + (1'h1)))
                    begin
                      reg356 <= $unsigned({(forvar259[(1'h1):(1'h0)] ?
                              (~|forvar333) : (^forvar270))});
                      reg357 <= forvar325;
                    end
                  for (forvar358 = (1'h0); (forvar358 < (2'h2)); forvar358 = (forvar358 + (1'h1)))
                    begin
                      reg359 <= $signed($unsigned($signed({forvar291})));
                      reg360 <= {reg307[(3'h5):(2'h3)]};
                      reg361 <= ($unsigned($signed($signed((8'h9c)))) ?
                          (&$unsigned(reg256[(1'h1):(1'h0)])) : $unsigned((-$unsigned(forvar318))));
                    end
                  if ((&($unsigned(wire316) >>> $signed(reg309[(4'hb):(3'h7)]))))
                    begin
                      reg362 <= $signed((reg285[(3'h4):(2'h2)] ?
                          (~&(reg319 - forvar238)) : (^$unsigned(reg233))));
                    end
                  else
                    begin
                      reg362 <= $unsigned($unsigned((reg360 ?
                          (!forvar220) : $signed((8'hb8)))));
                      reg363 <= $unsigned((reg278[(1'h1):(1'h1)] ?
                          ($unsigned(forvar310) ^~ $unsigned((8'ha7))) : $unsigned({reg327})));
                      reg364 <= ($unsigned({{reg265}}) && $unsigned(((reg266 > reg342) >> forvar260)));
                    end
                end
            end
          reg365 <= reg363;
        end
      else
        begin
          for (forvar340 = (1'h0); (forvar340 < (1'h0)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 <= $signed((|($signed(forvar278) ?
                  {(8'ha0)} : (|reg342))));
              for (forvar342 = (1'h0); (forvar342 < (2'h3)); forvar342 = (forvar342 + (1'h1)))
                begin
                  reg343 <= (reg218 >>> ($signed((reg317 > forvar340)) ?
                      forvar354[(1'h0):(1'h0)] : reg221[(4'ha):(3'h6)]));
                end
            end
          if (reg233[(4'hb):(3'h4)])
            begin
              for (forvar344 = (1'h0); (forvar344 < (1'h1)); forvar344 = (forvar344 + (1'h1)))
                begin
                  for (forvar345 = (1'h0); (forvar345 < (2'h2)); forvar345 = (forvar345 + (1'h1)))
                    begin
                      reg346 <= reg298[(2'h2):(1'h0)];
                      reg347 <= $signed($unsigned(reg224));
                      reg348 <= ((-({reg292} <<< ((8'h9e) != forvar350))) >> reg266[(4'h9):(2'h3)]);
                      reg349 <= reg225[(3'h4):(1'h1)];
                    end
                end
            end
          else
            begin
              reg344 <= (($unsigned(reg348[(1'h1):(1'h0)]) ?
                  $unsigned($signed(reg243)) : ($unsigned(reg258) ?
                      forvar259[(1'h1):(1'h0)] : (reg360 ?
                          reg346 : reg348))) && (reg325[(4'hc):(2'h2)] || $unsigned($signed((8'hba)))));
              if (wire212)
                begin
                  if (((!$signed(reg278)) & {$unsigned(forvar325)}))
                    begin
                      reg345 <= reg241[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg345 <= (^~{reg238});
                    end
                end
              else
                begin
                  reg345 <= $unsigned($signed($unsigned((^~(8'ha2)))));
                  for (forvar346 = (1'h0); (forvar346 < (2'h2)); forvar346 = (forvar346 + (1'h1)))
                    begin
                      reg347 <= ($unsigned(reg338[(1'h1):(1'h0)]) - reg224[(2'h3):(2'h3)]);
                    end
                end
            end
          for (forvar350 = (1'h0); (forvar350 < (2'h3)); forvar350 = (forvar350 + (1'h1)))
            begin
              if ($unsigned(reg268))
                begin
                  for (forvar351 = (1'h0); (forvar351 < (2'h3)); forvar351 = (forvar351 + (1'h1)))
                    begin
                      reg352 <= $unsigned({(^~((8'hb8) ?
                              forvar254 : forvar222))});
                      reg353 <= ($unsigned((reg357[(3'h7):(2'h3)] > (~&forvar228))) ?
                          ({forvar325[(1'h0):(1'h0)]} ?
                              (^(forvar340 ?
                                  reg353 : reg257)) : ($unsigned((8'hb9)) + (forvar274 & reg359))) : (^~(&reg305)));
                      reg354 <= $unsigned((~&((reg325 <<< (8'hb8)) < $unsigned((8'ha8)))));
                      reg355 <= {$unsigned((+forvar237[(4'hd):(3'h6)]))};
                    end
                end
              else
                begin
                  for (forvar351 = (1'h0); (forvar351 < (2'h3)); forvar351 = (forvar351 + (1'h1)))
                    begin
                      reg352 <= ($signed(reg360[(3'h4):(1'h0)]) ?
                          {reg343} : (!(forvar277 ?
                              $unsigned(forvar302) : $unsigned((8'h9e)))));
                      reg353 <= (~^forvar350);
                      reg354 <= (~(~&{(reg308 ^ reg339)}));
                    end
                  for (forvar355 = (1'h0); (forvar355 < (2'h3)); forvar355 = (forvar355 + (1'h1)))
                    begin
                      reg356 <= ($unsigned($signed(((8'hb6) > reg229))) ?
                          $signed(($unsigned((8'ha6)) ?
                              $signed(forvar240) : $signed(reg357))) : (~&(8'hb4)));
                      reg357 <= $unsigned(reg230[(2'h2):(2'h2)]);
                    end
                end
              if ($signed($signed((^~(forvar302 ? reg303 : forvar306)))))
                begin
                  reg358 <= $unsigned(($unsigned((forvar270 ?
                      reg332 : reg328)) <= {(~&reg232)}));
                  reg359 <= $signed((^~$signed((~reg250))));
                  for (forvar360 = (1'h0); (forvar360 < (2'h3)); forvar360 = (forvar360 + (1'h1)))
                    begin
                      reg361 <= forvar355[(3'h6):(1'h1)];
                      reg362 <= reg246[(2'h2):(2'h2)];
                      reg363 <= ($unsigned((^~forvar340)) ?
                          (($signed(reg328) - $signed(forvar302)) > wire316[(4'h8):(3'h7)]) : reg332[(1'h0):(1'h0)]);
                      reg364 <= (reg361[(4'ha):(1'h0)] ^ forvar222[(2'h2):(1'h0)]);
                    end
                end
              else
                begin
                  if (((reg345 * (|$signed(reg313))) ^ ({$signed((8'hb2))} != {(!(8'hb0))})))
                    begin
                      reg358 <= reg253[(1'h1):(1'h0)];
                      reg359 <= ($unsigned(reg274) ? (&reg338) : wire315);
                    end
                  else
                    begin
                      reg358 <= $unsigned(reg260[(3'h7):(3'h6)]);
                      reg359 <= (~(((reg332 & reg347) > (forvar219 < reg270)) ?
                          $signed((^forvar270)) : ((reg327 || reg300) ?
                              ((8'h9c) ^~ reg341) : $signed(reg338))));
                    end
                  for (forvar360 = (1'h0); (forvar360 < (2'h3)); forvar360 = (forvar360 + (1'h1)))
                    begin
                      reg361 <= ((($signed((8'had)) ?
                              (reg324 ? reg235 : reg241) : (^forvar341)) ?
                          $signed($signed(forvar220)) : (+(reg240 >> reg267))) << (|{(~&reg350)}));
                      reg362 <= reg340;
                      reg363 <= reg229[(4'hf):(4'h9)];
                      reg364 <= ($unsigned({(~&reg227)}) ?
                          $unsigned(wire316[(4'ha):(4'h8)]) : {{$unsigned((8'hb7))}});
                    end
                end
              for (forvar365 = (1'h0); (forvar365 < (1'h1)); forvar365 = (forvar365 + (1'h1)))
                begin
                  reg366 <= reg361;
                end
              if ((reg355 ?
                  ((~(~^reg348)) ?
                      ((reg361 ? (8'had) : forvar283) ?
                          (reg225 ?
                              (8'ha7) : (8'hb6)) : $unsigned((8'hb4))) : ((forvar301 ?
                              reg257 : reg341) ?
                          (reg325 ? reg275 : (8'hb1)) : {wire217})) : wire314))
                begin
                  reg367 <= (({$signed(reg336)} ?
                          $unsigned($signed(reg232)) : (reg275[(2'h3):(1'h1)] == $unsigned(reg277))) ?
                      (reg259[(3'h6):(2'h3)] >= ({reg362} + {reg360})) : ((forvar345 < $signed(forvar358)) ?
                          {$unsigned(forvar285)} : reg227));
                  for (forvar368 = (1'h0); (forvar368 < (2'h2)); forvar368 = (forvar368 + (1'h1)))
                    begin
                      reg369 <= ((((-reg284) ?
                              $signed(reg274) : $signed(forvar310)) && ({reg284} >= (^forvar270))) ?
                          $unsigned($unsigned($unsigned(reg363))) : ($signed({(8'hb9)}) - $unsigned((forvar283 <<< (8'hb5)))));
                      reg370 <= reg336;
                    end
                  if ((^$signed(reg328)))
                    begin
                      reg371 <= $unsigned(($signed((reg354 ?
                              forvar333 : reg309)) ?
                          ($unsigned(reg241) ?
                              (reg248 ?
                                  reg226 : reg266) : $unsigned(reg356)) : {forvar365}));
                    end
                  else
                    begin
                      reg371 <= $signed($unsigned(forvar302[(1'h0):(1'h0)]));
                      reg372 <= (!$unsigned(((8'hb2) ?
                          (wire314 ? reg308 : reg317) : $signed(wire212))));
                      reg373 <= forvar261;
                      reg374 <= (8'hb0);
                    end
                end
              else
                begin
                  if ((^(reg261 >> {(reg238 ? reg355 : reg370)})))
                    begin
                      reg367 <= reg262[(2'h3):(1'h1)];
                      reg368 <= (reg227 <= $signed($signed(reg360)));
                      reg369 <= {reg322[(4'ha):(3'h6)]};
                    end
                  else
                    begin
                      reg367 <= ($unsigned((+((8'h9e) ~^ reg351))) & forvar355[(4'hd):(3'h7)]);
                      reg368 <= reg342[(4'h8):(3'h7)];
                      reg369 <= ($unsigned((^(8'hab))) ?
                          reg329[(1'h1):(1'h0)] : $unsigned(reg244));
                    end
                  if (({((reg262 ? reg339 : (8'hba)) ?
                          (^~forvar255) : reg330)} >= $signed($unsigned(reg343[(1'h0):(1'h0)]))))
                    begin
                      reg370 <= (($signed(forvar283) ? reg348 : reg335) ?
                          $signed((reg322 == (8'hb3))) : reg371[(1'h0):(1'h0)]);
                      reg371 <= $signed($unsigned(((wire212 ?
                          reg325 : reg235) & $unsigned(wire217))));
                      reg372 <= $signed($signed((!(reg373 ? reg224 : reg295))));
                      reg373 <= $signed(((forvar333 ?
                          (reg274 ?
                              forvar365 : reg290) : $signed(reg351)) - ((~|reg240) ?
                          (&reg304) : (~&reg286))));
                    end
                  else
                    begin
                      reg370 <= $signed($signed(((reg354 ? (8'hac) : reg359) ?
                          reg343 : reg260[(3'h6):(1'h0)])));
                      reg371 <= forvar310;
                      reg372 <= ($unsigned(($unsigned(reg257) ?
                              reg349[(2'h3):(2'h2)] : reg281)) ?
                          forvar347[(3'h5):(2'h2)] : (|reg354));
                      reg373 <= $signed(((&{wire216}) ?
                          (~(~|reg343)) : $signed(reg370)));
                    end
                end
            end
        end
      if (reg333[(1'h1):(1'h0)])
        begin
          for (forvar375 = (1'h0); (forvar375 < (2'h3)); forvar375 = (forvar375 + (1'h1)))
            begin
              for (forvar376 = (1'h0); (forvar376 < (1'h0)); forvar376 = (forvar376 + (1'h1)))
                begin
                  if (reg319[(3'h5):(3'h4)])
                    begin
                      reg377 <= (-(+forvar340[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg377 <= (!$unsigned($signed(((8'hb0) ?
                          reg365 : forvar347))));
                      reg378 <= reg266;
                      reg379 <= $signed(reg364);
                      reg380 <= forvar228[(4'h8):(1'h0)];
                    end
                  reg381 <= forvar264[(2'h3):(1'h1)];
                end
              if ($signed($unsigned((8'ha6))))
                begin
                  reg382 <= reg267[(2'h3):(1'h1)];
                  for (forvar383 = (1'h0); (forvar383 < (1'h1)); forvar383 = (forvar383 + (1'h1)))
                    begin
                      reg384 <= reg363;
                      reg385 <= (~((8'h9e) >>> {(forvar358 == forvar383)}));
                      reg386 <= $unsigned(((~^(~|forvar252)) || reg264[(1'h1):(1'h1)]));
                      reg387 <= ($unsigned(reg358[(4'h9):(2'h3)]) >= $signed(forvar368[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar382 = (1'h0); (forvar382 < (2'h3)); forvar382 = (forvar382 + (1'h1)))
                    begin
                      reg383 <= {reg294};
                      reg384 <= (~(~$unsigned($unsigned((8'ha4)))));
                      reg385 <= (($unsigned((reg232 < forvar296)) ?
                              forvar368[(2'h2):(1'h1)] : ($unsigned(reg384) ?
                                  $unsigned(forvar252) : reg346[(4'h9):(3'h6)])) ?
                          reg285[(3'h4):(1'h0)] : $signed((((8'hb0) & (8'ha6)) > $signed(reg342))));
                    end
                  for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
                    begin
                      reg387 <= (8'hb6);
                      reg388 <= reg280[(3'h5):(1'h1)];
                    end
                end
              for (forvar389 = (1'h0); (forvar389 < (2'h3)); forvar389 = (forvar389 + (1'h1)))
                begin
                  reg390 <= reg307[(2'h2):(2'h2)];
                  for (forvar391 = (1'h0); (forvar391 < (2'h2)); forvar391 = (forvar391 + (1'h1)))
                    begin
                      reg392 <= ($signed(($unsigned(forvar351) > {reg378})) ^ forvar333[(4'ha):(4'h9)]);
                      reg393 <= reg382[(4'ha):(4'h9)];
                    end
                  reg394 <= reg243[(3'h4):(2'h2)];
                end
            end
        end
      else
        begin
          for (forvar375 = (1'h0); (forvar375 < (2'h3)); forvar375 = (forvar375 + (1'h1)))
            begin
              if (reg258)
                begin
                  if ($unsigned({reg248[(4'hc):(2'h3)]}))
                    begin
                      reg376 <= forvar278;
                      reg377 <= (reg289 >> ((^~(reg297 ? reg374 : forvar333)) ?
                          $unsigned((~&forvar340)) : {(~^forvar382)}));
                      reg378 <= (^reg299);
                    end
                  else
                    begin
                      reg376 <= $signed((reg362[(1'h0):(1'h0)] ?
                          (forvar342 >>> (~(8'ha9))) : ($signed(reg348) > (~|reg245))));
                    end
                  if ((((|(8'ha7)) ?
                          $unsigned(((8'haa) ?
                              forvar288 : (8'hb8))) : forvar375[(3'h7):(2'h2)]) ?
                      forvar391 : $signed((reg322 | reg383[(4'hd):(4'ha)]))))
                    begin
                      reg379 <= (^~(~{$signed((8'ha8))}));
                    end
                  else
                    begin
                      reg379 <= (~$unsigned($unsigned(forvar276[(1'h0):(1'h0)])));
                    end
                end
              else
                begin
                  if ({($unsigned($unsigned(reg324)) < ($signed(reg390) ?
                          ((8'ha0) == reg250) : reg263[(2'h3):(2'h3)]))})
                    begin
                      reg376 <= reg298[(1'h0):(1'h0)];
                      reg377 <= (~$unsigned((~^forvar274)));
                      reg378 <= forvar355;
                    end
                  else
                    begin
                      reg376 <= (~(~&(reg239 & {reg286})));
                      reg377 <= (forvar342[(3'h7):(2'h3)] ?
                          forvar237[(4'ha):(1'h0)] : ((+$unsigned((8'hb7))) ?
                              {forvar344[(4'he):(4'h9)]} : ((~&reg243) ~^ forvar278)));
                      reg378 <= (^~({(reg277 | (8'ha1))} ?
                          (forvar265 ?
                              $unsigned(forvar386) : forvar347[(1'h0):(1'h0)]) : reg349));
                    end
                  for (forvar379 = (1'h0); (forvar379 < (2'h2)); forvar379 = (forvar379 + (1'h1)))
                    begin
                      reg380 <= ((8'hb6) >= reg241);
                      reg381 <= (($signed($signed(reg370)) * wire213[(3'h7):(2'h3)]) ?
                          (wire316 ?
                              reg368[(1'h0):(1'h0)] : ($unsigned(reg260) <= {reg299})) : ({reg363} ?
                              reg371 : (reg390 ^~ $signed(forvar355))));
                      reg382 <= ((^$signed(forvar296[(1'h1):(1'h0)])) ?
                          forvar383[(2'h3):(2'h3)] : ($unsigned(((8'ha9) <= forvar383)) ?
                              forvar260[(3'h4):(2'h2)] : reg319));
                      reg383 <= (reg304 >> {({reg327} ^ (reg276 | (8'hb9)))});
                    end
                  if ((&(reg355[(4'h8):(3'h4)] != $signed(reg328[(3'h6):(1'h1)]))))
                    begin
                      reg384 <= $signed({((!reg359) << reg273)});
                      reg385 <= reg354;
                      reg386 <= {reg308};
                    end
                  else
                    begin
                      reg384 <= reg246[(1'h0):(1'h0)];
                    end
                end
              for (forvar387 = (1'h0); (forvar387 < (2'h2)); forvar387 = (forvar387 + (1'h1)))
                begin
                  for (forvar388 = (1'h0); (forvar388 < (2'h3)); forvar388 = (forvar388 + (1'h1)))
                    begin
                      reg389 <= (($unsigned($unsigned((8'had))) ?
                          ($unsigned(reg344) >>> (-forvar264)) : forvar228) == $signed($signed(reg269)));
                      reg390 <= (8'hb7);
                    end
                  for (forvar391 = (1'h0); (forvar391 < (2'h3)); forvar391 = (forvar391 + (1'h1)))
                    begin
                      reg392 <= ($unsigned(forvar274) ?
                          (^~forvar318) : (~&(!$signed(forvar375))));
                      reg393 <= ((($signed(reg334) >= (reg353 <<< reg323)) * reg380) ?
                          ((reg225 >= reg298[(2'h2):(1'h0)]) * forvar264) : {forvar278[(2'h2):(1'h0)]});
                      reg394 <= (forvar279[(3'h5):(2'h3)] & ($signed({reg345}) ?
                          ($unsigned(reg271) | $signed(forvar288)) : $signed(((8'had) ?
                              reg251 : (8'ha7)))));
                    end
                  if ((&reg351[(2'h2):(2'h2)]))
                    begin
                      reg395 <= (|reg354[(1'h1):(1'h0)]);
                      reg396 <= ($signed($signed((!(8'hb6)))) ~^ (8'ha9));
                      reg397 <= reg264[(1'h0):(1'h0)];
                      reg398 <= ((forvar329[(3'h4):(1'h0)] ^ $signed($signed(forvar375))) ?
                          $signed((-$unsigned((8'hb1)))) : ($signed((forvar341 << reg263)) * (forvar333[(4'h8):(3'h7)] | $signed((8'ha6)))));
                    end
                  else
                    begin
                      reg395 <= $signed(($unsigned($unsigned(reg335)) * $signed(reg309[(4'hb):(3'h4)])));
                      reg396 <= ((^~$unsigned($signed(reg238))) ~^ ((reg395[(2'h3):(2'h3)] ?
                          (forvar261 * forvar297) : (reg321 <<< reg230)) >>> reg246[(1'h0):(1'h0)]));
                      reg397 <= {(|$unsigned($signed(forvar348)))};
                      reg398 <= reg395;
                    end
                  for (forvar399 = (1'h0); (forvar399 < (1'h1)); forvar399 = (forvar399 + (1'h1)))
                    begin
                      reg400 <= $signed({$signed(reg299[(4'he):(1'h1)])});
                      reg401 <= ((~^reg338[(2'h2):(1'h1)]) ?
                          (~|(^~(reg241 >= reg372))) : ({$signed(forvar238)} < {reg342[(3'h6):(3'h4)]}));
                      reg402 <= (reg381[(1'h1):(1'h0)] ?
                          $signed(((^~forvar291) ?
                              $unsigned(reg242) : {forvar320})) : reg240);
                    end
                end
              for (forvar403 = (1'h0); (forvar403 < (2'h2)); forvar403 = (forvar403 + (1'h1)))
                begin
                  reg404 <= reg385;
                  for (forvar405 = (1'h0); (forvar405 < (1'h1)); forvar405 = (forvar405 + (1'h1)))
                    begin
                      reg406 <= $unsigned({($unsigned(forvar219) ?
                              {(8'hb4)} : (reg297 - forvar273))});
                    end
                  for (forvar407 = (1'h0); (forvar407 < (2'h3)); forvar407 = (forvar407 + (1'h1)))
                    begin
                      reg408 <= $unsigned(reg368[(1'h1):(1'h1)]);
                      reg409 <= (reg229 ~^ (~|$signed((reg319 ^ reg382))));
                    end
                end
              for (forvar410 = (1'h0); (forvar410 < (1'h1)); forvar410 = (forvar410 + (1'h1)))
                begin
                  if ($signed(reg323[(1'h1):(1'h1)]))
                    begin
                      reg411 <= reg392;
                    end
                  else
                    begin
                      reg411 <= (~|$signed(reg400));
                      reg412 <= ({$signed((+reg275))} > forvar274);
                    end
                  if ($signed(((^~{forvar265}) | ($unsigned(reg408) ?
                      $signed(reg317) : (forvar330 == reg307)))))
                    begin
                      reg413 <= (-$unsigned(forvar261[(4'hc):(4'hc)]));
                      reg414 <= (reg368 ~^ $signed((&(reg327 >>> reg342))));
                      reg415 <= wire216;
                    end
                  else
                    begin
                      reg413 <= $unsigned((8'hac));
                      reg414 <= (((-(forvar351 ? reg286 : forvar261)) ?
                          (-$signed(reg245)) : ($unsigned(reg236) < (reg387 ?
                              (8'h9e) : reg303))) - (+(~|forvar375[(4'h9):(4'h8)])));
                    end
                  if (forvar238)
                    begin
                      reg416 <= (&{$unsigned($signed(forvar387))});
                      reg417 <= (~^reg317[(1'h1):(1'h1)]);
                      reg418 <= $signed(reg359[(3'h5):(1'h1)]);
                    end
                  else
                    begin
                      reg416 <= wire212[(3'h5):(1'h1)];
                      reg417 <= ($unsigned($signed((forvar296 < (8'h9d)))) ?
                          $signed(((reg221 ?
                              wire216 : reg328) ^ $signed(reg331))) : reg382);
                      reg418 <= ($signed($unsigned(((8'haf) ?
                              forvar389 : reg284))) ?
                          $signed(reg341) : forvar222);
                    end
                  reg419 <= forvar346[(3'h7):(2'h2)];
                end
            end
          if (reg303)
            begin
              if ({(forvar249[(2'h2):(2'h2)] ?
                      $signed({forvar344}) : $unsigned($signed(reg273)))})
                begin
                  if ({$unsigned(((~&forvar297) * (reg295 ?
                          forvar347 : (8'ha8))))})
                    begin
                      reg420 <= {reg393};
                      reg421 <= forvar291;
                      reg422 <= {(^reg376[(3'h5):(3'h4)])};
                      reg423 <= (~|reg267[(3'h5):(1'h1)]);
                    end
                  else
                    begin
                      reg420 <= (wire217[(2'h3):(2'h3)] + reg379[(4'h8):(2'h2)]);
                      reg421 <= reg383[(1'h0):(1'h0)];
                      reg422 <= reg300;
                      reg423 <= {(forvar301[(1'h0):(1'h0)] < (8'hb0))};
                    end
                  if (reg341)
                    begin
                      reg424 <= $signed(((^~$signed(forvar260)) && {(reg416 <<< reg250)}));
                      reg425 <= $unsigned(reg225[(4'ha):(3'h5)]);
                      reg426 <= ($signed(reg406[(3'h5):(1'h0)]) ?
                          reg253[(3'h4):(2'h3)] : reg234);
                      reg427 <= (~(&forvar254[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg424 <= $signed($signed((reg289 >= (forvar330 ?
                          wire212 : forvar388))));
                      reg425 <= forvar342[(2'h2):(1'h1)];
                    end
                  for (forvar428 = (1'h0); (forvar428 < (2'h2)); forvar428 = (forvar428 + (1'h1)))
                    begin
                      reg429 <= {($unsigned((reg246 <= forvar219)) <= $signed((&reg360)))};
                      reg430 <= (^~(forvar382 ?
                          $signed(reg280) : (^$signed(reg387))));
                      reg431 <= $signed((+((8'hb9) ?
                          $unsigned(reg412) : (+forvar344))));
                      reg432 <= $signed($unsigned((~|(reg335 ?
                          forvar273 : reg325))));
                    end
                end
              else
                begin
                  if ({(((|reg263) || wire315) * reg236)})
                    begin
                      reg420 <= $unsigned(forvar382[(4'h8):(1'h1)]);
                    end
                  else
                    begin
                      reg420 <= $unsigned(reg234);
                      reg421 <= reg419;
                      reg422 <= (($signed($unsigned(reg354)) ?
                              (reg334 ?
                                  $unsigned((8'haa)) : (reg235 * reg394)) : ((forvar260 ?
                                      reg430 : reg422) ?
                                  {reg348} : {reg262})) ?
                          forvar220[(2'h2):(1'h1)] : reg323[(2'h2):(2'h2)]);
                    end
                  for (forvar423 = (1'h0); (forvar423 < (1'h1)); forvar423 = (forvar423 + (1'h1)))
                    begin
                      reg424 <= $unsigned((({forvar325} ?
                          (reg343 ~^ reg294) : reg423) * ($unsigned(reg413) + ((8'hba) < forvar265))));
                      reg425 <= (reg258[(3'h4):(3'h4)] ?
                          ($signed((~(8'ha0))) ?
                              (~&reg224[(2'h3):(1'h1)]) : $signed((forvar291 == reg415))) : $unsigned($signed(forvar386[(1'h0):(1'h0)])));
                      reg426 <= $unsigned(reg300);
                    end
                  if (($unsigned(((~^reg271) ?
                          $unsigned((8'h9c)) : forvar368[(2'h3):(2'h2)])) ?
                      (&(reg413[(4'hb):(4'hb)] & $signed(reg304))) : (((reg262 != reg326) >> reg283[(1'h0):(1'h0)]) ?
                          ($unsigned(reg384) == (&reg266)) : $unsigned(forvar347[(2'h2):(1'h0)]))))
                    begin
                      reg427 <= forvar261[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg427 <= $unsigned((~&$unsigned((^~reg330))));
                      reg428 <= (+reg402[(2'h2):(1'h1)]);
                      reg429 <= (+$unsigned({$unsigned(reg352)}));
                    end
                  for (forvar430 = (1'h0); (forvar430 < (1'h1)); forvar430 = (forvar430 + (1'h1)))
                    begin
                      reg431 <= {(!reg280[(4'he):(1'h1)])};
                      reg432 <= reg275[(2'h3):(2'h3)];
                      reg433 <= (^{$signed(reg232)});
                    end
                end
              reg434 <= ((((reg342 >= reg387) ?
                      $signed(reg280) : $unsigned(reg347)) & ((forvar354 ?
                          reg247 : (8'hba)) ?
                      forvar259[(1'h1):(1'h0)] : (forvar285 ?
                          forvar329 : reg406))) ?
                  reg278 : ($signed(forvar382[(4'ha):(3'h7)]) ?
                      reg427 : $signed($unsigned(reg245))));
              for (forvar435 = (1'h0); (forvar435 < (2'h2)); forvar435 = (forvar435 + (1'h1)))
                begin
                  for (forvar436 = (1'h0); (forvar436 < (2'h2)); forvar436 = (forvar436 + (1'h1)))
                    begin
                      reg437 <= (($unsigned(((8'hb8) + reg247)) ^~ (~$unsigned(reg312))) ?
                          (!reg380[(1'h0):(1'h0)]) : {reg366});
                      reg438 <= (forvar350 ?
                          reg277[(1'h0):(1'h0)] : ($unsigned({reg270}) << {$unsigned(reg334)}));
                      reg439 <= (-(-$unsigned($signed(reg234))));
                      reg440 <= ($signed($unsigned((forvar258 ^ reg432))) >> reg344);
                    end
                end
            end
          else
            begin
              if ($signed($unsigned(forvar325[(4'h9):(4'h9)])))
                begin
                  if ((~^{forvar410[(1'h0):(1'h0)]}))
                    begin
                      reg420 <= reg371[(4'hc):(3'h7)];
                      reg421 <= {$signed(wire213[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg420 <= {(8'ha3)};
                    end
                  if (forvar237[(4'hd):(1'h0)])
                    begin
                      reg422 <= $signed((($signed(reg273) ?
                          forvar391[(1'h1):(1'h0)] : (reg374 ^ reg374)) > $unsigned(((8'hb9) != reg432))));
                      reg423 <= ($signed(forvar278) >= (((forvar387 != forvar405) ?
                          reg263 : (reg426 ? reg226 : reg365)) | ((forvar325 ?
                          reg404 : reg383) < ((8'hb2) > reg292))));
                    end
                  else
                    begin
                      reg422 <= $signed($unsigned(((~reg439) ?
                          (reg282 > reg294) : (reg409 ? (8'hb8) : reg388))));
                      reg423 <= $unsigned($signed(((reg271 || reg341) ?
                          $signed(reg380) : ((8'hb9) ? reg321 : reg411))));
                      reg424 <= (|((8'hb8) << forvar254));
                    end
                  for (forvar425 = (1'h0); (forvar425 < (2'h2)); forvar425 = (forvar425 + (1'h1)))
                    begin
                      reg426 <= (^~((~|{(8'hb9)}) ?
                          ($unsigned((8'hb9)) ?
                              forvar259 : {wire316}) : $unsigned(reg386[(2'h2):(1'h0)])));
                      reg427 <= reg267[(2'h2):(2'h2)];
                    end
                  if ({$signed((forvar277 ?
                          $signed(reg242) : (reg267 ? wire214 : wire215)))})
                    begin
                      reg428 <= reg402[(2'h2):(2'h2)];
                      reg429 <= $unsigned(reg419[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg428 <= reg232;
                    end
                end
              else
                begin
                  for (forvar420 = (1'h0); (forvar420 < (2'h3)); forvar420 = (forvar420 + (1'h1)))
                    begin
                      reg421 <= reg284[(4'h9):(3'h4)];
                    end
                  reg422 <= ($unsigned((~|(8'ha1))) ?
                      reg234[(1'h1):(1'h0)] : ((forvar265[(2'h3):(1'h0)] >> (reg266 + forvar355)) && {forvar428[(3'h4):(2'h3)]}));
                  for (forvar423 = (1'h0); (forvar423 < (1'h1)); forvar423 = (forvar423 + (1'h1)))
                    begin
                      reg424 <= $unsigned($signed(reg226[(3'h4):(2'h2)]));
                    end
                  reg425 <= $signed(reg245[(2'h3):(2'h2)]);
                end
            end
          reg441 <= (reg394[(1'h1):(1'h1)] ?
              $signed(((8'hae) - (reg358 ?
                  reg388 : reg372))) : reg287[(2'h2):(1'h0)]);
          reg442 <= (forvar405 ?
              ($signed({(8'hb3)}) < reg387[(2'h2):(1'h0)]) : (forvar238[(3'h6):(2'h3)] ?
                  $unsigned(reg412) : $unsigned((8'hb7))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar443 = (1'h0); (forvar443 < (1'h0)); forvar443 = (forvar443 + (1'h1)))
        begin
          reg444 <= reg309;
          for (forvar445 = (1'h0); (forvar445 < (2'h3)); forvar445 = (forvar445 + (1'h1)))
            begin
              if ($signed(reg327))
                begin
                  if ($unsigned($unsigned((^~$signed(forvar297)))))
                    begin
                      reg446 <= ($signed({{forvar278}}) < {$signed((~&reg250))});
                      reg447 <= ((~^reg414[(1'h0):(1'h0)]) && $unsigned(((~^(8'ha3)) ^~ (reg390 < forvar277))));
                      reg448 <= ((~|$unsigned(forvar436)) >>> forvar355);
                    end
                  else
                    begin
                      reg446 <= reg263;
                    end
                end
              else
                begin
                  if ($unsigned((((reg231 ^~ forvar350) ?
                          $signed(reg392) : forvar342) ?
                      $unsigned((+reg409)) : (^~(|reg350)))))
                    begin
                      reg446 <= reg295;
                      reg447 <= {(|(~reg333))};
                    end
                  else
                    begin
                      reg446 <= {(&forvar420)};
                    end
                  if (reg233)
                    begin
                      reg448 <= (((!(reg327 ? reg385 : reg411)) ?
                              reg409 : $signed($signed(reg236))) ?
                          (|$unsigned($signed((8'hb5)))) : ($signed($unsigned(reg283)) >> forvar436));
                      reg449 <= reg434;
                      reg450 <= {($signed((reg369 + forvar273)) ?
                              (reg324 || wire214) : reg371)};
                    end
                  else
                    begin
                      reg448 <= reg380[(4'hc):(1'h0)];
                      reg449 <= wire316;
                    end
                  for (forvar451 = (1'h0); (forvar451 < (1'h1)); forvar451 = (forvar451 + (1'h1)))
                    begin
                      reg452 <= $unsigned(($signed($unsigned(forvar383)) ?
                          reg360 : ((reg366 ? reg230 : forvar360) ?
                              (^~reg376) : (+forvar238))));
                    end
                  for (forvar453 = (1'h0); (forvar453 < (2'h3)); forvar453 = (forvar453 + (1'h1)))
                    begin
                      reg454 <= (8'hb8);
                      reg455 <= $unsigned((!$unsigned((forvar264 - reg422))));
                      reg456 <= {forvar220};
                    end
                end
              if ($unsigned((^~(&reg371))))
                begin
                  reg457 <= ($unsigned((reg427 ^ $unsigned(forvar342))) ?
                      (^$unsigned(forvar285)) : $unsigned(reg416[(3'h5):(2'h2)]));
                end
              else
                begin
                  for (forvar457 = (1'h0); (forvar457 < (2'h2)); forvar457 = (forvar457 + (1'h1)))
                    begin
                      reg458 <= reg398;
                      reg459 <= ((reg353[(3'h6):(2'h3)] == $unsigned(reg413[(2'h3):(2'h2)])) ?
                          (8'h9f) : (+reg373[(3'h6):(2'h3)]));
                      reg460 <= forvar320;
                      reg461 <= (forvar351 ?
                          reg458[(4'ha):(1'h0)] : reg372[(4'hd):(4'hb)]);
                    end
                  for (forvar462 = (1'h0); (forvar462 < (2'h2)); forvar462 = (forvar462 + (1'h1)))
                    begin
                      reg463 <= (((forvar276[(3'h4):(1'h1)] >= (reg336 >> forvar428)) ?
                              reg308[(1'h1):(1'h1)] : (~|$signed(reg360))) ?
                          forvar410[(1'h0):(1'h0)] : reg416);
                      reg464 <= $unsigned($signed({(~&reg269)}));
                      reg465 <= (8'hab);
                      reg466 <= reg336[(2'h2):(1'h0)];
                    end
                  reg467 <= forvar254[(4'h9):(1'h0)];
                  reg468 <= (&forvar276);
                end
              reg469 <= (8'haf);
            end
          if ((+$signed(((~|forvar407) >>> reg236))))
            begin
              if (reg456[(2'h3):(2'h3)])
                begin
                  for (forvar470 = (1'h0); (forvar470 < (2'h2)); forvar470 = (forvar470 + (1'h1)))
                    begin
                      reg471 <= ((^reg259) || ({reg344} ?
                          (reg279[(1'h0):(1'h0)] < (wire314 <= forvar297)) : (-$unsigned(reg231))));
                    end
                  if (forvar259)
                    begin
                      reg472 <= (^$signed($unsigned(reg275)));
                      reg473 <= reg269[(3'h7):(3'h4)];
                      reg474 <= $signed(($unsigned(forvar323) ?
                          reg356 : $signed({reg398})));
                      reg475 <= forvar383[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg472 <= (&(~$signed((reg331 << reg464))));
                      reg473 <= reg371[(2'h3):(2'h3)];
                      reg474 <= (forvar259[(1'h1):(1'h0)] | $unsigned(((^reg303) && (reg472 & forvar274))));
                      reg475 <= (forvar302 ? forvar358[(1'h0):(1'h0)] : reg311);
                    end
                  if ($unsigned($unsigned($signed(reg231))))
                    begin
                      reg476 <= (($signed($signed(reg274)) ?
                              (~|reg283[(2'h3):(1'h1)]) : (!(reg457 ?
                                  (8'haa) : reg363))) ?
                          (($unsigned((8'h9d)) & (reg420 ?
                              (8'ha0) : forvar443)) == $unsigned($unsigned(reg276))) : ((^(|(8'ha2))) + ((reg457 << forvar462) ?
                              reg259 : {(8'hae)})));
                    end
                  else
                    begin
                      reg476 <= reg331[(3'h4):(2'h2)];
                      reg477 <= {$signed($unsigned((reg411 ~^ forvar410)))};
                      reg478 <= (8'hb4);
                      reg479 <= $signed(((forvar462 ?
                          forvar320[(2'h3):(1'h0)] : reg461) <<< {reg230[(2'h3):(1'h1)]}));
                    end
                  if (($signed($signed(reg469[(1'h0):(1'h0)])) < ($signed($signed(reg357)) + ($unsigned((8'ha9)) ?
                      (forvar301 <= reg341) : $signed((8'ha4))))))
                    begin
                      reg480 <= reg434[(3'h5):(2'h3)];
                      reg481 <= $unsigned(($signed($signed(reg384)) ?
                          reg243[(1'h1):(1'h0)] : (reg348[(2'h3):(1'h0)] > reg394[(1'h0):(1'h0)])));
                      reg482 <= ($unsigned(forvar354) ?
                          (^(8'hb3)) : reg430[(4'h8):(2'h2)]);
                      reg483 <= (~&(($unsigned(reg357) ?
                              (~^(8'hb5)) : forvar360) ?
                          $signed({wire216}) : {reg320}));
                    end
                  else
                    begin
                      reg480 <= ((+reg245[(1'h1):(1'h0)]) ?
                          $signed($unsigned((8'h9f))) : reg279[(4'ha):(3'h7)]);
                      reg481 <= (^~{$signed($signed((8'ha5)))});
                      reg482 <= {$unsigned($unsigned(reg479))};
                    end
                end
              else
                begin
                  for (forvar470 = (1'h0); (forvar470 < (2'h3)); forvar470 = (forvar470 + (1'h1)))
                    begin
                      reg471 <= forvar425[(2'h3):(1'h0)];
                      reg472 <= (~|(((^~forvar240) ?
                              {reg345} : ((8'ha4) + reg408)) ?
                          (^(~^reg387)) : (|(reg469 ? (8'hb8) : forvar383))));
                      reg473 <= reg238;
                      reg474 <= ((!reg298) << $signed(((reg464 ^~ (8'hae)) ?
                          (reg259 ? reg317 : reg253) : (reg266 < forvar320))));
                    end
                  if ({({$unsigned(reg401)} ?
                          ((reg377 ?
                              (8'haa) : reg481) == (reg362 ~^ forvar291)) : forvar296[(4'ha):(4'ha)])})
                    begin
                      reg475 <= $signed(reg335[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg475 <= reg257;
                      reg476 <= reg221[(3'h5):(2'h3)];
                      reg477 <= (~&$signed({forvar350[(2'h3):(2'h2)]}));
                      reg478 <= (reg303 == ($unsigned((+reg395)) ?
                          ((forvar272 ?
                              reg263 : forvar219) | forvar252[(2'h3):(1'h1)]) : forvar405));
                    end
                end
              if ((forvar368[(1'h0):(1'h0)] || $signed({reg326[(4'h8):(3'h5)]})))
                begin
                  for (forvar484 = (1'h0); (forvar484 < (1'h0)); forvar484 = (forvar484 + (1'h1)))
                    begin
                      reg485 <= (~^((reg414 ?
                          (~|reg372) : (reg230 ?
                              reg312 : reg325)) > ($signed(reg331) ^~ (|reg466))));
                    end
                  if (reg320[(1'h1):(1'h0)])
                    begin
                      reg486 <= (+reg246[(1'h1):(1'h0)]);
                      reg487 <= $signed($signed(($unsigned(forvar238) ?
                          ((8'hb5) ? reg408 : reg247) : (reg440 ?
                              reg346 : (8'hb7)))));
                      reg488 <= $signed($signed({reg262}));
                      reg489 <= forvar391[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg486 <= {reg312};
                    end
                  reg490 <= {{((reg239 <= reg486) ?
                              (8'h9d) : $signed(reg334))}};
                end
              else
                begin
                  for (forvar484 = (1'h0); (forvar484 < (1'h0)); forvar484 = (forvar484 + (1'h1)))
                    begin
                      reg485 <= ($unsigned(reg474) > $signed((~&$signed(reg408))));
                    end
                  for (forvar486 = (1'h0); (forvar486 < (2'h3)); forvar486 = (forvar486 + (1'h1)))
                    begin
                      reg487 <= (~$signed($unsigned($unsigned((8'h9c)))));
                      reg488 <= (({reg478} ?
                              $unsigned(reg483) : $signed((~forvar420))) ?
                          (-(8'hba)) : (reg395[(1'h0):(1'h0)] ?
                              reg328[(4'h9):(4'h8)] : (!reg239)));
                      reg489 <= reg416;
                    end
                end
              reg491 <= ((~(~&(reg411 ? reg234 : (8'hae)))) ?
                  reg430 : $unsigned({{forvar261}}));
              reg492 <= forvar389[(3'h5):(1'h0)];
            end
          else
            begin
              for (forvar470 = (1'h0); (forvar470 < (1'h0)); forvar470 = (forvar470 + (1'h1)))
                begin
                  for (forvar471 = (1'h0); (forvar471 < (2'h2)); forvar471 = (forvar471 + (1'h1)))
                    begin
                      reg472 <= reg479;
                    end
                  for (forvar473 = (1'h0); (forvar473 < (1'h0)); forvar473 = (forvar473 + (1'h1)))
                    begin
                      reg474 <= $signed(({(reg264 >>> forvar410)} ?
                          {$unsigned(reg312)} : (8'h9d)));
                    end
                end
              for (forvar475 = (1'h0); (forvar475 < (2'h2)); forvar475 = (forvar475 + (1'h1)))
                begin
                  reg476 <= forvar252[(2'h2):(1'h1)];
                  for (forvar477 = (1'h0); (forvar477 < (1'h1)); forvar477 = (forvar477 + (1'h1)))
                    begin
                      reg478 <= (reg441 ?
                          {((~|reg239) & (+forvar252))} : ((^~(forvar341 * reg251)) * (reg271[(3'h4):(1'h1)] | $unsigned(reg262))));
                      reg479 <= (reg430[(3'h6):(1'h1)] ?
                          (($unsigned(reg323) + $unsigned(forvar306)) ?
                              $unsigned($unsigned(reg437)) : ({reg439} ?
                                  $unsigned(reg279) : reg433)) : ({(8'hb3)} != $signed((reg284 ?
                              reg241 : reg459))));
                      reg480 <= {reg421};
                    end
                  if (reg278)
                    begin
                      reg481 <= (|$signed(reg322));
                      reg482 <= forvar329;
                    end
                  else
                    begin
                      reg481 <= reg388[(2'h3):(1'h0)];
                    end
                  for (forvar483 = (1'h0); (forvar483 < (1'h0)); forvar483 = (forvar483 + (1'h1)))
                    begin
                      reg484 <= ($unsigned(forvar365[(1'h1):(1'h1)]) | $signed({$signed(reg258)}));
                      reg485 <= $signed(((~(8'ha8)) ?
                          reg385[(4'hf):(1'h1)] : (+reg251[(4'h8):(3'h7)])));
                      reg486 <= reg227;
                      reg487 <= $signed($unsigned((((8'hb0) << reg319) ?
                          (reg396 ? forvar272 : (8'ha3)) : {forvar430})));
                    end
                end
            end
        end
      for (forvar493 = (1'h0); (forvar493 < (1'h0)); forvar493 = (forvar493 + (1'h1)))
        begin
          if ({{$unsigned((reg385 >> reg457))}})
            begin
              reg494 <= {$signed(((forvar445 ^ (8'hba)) >>> $signed(reg263)))};
            end
          else
            begin
              for (forvar494 = (1'h0); (forvar494 < (1'h0)); forvar494 = (forvar494 + (1'h1)))
                begin
                  if (reg393)
                    begin
                      reg495 <= (($signed((reg293 >>> reg342)) ?
                              reg366[(2'h2):(1'h0)] : ($unsigned(forvar405) || (8'hb7))) ?
                          forvar462[(1'h1):(1'h0)] : (&(!(~&forvar382))));
                      reg496 <= $signed((reg439[(4'hd):(4'hc)] ?
                          {((8'hae) ?
                                  reg440 : reg427)} : $unsigned((^~forvar443))));
                      reg497 <= (~&reg472);
                      reg498 <= (|{(-((8'ha3) ? reg347 : reg477))});
                    end
                  else
                    begin
                      reg495 <= reg330[(4'ha):(1'h1)];
                    end
                  reg499 <= forvar301;
                end
              for (forvar500 = (1'h0); (forvar500 < (1'h1)); forvar500 = (forvar500 + (1'h1)))
                begin
                  if ($signed((reg279 ~^ $signed((reg283 ? reg269 : (8'ha7))))))
                    begin
                      reg501 <= reg290;
                      reg502 <= (reg433 + reg241);
                    end
                  else
                    begin
                      reg501 <= reg277;
                      reg502 <= reg368;
                    end
                  for (forvar503 = (1'h0); (forvar503 < (2'h2)); forvar503 = (forvar503 + (1'h1)))
                    begin
                      reg504 <= $signed(($unsigned({reg267}) ?
                          (&(~^reg300)) : ($signed((8'hae)) ?
                              reg502[(4'hf):(4'hb)] : $signed(reg370))));
                      reg505 <= $unsigned((reg406[(2'h2):(2'h2)] ?
                          (-(reg440 ^~ reg264)) : (~forvar254[(1'h0):(1'h0)])));
                    end
                end
              if (((reg225[(4'ha):(2'h3)] * ((reg502 >> reg458) - $signed(reg415))) ?
                  (forvar453 != {forvar240[(1'h1):(1'h0)]}) : ((reg281 >= {reg454}) ~^ $signed((^~forvar238)))))
                begin
                  if (reg388[(2'h3):(2'h3)])
                    begin
                      reg506 <= reg250;
                      reg507 <= ((forvar360[(1'h1):(1'h1)] && (|forvar430)) ?
                          (+reg373[(3'h7):(3'h5)]) : $signed(((reg346 ^~ reg487) + forvar301)));
                      reg508 <= reg334[(3'h5):(3'h4)];
                      reg509 <= ($unsigned(($signed(forvar389) ?
                              reg434 : $unsigned((8'ha5)))) ?
                          $unsigned((~&reg418[(3'h4):(3'h4)])) : $unsigned(reg240[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg506 <= ({$unsigned((^reg468))} ?
                          (^~(8'hb7)) : {$unsigned((reg384 ?
                                  reg498 : reg456))});
                      reg507 <= ($signed(forvar445) << $signed((reg473[(1'h0):(1'h0)] ?
                          $unsigned(reg452) : $signed(forvar403))));
                    end
                  for (forvar510 = (1'h0); (forvar510 < (1'h1)); forvar510 = (forvar510 + (1'h1)))
                    begin
                      reg511 <= $signed($unsigned($unsigned((reg324 != forvar222))));
                      reg512 <= (^~(((forvar453 <<< forvar237) << (reg325 <<< reg349)) == (^(~|reg440))));
                      reg513 <= (~&{$signed(reg241)});
                    end
                  for (forvar514 = (1'h0); (forvar514 < (1'h1)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= $unsigned($signed(reg317[(3'h5):(2'h3)]));
                    end
                  if ($unsigned((reg230[(1'h0):(1'h0)] ?
                      (reg465[(1'h1):(1'h1)] ^~ $signed(forvar462)) : (8'ha4))))
                    begin
                      reg516 <= (~|{reg304});
                    end
                  else
                    begin
                      reg516 <= ($signed((~|{forvar270})) && $unsigned($signed((~^reg238))));
                      reg517 <= forvar443[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar506 = (1'h0); (forvar506 < (1'h1)); forvar506 = (forvar506 + (1'h1)))
                    begin
                      reg507 <= reg235;
                      reg508 <= reg476[(3'h4):(1'h1)];
                    end
                  for (forvar509 = (1'h0); (forvar509 < (2'h3)); forvar509 = (forvar509 + (1'h1)))
                    begin
                      reg510 <= $unsigned(reg516[(3'h4):(2'h3)]);
                      reg511 <= (($unsigned((reg388 ?
                              (8'haf) : reg339)) ^~ ($signed(reg417) ?
                              ((8'ha0) >> (8'hb8)) : $unsigned(reg469))) ?
                          ((((8'h9e) ?
                              forvar259 : forvar325) < (~reg348)) & (!$signed(forvar252))) : $unsigned((~&reg274)));
                    end
                  if ((8'hb3))
                    begin
                      reg512 <= $unsigned((|(!forvar484)));
                      reg513 <= reg373[(3'h4):(2'h3)];
                      reg514 <= reg344;
                      reg515 <= forvar509;
                    end
                  else
                    begin
                      reg512 <= (reg243 ?
                          (($signed((8'ha2)) | (forvar273 <<< (8'hb9))) ?
                              $unsigned(((8'ha0) ?
                                  forvar486 : forvar345)) : {reg488}) : $signed(reg421));
                    end
                end
            end
          if ((reg241 || (~|(~&$signed(reg431)))))
            begin
              if ((($signed($signed((8'ha8))) ?
                      $unsigned((forvar389 ?
                          reg477 : reg467)) : (~^(^forvar329))) ?
                  $signed((reg389[(3'h5):(2'h3)] < (&reg245))) : $unsigned(forvar237)))
                begin
                  if (reg427)
                    begin
                      reg518 <= reg444[(4'hc):(2'h2)];
                      reg519 <= $signed((~(&$signed(reg330))));
                      reg520 <= (reg438 ?
                          ({$unsigned(reg326)} ?
                              {reg440} : $signed(reg332[(2'h3):(2'h3)])) : $unsigned((|$unsigned(reg353))));
                    end
                  else
                    begin
                      reg518 <= (((!(^forvar228)) <<< ({(8'ha6)} & (reg487 > reg502))) ?
                          reg274[(5'h10):(4'ha)] : (~($unsigned(reg368) ^~ (reg286 ?
                              (8'hac) : reg335))));
                      reg519 <= {(~(reg483[(1'h0):(1'h0)] ?
                              (reg424 || reg430) : reg243[(1'h0):(1'h0)]))};
                    end
                end
              else
                begin
                  reg518 <= (~^($signed((-reg377)) | $signed({forvar323})));
                  if ((&(({reg259} ? (reg505 | reg262) : $unsigned(forvar341)) ?
                      reg492 : (8'hb0))))
                    begin
                      reg519 <= ((^~$signed(reg364[(3'h5):(3'h5)])) ?
                          reg478 : reg229);
                      reg520 <= (8'hb1);
                      reg521 <= forvar360;
                      reg522 <= reg473[(4'h9):(3'h5)];
                    end
                  else
                    begin
                      reg519 <= $signed($signed($unsigned(reg400)));
                      reg520 <= (^~$unsigned((&$unsigned(reg459))));
                      reg521 <= (reg345 ?
                          reg442 : $signed($unsigned((-reg476))));
                    end
                  reg523 <= reg242[(4'ha):(3'h4)];
                end
              for (forvar524 = (1'h0); (forvar524 < (2'h3)); forvar524 = (forvar524 + (1'h1)))
                begin
                  if ({reg521[(2'h2):(2'h2)]})
                    begin
                      reg525 <= {$signed($signed(reg446[(1'h0):(1'h0)]))};
                      reg526 <= {(reg406 ?
                              (reg390 ?
                                  (forvar484 ?
                                      reg340 : (8'hba)) : (~&wire214)) : (8'h9e))};
                      reg527 <= $unsigned(reg242[(4'he):(1'h1)]);
                      reg528 <= $signed((8'ha8));
                    end
                  else
                    begin
                      reg525 <= ((($signed(reg251) - (reg253 * reg260)) >> $signed({forvar368})) ?
                          reg415 : (~({reg383} ? (8'ha7) : (~^wire316))));
                      reg526 <= (^~reg253[(3'h4):(2'h2)]);
                      reg527 <= ($unsigned((~&(8'hab))) >>> $signed(($signed(reg433) ?
                          (^reg225) : reg406)));
                    end
                  for (forvar529 = (1'h0); (forvar529 < (1'h0)); forvar529 = (forvar529 + (1'h1)))
                    begin
                      reg530 <= ((forvar403 & (8'hac)) && (forvar420[(4'h8):(2'h2)] ^ (~(reg406 >= forvar514))));
                    end
                  for (forvar531 = (1'h0); (forvar531 < (2'h3)); forvar531 = (forvar531 + (1'h1)))
                    begin
                      reg532 <= forvar383[(3'h4):(2'h3)];
                      reg533 <= {$unsigned(reg421)};
                      reg534 <= reg265[(1'h1):(1'h0)];
                      reg535 <= reg381;
                    end
                end
            end
          else
            begin
              if (forvar302)
                begin
                  if (($unsigned(reg377) - ((&(reg340 ? (8'had) : reg313)) ?
                      forvar375 : (((8'hb9) < forvar310) ?
                          (8'ha2) : (reg338 ? reg350 : reg242)))))
                    begin
                      reg518 <= (reg245 ?
                          reg519[(2'h2):(2'h2)] : forvar301[(1'h1):(1'h0)]);
                      reg519 <= forvar451[(1'h0):(1'h0)];
                      reg520 <= forvar423;
                    end
                  else
                    begin
                      reg518 <= {($unsigned($unsigned(reg256)) || $unsigned((reg534 ?
                              reg471 : reg413)))};
                      reg519 <= $signed((((8'h9d) | {forvar531}) ?
                          (reg239[(3'h6):(1'h0)] ?
                              (~&(8'ha1)) : reg488[(2'h3):(1'h1)]) : {$signed(reg298)}));
                    end
                  for (forvar521 = (1'h0); (forvar521 < (1'h0)); forvar521 = (forvar521 + (1'h1)))
                    begin
                      reg522 <= reg527;
                      reg523 <= {$unsigned((reg447[(2'h3):(2'h3)] || reg265))};
                      reg524 <= forvar252;
                    end
                  for (forvar525 = (1'h0); (forvar525 < (2'h2)); forvar525 = (forvar525 + (1'h1)))
                    begin
                      reg526 <= reg528[(1'h1):(1'h0)];
                    end
                  for (forvar527 = (1'h0); (forvar527 < (2'h3)); forvar527 = (forvar527 + (1'h1)))
                    begin
                      reg528 <= $unsigned($signed((reg411[(2'h3):(2'h3)] != reg454)));
                      reg529 <= $signed((reg335[(3'h5):(1'h0)] ?
                          (-((8'hba) ? reg428 : reg527)) : ($unsigned(reg534) ?
                              $unsigned(forvar423) : {reg452})));
                      reg530 <= $signed($unsigned((((8'hb0) ?
                          reg372 : forvar425) >> (reg336 ? reg487 : reg508))));
                    end
                end
              else
                begin
                  if ({(!(reg317[(1'h0):(1'h0)] ?
                          (&reg507) : $signed(wire212)))})
                    begin
                      reg518 <= reg259;
                      reg519 <= $signed(((&$signed(reg334)) ?
                          $signed(reg319[(2'h2):(2'h2)]) : $signed((reg534 ?
                              (8'haf) : reg366))));
                    end
                  else
                    begin
                      reg518 <= (-$unsigned($signed($signed(wire213))));
                    end
                  reg520 <= $unsigned((($signed((8'h9f)) ?
                      ((8'h9f) && (8'hb9)) : {reg393}) && (-{reg342})));
                  if (reg281[(2'h3):(2'h2)])
                    begin
                      reg521 <= (~^$signed((^~forvar477[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg521 <= reg463[(2'h3):(1'h0)];
                      reg522 <= reg430[(4'hd):(4'hc)];
                    end
                end
              for (forvar531 = (1'h0); (forvar531 < (1'h1)); forvar531 = (forvar531 + (1'h1)))
                begin
                  if ((~|reg378))
                    begin
                      reg532 <= $unsigned(reg369[(4'hb):(4'hb)]);
                    end
                  else
                    begin
                      reg532 <= reg251;
                      reg533 <= reg337;
                      reg534 <= $unsigned($signed($signed((forvar514 << reg376))));
                    end
                  for (forvar535 = (1'h0); (forvar535 < (2'h2)); forvar535 = (forvar535 + (1'h1)))
                    begin
                      reg536 <= $signed((forvar445 - $signed(reg357[(3'h5):(3'h5)])));
                      reg537 <= $signed(wire216);
                    end
                  for (forvar538 = (1'h0); (forvar538 < (2'h2)); forvar538 = (forvar538 + (1'h1)))
                    begin
                      reg539 <= (8'ha9);
                      reg540 <= ((|$signed((forvar382 ?
                          reg535 : reg484))) >> {(~reg497)});
                      reg541 <= (8'hb6);
                    end
                end
              for (forvar542 = (1'h0); (forvar542 < (2'h2)); forvar542 = (forvar542 + (1'h1)))
                begin
                  if (forvar423[(2'h2):(2'h2)])
                    begin
                      reg543 <= reg348[(2'h3):(1'h1)];
                      reg544 <= reg521[(2'h3):(1'h1)];
                      reg545 <= $signed(forvar423[(4'h9):(3'h5)]);
                    end
                  else
                    begin
                      reg543 <= $unsigned(reg295);
                      reg544 <= reg502[(3'h6):(3'h6)];
                    end
                  for (forvar546 = (1'h0); (forvar546 < (1'h1)); forvar546 = (forvar546 + (1'h1)))
                    begin
                      reg547 <= (reg374 ? reg423 : (&(-(~|reg358))));
                      reg548 <= ($signed((8'hb7)) ?
                          (&reg394[(1'h0):(1'h0)]) : (!($unsigned((8'ha6)) ?
                              $unsigned(reg325) : {reg392})));
                    end
                end
            end
          for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
            begin
              for (forvar550 = (1'h0); (forvar550 < (1'h0)); forvar550 = (forvar550 + (1'h1)))
                begin
                  for (forvar551 = (1'h0); (forvar551 < (2'h3)); forvar551 = (forvar551 + (1'h1)))
                    begin
                      reg552 <= $signed($signed($unsigned({(8'ha0)})));
                      reg553 <= forvar471;
                    end
                end
              if ($signed((((forvar260 ? reg330 : reg329) ?
                      reg455[(3'h6):(3'h4)] : (reg353 <<< reg334)) ?
                  (~&reg330) : ($unsigned(forvar551) ? (|(8'ha4)) : {reg240}))))
                begin
                  if (($unsigned((^$unsigned((8'haf)))) > {reg251[(2'h2):(1'h1)]}))
                    begin
                      reg554 <= (($signed((forvar350 ? reg505 : forvar428)) ?
                              ($unsigned(reg242) <<< $signed(forvar260)) : $signed($signed(forvar386))) ?
                          (~((reg256 ?
                              reg259 : reg504) | reg346)) : $signed((^~reg221)));
                    end
                  else
                    begin
                      reg554 <= {((reg266[(3'h6):(2'h2)] ?
                                  (+reg341) : forvar354[(1'h1):(1'h0)]) ?
                              (+$signed((8'hb5))) : ((reg236 < reg364) ?
                                  reg327[(1'h1):(1'h1)] : {(8'haf)}))};
                      reg555 <= reg287;
                    end
                  reg556 <= ({$signed($signed((8'ha4)))} || $unsigned(($unsigned(reg323) ^~ ((8'ha8) ?
                      reg529 : (8'hb2)))));
                  if (($unsigned((reg382 ?
                      (8'hae) : (8'ha8))) >> {reg487[(4'hb):(1'h1)]}))
                    begin
                      reg557 <= reg467;
                      reg558 <= (~&(!(reg374[(4'hf):(1'h1)] >= (~|reg523))));
                      reg559 <= {$unsigned($signed($unsigned(forvar403)))};
                      reg560 <= reg456[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg557 <= $unsigned((reg246 ?
                          $unsigned((|reg384)) : {$unsigned((8'hb8))}));
                      reg558 <= forvar277[(4'hb):(2'h3)];
                      reg559 <= $signed($unsigned((8'had)));
                    end
                  for (forvar561 = (1'h0); (forvar561 < (2'h2)); forvar561 = (forvar561 + (1'h1)))
                    begin
                      reg562 <= ($signed(reg322) < {$signed($signed(reg404))});
                      reg563 <= forvar344[(3'h6):(3'h6)];
                    end
                end
              else
                begin
                  for (forvar554 = (1'h0); (forvar554 < (2'h2)); forvar554 = (forvar554 + (1'h1)))
                    begin
                      reg555 <= $signed({reg307});
                    end
                  for (forvar556 = (1'h0); (forvar556 < (1'h0)); forvar556 = (forvar556 + (1'h1)))
                    begin
                      reg557 <= ($signed((&(forvar503 ?
                          forvar272 : reg483))) > ($signed($signed(reg294)) ?
                          ((reg420 >> reg380) ?
                              ((8'haa) ? (8'ha4) : reg367) : (reg263 ?
                                  reg499 : reg352)) : $unsigned($unsigned(forvar340))));
                      reg558 <= (~^(+($unsigned(reg362) ?
                          forvar484[(3'h6):(2'h2)] : reg349)));
                    end
                  reg559 <= (~^$signed(($signed(reg253) ?
                      reg338 : $unsigned(reg250))));
                end
            end
        end
    end
  assign wire564 = (($unsigned((&reg371)) >>> {(~&(8'h9e))}) ?
                       (+($unsigned(reg467) * $unsigned(reg423))) : forvar445);
  assign wire565 = {(^($unsigned(forvar342) ?
                           {reg490} : reg280[(1'h0):(1'h0)]))};
  assign wire566 = {$unsigned((!reg545))};
  assign wire567 = ($signed($unsigned(reg465[(2'h2):(2'h2)])) ?
                       (reg367 & (((8'haa) ? reg512 : reg421) ?
                           forvar341 : reg446)) : $signed(reg506[(1'h0):(1'h0)]));
  assign wire568 = ($signed($signed($signed(reg350))) | $signed(($unsigned(wire217) ~^ $signed((8'hb2)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module641
#( parameter param4145 = (({(^(8'hac))} ? (((8'hb8) ? (8'ha3) : (8'hb8)) || {(8'hab)}) : {(^(8'haf))}) > ((((8'ha4) ? (8'ha0) : (8'hb6)) ? {(8'hb5)} : ((8'hab) << (8'hb4))) > ((~(8'ha0)) ? ((8'ha1) ? (8'ha6) : (8'hb1)) : ((8'h9e) >>> (8'hb6))))) )
(y, clk, wire645, wire644, wire643, wire642);
  output wire [(32'ha33):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire645;
  input wire [(4'h8):(1'h0)] wire644;
  input wire [(4'he):(1'h0)] wire643;
  input wire signed [(4'h8):(1'h0)] wire642;
  wire signed [(4'he):(1'h0)] wire4144;
  wire signed [(4'hd):(1'h0)] wire4143;
  reg signed [(4'hc):(1'h0)] reg4142 = (1'h0);
  reg [(3'h5):(1'h0)] reg4122 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4119 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4117 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4116 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4112 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4111 = (1'h0);
  reg [(4'hf):(1'h0)] reg4110 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4108 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4106 = (1'h0);
  reg [(3'h7):(1'h0)] reg4105 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4102 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4099 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4095 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4092 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4088 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4141 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4140 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4127 = (1'h0);
  reg [(4'h9):(1'h0)] reg4139 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4138 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4137 = (1'h0);
  reg [(3'h4):(1'h0)] reg4136 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4135 = (1'h0);
  reg [(4'ha):(1'h0)] reg4134 = (1'h0);
  reg [(4'hc):(1'h0)] reg4133 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4132 = (1'h0);
  reg [(2'h2):(1'h0)] reg4131 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4130 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4129 = (1'h0);
  reg [(4'h9):(1'h0)] reg4128 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4127 = (1'h0);
  reg [(4'h8):(1'h0)] reg4126 = (1'h0);
  reg [(2'h2):(1'h0)] reg4125 = (1'h0);
  reg [(4'he):(1'h0)] reg4124 = (1'h0);
  reg [(3'h4):(1'h0)] reg4123 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4122 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4121 = (1'h0);
  reg [(4'hc):(1'h0)] reg4120 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4119 = (1'h0);
  reg [(3'h7):(1'h0)] reg4118 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4117 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4116 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4115 = (1'h0);
  reg [(3'h6):(1'h0)] reg4114 = (1'h0);
  reg [(3'h7):(1'h0)] reg4113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4112 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4111 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4110 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4109 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4108 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4107 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4106 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4105 = (1'h0);
  reg [(4'ha):(1'h0)] reg4104 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4103 = (1'h0);
  reg [(4'hc):(1'h0)] reg4102 = (1'h0);
  reg [(3'h7):(1'h0)] reg4101 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4089 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4100 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4099 = (1'h0);
  reg [(3'h7):(1'h0)] reg4098 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4097 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4096 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4095 = (1'h0);
  reg [(3'h6):(1'h0)] reg4094 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4093 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4092 = (1'h0);
  reg [(4'he):(1'h0)] reg4091 = (1'h0);
  reg [(2'h2):(1'h0)] reg4090 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4089 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4088 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4087 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire4086;
  reg signed [(3'h6):(1'h0)] reg4085 = (1'h0);
  reg [(3'h5):(1'h0)] reg4084 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4083 = (1'h0);
  reg [(4'hb):(1'h0)] reg4082 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4081 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4078 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4080 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4079 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4078 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4077 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4076 = (1'h0);
  reg [(4'hc):(1'h0)] reg4075 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4074 = (1'h0);
  reg [(4'he):(1'h0)] reg4073 = (1'h0);
  reg [(4'h8):(1'h0)] reg4072 = (1'h0);
  reg [(4'h9):(1'h0)] reg4071 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4070 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4069 = (1'h0);
  reg [(4'hc):(1'h0)] reg4065 = (1'h0);
  reg [(2'h2):(1'h0)] reg4068 = (1'h0);
  reg [(4'ha):(1'h0)] reg4067 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4066 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4065 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4064 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4063 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4062 = (1'h0);
  reg [(3'h6):(1'h0)] reg4061 = (1'h0);
  reg [(4'ha):(1'h0)] reg4060 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4059 = (1'h0);
  reg [(3'h5):(1'h0)] reg4058 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4054 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4051 = (1'h0);
  reg [(3'h6):(1'h0)] reg4050 = (1'h0);
  reg [(4'h9):(1'h0)] reg4057 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4056 = (1'h0);
  reg [(4'hb):(1'h0)] reg4055 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4054 = (1'h0);
  reg [(4'h9):(1'h0)] reg4053 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4052 = (1'h0);
  reg [(4'hd):(1'h0)] reg4051 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4050 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4049 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4048 = (1'h0);
  reg [(4'he):(1'h0)] forvar4047 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4046 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4036 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4030 = (1'h0);
  reg [(4'h8):(1'h0)] reg4025 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4024 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4022 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4018 = (1'h0);
  reg [(2'h3):(1'h0)] reg4045 = (1'h0);
  reg [(4'h9):(1'h0)] reg4044 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4043 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4042 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4041 = (1'h0);
  reg [(3'h4):(1'h0)] reg4040 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4039 = (1'h0);
  reg [(3'h4):(1'h0)] reg4038 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4037 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4036 = (1'h0);
  reg [(4'h9):(1'h0)] reg4035 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4034 = (1'h0);
  reg [(3'h7):(1'h0)] reg4033 = (1'h0);
  reg [(4'h8):(1'h0)] reg4032 = (1'h0);
  reg [(3'h6):(1'h0)] reg4031 = (1'h0);
  reg [(4'he):(1'h0)] forvar4030 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4029 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4028 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4027 = (1'h0);
  reg [(5'h10):(1'h0)] reg4026 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4025 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4024 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4020 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4023 = (1'h0);
  reg [(4'hc):(1'h0)] reg4022 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4021 = (1'h0);
  reg [(4'hf):(1'h0)] reg4020 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4019 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4018 = (1'h0);
  reg [(4'hf):(1'h0)] reg4017 = (1'h0);
  reg [(4'ha):(1'h0)] reg4016 = (1'h0);
  reg [(3'h4):(1'h0)] reg4015 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4012 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4011 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4009 = (1'h0);
  reg [(5'h10):(1'h0)] reg4014 = (1'h0);
  reg [(3'h6):(1'h0)] reg4013 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4012 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4011 = (1'h0);
  reg [(2'h2):(1'h0)] reg4010 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4009 = (1'h0);
  reg [(4'hb):(1'h0)] reg4005 = (1'h0);
  reg [(4'h9):(1'h0)] reg4008 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4007 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4006 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4005 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4004 = (1'h0);
  reg [(3'h4):(1'h0)] reg4001 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4003 = (1'h0);
  reg [(4'hf):(1'h0)] reg4002 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4001 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4000 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3999 = (1'h0);
  wire [(4'hf):(1'h0)] wire3998;
  wire [(4'hc):(1'h0)] wire3996;
  wire signed [(4'he):(1'h0)] wire1056;
  wire [(4'he):(1'h0)] wire646;
  wire [(4'ha):(1'h0)] wire1058;
  reg [(4'ha):(1'h0)] forvar1059 = (1'h0);
  reg [(4'hd):(1'h0)] reg1060 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1060 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1061 = (1'h0);
  reg [(3'h6):(1'h0)] reg1062 = (1'h0);
  reg [(4'h8):(1'h0)] reg1063 = (1'h0);
  reg [(4'hb):(1'h0)] reg1064 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1065 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1066 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1067 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1068 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1069 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1070 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1071 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1072 = (1'h0);
  reg [(4'ha):(1'h0)] reg1073 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1074 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1070 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1075 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1076 = (1'h0);
  reg [(4'he):(1'h0)] reg1077 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1078 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1079 = (1'h0);
  reg [(4'hc):(1'h0)] reg1080 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1081 = (1'h0);
  reg [(4'h8):(1'h0)] reg1082 = (1'h0);
  reg [(2'h2):(1'h0)] reg1083 = (1'h0);
  reg [(4'hc):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1085 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1086 = (1'h0);
  reg [(3'h6):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1088 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1089 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1090 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1091 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1092 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1093 = (1'h0);
  reg [(3'h4):(1'h0)] reg1094 = (1'h0);
  reg [(4'he):(1'h0)] forvar1095 = (1'h0);
  reg [(4'hb):(1'h0)] reg1096 = (1'h0);
  reg [(4'hc):(1'h0)] reg1097 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1098 = (1'h0);
  reg [(5'h10):(1'h0)] reg1099 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1100 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1101 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1102 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1103 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1104 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1105 = (1'h0);
  reg [(3'h4):(1'h0)] reg1106 = (1'h0);
  reg [(4'hd):(1'h0)] reg1107 = (1'h0);
  reg [(3'h5):(1'h0)] reg1108 = (1'h0);
  reg [(4'hc):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1110 = (1'h0);
  reg [(3'h5):(1'h0)] reg1111 = (1'h0);
  reg [(4'hf):(1'h0)] reg1112 = (1'h0);
  reg [(4'h8):(1'h0)] reg1113 = (1'h0);
  reg [(4'hb):(1'h0)] reg1114 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1103 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1104 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1105 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1107 = (1'h0);
  reg [(4'he):(1'h0)] forvar1115 = (1'h0);
  reg [(3'h4):(1'h0)] reg1116 = (1'h0);
  reg [(2'h2):(1'h0)] reg1117 = (1'h0);
  reg [(4'h8):(1'h0)] reg1118 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1119 = (1'h0);
  reg [(3'h6):(1'h0)] reg1120 = (1'h0);
  reg [(4'hd):(1'h0)] reg1121 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1122 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1123 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1124 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1125 = (1'h0);
  reg [(4'hf):(1'h0)] reg1126 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1127 = (1'h0);
  reg [(3'h6):(1'h0)] reg1128 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1129 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1130 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1131 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1132 = (1'h0);
  reg [(4'ha):(1'h0)] reg1133 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1134 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1135 = (1'h0);
  reg [(4'he):(1'h0)] reg1136 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1137 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1138 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1139 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1141 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1142 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1143 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1144 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1145 = (1'h0);
  reg [(4'ha):(1'h0)] reg1146 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1147 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1148 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1149 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1150 = (1'h0);
  reg [(2'h2):(1'h0)] reg1151 = (1'h0);
  wire [(5'h10):(1'h0)] wire1152;
  wire [(4'hd):(1'h0)] wire3994;
  assign y = {wire4144,
                 wire4143,
                 reg4142,
                 reg4122,
                 reg4119,
                 forvar4117,
                 forvar4116,
                 forvar4112,
                 forvar4111,
                 reg4110,
                 reg4108,
                 forvar4106,
                 reg4105,
                 forvar4102,
                 forvar4099,
                 forvar4095,
                 forvar4092,
                 reg4088,
                 reg4141,
                 reg4140,
                 reg4127,
                 reg4139,
                 reg4138,
                 reg4137,
                 reg4136,
                 forvar4135,
                 reg4134,
                 reg4133,
                 forvar4132,
                 reg4131,
                 reg4130,
                 reg4129,
                 reg4128,
                 forvar4127,
                 reg4126,
                 reg4125,
                 reg4124,
                 reg4123,
                 forvar4122,
                 reg4121,
                 reg4120,
                 forvar4119,
                 reg4118,
                 reg4117,
                 reg4116,
                 reg4115,
                 reg4114,
                 reg4113,
                 reg4112,
                 reg4111,
                 forvar4110,
                 reg4109,
                 forvar4108,
                 reg4107,
                 reg4106,
                 forvar4105,
                 reg4104,
                 reg4103,
                 reg4102,
                 reg4101,
                 reg4089,
                 reg4100,
                 reg4099,
                 reg4098,
                 forvar4097,
                 reg4096,
                 reg4095,
                 reg4094,
                 reg4093,
                 reg4092,
                 reg4091,
                 reg4090,
                 forvar4089,
                 forvar4088,
                 reg4087,
                 wire4086,
                 reg4085,
                 reg4084,
                 reg4083,
                 reg4082,
                 reg4081,
                 forvar4078,
                 reg4080,
                 reg4079,
                 reg4078,
                 reg4077,
                 reg4076,
                 reg4075,
                 reg4074,
                 reg4073,
                 reg4072,
                 reg4071,
                 reg4070,
                 forvar4069,
                 reg4065,
                 reg4068,
                 reg4067,
                 reg4066,
                 forvar4065,
                 reg4064,
                 reg4063,
                 reg4062,
                 reg4061,
                 reg4060,
                 reg4059,
                 reg4058,
                 reg4054,
                 forvar4051,
                 reg4050,
                 reg4057,
                 reg4056,
                 reg4055,
                 forvar4054,
                 reg4053,
                 reg4052,
                 reg4051,
                 forvar4050,
                 reg4049,
                 forvar4048,
                 forvar4047,
                 forvar4046,
                 reg4036,
                 reg4030,
                 reg4025,
                 forvar4024,
                 forvar4022,
                 forvar4018,
                 reg4045,
                 reg4044,
                 reg4043,
                 reg4042,
                 forvar4041,
                 reg4040,
                 reg4039,
                 reg4038,
                 reg4037,
                 forvar4036,
                 reg4035,
                 reg4034,
                 reg4033,
                 reg4032,
                 reg4031,
                 forvar4030,
                 forvar4029,
                 reg4028,
                 reg4027,
                 reg4026,
                 forvar4025,
                 reg4024,
                 forvar4020,
                 reg4023,
                 reg4022,
                 reg4021,
                 reg4020,
                 reg4019,
                 reg4018,
                 reg4017,
                 reg4016,
                 reg4015,
                 reg4012,
                 forvar4011,
                 forvar4009,
                 reg4014,
                 reg4013,
                 forvar4012,
                 reg4011,
                 reg4010,
                 reg4009,
                 reg4005,
                 reg4008,
                 reg4007,
                 reg4006,
                 forvar4005,
                 reg4004,
                 reg4001,
                 reg4003,
                 reg4002,
                 forvar4001,
                 forvar4000,
                 forvar3999,
                 wire3998,
                 wire3996,
                 wire1056,
                 wire646,
                 wire1058,
                 forvar1059,
                 reg1060,
                 forvar1060,
                 reg1061,
                 reg1062,
                 reg1063,
                 reg1064,
                 reg1065,
                 reg1066,
                 reg1067,
                 reg1068,
                 forvar1069,
                 forvar1070,
                 reg1071,
                 reg1072,
                 reg1073,
                 reg1074,
                 reg1070,
                 forvar1075,
                 reg1076,
                 reg1077,
                 reg1078,
                 forvar1079,
                 reg1080,
                 reg1081,
                 reg1082,
                 reg1083,
                 reg1084,
                 reg1085,
                 reg1086,
                 reg1087,
                 reg1088,
                 reg1089,
                 forvar1090,
                 forvar1091,
                 forvar1092,
                 reg1093,
                 reg1094,
                 forvar1095,
                 reg1096,
                 reg1097,
                 reg1098,
                 reg1099,
                 reg1100,
                 reg1101,
                 forvar1102,
                 reg1103,
                 forvar1104,
                 reg1105,
                 reg1106,
                 reg1107,
                 reg1108,
                 reg1109,
                 reg1110,
                 reg1111,
                 reg1112,
                 reg1113,
                 reg1114,
                 forvar1103,
                 reg1104,
                 forvar1105,
                 forvar1107,
                 forvar1115,
                 reg1116,
                 reg1117,
                 reg1118,
                 forvar1119,
                 reg1120,
                 reg1121,
                 forvar1122,
                 reg1123,
                 reg1124,
                 reg1125,
                 reg1126,
                 reg1127,
                 reg1128,
                 reg1129,
                 forvar1130,
                 forvar1131,
                 forvar1132,
                 reg1133,
                 reg1134,
                 reg1135,
                 reg1136,
                 reg1137,
                 forvar1138,
                 reg1139,
                 reg1140,
                 reg1141,
                 forvar1142,
                 reg1143,
                 reg1144,
                 forvar1145,
                 reg1146,
                 reg1147,
                 reg1148,
                 reg1149,
                 reg1150,
                 reg1151,
                 wire1152,
                 wire3994,
                 (1'h0)};
  assign wire646 = ($signed(($signed(wire645) * (wire645 > wire643))) ?
                       wire642[(3'h6):(2'h3)] : wire643);
  module647 modinst1057 (.clk(clk), .wire649(wire646), .wire648(wire643), .wire650(wire644), .wire652(wire642), .y(wire1056), .wire651(wire645));
  assign wire1058 = wire1056[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar1059 = (1'h0); (forvar1059 < (1'h0)); forvar1059 = (forvar1059 + (1'h1)))
        begin
          if ($signed(($unsigned((-(8'h9f))) >= (wire1058[(3'h7):(2'h2)] << {wire1058}))))
            begin
              reg1060 <= wire646[(3'h4):(2'h3)];
            end
          else
            begin
              for (forvar1060 = (1'h0); (forvar1060 < (1'h1)); forvar1060 = (forvar1060 + (1'h1)))
                begin
                  if ($signed(wire646))
                    begin
                      reg1061 <= $unsigned(({$signed((8'hb3))} ~^ (wire643[(1'h1):(1'h0)] ?
                          (wire643 ? wire642 : wire645) : $unsigned(reg1060))));
                      reg1062 <= (wire1056 ^~ $unsigned($unsigned($signed(wire1056))));
                      reg1063 <= (!reg1060);
                      reg1064 <= (((forvar1059 && $unsigned(wire643)) ?
                              $signed((~&wire644)) : wire645[(1'h0):(1'h0)]) ?
                          {($unsigned(reg1061) ?
                                  (reg1063 - wire646) : (reg1061 ?
                                      wire643 : (8'hab)))} : (8'ha2));
                    end
                  else
                    begin
                      reg1061 <= (8'hb7);
                    end
                  if (($unsigned($unsigned((-reg1063))) ?
                      (+forvar1059) : wire1056))
                    begin
                      reg1065 <= (~^$unsigned(forvar1059[(1'h0):(1'h0)]));
                      reg1066 <= $unsigned((8'ha3));
                      reg1067 <= $unsigned($unsigned(reg1066));
                    end
                  else
                    begin
                      reg1065 <= reg1064;
                    end
                end
              reg1068 <= (~^(|{$unsigned((8'h9f))}));
            end
          for (forvar1069 = (1'h0); (forvar1069 < (1'h1)); forvar1069 = (forvar1069 + (1'h1)))
            begin
              if ((~forvar1059))
                begin
                  for (forvar1070 = (1'h0); (forvar1070 < (2'h2)); forvar1070 = (forvar1070 + (1'h1)))
                    begin
                      reg1071 <= $signed(reg1066);
                    end
                  if ({(($unsigned(wire644) >> wire642[(3'h4):(1'h1)]) ?
                          (8'ha1) : reg1062)})
                    begin
                      reg1072 <= $signed((~|reg1067[(2'h3):(2'h3)]));
                      reg1073 <= reg1061[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg1072 <= $unsigned((8'hb3));
                      reg1073 <= (8'hab);
                      reg1074 <= reg1073[(3'h4):(2'h3)];
                    end
                end
              else
                begin
                  if ((|$signed($signed({forvar1059}))))
                    begin
                      reg1070 <= {($signed(reg1068) ?
                              (&(^~reg1061)) : ($unsigned(wire645) ?
                                  (wire643 >> forvar1059) : {wire643}))};
                      reg1071 <= reg1070;
                      reg1072 <= ((^~((wire646 + reg1072) ?
                          (reg1073 ?
                              reg1072 : forvar1069) : (-wire646))) ^ (^~reg1062[(3'h4):(3'h4)]));
                    end
                  else
                    begin
                      reg1070 <= (-($signed(forvar1060) > ((&reg1073) ?
                          forvar1070[(1'h0):(1'h0)] : wire645)));
                      reg1071 <= $signed(forvar1059);
                    end
                end
              for (forvar1075 = (1'h0); (forvar1075 < (1'h1)); forvar1075 = (forvar1075 + (1'h1)))
                begin
                  if (((~|($unsigned(wire1058) <= ((8'hb5) ?
                          reg1066 : forvar1059))) ?
                      $signed($signed(forvar1070)) : reg1073[(2'h2):(1'h1)]))
                    begin
                      reg1076 <= wire1056[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1076 <= (+(reg1062 > ({wire644} * $unsigned(wire643))));
                      reg1077 <= ($signed($signed(((8'h9e) ?
                              (8'hae) : reg1076))) ?
                          reg1068 : {forvar1059});
                    end
                  if ($unsigned({reg1071[(3'h5):(2'h3)]}))
                    begin
                      reg1078 <= forvar1075[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg1078 <= ($signed($unsigned($unsigned(wire1056))) & (^(&(~&reg1073))));
                    end
                end
              for (forvar1079 = (1'h0); (forvar1079 < (1'h1)); forvar1079 = (forvar1079 + (1'h1)))
                begin
                  if ({reg1063})
                    begin
                      reg1080 <= $signed($unsigned($signed((reg1062 ?
                          reg1065 : reg1067))));
                      reg1081 <= forvar1070;
                      reg1082 <= reg1081[(4'hc):(1'h0)];
                      reg1083 <= (~^$unsigned((8'h9c)));
                    end
                  else
                    begin
                      reg1080 <= reg1062;
                      reg1081 <= reg1065[(1'h1):(1'h0)];
                      reg1082 <= $signed(reg1071[(1'h0):(1'h0)]);
                      reg1083 <= $unsigned($signed((-$unsigned(reg1068))));
                    end
                  if (reg1065[(1'h1):(1'h0)])
                    begin
                      reg1084 <= (^{((forvar1059 ? reg1074 : reg1063) ?
                              (reg1068 > forvar1069) : (reg1074 ?
                                  (8'h9e) : forvar1079))});
                      reg1085 <= $unsigned(((|((8'had) ? reg1072 : (8'h9c))) ?
                          (8'hb4) : ({reg1072} >>> (~^wire645))));
                    end
                  else
                    begin
                      reg1084 <= (~|$signed((reg1077[(3'h7):(1'h0)] ^~ (8'hb6))));
                      reg1085 <= $unsigned(($signed($unsigned(reg1078)) ?
                          ((^reg1085) * $signed(reg1081)) : ((8'hb8) ?
                              $signed(forvar1059) : (reg1070 != reg1078))));
                    end
                  if (($signed((~reg1061[(4'hb):(4'h8)])) ?
                      $signed(((&(8'had)) ?
                          (!wire645) : reg1076[(2'h2):(1'h1)])) : ((~&(~^reg1071)) >> ((forvar1069 ?
                          reg1074 : wire644) ^ reg1064))))
                    begin
                      reg1086 <= $unsigned($unsigned(forvar1069[(3'h5):(3'h4)]));
                      reg1087 <= ($signed(reg1086) ?
                          $signed((^~{reg1073})) : (!(|forvar1070)));
                      reg1088 <= reg1070[(2'h3):(1'h1)];
                      reg1089 <= $signed({(reg1062[(3'h4):(1'h0)] ?
                              (reg1084 ? (8'had) : (8'h9d)) : {(8'haf)})});
                    end
                  else
                    begin
                      reg1086 <= ({reg1083} ?
                          (forvar1075 ?
                              (^~(reg1061 + (8'ha4))) : (~&$unsigned(wire646))) : reg1062[(3'h4):(2'h2)]);
                      reg1087 <= $signed(((!(wire646 ? reg1062 : (8'h9c))) ?
                          $unsigned(((8'haf) < reg1064)) : forvar1070[(2'h3):(1'h0)]));
                      reg1088 <= reg1068[(3'h5):(2'h2)];
                      reg1089 <= $unsigned(({(-reg1066)} <<< (wire644[(1'h0):(1'h0)] ?
                          (reg1063 << wire644) : $unsigned(reg1067))));
                    end
                end
            end
          for (forvar1090 = (1'h0); (forvar1090 < (2'h3)); forvar1090 = (forvar1090 + (1'h1)))
            begin
              for (forvar1091 = (1'h0); (forvar1091 < (2'h3)); forvar1091 = (forvar1091 + (1'h1)))
                begin
                  for (forvar1092 = (1'h0); (forvar1092 < (2'h3)); forvar1092 = (forvar1092 + (1'h1)))
                    begin
                      reg1093 <= reg1071;
                      reg1094 <= (~^forvar1075[(1'h0):(1'h0)]);
                    end
                  for (forvar1095 = (1'h0); (forvar1095 < (2'h2)); forvar1095 = (forvar1095 + (1'h1)))
                    begin
                      reg1096 <= (((|(wire1056 ? (8'ha9) : wire643)) ?
                          $unsigned(forvar1095) : ({reg1078} ^~ (~^reg1089))) ^ $signed($signed((~^forvar1091))));
                    end
                  if ($signed(reg1089))
                    begin
                      reg1097 <= ($unsigned((~&reg1080[(3'h7):(3'h4)])) ?
                          (forvar1069[(3'h6):(3'h5)] ?
                              reg1096[(4'hb):(3'h7)] : $signed((8'ha7))) : reg1067);
                      reg1098 <= reg1081;
                      reg1099 <= $unsigned(reg1088[(4'h8):(3'h7)]);
                      reg1100 <= reg1098;
                    end
                  else
                    begin
                      reg1097 <= reg1097[(3'h7):(3'h4)];
                      reg1098 <= reg1064[(1'h0):(1'h0)];
                      reg1099 <= reg1063[(3'h4):(2'h2)];
                      reg1100 <= {(^$unsigned(reg1067[(2'h3):(2'h3)]))};
                    end
                  reg1101 <= $unsigned(wire1056);
                end
            end
        end
      for (forvar1102 = (1'h0); (forvar1102 < (1'h0)); forvar1102 = (forvar1102 + (1'h1)))
        begin
          if (reg1074[(1'h1):(1'h0)])
            begin
              reg1103 <= wire646;
              for (forvar1104 = (1'h0); (forvar1104 < (1'h1)); forvar1104 = (forvar1104 + (1'h1)))
                begin
                  if ($unsigned(reg1100))
                    begin
                      reg1105 <= $signed(forvar1060);
                    end
                  else
                    begin
                      reg1105 <= {$signed({(forvar1075 * forvar1090)})};
                      reg1106 <= $signed((&$unsigned($unsigned(reg1068))));
                      reg1107 <= {forvar1090[(4'h9):(3'h4)]};
                      reg1108 <= $unsigned(forvar1104);
                    end
                  if ((((forvar1095 > (~|reg1105)) ?
                          ($unsigned(reg1105) && (reg1107 == forvar1059)) : reg1101) ?
                      (reg1093 ? forvar1092 : (|$unsigned(reg1107))) : reg1077))
                    begin
                      reg1109 <= $unsigned($unsigned(reg1101));
                      reg1110 <= {($signed((^reg1080)) ?
                              (^~reg1086) : ({reg1074} && $unsigned(reg1097)))};
                      reg1111 <= reg1107;
                    end
                  else
                    begin
                      reg1109 <= forvar1075[(1'h1):(1'h1)];
                    end
                  if (reg1062)
                    begin
                      reg1112 <= $unsigned(forvar1059);
                      reg1113 <= (&{$signed(((8'hba) ? reg1082 : reg1072))});
                      reg1114 <= (8'h9c);
                    end
                  else
                    begin
                      reg1112 <= ($unsigned((forvar1070[(3'h4):(1'h1)] ?
                              {reg1071} : $signed((8'haa)))) ?
                          {$signed($signed(reg1066))} : reg1093);
                      reg1113 <= reg1081;
                      reg1114 <= ((~^(+wire643[(4'h8):(3'h7)])) ?
                          ((reg1106[(1'h1):(1'h1)] == (wire643 < reg1096)) << {(~^forvar1095)}) : (~&(reg1113 <<< (~&(8'haf)))));
                    end
                end
            end
          else
            begin
              for (forvar1103 = (1'h0); (forvar1103 < (2'h2)); forvar1103 = (forvar1103 + (1'h1)))
                begin
                  reg1104 <= reg1088;
                end
              if ($unsigned(reg1062))
                begin
                  for (forvar1105 = (1'h0); (forvar1105 < (2'h3)); forvar1105 = (forvar1105 + (1'h1)))
                    begin
                      reg1106 <= ((reg1080 & ((8'ha9) != (forvar1103 | reg1089))) ?
                          ($signed($signed(reg1093)) ?
                              (forvar1079 <<< {forvar1075}) : wire646[(3'h5):(3'h4)]) : ($unsigned(forvar1091) - forvar1091));
                    end
                  for (forvar1107 = (1'h0); (forvar1107 < (1'h0)); forvar1107 = (forvar1107 + (1'h1)))
                    begin
                      reg1108 <= ((~&$signed($signed(reg1083))) >= (((!forvar1059) > $signed(reg1098)) << reg1072[(3'h4):(2'h3)]));
                      reg1109 <= $signed((+forvar1102));
                      reg1110 <= {({(reg1109 > reg1113)} ?
                              ({reg1063} ?
                                  (reg1081 ~^ reg1082) : reg1107) : (&$unsigned(reg1110)))};
                      reg1111 <= {$signed((-$unsigned(reg1070)))};
                    end
                  if ((&reg1078[(4'h9):(3'h7)]))
                    begin
                      reg1112 <= {({(wire643 ~^ reg1113)} | ({(8'hb0)} ?
                              reg1061 : (reg1064 ? reg1060 : reg1098)))};
                      reg1113 <= reg1101;
                      reg1114 <= (forvar1107[(2'h2):(2'h2)] * $signed(((reg1097 ?
                          forvar1075 : reg1082) == reg1063[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg1112 <= forvar1107[(3'h4):(2'h2)];
                      reg1113 <= {$unsigned(forvar1104)};
                      reg1114 <= {{(reg1071 ?
                                  (~^wire646) : $unsigned(wire1058))}};
                    end
                  for (forvar1115 = (1'h0); (forvar1115 < (1'h0)); forvar1115 = (forvar1115 + (1'h1)))
                    begin
                      reg1116 <= (8'h9d);
                      reg1117 <= wire646[(2'h2):(2'h2)];
                      reg1118 <= $signed(reg1061[(2'h3):(1'h0)]);
                    end
                end
              else
                begin
                  reg1105 <= forvar1105[(2'h2):(2'h2)];
                end
              for (forvar1119 = (1'h0); (forvar1119 < (2'h3)); forvar1119 = (forvar1119 + (1'h1)))
                begin
                  reg1120 <= forvar1059;
                  reg1121 <= ($unsigned({$signed(forvar1060)}) != (reg1073 ?
                      forvar1069 : forvar1119));
                end
              for (forvar1122 = (1'h0); (forvar1122 < (1'h1)); forvar1122 = (forvar1122 + (1'h1)))
                begin
                  if (($unsigned(wire1056) ?
                      $unsigned(reg1081) : {$signed($signed(forvar1104))}))
                    begin
                      reg1123 <= (reg1078 ?
                          ((~wire1056) ~^ ((forvar1070 ? reg1088 : reg1116) ?
                              $signed(forvar1122) : reg1080)) : $signed(reg1078[(4'h8):(3'h5)]));
                    end
                  else
                    begin
                      reg1123 <= (^forvar1102[(3'h4):(1'h0)]);
                      reg1124 <= $signed($unsigned(reg1106));
                      reg1125 <= reg1068[(3'h5):(2'h3)];
                    end
                  if ((8'hb0))
                    begin
                      reg1126 <= reg1062[(3'h5):(1'h0)];
                      reg1127 <= {(((reg1083 ? reg1084 : reg1116) ?
                              (forvar1090 == reg1072) : $signed(wire644)) >= $signed((reg1089 ?
                              (8'hab) : reg1088)))};
                    end
                  else
                    begin
                      reg1126 <= ((($unsigned(reg1105) << (forvar1115 ?
                              reg1120 : reg1070)) ?
                          {{reg1064}} : reg1121[(3'h4):(1'h1)]) | $unsigned({$unsigned(forvar1119)}));
                      reg1127 <= $signed(($signed((reg1082 < (8'ha3))) >= $signed($unsigned(forvar1095))));
                      reg1128 <= ((~^$unsigned(reg1073)) ?
                          {$signed((~reg1127))} : reg1074);
                      reg1129 <= reg1117[(1'h1):(1'h0)];
                    end
                end
            end
          for (forvar1130 = (1'h0); (forvar1130 < (1'h1)); forvar1130 = (forvar1130 + (1'h1)))
            begin
              for (forvar1131 = (1'h0); (forvar1131 < (2'h2)); forvar1131 = (forvar1131 + (1'h1)))
                begin
                  for (forvar1132 = (1'h0); (forvar1132 < (1'h0)); forvar1132 = (forvar1132 + (1'h1)))
                    begin
                      reg1133 <= reg1128[(1'h1):(1'h1)];
                    end
                  if ((~&{(~^$signed(reg1080))}))
                    begin
                      reg1134 <= (|$signed($signed($unsigned(reg1113))));
                      reg1135 <= {reg1120[(3'h6):(3'h4)]};
                      reg1136 <= reg1129[(2'h3):(1'h0)];
                      reg1137 <= wire643[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg1134 <= $unsigned(((forvar1107[(1'h0):(1'h0)] ?
                          (reg1114 & reg1100) : (-reg1089)) ~^ wire1056[(4'h8):(2'h2)]));
                    end
                  for (forvar1138 = (1'h0); (forvar1138 < (1'h1)); forvar1138 = (forvar1138 + (1'h1)))
                    begin
                      reg1139 <= ($unsigned(reg1129[(3'h5):(1'h1)]) <= (((reg1068 <= forvar1090) ?
                          forvar1105 : (reg1080 ?
                              reg1084 : reg1087)) ^~ $signed((reg1078 >> reg1062))));
                      reg1140 <= ((reg1127 ?
                              {$signed((8'had))} : $signed(reg1124)) ?
                          (&($unsigned(reg1127) ?
                              (reg1113 ?
                                  reg1121 : forvar1079) : (+wire645))) : (~|(8'h9e)));
                      reg1141 <= {(~|reg1112)};
                    end
                end
              for (forvar1142 = (1'h0); (forvar1142 < (1'h0)); forvar1142 = (forvar1142 + (1'h1)))
                begin
                  reg1143 <= $unsigned((~$signed($signed(reg1082))));
                  reg1144 <= reg1125;
                  for (forvar1145 = (1'h0); (forvar1145 < (1'h0)); forvar1145 = (forvar1145 + (1'h1)))
                    begin
                      reg1146 <= $unsigned((reg1071[(2'h2):(2'h2)] ?
                          {$signed(reg1141)} : ((reg1110 ?
                              reg1067 : (8'hb8)) == $signed(reg1093))));
                      reg1147 <= $signed(((reg1128 ?
                          (forvar1059 ^ (8'hb9)) : {(8'haa)}) * $signed({reg1124})));
                      reg1148 <= $unsigned((reg1068 ?
                          forvar1075 : {$signed(reg1121)}));
                      reg1149 <= (~&reg1084);
                    end
                end
            end
          reg1150 <= forvar1070[(2'h3):(1'h1)];
        end
      reg1151 <= forvar1104;
    end
  assign wire1152 = {$unsigned((reg1100 ?
                            (reg1074 ?
                                reg1114 : forvar1102) : forvar1132[(3'h4):(1'h0)]))};
  module1153 modinst3995 (wire3994, clk, reg1126, forvar1090, reg1107, reg1099, forvar1132);
  module2367 modinst3997 (.y(wire3996), .wire2371(reg1063), .wire2369(reg1099), .clk(clk), .wire2368(reg1149), .wire2370(reg1127));
  assign wire3998 = $unsigned(reg1065[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar3999 = (1'h0); (forvar3999 < (2'h3)); forvar3999 = (forvar3999 + (1'h1)))
        begin
          if ((-($signed((!(8'ha8))) * $unsigned($unsigned(reg1144)))))
            begin
              for (forvar4000 = (1'h0); (forvar4000 < (1'h1)); forvar4000 = (forvar4000 + (1'h1)))
                begin
                  for (forvar4001 = (1'h0); (forvar4001 < (2'h3)); forvar4001 = (forvar4001 + (1'h1)))
                    begin
                      reg4002 <= forvar1119[(2'h2):(2'h2)];
                    end
                  reg4003 <= forvar1103[(4'h9):(3'h7)];
                end
            end
          else
            begin
              for (forvar4000 = (1'h0); (forvar4000 < (2'h3)); forvar4000 = (forvar4000 + (1'h1)))
                begin
                  if ((forvar1105[(2'h3):(2'h2)] <= (8'haf)))
                    begin
                      reg4001 <= ($unsigned(wire1056[(3'h5):(2'h3)]) ?
                          (8'hba) : reg1073[(2'h2):(2'h2)]);
                      reg4002 <= {{reg1084}};
                      reg4003 <= (+$unsigned(((forvar1090 ?
                          (8'h9e) : reg1063) | (+reg1103))));
                    end
                  else
                    begin
                      reg4001 <= reg1150;
                      reg4002 <= $signed($unsigned(((forvar1105 ?
                          reg1103 : reg1116) <= $unsigned(forvar1103))));
                      reg4003 <= ($signed({forvar1107}) + forvar1145[(3'h4):(3'h4)]);
                    end
                  reg4004 <= $unsigned($signed(reg1127[(2'h3):(2'h2)]));
                end
              if ((^~reg1060))
                begin
                  for (forvar4005 = (1'h0); (forvar4005 < (2'h2)); forvar4005 = (forvar4005 + (1'h1)))
                    begin
                      reg4006 <= (&reg1121[(1'h1):(1'h0)]);
                      reg4007 <= ($unsigned(($signed(reg1070) ?
                              $signed(reg1136) : forvar1091[(4'h9):(4'h8)])) ?
                          {reg1118} : $unsigned(reg1147));
                    end
                  reg4008 <= $signed((-(8'hb4)));
                end
              else
                begin
                  if ((~|wire3996[(3'h5):(3'h4)]))
                    begin
                      reg4005 <= wire1152;
                    end
                  else
                    begin
                      reg4005 <= ($signed(reg1111) ?
                          (reg1112[(4'he):(2'h2)] << (|(wire3994 ?
                              reg1151 : reg1100))) : reg1124);
                      reg4006 <= ({$signed((!wire3994))} >= (~|(+(forvar1069 << reg4002))));
                      reg4007 <= reg1068;
                    end
                end
              if ((8'haf))
                begin
                  if ($signed(reg1112))
                    begin
                      reg4009 <= {reg1148};
                      reg4010 <= (!$signed($unsigned(reg1136[(3'h6):(3'h4)])));
                    end
                  else
                    begin
                      reg4009 <= (wire643 ?
                          (((forvar1079 ? reg4003 : reg1128) ?
                                  reg1135 : (forvar1132 && reg1068)) ?
                              ((-forvar1079) ?
                                  $signed(reg4001) : (!forvar4005)) : forvar1104) : (-forvar1103));
                      reg4010 <= $unsigned((reg4004[(1'h0):(1'h0)] << ((forvar1102 >> (8'ha3)) <<< $unsigned(forvar1075))));
                      reg4011 <= $signed({({reg1082} || reg1085)});
                    end
                  for (forvar4012 = (1'h0); (forvar4012 < (1'h0)); forvar4012 = (forvar4012 + (1'h1)))
                    begin
                      reg4013 <= ({wire644} <= (($unsigned(reg1110) - (~reg4006)) ?
                          $signed($unsigned(forvar4000)) : ((|(8'ha2)) ?
                              $signed(forvar1069) : {(8'ha6)})));
                      reg4014 <= $signed($signed(reg1088[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  for (forvar4009 = (1'h0); (forvar4009 < (1'h0)); forvar4009 = (forvar4009 + (1'h1)))
                    begin
                      reg4010 <= reg1151;
                    end
                  for (forvar4011 = (1'h0); (forvar4011 < (2'h2)); forvar4011 = (forvar4011 + (1'h1)))
                    begin
                      reg4012 <= $signed((((forvar4001 ?
                          (8'h9f) : reg1108) >> reg4007[(1'h1):(1'h1)]) != reg1114[(4'h8):(2'h3)]));
                      reg4013 <= $signed((~&reg1120));
                    end
                  if (reg1068)
                    begin
                      reg4014 <= forvar1107;
                      reg4015 <= {forvar1059};
                    end
                  else
                    begin
                      reg4014 <= (({$unsigned(wire3996)} ?
                              (reg4008 ?
                                  reg1148[(2'h2):(1'h0)] : (reg1134 * wire642)) : $unsigned((reg1147 ^~ wire645))) ?
                          (({reg1137} ?
                              ((8'hb8) & forvar4011) : (forvar1107 >= reg4011)) <<< reg1077[(4'h8):(2'h2)]) : reg1110[(3'h5):(3'h4)]);
                      reg4015 <= forvar1122[(2'h2):(1'h1)];
                      reg4016 <= (~(^$signed((reg4015 || (8'hb4)))));
                      reg4017 <= $signed({$unsigned((reg1124 <<< reg1063))});
                    end
                end
            end
          if ({((^~(~^reg1147)) ?
                  ($unsigned(reg1146) ?
                      (reg1121 ~^ reg1107) : $unsigned(wire643)) : {(reg1085 ?
                          reg1108 : reg1126)})})
            begin
              if ($unsigned({(forvar1115 | forvar1070)}))
                begin
                  if (($unsigned($signed(reg4014[(1'h1):(1'h0)])) ?
                      reg1099 : $unsigned((^~{(8'hab)}))))
                    begin
                      reg4018 <= forvar4012[(1'h1):(1'h0)];
                      reg4019 <= reg4018;
                      reg4020 <= forvar1075;
                      reg4021 <= $signed(forvar1070[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg4018 <= forvar1090;
                      reg4019 <= ($unsigned(reg1068[(3'h5):(3'h4)]) ?
                          (reg1149 == {forvar1142}) : (-$unsigned((^~reg4009))));
                    end
                  if (reg1103)
                    begin
                      reg4022 <= $signed($unsigned({((8'hb1) ^ reg4021)}));
                    end
                  else
                    begin
                      reg4022 <= (&(reg1099[(4'hc):(1'h0)] == {(reg1105 ?
                              forvar1070 : reg1073)}));
                      reg4023 <= $signed(reg1101[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  if (forvar1131[(3'h7):(3'h6)])
                    begin
                      reg4018 <= (forvar4009[(1'h0):(1'h0)] ?
                          {$unsigned(reg1117)} : $unsigned(({reg1120} ?
                              {reg1149} : (reg1114 ? reg1150 : reg4016))));
                    end
                  else
                    begin
                      reg4018 <= (({(|(8'hb7))} ?
                              (reg1077 > ((8'hb3) ?
                                  reg4017 : forvar1142)) : (~^$unsigned(reg1113))) ?
                          (wire644[(3'h6):(2'h3)] ?
                              wire3996[(2'h3):(1'h1)] : $signed(reg1124[(1'h1):(1'h0)])) : $unsigned(forvar4000));
                      reg4019 <= $signed((~reg1063));
                    end
                  for (forvar4020 = (1'h0); (forvar4020 < (1'h1)); forvar4020 = (forvar4020 + (1'h1)))
                    begin
                      reg4021 <= reg1141[(4'h8):(3'h7)];
                      reg4022 <= $unsigned($unsigned($signed($signed(reg1127))));
                      reg4023 <= $unsigned($unsigned($signed($unsigned(reg1150))));
                      reg4024 <= $unsigned($unsigned($signed((reg1066 - reg1067))));
                    end
                  for (forvar4025 = (1'h0); (forvar4025 < (1'h0)); forvar4025 = (forvar4025 + (1'h1)))
                    begin
                      reg4026 <= $signed((forvar4012[(1'h1):(1'h1)] ?
                          (~$signed(forvar1142)) : (8'h9f)));
                      reg4027 <= (|reg1147);
                      reg4028 <= (~&$unsigned((|reg1116[(1'h0):(1'h0)])));
                    end
                end
              for (forvar4029 = (1'h0); (forvar4029 < (1'h0)); forvar4029 = (forvar4029 + (1'h1)))
                begin
                  for (forvar4030 = (1'h0); (forvar4030 < (1'h1)); forvar4030 = (forvar4030 + (1'h1)))
                    begin
                      reg4031 <= wire3996[(3'h4):(2'h3)];
                      reg4032 <= (~$unsigned(($signed((8'hb8)) & (forvar4025 ?
                          forvar1092 : wire1056))));
                      reg4033 <= $signed(reg1088);
                      reg4034 <= reg1078[(2'h3):(2'h3)];
                    end
                end
              reg4035 <= reg1137;
              for (forvar4036 = (1'h0); (forvar4036 < (1'h1)); forvar4036 = (forvar4036 + (1'h1)))
                begin
                  if ($signed(((^{reg4002}) ^~ (8'hba))))
                    begin
                      reg4037 <= wire1056;
                      reg4038 <= $signed($unsigned(($unsigned(reg1064) << reg4037[(4'h8):(1'h1)])));
                      reg4039 <= (reg1114 ?
                          (~&reg1151[(2'h2):(1'h0)]) : reg4019);
                      reg4040 <= ((!(wire3994 ?
                          (&reg1070) : wire642[(3'h5):(1'h1)])) == forvar1091);
                    end
                  else
                    begin
                      reg4037 <= (8'hab);
                      reg4038 <= (-($signed(wire642[(2'h2):(1'h0)]) >= forvar1090[(4'h9):(4'h8)]));
                      reg4039 <= $unsigned((^~$signed($signed(forvar4020))));
                      reg4040 <= $signed((&reg4002[(3'h7):(3'h6)]));
                    end
                  for (forvar4041 = (1'h0); (forvar4041 < (2'h3)); forvar4041 = (forvar4041 + (1'h1)))
                    begin
                      reg4042 <= reg1126[(3'h5):(1'h0)];
                      reg4043 <= (+reg1062);
                      reg4044 <= $signed(reg1107);
                    end
                  reg4045 <= $unsigned((~|$signed(reg1109)));
                end
            end
          else
            begin
              for (forvar4018 = (1'h0); (forvar4018 < (2'h3)); forvar4018 = (forvar4018 + (1'h1)))
                begin
                  reg4019 <= $unsigned((reg1070 ^~ $signed((reg4014 ?
                      reg1143 : (8'hb5)))));
                end
              for (forvar4020 = (1'h0); (forvar4020 < (1'h1)); forvar4020 = (forvar4020 + (1'h1)))
                begin
                  reg4021 <= $signed((((reg1073 <<< forvar1105) ?
                          (reg1085 * forvar4001) : {reg1113}) ?
                      $signed(reg4018) : reg1143[(4'h8):(4'h8)]));
                  for (forvar4022 = (1'h0); (forvar4022 < (2'h2)); forvar4022 = (forvar4022 + (1'h1)))
                    begin
                      reg4023 <= (forvar3999[(1'h0):(1'h0)] & reg4027);
                    end
                end
              for (forvar4024 = (1'h0); (forvar4024 < (1'h1)); forvar4024 = (forvar4024 + (1'h1)))
                begin
                  if (($unsigned((8'haa)) ?
                      ((^reg1088) <= reg4023) : (~^(reg1073[(1'h1):(1'h1)] ?
                          forvar4000 : (reg1149 + reg4010)))))
                    begin
                      reg4025 <= ({{$signed(forvar4000)}} << $signed((|((8'hba) << forvar1105))));
                      reg4026 <= reg4031;
                      reg4027 <= $unsigned(forvar1145[(4'h8):(1'h1)]);
                    end
                  else
                    begin
                      reg4025 <= (($signed(forvar1092[(3'h5):(1'h1)]) ?
                              reg1108 : $signed(((8'hb2) ^ reg4034))) ?
                          {reg1120} : ({(|reg4004)} ?
                              $signed($signed(reg1150)) : $signed({forvar4018})));
                      reg4026 <= (reg4020 ^ forvar4036);
                      reg4027 <= $unsigned((($signed(reg4039) ?
                              wire3998 : forvar4036[(2'h2):(2'h2)]) ?
                          $unsigned(forvar4029) : $unsigned((forvar1104 ?
                              reg4025 : reg4008))));
                      reg4028 <= (reg4001 >> $unsigned($signed(((8'ha2) - reg1074))));
                    end
                  for (forvar4029 = (1'h0); (forvar4029 < (2'h3)); forvar4029 = (forvar4029 + (1'h1)))
                    begin
                      reg4030 <= ($unsigned($unsigned(reg1147)) ?
                          reg1078 : (-(|(forvar4011 != reg1084))));
                      reg4031 <= $signed(({{(8'hb4)}} ?
                          reg4021 : reg4012[(1'h1):(1'h1)]));
                    end
                  if ((reg4005 ?
                      (-(~reg4010[(1'h0):(1'h0)])) : (+$signed((reg1151 | reg4031)))))
                    begin
                      reg4032 <= reg1081;
                    end
                  else
                    begin
                      reg4032 <= (forvar1119[(1'h0):(1'h0)] ?
                          ($unsigned(reg1099) || reg4040) : (reg1087[(3'h4):(1'h0)] ?
                              ((&forvar4036) != $unsigned(forvar1105)) : $unsigned(forvar1130)));
                      reg4033 <= $unsigned(($unsigned((reg1078 == (8'h9d))) ?
                          ($unsigned(forvar1105) != $unsigned(reg1127)) : $unsigned((reg1121 ?
                              reg1067 : reg4045))));
                      reg4034 <= ($signed((-reg1104[(1'h1):(1'h0)])) ^ $unsigned(({forvar4029} ?
                          (forvar1069 ?
                              reg4015 : reg1060) : (forvar4005 >> reg1094))));
                      reg4035 <= $signed((8'ha9));
                    end
                end
              reg4036 <= $signed($signed(((~&(8'hb6)) ?
                  ((8'hb0) ? reg4022 : forvar1102) : (reg4037 > (8'hba)))));
            end
          for (forvar4046 = (1'h0); (forvar4046 < (2'h3)); forvar4046 = (forvar4046 + (1'h1)))
            begin
              for (forvar4047 = (1'h0); (forvar4047 < (2'h3)); forvar4047 = (forvar4047 + (1'h1)))
                begin
                  for (forvar4048 = (1'h0); (forvar4048 < (2'h2)); forvar4048 = (forvar4048 + (1'h1)))
                    begin
                      reg4049 <= (^($unsigned($signed(reg4022)) == (-forvar4005)));
                    end
                end
              if (($unsigned({$unsigned(reg1107)}) ?
                  (((reg4007 ? forvar1069 : reg1084) | {reg4049}) ?
                      (reg1120[(3'h4):(2'h3)] ?
                          $signed(reg1149) : $signed(forvar4020)) : {wire3998}) : ($signed(reg4010[(1'h0):(1'h0)]) ?
                      reg4011[(2'h3):(2'h3)] : $unsigned({reg1078}))))
                begin
                  for (forvar4050 = (1'h0); (forvar4050 < (2'h2)); forvar4050 = (forvar4050 + (1'h1)))
                    begin
                      reg4051 <= $signed($unsigned($unsigned(reg1126)));
                    end
                  if ($unsigned({((reg1136 ? reg1073 : reg1135) ?
                          $signed(reg1150) : (reg1112 ?
                              forvar1132 : forvar3999))}))
                    begin
                      reg4052 <= (({reg1141} << $signed(((8'ha3) | reg4009))) ?
                          forvar4029[(1'h0):(1'h0)] : (reg1088 ?
                              $unsigned({reg4021}) : (|reg4025)));
                    end
                  else
                    begin
                      reg4052 <= $signed(($unsigned((8'h9c)) ?
                          $signed((^~(8'hb8))) : reg4052));
                      reg4053 <= $signed($unsigned((reg1150[(3'h5):(1'h1)] == (reg4021 ?
                          reg1066 : reg1133))));
                    end
                  for (forvar4054 = (1'h0); (forvar4054 < (2'h2)); forvar4054 = (forvar4054 + (1'h1)))
                    begin
                      reg4055 <= reg1116;
                      reg4056 <= $signed(forvar1095[(4'h9):(2'h2)]);
                    end
                  reg4057 <= reg1088[(4'ha):(1'h1)];
                end
              else
                begin
                  reg4050 <= $signed($unsigned(reg1124));
                  for (forvar4051 = (1'h0); (forvar4051 < (1'h0)); forvar4051 = (forvar4051 + (1'h1)))
                    begin
                      reg4052 <= $unsigned($signed((reg1086 ?
                          (reg4044 ?
                              reg1074 : reg1105) : reg1139[(2'h2):(1'h1)])));
                      reg4053 <= $signed({(8'hb2)});
                      reg4054 <= $unsigned($signed(((reg4013 >> reg4052) ?
                          $signed(reg1105) : (-forvar4018))));
                      reg4055 <= (^reg1109);
                    end
                  if ($unsigned($signed(reg1065)))
                    begin
                      reg4056 <= $signed(forvar1070[(3'h5):(3'h4)]);
                      reg4057 <= ($signed({reg1140}) ?
                          {($unsigned(reg1105) ?
                                  ((8'haf) ? reg4027 : reg4025) : ((8'hb7) ?
                                      reg1133 : reg4039))} : {wire646});
                      reg4058 <= (reg4017[(4'ha):(3'h4)] <<< reg1127[(3'h6):(1'h1)]);
                    end
                  else
                    begin
                      reg4056 <= reg4015[(2'h2):(1'h1)];
                      reg4057 <= reg4042[(2'h2):(2'h2)];
                      reg4058 <= ((8'h9c) <= reg1133);
                      reg4059 <= (8'hb5);
                    end
                  if (reg4003)
                    begin
                      reg4060 <= $signed($unsigned(($signed(forvar4030) || (reg1120 ?
                          (8'hba) : reg4028))));
                    end
                  else
                    begin
                      reg4060 <= ((reg4055 >>> {reg4009}) ?
                          $unsigned($unsigned((reg1099 >> (8'ha5)))) : $unsigned((((8'h9e) ?
                              reg1108 : reg4011) << (|(8'hac)))));
                      reg4061 <= ({reg4043} ?
                          (8'hac) : (reg1066 ^ (|(reg4044 ?
                              forvar1145 : (8'ha4)))));
                      reg4062 <= (reg1100 << reg4014[(3'h6):(3'h4)]);
                      reg4063 <= reg1096;
                    end
                end
              if ($unsigned(reg1121[(4'h9):(3'h4)]))
                begin
                  reg4064 <= ($signed((!(~&(8'hb0)))) ?
                      $unsigned(({wire3994} ?
                          reg1098[(4'h8):(1'h1)] : $signed(reg4023))) : reg4053[(4'h8):(1'h0)]);
                  for (forvar4065 = (1'h0); (forvar4065 < (2'h3)); forvar4065 = (forvar4065 + (1'h1)))
                    begin
                      reg4066 <= ((+reg4038) ? {(+reg1076)} : forvar4005);
                      reg4067 <= $unsigned((reg4049 ?
                          reg4022 : $signed($signed(reg1116))));
                      reg4068 <= forvar1079;
                    end
                end
              else
                begin
                  reg4064 <= $signed((reg4056 >= reg4028[(3'h7):(2'h2)]));
                  if ((forvar1079 ?
                      wire3994[(1'h0):(1'h0)] : $signed(({(8'h9f)} ?
                          reg1093 : {reg1117}))))
                    begin
                      reg4065 <= (({(+reg1073)} ?
                              ($unsigned(reg4008) ?
                                  (forvar4065 ?
                                      reg1137 : reg4024) : (~&wire3996)) : ($unsigned(wire643) ?
                                  (reg4020 != (8'h9e)) : $unsigned(reg4054))) ?
                          $signed(((&reg4028) ?
                              (reg1125 || (8'ha1)) : $signed(reg4033))) : (^~((forvar1104 ?
                              forvar4029 : reg4059) > $unsigned(reg1081))));
                      reg4066 <= {((~&$unsigned(reg1134)) - ($signed(wire642) ?
                              (|forvar1122) : reg1108[(1'h1):(1'h1)]))};
                      reg4067 <= (8'ha2);
                      reg4068 <= (~|reg1113[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg4065 <= $unsigned($unsigned(({forvar1059} ?
                          reg4057[(2'h2):(1'h1)] : (reg1129 >= wire3998))));
                      reg4066 <= ($unsigned(({reg1137} ?
                              $unsigned(forvar1090) : (~^(8'hb4)))) ?
                          ($signed((reg1133 >= reg1140)) ?
                              (|(forvar4000 * reg1120)) : reg4031[(3'h6):(1'h0)]) : (^forvar1075[(2'h3):(2'h3)]));
                      reg4067 <= (8'ha9);
                      reg4068 <= forvar4009;
                    end
                  for (forvar4069 = (1'h0); (forvar4069 < (2'h2)); forvar4069 = (forvar4069 + (1'h1)))
                    begin
                      reg4070 <= $signed((reg1086 ?
                          (reg1078 ~^ $unsigned(reg4027)) : ($unsigned(wire644) & forvar1119[(1'h1):(1'h1)])));
                      reg4071 <= $signed($unsigned(((8'hb1) ?
                          $signed(forvar1091) : forvar1130[(4'ha):(1'h1)])));
                      reg4072 <= $unsigned({(((8'ha9) ?
                              reg4016 : reg4008) != $unsigned(reg1104))});
                      reg4073 <= reg1073;
                    end
                  if (((forvar1142[(2'h2):(1'h0)] >> {forvar4047}) ^~ $signed(((forvar1079 | forvar1122) & {(8'ha7)}))))
                    begin
                      reg4074 <= {((|reg1108[(1'h1):(1'h1)]) ?
                              (-$unsigned(reg4066)) : ($signed(reg4035) ?
                                  $unsigned(forvar4022) : reg1120[(3'h4):(1'h1)]))};
                      reg4075 <= reg4072[(3'h7):(3'h5)];
                      reg4076 <= $unsigned(forvar4048[(1'h0):(1'h0)]);
                      reg4077 <= reg4025[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg4074 <= (((8'ha5) ?
                              $unsigned($unsigned((8'ha2))) : ($signed(reg4004) ?
                                  {reg1087} : reg1077)) ?
                          $signed((~&$unsigned(forvar4011))) : $unsigned({(reg1151 ?
                                  reg4045 : forvar1090)}));
                      reg4075 <= (reg4062 <= forvar1079);
                      reg4076 <= reg4007[(4'hc):(3'h7)];
                    end
                end
              if (($unsigned((&forvar1131)) & $unsigned(((reg4058 <<< (8'ha7)) ?
                  (reg1107 ? reg1070 : reg4054) : $signed(reg1123)))))
                begin
                  if (($unsigned($unsigned((reg1121 <= reg1063))) ?
                      $signed(({reg4038} ?
                          (reg1111 ?
                              reg1066 : reg1113) : (reg4017 <= reg1080))) : {$unsigned(reg1134[(3'h5):(2'h2)])}))
                    begin
                      reg4078 <= $signed((~|((forvar1105 & reg1087) ?
                          (wire646 ? reg1111 : reg4017) : $signed(reg4035))));
                      reg4079 <= reg1134;
                    end
                  else
                    begin
                      reg4078 <= $signed(reg4039[(3'h4):(1'h1)]);
                      reg4079 <= {((~$signed(wire3996)) << forvar4012)};
                      reg4080 <= (reg4001 ?
                          $unsigned(((wire1152 != (8'ha0)) + $unsigned(wire3996))) : ((^(~^(8'hb0))) <<< reg4074[(2'h3):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar4078 = (1'h0); (forvar4078 < (2'h2)); forvar4078 = (forvar4078 + (1'h1)))
                    begin
                      reg4079 <= $unsigned((^~forvar1122));
                      reg4080 <= reg1084;
                    end
                  reg4081 <= reg4068;
                  if ($signed((^$signed($signed(reg4025)))))
                    begin
                      reg4082 <= {(^~$unsigned((reg4026 ? reg4020 : (8'hba))))};
                      reg4083 <= $signed($signed(reg1141));
                      reg4084 <= ({$signed((reg4073 ? (8'haa) : reg1088))} ?
                          (^~{reg1120}) : {reg1143[(3'h5):(3'h5)]});
                      reg4085 <= wire642[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg4082 <= ((reg4032[(1'h1):(1'h0)] ?
                              reg1134[(2'h2):(1'h0)] : {(~&reg1093)}) ?
                          {($unsigned(reg1061) | reg4061)} : (reg4037 ?
                              (reg1068 ?
                                  reg1068[(1'h1):(1'h1)] : ((8'hb4) ?
                                      (8'ha3) : (8'haa))) : reg1128));
                      reg4083 <= ((^~(~^(reg4001 ? reg4039 : forvar1105))) ?
                          (wire3996 ?
                              reg4031[(2'h3):(1'h1)] : $unsigned($signed(reg4032))) : (~|wire644[(1'h1):(1'h0)]));
                      reg4084 <= reg4003;
                      reg4085 <= $unsigned(reg4001);
                    end
                end
            end
        end
    end
  assign wire4086 = reg4055[(4'ha):(4'h9)];
  always
    @(posedge clk) begin
      reg4087 <= (reg4033 == reg1123);
      if ((8'h9d))
        begin
          for (forvar4088 = (1'h0); (forvar4088 < (2'h2)); forvar4088 = (forvar4088 + (1'h1)))
            begin
              if (reg1084[(3'h7):(3'h4)])
                begin
                  for (forvar4089 = (1'h0); (forvar4089 < (2'h3)); forvar4089 = (forvar4089 + (1'h1)))
                    begin
                      reg4090 <= $unsigned(reg4052[(3'h6):(3'h4)]);
                      reg4091 <= $signed($unsigned((^$signed(reg4050))));
                      reg4092 <= (reg4012[(3'h4):(1'h0)] ?
                          {reg1141[(2'h3):(2'h3)]} : reg1121);
                      reg4093 <= (($signed((reg1081 - reg4024)) + (^~(8'ha8))) ?
                          reg1136 : reg1083[(1'h0):(1'h0)]);
                    end
                  if ($unsigned(reg1066))
                    begin
                      reg4094 <= $signed(forvar1079[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg4094 <= (~&(8'ha4));
                      reg4095 <= (~|$unsigned(($unsigned(reg4075) < $unsigned(reg1112))));
                      reg4096 <= ($unsigned({$signed(wire1152)}) ?
                          (($unsigned(reg1127) ?
                                  (forvar4065 ?
                                      reg4057 : reg1060) : {reg4015}) ?
                              reg1134 : (~(+reg4076))) : reg4031[(2'h2):(1'h1)]);
                    end
                  for (forvar4097 = (1'h0); (forvar4097 < (1'h1)); forvar4097 = (forvar4097 + (1'h1)))
                    begin
                      reg4098 <= ((8'h9d) > $signed(($signed(reg1110) ^~ (~(8'hb5)))));
                      reg4099 <= {(($signed((8'hb5)) ?
                              (reg1139 ?
                                  reg4031 : reg1084) : {reg4095}) < reg4026)};
                      reg4100 <= $signed((reg4042[(1'h0):(1'h0)] ?
                          (reg1074 <= (~wire646)) : forvar4069));
                    end
                end
              else
                begin
                  if ((8'hb1))
                    begin
                      reg4089 <= $signed((~&reg4067));
                    end
                  else
                    begin
                      reg4089 <= $signed((~$signed({reg4032})));
                    end
                end
              if (((reg1137 ?
                      $signed($signed(reg4008)) : (&(forvar4005 <<< reg4030))) ?
                  reg4052[(3'h5):(2'h3)] : $unsigned((reg1082[(4'h8):(2'h3)] ?
                      (reg4039 ? (8'ha7) : reg1151) : ((8'hab) <<< reg4011)))))
                begin
                  if ((reg4078[(4'h9):(3'h4)] ?
                      ((+(reg1078 * forvar1069)) ?
                          $signed((reg4063 | reg1146)) : $unsigned(forvar4009)) : (((reg4055 ?
                              reg4100 : forvar4022) ~^ (reg4093 ?
                              reg4078 : reg4067)) ?
                          (!$unsigned(forvar1079)) : reg1088)))
                    begin
                      reg4101 <= wire644[(3'h4):(3'h4)];
                      reg4102 <= $signed(reg4038);
                      reg4103 <= $signed(($signed($unsigned(reg1112)) ~^ ((reg4034 >= reg4053) ?
                          (reg4062 & reg1143) : (~forvar1069))));
                      reg4104 <= wire3996[(3'h6):(3'h6)];
                    end
                  else
                    begin
                      reg4101 <= (reg4054[(3'h4):(2'h3)] | $signed({(reg1112 ?
                              reg1078 : (8'ha7))}));
                    end
                  for (forvar4105 = (1'h0); (forvar4105 < (2'h2)); forvar4105 = (forvar4105 + (1'h1)))
                    begin
                      reg4106 <= (reg1066[(1'h0):(1'h0)] + reg4021[(3'h4):(2'h2)]);
                    end
                  reg4107 <= ($unsigned((+reg1105[(2'h3):(1'h0)])) ?
                      ($signed((reg1065 != reg4098)) <<< (|reg4077)) : (-((reg4062 ?
                          (8'hb9) : forvar1142) <<< (forvar1103 ?
                          (8'hab) : forvar4000))));
                  for (forvar4108 = (1'h0); (forvar4108 < (2'h2)); forvar4108 = (forvar4108 + (1'h1)))
                    begin
                      reg4109 <= reg4045[(2'h3):(1'h0)];
                    end
                end
              else
                begin
                  reg4101 <= $signed(reg4082);
                end
              for (forvar4110 = (1'h0); (forvar4110 < (1'h1)); forvar4110 = (forvar4110 + (1'h1)))
                begin
                  if (wire3998[(3'h4):(2'h3)])
                    begin
                      reg4111 <= $unsigned(wire3994);
                      reg4112 <= ($unsigned($signed(((8'ha9) ?
                          reg1073 : forvar4005))) ^ (~|(reg4045[(2'h2):(1'h1)] ?
                          ((8'hb1) ? (8'hb4) : forvar1131) : {(8'hab)})));
                      reg4113 <= $unsigned($unsigned(({reg4066} ?
                          forvar4024 : $signed(reg1140))));
                      reg4114 <= $unsigned($unsigned(($unsigned(reg1151) & (reg4036 ?
                          reg4080 : forvar4001))));
                    end
                  else
                    begin
                      reg4111 <= ($unsigned(((reg1135 ? forvar1060 : reg4034) ?
                              (reg4057 ? (8'h9e) : wire3994) : (-reg1143))) ?
                          (|{$unsigned(forvar1142)}) : ({$unsigned(reg1112)} && $unsigned(forvar1131)));
                    end
                  if ($unsigned(reg4030[(1'h0):(1'h0)]))
                    begin
                      reg4115 <= $signed($unsigned(reg1063[(4'h8):(2'h2)]));
                    end
                  else
                    begin
                      reg4115 <= (reg4004 & $signed(forvar1092[(4'h8):(4'h8)]));
                      reg4116 <= reg4028[(3'h6):(3'h5)];
                      reg4117 <= {(~^{reg4068[(2'h2):(1'h1)]})};
                      reg4118 <= {reg1128[(2'h3):(2'h3)]};
                    end
                  for (forvar4119 = (1'h0); (forvar4119 < (2'h3)); forvar4119 = (forvar4119 + (1'h1)))
                    begin
                      reg4120 <= (8'ha4);
                    end
                end
            end
          reg4121 <= $signed((~|({reg4082} ^ {forvar4050})));
          for (forvar4122 = (1'h0); (forvar4122 < (2'h3)); forvar4122 = (forvar4122 + (1'h1)))
            begin
              if (reg4082)
                begin
                  if (reg1124)
                    begin
                      reg4123 <= $signed($signed($signed(forvar1131[(3'h7):(1'h0)])));
                      reg4124 <= reg4027[(2'h2):(2'h2)];
                      reg4125 <= $unsigned((reg4014[(3'h5):(1'h1)] ?
                          reg4117 : reg4044[(4'h9):(1'h0)]));
                      reg4126 <= $unsigned($unsigned((~&(~&(8'ha8)))));
                    end
                  else
                    begin
                      reg4123 <= reg4012;
                      reg4124 <= $unsigned((|(&$unsigned(reg1099))));
                    end
                  for (forvar4127 = (1'h0); (forvar4127 < (2'h2)); forvar4127 = (forvar4127 + (1'h1)))
                    begin
                      reg4128 <= (~&(|(|(|reg1080))));
                      reg4129 <= {($signed((~^reg4051)) ?
                              reg1128 : reg4126[(2'h3):(2'h3)])};
                      reg4130 <= (8'h9e);
                      reg4131 <= $unsigned((~reg4027[(1'h0):(1'h0)]));
                    end
                  for (forvar4132 = (1'h0); (forvar4132 < (2'h3)); forvar4132 = (forvar4132 + (1'h1)))
                    begin
                      reg4133 <= {$signed({(^forvar4024)})};
                      reg4134 <= (reg4115[(3'h6):(2'h3)] ?
                          forvar4097[(2'h2):(2'h2)] : reg4044[(1'h1):(1'h1)]);
                    end
                  for (forvar4135 = (1'h0); (forvar4135 < (1'h0)); forvar4135 = (forvar4135 + (1'h1)))
                    begin
                      reg4136 <= wire643;
                      reg4137 <= $signed((($signed(reg4084) * reg4123[(2'h3):(1'h1)]) ?
                          reg4099[(3'h6):(1'h0)] : (~^$unsigned(reg1111))));
                      reg4138 <= reg1143[(1'h1):(1'h0)];
                      reg4139 <= $unsigned($unsigned(reg4102[(4'h9):(2'h2)]));
                    end
                end
              else
                begin
                  if (((^forvar1059[(4'ha):(3'h7)]) ?
                      reg4116[(2'h2):(1'h0)] : $unsigned((reg1088[(2'h3):(1'h1)] ?
                          (forvar4000 && reg4099) : $signed(reg4031)))))
                    begin
                      reg4123 <= reg1141;
                      reg4124 <= (!$signed(((forvar1092 || forvar1119) >= $signed(forvar4119))));
                      reg4125 <= (reg1083 ?
                          (($signed(reg1083) ^ $signed(reg4078)) ?
                              $signed($signed((8'hb3))) : forvar4105) : {$signed($unsigned(reg4068))});
                    end
                  else
                    begin
                      reg4123 <= reg4115;
                      reg4124 <= reg1129[(3'h5):(2'h3)];
                    end
                  if (reg1123[(2'h2):(1'h0)])
                    begin
                      reg4126 <= $signed(($signed($unsigned((8'ha0))) ?
                          wire643[(2'h2):(1'h0)] : $unsigned({(8'hb3)})));
                      reg4127 <= ($signed(reg4008) ?
                          (8'hb7) : reg4010[(1'h0):(1'h0)]);
                      reg4128 <= $signed(wire1058[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg4126 <= (~^$signed($unsigned((reg1086 ?
                          reg1101 : forvar4000))));
                      reg4127 <= ($unsigned(reg4033[(3'h7):(1'h0)]) ~^ $signed($signed(forvar4005)));
                      reg4128 <= forvar1092[(1'h0):(1'h0)];
                    end
                  if ((~&(reg4035[(2'h2):(1'h1)] || (~|$unsigned(reg4074)))))
                    begin
                      reg4129 <= wire644[(4'h8):(2'h3)];
                      reg4130 <= reg4098[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg4129 <= ({reg4113[(2'h3):(2'h3)]} ?
                          $unsigned(((8'hb3) <= (~|(8'ha3)))) : reg4036);
                    end
                end
              reg4140 <= reg4129;
              reg4141 <= {$unsigned($unsigned($signed(wire645)))};
            end
        end
      else
        begin
          if ((~(~|(~|(!wire3996)))))
            begin
              reg4088 <= {$signed(((wire642 >>> reg4013) == (forvar4005 ?
                      reg4053 : reg4117)))};
              if (reg4087[(3'h5):(2'h3)])
                begin
                  for (forvar4089 = (1'h0); (forvar4089 < (1'h0)); forvar4089 = (forvar4089 + (1'h1)))
                    begin
                      reg4090 <= (reg4066[(4'ha):(3'h7)] ?
                          reg4003[(2'h3):(1'h1)] : (~|{reg4136[(2'h2):(2'h2)]}));
                      reg4091 <= forvar4097[(1'h0):(1'h0)];
                    end
                  for (forvar4092 = (1'h0); (forvar4092 < (1'h0)); forvar4092 = (forvar4092 + (1'h1)))
                    begin
                      reg4093 <= {$unsigned(((~forvar4135) >> reg4006))};
                    end
                end
              else
                begin
                  for (forvar4089 = (1'h0); (forvar4089 < (2'h2)); forvar4089 = (forvar4089 + (1'h1)))
                    begin
                      reg4090 <= $unsigned($signed(reg4051));
                    end
                  reg4091 <= $unsigned($unsigned(({reg4092} >> (reg1149 ?
                      reg4101 : (8'ha7)))));
                  if ($unsigned($signed((&$unsigned(reg1085)))))
                    begin
                      reg4092 <= reg4075[(3'h7):(3'h6)];
                    end
                  else
                    begin
                      reg4092 <= {(-((reg1136 ?
                              reg1099 : reg4102) | (|reg4123)))};
                      reg4093 <= ($signed($unsigned((reg1151 ?
                              reg4131 : reg4059))) ?
                          $signed($unsigned((8'hb6))) : (!$signed({forvar4001})));
                      reg4094 <= forvar4001[(3'h5):(3'h4)];
                    end
                  for (forvar4095 = (1'h0); (forvar4095 < (1'h0)); forvar4095 = (forvar4095 + (1'h1)))
                    begin
                      reg4096 <= reg4011;
                    end
                end
              for (forvar4097 = (1'h0); (forvar4097 < (1'h0)); forvar4097 = (forvar4097 + (1'h1)))
                begin
                  reg4098 <= $unsigned((((forvar4030 > (8'hb1)) ?
                          reg1144 : ((8'hb2) & reg4111)) ?
                      (~wire3994[(4'hc):(3'h6)]) : $unsigned(forvar1122)));
                  for (forvar4099 = (1'h0); (forvar4099 < (2'h3)); forvar4099 = (forvar4099 + (1'h1)))
                    begin
                      reg4100 <= (reg4117[(1'h0):(1'h0)] ^ ($unsigned({(8'hae)}) ?
                          (8'hb1) : $signed((reg1111 ? reg1104 : (8'hac)))));
                      reg4101 <= {(forvar1060 ^ ((reg4081 ?
                                  reg4087 : forvar4110) ?
                              ((8'hba) && (8'hb6)) : (reg4061 <= (8'h9e))))};
                    end
                  for (forvar4102 = (1'h0); (forvar4102 < (2'h2)); forvar4102 = (forvar4102 + (1'h1)))
                    begin
                      reg4103 <= reg1151[(2'h2):(2'h2)];
                      reg4104 <= $signed($unsigned((reg4018[(2'h2):(1'h0)] == reg4114)));
                      reg4105 <= $signed((reg4137[(3'h7):(3'h5)] ?
                          $signed(reg1103) : (-$signed(reg4099))));
                    end
                  for (forvar4106 = (1'h0); (forvar4106 < (1'h1)); forvar4106 = (forvar4106 + (1'h1)))
                    begin
                      reg4107 <= (reg1134 ?
                          reg4043 : $signed(reg1108[(2'h3):(1'h0)]));
                      reg4108 <= (|(reg4009 ?
                          ((reg4136 != forvar4089) || reg1100) : $unsigned({(8'hb3)})));
                      reg4109 <= reg4121;
                    end
                end
            end
          else
            begin
              for (forvar4088 = (1'h0); (forvar4088 < (1'h1)); forvar4088 = (forvar4088 + (1'h1)))
                begin
                  reg4089 <= ($unsigned(reg1111) | reg4103[(4'hd):(2'h3)]);
                end
            end
          reg4110 <= forvar4005[(3'h4):(2'h2)];
          for (forvar4111 = (1'h0); (forvar4111 < (1'h0)); forvar4111 = (forvar4111 + (1'h1)))
            begin
              for (forvar4112 = (1'h0); (forvar4112 < (1'h1)); forvar4112 = (forvar4112 + (1'h1)))
                begin
                  if (((~|{forvar4041}) ?
                      $signed(((reg4089 || reg1118) ^~ $signed(reg1105))) : (+((wire644 >= forvar1104) != reg4101))))
                    begin
                      reg4113 <= $signed({reg4037});
                      reg4114 <= (8'hb5);
                      reg4115 <= (((+(^~(8'h9f))) << $unsigned({reg4001})) ?
                          ((reg1108 ^~ (forvar4088 ^ (8'hb9))) ?
                              (~|$unsigned(reg1112)) : $unsigned((reg4014 <<< reg4077))) : $unsigned(wire1152));
                    end
                  else
                    begin
                      reg4113 <= reg4095[(4'h8):(2'h2)];
                      reg4114 <= ((($signed(reg4050) <= $unsigned(reg1078)) ?
                              $unsigned((reg4014 || reg1104)) : reg1143[(4'hc):(4'hc)]) ?
                          reg4103 : $signed(((~reg1141) || $unsigned((8'hb2)))));
                    end
                end
              for (forvar4116 = (1'h0); (forvar4116 < (2'h2)); forvar4116 = (forvar4116 + (1'h1)))
                begin
                  for (forvar4117 = (1'h0); (forvar4117 < (2'h3)); forvar4117 = (forvar4117 + (1'h1)))
                    begin
                      reg4118 <= $signed({(forvar1115 ?
                              $signed(reg4034) : reg4004)});
                      reg4119 <= $signed($signed((-reg1134[(3'h7):(2'h2)])));
                      reg4120 <= ((^wire646[(4'hb):(3'h6)]) ?
                          ($unsigned((reg4136 * (8'haf))) & (forvar1103 ?
                              reg4095 : (reg4064 == (8'had)))) : {$unsigned($signed(reg4030))});
                    end
                  if ($unsigned(forvar4122[(1'h1):(1'h1)]))
                    begin
                      reg4121 <= (~^forvar4069[(4'h9):(1'h0)]);
                      reg4122 <= forvar4099[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg4121 <= ((~^(~|(~forvar1092))) ?
                          reg1085[(3'h7):(3'h7)] : $unsigned((~(8'had))));
                    end
                end
              reg4123 <= $signed($signed({$signed((8'had))}));
              reg4124 <= $signed(({reg4094} != (8'hb7)));
            end
          reg4125 <= (reg4040 ? $signed({reg1137}) : reg1106);
        end
      reg4142 <= ($unsigned({forvar1122}) | reg4093);
    end
  assign wire4143 = ($signed((reg1150 ?
                        (^forvar1104) : (8'ha0))) ~^ {reg4019[(2'h2):(2'h2)]});
  assign wire4144 = $unsigned(reg1113[(1'h0):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1153
#( parameter param3993 = ((({(8'hb5)} << {(8'haa)}) ? (((8'haa) != (8'hab)) ? ((8'hb9) ? (8'h9f) : (8'haa)) : (|(8'h9e))) : (~&((8'hb0) ? (8'h9e) : (8'ha5)))) ? ((^(~|(8'ha3))) - ((~(8'h9e)) & ((8'haf) && (8'ha2)))) : (!(~^((8'ha9) ? (8'ha5) : (8'hb6))))) )
(y, clk, wire1158, wire1157, wire1156, wire1155, wire1154);
  output wire [(32'hf8b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire1158;
  input wire signed [(4'hf):(1'h0)] wire1157;
  input wire signed [(4'hd):(1'h0)] wire1156;
  input wire [(5'h10):(1'h0)] wire1155;
  input wire [(4'hb):(1'h0)] wire1154;
  wire [(4'hc):(1'h0)] wire3992;
  reg [(4'he):(1'h0)] reg3991 = (1'h0);
  reg [(4'he):(1'h0)] reg3990 = (1'h0);
  reg [(2'h2):(1'h0)] reg3989 = (1'h0);
  reg [(4'he):(1'h0)] reg3988 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3987 = (1'h0);
  reg [(4'hd):(1'h0)] reg3986 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3985 = (1'h0);
  reg [(4'h9):(1'h0)] reg3984 = (1'h0);
  reg [(3'h7):(1'h0)] reg3983 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3982 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3981 = (1'h0);
  reg [(4'he):(1'h0)] forvar3980 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3975 = (1'h0);
  reg [(4'he):(1'h0)] reg3979 = (1'h0);
  reg [(4'h9):(1'h0)] reg3978 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3977 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3976 = (1'h0);
  reg [(4'hf):(1'h0)] reg3975 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3974 = (1'h0);
  reg [(4'ha):(1'h0)] reg3973 = (1'h0);
  reg [(4'he):(1'h0)] reg3972 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3971 = (1'h0);
  reg [(4'he):(1'h0)] reg3970 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3969 = (1'h0);
  reg [(3'h5):(1'h0)] reg3968 = (1'h0);
  reg [(3'h6):(1'h0)] reg3967 = (1'h0);
  reg [(4'hf):(1'h0)] reg3966 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3965 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3964 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3963 = (1'h0);
  reg [(4'hf):(1'h0)] reg3962 = (1'h0);
  reg [(2'h3):(1'h0)] reg3961 = (1'h0);
  reg [(3'h6):(1'h0)] reg3960 = (1'h0);
  reg [(5'h10):(1'h0)] reg3959 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3958 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3957 = (1'h0);
  reg [(5'h10):(1'h0)] reg3956 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3955 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3954 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3953 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3952 = (1'h0);
  reg [(4'hc):(1'h0)] reg3951 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3950 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3949 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3948 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3947 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3946 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3945 = (1'h0);
  reg [(3'h7):(1'h0)] reg3944 = (1'h0);
  reg [(3'h4):(1'h0)] reg3943 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3942 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3941 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3940 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3939 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3887 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3886 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3879 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3882 = (1'h0);
  reg [(2'h3):(1'h0)] reg3877 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3874 = (1'h0);
  reg [(3'h7):(1'h0)] reg3873 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3872 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3869 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3868 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3865 = (1'h0);
  reg [(4'hc):(1'h0)] reg3863 = (1'h0);
  reg [(4'hd):(1'h0)] reg3938 = (1'h0);
  reg [(2'h3):(1'h0)] reg3937 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3936 = (1'h0);
  reg [(2'h3):(1'h0)] reg3935 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3934 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3933 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3932 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3931 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3930 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3929 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3928 = (1'h0);
  reg [(2'h3):(1'h0)] reg3927 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3926 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3922 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3921 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3925 = (1'h0);
  reg [(3'h7):(1'h0)] reg3924 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3923 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3922 = (1'h0);
  reg [(4'hd):(1'h0)] reg3921 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3920 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3919 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3918 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3917 = (1'h0);
  reg [(3'h6):(1'h0)] reg3916 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3915 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3914 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3913 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3912 = (1'h0);
  reg [(4'he):(1'h0)] reg3911 = (1'h0);
  reg [(4'hd):(1'h0)] reg3910 = (1'h0);
  reg [(4'he):(1'h0)] reg3909 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3908 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3907 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3906 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3905 = (1'h0);
  reg [(2'h2):(1'h0)] reg3904 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3903 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3902 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3901 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3900 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3899 = (1'h0);
  reg [(4'ha):(1'h0)] reg3898 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3897 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3896 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3895 = (1'h0);
  reg [(4'hf):(1'h0)] reg3894 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3893 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3892 = (1'h0);
  reg [(4'he):(1'h0)] reg3891 = (1'h0);
  reg [(3'h4):(1'h0)] reg3890 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3889 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3888 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3887 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3886 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3885 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3880 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3884 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3883 = (1'h0);
  reg [(2'h3):(1'h0)] reg3882 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3881 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3880 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3879 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3878 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3877 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3876 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3875 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3874 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3873 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3872 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3871 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3870 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3869 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3868 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3867 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3866 = (1'h0);
  reg [(4'h8):(1'h0)] reg3865 = (1'h0);
  reg [(4'hc):(1'h0)] reg3864 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3863 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3862 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3861 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3855 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3853 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3850 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3849 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3842 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3838 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3860 = (1'h0);
  reg [(4'he):(1'h0)] reg3859 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3858 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3857 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3856 = (1'h0);
  reg [(2'h3):(1'h0)] reg3855 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3854 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3853 = (1'h0);
  reg [(5'h10):(1'h0)] reg3852 = (1'h0);
  reg [(2'h3):(1'h0)] reg3851 = (1'h0);
  reg [(4'hf):(1'h0)] reg3850 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3849 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3848 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3847 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3843 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3847 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3846 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3845 = (1'h0);
  reg [(2'h3):(1'h0)] reg3844 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3843 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3841 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3837 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3836 = (1'h0);
  reg [(4'hc):(1'h0)] reg3842 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3841 = (1'h0);
  reg [(3'h5):(1'h0)] reg3840 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3839 = (1'h0);
  reg [(4'hb):(1'h0)] reg3838 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3837 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3836 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire3835;
  reg [(5'h10):(1'h0)] reg3834 = (1'h0);
  reg [(2'h3):(1'h0)] reg3833 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3832 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3824 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3821 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3819 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3818 = (1'h0);
  reg [(4'h9):(1'h0)] reg3831 = (1'h0);
  reg [(4'ha):(1'h0)] reg3830 = (1'h0);
  reg [(3'h4):(1'h0)] reg3829 = (1'h0);
  reg [(4'hc):(1'h0)] reg3828 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3827 = (1'h0);
  reg [(4'hc):(1'h0)] reg3826 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3825 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3824 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3823 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3822 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3821 = (1'h0);
  reg [(5'h10):(1'h0)] reg3820 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3819 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3818 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3817 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3816 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3815 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3814 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3813 = (1'h0);
  reg [(4'h9):(1'h0)] reg3812 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3811 = (1'h0);
  reg [(5'h10):(1'h0)] reg3810 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3809 = (1'h0);
  reg [(4'hf):(1'h0)] reg3808 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3807 = (1'h0);
  reg [(4'hf):(1'h0)] reg3806 = (1'h0);
  reg [(2'h2):(1'h0)] reg3805 = (1'h0);
  reg [(5'h10):(1'h0)] reg3804 = (1'h0);
  reg [(4'hc):(1'h0)] reg3803 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3802 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3801 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3801 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3800 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3799 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3798 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3797 = (1'h0);
  reg [(3'h4):(1'h0)] reg3796 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3795 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3794 = (1'h0);
  reg [(4'h9):(1'h0)] reg3793 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3792 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3791 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3790 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3789 = (1'h0);
  reg [(2'h3):(1'h0)] reg3788 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3787 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3786 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3785 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3784 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3783 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3782 = (1'h0);
  reg [(4'h8):(1'h0)] reg3781 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3780 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3779 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3778 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3777 = (1'h0);
  reg [(4'h9):(1'h0)] reg3776 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3775 = (1'h0);
  reg [(4'h9):(1'h0)] reg3774 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3773 = (1'h0);
  reg [(4'h8):(1'h0)] reg3772 = (1'h0);
  reg [(3'h6):(1'h0)] reg3771 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3770 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3769 = (1'h0);
  reg [(4'h8):(1'h0)] reg3768 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3767 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3766 = (1'h0);
  reg [(4'h8):(1'h0)] reg3765 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3764 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3763 = (1'h0);
  reg [(4'he):(1'h0)] reg3762 = (1'h0);
  reg [(2'h2):(1'h0)] reg3761 = (1'h0);
  reg [(3'h6):(1'h0)] reg3760 = (1'h0);
  reg [(4'hd):(1'h0)] reg3759 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3758 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3757 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3756 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3755 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3753 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3752 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3754 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3753 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3752 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3751 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3750 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3717 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3716 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3749 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3748 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3747 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3746 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3745 = (1'h0);
  reg [(3'h6):(1'h0)] reg3744 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3743 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3742 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3741 = (1'h0);
  reg [(3'h5):(1'h0)] reg3740 = (1'h0);
  reg [(4'hc):(1'h0)] reg3739 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3738 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3737 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3736 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3735 = (1'h0);
  reg [(3'h6):(1'h0)] reg3734 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3733 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3732 = (1'h0);
  reg [(2'h3):(1'h0)] reg3731 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3730 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3729 = (1'h0);
  reg [(4'hf):(1'h0)] reg3728 = (1'h0);
  reg [(2'h2):(1'h0)] reg3727 = (1'h0);
  reg [(2'h2):(1'h0)] reg3726 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3725 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3724 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3723 = (1'h0);
  reg [(3'h5):(1'h0)] reg3722 = (1'h0);
  reg [(4'hc):(1'h0)] reg3721 = (1'h0);
  reg [(4'hc):(1'h0)] reg3720 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3719 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3718 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3717 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3716 = (1'h0);
  reg [(4'h9):(1'h0)] reg3715 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3714 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3673 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3670 = (1'h0);
  reg [(4'he):(1'h0)] forvar3666 = (1'h0);
  reg [(4'ha):(1'h0)] reg3663 = (1'h0);
  reg [(2'h2):(1'h0)] reg3659 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3657 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3656 = (1'h0);
  reg [(4'hc):(1'h0)] reg3655 = (1'h0);
  reg [(3'h7):(1'h0)] reg3650 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3647 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3646 = (1'h0);
  reg [(3'h6):(1'h0)] reg3642 = (1'h0);
  reg [(3'h6):(1'h0)] reg3644 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3707 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3704 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3700 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3696 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3713 = (1'h0);
  reg [(2'h2):(1'h0)] reg3712 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3711 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3710 = (1'h0);
  reg [(3'h5):(1'h0)] reg3709 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3708 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3707 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3706 = (1'h0);
  reg [(4'ha):(1'h0)] reg3705 = (1'h0);
  reg [(4'hf):(1'h0)] reg3704 = (1'h0);
  reg [(4'h9):(1'h0)] reg3703 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3702 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3701 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3700 = (1'h0);
  reg [(4'he):(1'h0)] reg3699 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3698 = (1'h0);
  reg [(2'h3):(1'h0)] reg3697 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3696 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3695 = (1'h0);
  reg [(3'h4):(1'h0)] reg3694 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3693 = (1'h0);
  reg [(4'he):(1'h0)] forvar3692 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3689 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3687 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3684 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3682 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3678 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3691 = (1'h0);
  reg [(3'h7):(1'h0)] reg3690 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3689 = (1'h0);
  reg [(4'ha):(1'h0)] reg3688 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3687 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3686 = (1'h0);
  reg [(4'h9):(1'h0)] reg3685 = (1'h0);
  reg [(2'h3):(1'h0)] reg3684 = (1'h0);
  reg [(5'h10):(1'h0)] reg3683 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3682 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3681 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3680 = (1'h0);
  reg [(5'h10):(1'h0)] reg3679 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3678 = (1'h0);
  reg [(2'h2):(1'h0)] reg3677 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3676 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3675 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3674 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3673 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3672 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3671 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3670 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3669 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3668 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3667 = (1'h0);
  reg [(4'hb):(1'h0)] reg3666 = (1'h0);
  reg [(4'he):(1'h0)] reg3665 = (1'h0);
  reg [(4'hf):(1'h0)] reg3664 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3663 = (1'h0);
  reg [(4'he):(1'h0)] forvar3662 = (1'h0);
  reg [(4'hb):(1'h0)] reg3661 = (1'h0);
  reg [(4'hc):(1'h0)] reg3660 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3659 = (1'h0);
  reg [(2'h2):(1'h0)] reg3658 = (1'h0);
  reg [(4'he):(1'h0)] forvar3657 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3656 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3655 = (1'h0);
  reg [(3'h7):(1'h0)] reg3654 = (1'h0);
  reg [(4'h8):(1'h0)] reg3653 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3652 = (1'h0);
  reg [(4'h9):(1'h0)] reg3651 = (1'h0);
  reg [(4'he):(1'h0)] forvar3650 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3649 = (1'h0);
  reg [(4'hf):(1'h0)] reg3648 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3647 = (1'h0);
  reg [(3'h6):(1'h0)] reg3646 = (1'h0);
  reg [(2'h2):(1'h0)] reg3645 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3644 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3643 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3642 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3641 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3640 = (1'h0);
  reg [(2'h2):(1'h0)] reg3639 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3638 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3637 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3636 = (1'h0);
  wire [(4'ha):(1'h0)] wire3634;
  wire signed [(4'h8):(1'h0)] wire3633;
  wire [(5'h10):(1'h0)] wire3365;
  wire signed [(2'h3):(1'h0)] wire2167;
  wire [(4'he):(1'h0)] wire2166;
  wire [(4'hf):(1'h0)] wire2165;
  wire [(4'hf):(1'h0)] wire2164;
  wire signed [(4'he):(1'h0)] wire2162;
  wire signed [(4'hb):(1'h0)] wire1159;
  wire signed [(4'h9):(1'h0)] wire3631;
  assign y = {wire3992,
                 reg3991,
                 reg3990,
                 reg3989,
                 reg3988,
                 reg3987,
                 reg3986,
                 reg3985,
                 reg3984,
                 reg3983,
                 forvar3982,
                 forvar3981,
                 forvar3980,
                 forvar3975,
                 reg3979,
                 reg3978,
                 reg3977,
                 reg3976,
                 reg3975,
                 reg3974,
                 reg3973,
                 reg3972,
                 forvar3971,
                 reg3970,
                 reg3969,
                 reg3968,
                 reg3967,
                 reg3966,
                 forvar3965,
                 forvar3964,
                 reg3963,
                 reg3962,
                 reg3961,
                 reg3960,
                 reg3959,
                 forvar3958,
                 reg3957,
                 reg3956,
                 reg3955,
                 forvar3954,
                 forvar3953,
                 reg3952,
                 reg3951,
                 reg3950,
                 forvar3949,
                 reg3948,
                 reg3947,
                 reg3946,
                 forvar3945,
                 reg3944,
                 reg3943,
                 reg3942,
                 reg3941,
                 forvar3940,
                 forvar3939,
                 reg3887,
                 reg3886,
                 forvar3879,
                 forvar3882,
                 reg3877,
                 forvar3874,
                 reg3873,
                 reg3872,
                 forvar3869,
                 reg3868,
                 forvar3865,
                 reg3863,
                 reg3938,
                 reg3937,
                 reg3936,
                 reg3935,
                 reg3934,
                 forvar3933,
                 reg3932,
                 reg3931,
                 reg3930,
                 forvar3929,
                 reg3928,
                 reg3927,
                 forvar3926,
                 reg3922,
                 forvar3921,
                 reg3925,
                 reg3924,
                 reg3923,
                 forvar3922,
                 reg3921,
                 forvar3920,
                 reg3919,
                 reg3918,
                 forvar3917,
                 reg3916,
                 reg3915,
                 reg3914,
                 reg3913,
                 forvar3912,
                 reg3911,
                 reg3910,
                 reg3909,
                 reg3908,
                 reg3907,
                 reg3906,
                 reg3905,
                 reg3904,
                 forvar3903,
                 reg3902,
                 reg3901,
                 forvar3900,
                 reg3899,
                 reg3898,
                 forvar3897,
                 reg3896,
                 reg3895,
                 reg3894,
                 reg3893,
                 forvar3892,
                 reg3891,
                 reg3890,
                 reg3889,
                 forvar3888,
                 forvar3887,
                 forvar3886,
                 reg3885,
                 reg3880,
                 reg3884,
                 reg3883,
                 reg3882,
                 reg3881,
                 forvar3880,
                 reg3879,
                 reg3878,
                 forvar3877,
                 reg3876,
                 reg3875,
                 reg3874,
                 forvar3873,
                 forvar3872,
                 reg3871,
                 reg3870,
                 reg3869,
                 forvar3868,
                 reg3867,
                 reg3866,
                 reg3865,
                 reg3864,
                 forvar3863,
                 forvar3862,
                 forvar3861,
                 forvar3855,
                 reg3853,
                 forvar3850,
                 forvar3849,
                 forvar3842,
                 forvar3838,
                 reg3860,
                 reg3859,
                 reg3858,
                 reg3857,
                 reg3856,
                 reg3855,
                 reg3854,
                 forvar3853,
                 reg3852,
                 reg3851,
                 reg3850,
                 reg3849,
                 forvar3848,
                 forvar3847,
                 forvar3843,
                 reg3847,
                 reg3846,
                 reg3845,
                 reg3844,
                 reg3843,
                 reg3841,
                 reg3837,
                 forvar3836,
                 reg3842,
                 forvar3841,
                 reg3840,
                 reg3839,
                 reg3838,
                 forvar3837,
                 reg3836,
                 wire3835,
                 reg3834,
                 reg3833,
                 reg3832,
                 forvar3824,
                 reg3821,
                 forvar3819,
                 reg3818,
                 reg3831,
                 reg3830,
                 reg3829,
                 reg3828,
                 forvar3827,
                 reg3826,
                 reg3825,
                 reg3824,
                 reg3823,
                 reg3822,
                 forvar3821,
                 reg3820,
                 reg3819,
                 forvar3818,
                 forvar3817,
                 reg3816,
                 reg3815,
                 forvar3814,
                 reg3813,
                 reg3812,
                 forvar3811,
                 reg3810,
                 reg3809,
                 reg3808,
                 reg3807,
                 reg3806,
                 reg3805,
                 reg3804,
                 reg3803,
                 forvar3802,
                 forvar3801,
                 reg3801,
                 forvar3800,
                 reg3799,
                 reg3798,
                 reg3797,
                 reg3796,
                 reg3795,
                 reg3794,
                 reg3793,
                 reg3792,
                 forvar3791,
                 reg3790,
                 forvar3789,
                 reg3788,
                 reg3787,
                 reg3786,
                 reg3785,
                 reg3784,
                 reg3783,
                 forvar3782,
                 reg3781,
                 forvar3780,
                 forvar3779,
                 forvar3778,
                 reg3777,
                 reg3776,
                 reg3775,
                 reg3774,
                 reg3773,
                 reg3772,
                 reg3771,
                 forvar3770,
                 reg3769,
                 reg3768,
                 reg3767,
                 reg3766,
                 reg3765,
                 forvar3764,
                 forvar3763,
                 reg3762,
                 reg3761,
                 reg3760,
                 reg3759,
                 reg3758,
                 reg3757,
                 reg3756,
                 forvar3755,
                 forvar3753,
                 reg3752,
                 reg3754,
                 reg3753,
                 forvar3752,
                 forvar3751,
                 reg3750,
                 reg3717,
                 reg3716,
                 reg3749,
                 reg3748,
                 reg3747,
                 forvar3746,
                 reg3745,
                 reg3744,
                 reg3743,
                 forvar3742,
                 reg3741,
                 reg3740,
                 reg3739,
                 reg3738,
                 forvar3737,
                 reg3736,
                 reg3735,
                 reg3734,
                 reg3733,
                 forvar3732,
                 reg3731,
                 reg3730,
                 reg3729,
                 reg3728,
                 reg3727,
                 reg3726,
                 reg3725,
                 forvar3724,
                 reg3723,
                 reg3722,
                 reg3721,
                 reg3720,
                 forvar3719,
                 reg3718,
                 forvar3717,
                 forvar3716,
                 reg3715,
                 forvar3714,
                 reg3673,
                 forvar3670,
                 forvar3666,
                 reg3663,
                 reg3659,
                 reg3657,
                 reg3656,
                 reg3655,
                 reg3650,
                 forvar3647,
                 forvar3646,
                 reg3642,
                 reg3644,
                 reg3707,
                 forvar3704,
                 forvar3700,
                 reg3696,
                 reg3713,
                 reg3712,
                 reg3711,
                 reg3710,
                 reg3709,
                 forvar3708,
                 forvar3707,
                 reg3706,
                 reg3705,
                 reg3704,
                 reg3703,
                 reg3702,
                 reg3701,
                 reg3700,
                 reg3699,
                 reg3698,
                 reg3697,
                 forvar3696,
                 reg3695,
                 reg3694,
                 forvar3693,
                 forvar3692,
                 reg3689,
                 reg3687,
                 forvar3684,
                 reg3682,
                 forvar3678,
                 reg3691,
                 reg3690,
                 forvar3689,
                 reg3688,
                 forvar3687,
                 reg3686,
                 reg3685,
                 reg3684,
                 reg3683,
                 forvar3682,
                 reg3681,
                 reg3680,
                 reg3679,
                 reg3678,
                 reg3677,
                 reg3676,
                 reg3675,
                 reg3674,
                 forvar3673,
                 reg3672,
                 reg3671,
                 reg3670,
                 reg3669,
                 reg3668,
                 reg3667,
                 reg3666,
                 reg3665,
                 reg3664,
                 forvar3663,
                 forvar3662,
                 reg3661,
                 reg3660,
                 forvar3659,
                 reg3658,
                 forvar3657,
                 forvar3656,
                 forvar3655,
                 reg3654,
                 reg3653,
                 reg3652,
                 reg3651,
                 forvar3650,
                 reg3649,
                 reg3648,
                 reg3647,
                 reg3646,
                 reg3645,
                 forvar3644,
                 reg3643,
                 forvar3642,
                 forvar3641,
                 reg3640,
                 reg3639,
                 forvar3638,
                 forvar3637,
                 forvar3636,
                 wire3634,
                 wire3633,
                 wire3365,
                 wire2167,
                 wire2166,
                 wire2165,
                 wire2164,
                 wire2162,
                 wire1159,
                 wire3631,
                 (1'h0)};
  assign wire1159 = (($unsigned({(8'h9d)}) - {(wire1157 == wire1154)}) <= ((|wire1157[(4'ha):(1'h0)]) ?
                        ((wire1157 ^~ wire1158) ?
                            (~&(8'hb2)) : {wire1156}) : $signed((-wire1154))));
  module1160 modinst2163 (wire2162, clk, wire1157, wire1155, wire1156, wire1159);
  assign wire2164 = wire1158[(2'h2):(2'h2)];
  assign wire2165 = (!$unsigned(wire1159));
  assign wire2166 = wire1156[(4'ha):(4'ha)];
  assign wire2167 = (($signed((wire1158 ?
                            wire2166 : wire1154)) + $signed(((8'haa) != wire1154))) ?
                        (^~$unsigned($signed(wire1154))) : ((~^(wire1159 <<< wire1155)) ?
                            (wire1159 ?
                                {wire1154} : (wire2162 + wire1159)) : $unsigned(wire2165[(1'h0):(1'h0)])));
  module2168 modinst3366 (.y(wire3365), .clk(clk), .wire2171(wire2162), .wire2170(wire1156), .wire2169(wire1154), .wire2173(wire2164), .wire2172(wire1158));
  module3367 modinst3632 (.wire3370(wire1157), .clk(clk), .y(wire3631), .wire3371(wire1155), .wire3368(wire2166), .wire3372(wire3365), .wire3369(wire1154));
  assign wire3633 = $unsigned($signed((-wire1157)));
  module2367 modinst3635 (.wire2369(wire1155), .clk(clk), .wire2368(wire2165), .y(wire3634), .wire2370(wire1158), .wire2371(wire1157));
  always
    @(posedge clk) begin
      for (forvar3636 = (1'h0); (forvar3636 < (1'h0)); forvar3636 = (forvar3636 + (1'h1)))
        begin
          for (forvar3637 = (1'h0); (forvar3637 < (2'h3)); forvar3637 = (forvar3637 + (1'h1)))
            begin
              for (forvar3638 = (1'h0); (forvar3638 < (1'h1)); forvar3638 = (forvar3638 + (1'h1)))
                begin
                  if (wire3365[(3'h5):(1'h0)])
                    begin
                      reg3639 <= (^($signed($unsigned(wire1155)) << (wire3634[(3'h6):(2'h3)] != {(8'hb4)})));
                      reg3640 <= (((-wire3634) ?
                              ((&wire3365) ~^ (wire1159 ?
                                  reg3639 : wire1158)) : {forvar3636}) ?
                          wire1159[(4'ha):(3'h4)] : (^forvar3636));
                    end
                  else
                    begin
                      reg3639 <= $signed((~&$signed($unsigned(wire2166))));
                      reg3640 <= (~(wire3634[(2'h3):(1'h0)] || ((|forvar3638) ?
                          (!wire2162) : $signed(reg3639))));
                    end
                end
            end
        end
      if ($unsigned((~^$signed((^~wire3633)))))
        begin
          for (forvar3641 = (1'h0); (forvar3641 < (2'h2)); forvar3641 = (forvar3641 + (1'h1)))
            begin
              for (forvar3642 = (1'h0); (forvar3642 < (2'h2)); forvar3642 = (forvar3642 + (1'h1)))
                begin
                  reg3643 <= $signed((($unsigned(wire1154) ?
                          wire1157[(4'hc):(3'h6)] : wire1157) ?
                      $unsigned(wire1157) : ((wire1157 ? reg3639 : forvar3637) ?
                          (~^wire2165) : $unsigned(reg3639))));
                  for (forvar3644 = (1'h0); (forvar3644 < (2'h2)); forvar3644 = (forvar3644 + (1'h1)))
                    begin
                      reg3645 <= $signed($signed(reg3639));
                    end
                  if ((+(&wire1158[(4'hd):(4'hd)])))
                    begin
                      reg3646 <= (wire2165 ^~ $unsigned((forvar3636 ?
                          (reg3645 & wire1155) : (~(8'hb6)))));
                      reg3647 <= $signed(reg3643[(4'hd):(4'hd)]);
                      reg3648 <= ((&((forvar3636 ? forvar3637 : (8'ha4)) ?
                              (wire3365 & wire1154) : (forvar3641 + wire1155))) ?
                          wire3631 : $signed(((wire1154 ? wire3631 : wire1156) ?
                              (forvar3641 ? wire3631 : wire2166) : (reg3646 ?
                                  reg3645 : reg3643))));
                      reg3649 <= ($unsigned($unsigned((~wire1154))) != $signed((^{wire3365})));
                    end
                  else
                    begin
                      reg3646 <= wire2165[(4'ha):(4'ha)];
                    end
                  for (forvar3650 = (1'h0); (forvar3650 < (2'h2)); forvar3650 = (forvar3650 + (1'h1)))
                    begin
                      reg3651 <= wire2162;
                      reg3652 <= wire3631;
                      reg3653 <= $signed(reg3649[(4'h9):(1'h1)]);
                      reg3654 <= $unsigned(wire2164);
                    end
                end
            end
          for (forvar3655 = (1'h0); (forvar3655 < (2'h2)); forvar3655 = (forvar3655 + (1'h1)))
            begin
              for (forvar3656 = (1'h0); (forvar3656 < (2'h3)); forvar3656 = (forvar3656 + (1'h1)))
                begin
                  for (forvar3657 = (1'h0); (forvar3657 < (2'h3)); forvar3657 = (forvar3657 + (1'h1)))
                    begin
                      reg3658 <= (8'ha3);
                    end
                  for (forvar3659 = (1'h0); (forvar3659 < (1'h1)); forvar3659 = (forvar3659 + (1'h1)))
                    begin
                      reg3660 <= $signed(forvar3655);
                      reg3661 <= (((~&$signed(reg3646)) - reg3658) ?
                          wire1159[(4'h8):(1'h1)] : ($signed((forvar3650 || (8'ha9))) * (-wire2165[(1'h1):(1'h0)])));
                    end
                end
              for (forvar3662 = (1'h0); (forvar3662 < (1'h1)); forvar3662 = (forvar3662 + (1'h1)))
                begin
                  for (forvar3663 = (1'h0); (forvar3663 < (2'h2)); forvar3663 = (forvar3663 + (1'h1)))
                    begin
                      reg3664 <= reg3653;
                      reg3665 <= ((wire2166[(3'h6):(2'h3)] <= (~&reg3639[(1'h0):(1'h0)])) <<< (forvar3656[(2'h2):(2'h2)] ?
                          $unsigned($unsigned((8'hb3))) : $unsigned({forvar3655})));
                      reg3666 <= (8'hb9);
                      reg3667 <= ($signed((reg3666 ?
                              reg3646 : $signed(wire2166))) ?
                          (^$unsigned($signed(forvar3644))) : $signed({(8'hba)}));
                    end
                  if ((((~&wire2162[(4'h8):(2'h2)]) ~^ ((8'haf) ?
                          reg3661[(2'h3):(2'h2)] : wire1159)) ?
                      reg3658[(2'h2):(2'h2)] : reg3639[(2'h2):(1'h0)]))
                    begin
                      reg3668 <= $signed(($unsigned(reg3640) * forvar3644));
                      reg3669 <= (&((((8'hba) >= wire2166) ^ (forvar3637 || forvar3644)) ?
                          $unsigned(wire1158) : (&(wire3631 <<< reg3667))));
                      reg3670 <= {$signed(reg3643[(3'h5):(3'h5)])};
                      reg3671 <= $unsigned($unsigned(wire1159));
                    end
                  else
                    begin
                      reg3668 <= $signed((($signed(reg3654) * reg3665[(1'h1):(1'h1)]) ~^ $signed((8'hba))));
                    end
                  reg3672 <= (($signed($signed(wire2164)) << ($signed(reg3647) ?
                      forvar3656 : reg3654[(2'h3):(1'h1)])) == ((reg3669[(2'h2):(2'h2)] ?
                      {reg3653} : $unsigned(forvar3656)) && forvar3637[(4'hc):(2'h3)]));
                  for (forvar3673 = (1'h0); (forvar3673 < (1'h0)); forvar3673 = (forvar3673 + (1'h1)))
                    begin
                      reg3674 <= (($signed(forvar3650[(2'h3):(2'h2)]) << $signed((wire2164 || wire1159))) < $unsigned($unsigned(reg3639[(1'h0):(1'h0)])));
                      reg3675 <= {$signed((!$unsigned(reg3646)))};
                      reg3676 <= reg3665[(4'hc):(4'h9)];
                      reg3677 <= ((~|$unsigned(reg3660)) ?
                          (((wire2165 ? reg3649 : reg3652) ?
                                  ((8'haa) ?
                                      (8'haf) : wire3633) : $unsigned(reg3658)) ?
                              ((forvar3657 < reg3676) ?
                                  (wire2166 ?
                                      reg3652 : reg3665) : wire1156[(3'h5):(2'h2)]) : ({wire3634} ?
                                  {reg3670} : ((8'ha7) ?
                                      (8'hae) : wire1158))) : {((wire1157 && reg3640) < {reg3646})});
                    end
                end
              if ((($unsigned(reg3676) ?
                      (forvar3659[(2'h2):(2'h2)] >> reg3652[(3'h7):(3'h6)]) : {(wire2166 ^ reg3649)}) ?
                  $unsigned(((reg3643 ? forvar3656 : reg3674) ?
                      (|reg3668) : (reg3666 <= reg3651))) : $unsigned({$signed(forvar3662)})))
                begin
                  if (forvar3657[(1'h1):(1'h0)])
                    begin
                      reg3678 <= (reg3667[(2'h2):(2'h2)] ?
                          (((|(8'haa)) ?
                              reg3665[(2'h3):(2'h2)] : $signed((8'had))) > $unsigned((reg3643 ?
                              (8'h9d) : reg3645))) : $unsigned(((forvar3637 ?
                                  forvar3663 : (8'hb5)) ?
                              $signed(reg3648) : $unsigned(reg3666))));
                      reg3679 <= (~^reg3643[(2'h3):(2'h3)]);
                      reg3680 <= $signed(reg3669[(1'h1):(1'h0)]);
                      reg3681 <= (-(($signed(reg3670) ?
                          (reg3647 ^~ (8'ha8)) : $unsigned(wire1155)) << (-$unsigned(reg3661))));
                    end
                  else
                    begin
                      reg3678 <= (({$signed(reg3639)} ?
                          (|(wire2167 ^ reg3680)) : $unsigned($unsigned((8'ha8)))) >= $unsigned($unsigned((reg3669 ?
                          wire3365 : forvar3656))));
                      reg3679 <= (^reg3660[(3'h5):(2'h3)]);
                    end
                  for (forvar3682 = (1'h0); (forvar3682 < (2'h3)); forvar3682 = (forvar3682 + (1'h1)))
                    begin
                      reg3683 <= {($unsigned(reg3676) ?
                              {$unsigned(reg3660)} : wire2166)};
                      reg3684 <= forvar3659[(2'h2):(2'h2)];
                      reg3685 <= (+reg3674);
                      reg3686 <= wire3633[(2'h2):(1'h1)];
                    end
                  for (forvar3687 = (1'h0); (forvar3687 < (1'h1)); forvar3687 = (forvar3687 + (1'h1)))
                    begin
                      reg3688 <= $unsigned((wire3631 ?
                          reg3668[(3'h5):(1'h0)] : (^~(-wire1154))));
                    end
                  for (forvar3689 = (1'h0); (forvar3689 < (1'h0)); forvar3689 = (forvar3689 + (1'h1)))
                    begin
                      reg3690 <= (-reg3680);
                      reg3691 <= ((({wire1157} >>> $unsigned(reg3681)) ^~ $signed(forvar3650)) ?
                          (($unsigned(reg3651) ?
                              {reg3652} : (!reg3667)) >> forvar3659[(1'h0):(1'h0)]) : reg3665);
                    end
                end
              else
                begin
                  for (forvar3678 = (1'h0); (forvar3678 < (1'h1)); forvar3678 = (forvar3678 + (1'h1)))
                    begin
                      reg3679 <= wire2164[(3'h5):(3'h5)];
                      reg3680 <= ((({wire3633} ?
                                  ((8'ha9) ? reg3661 : (8'ha7)) : wire3365) ?
                              $unsigned(wire3633[(3'h7):(2'h2)]) : ($signed(forvar3682) >= wire1155)) ?
                          $signed(((reg3668 ? (8'ha3) : wire1155) ?
                              reg3667 : (forvar3655 >> (8'ha0)))) : (-(!(reg3686 ?
                              reg3665 : wire2166))));
                      reg3681 <= ($signed($unsigned(reg3646)) ?
                          (reg3649[(3'h6):(3'h6)] ~^ $signed($unsigned(reg3645))) : ((8'haa) ^~ ((~^reg3680) ?
                              (reg3667 <= reg3680) : (~|forvar3682))));
                      reg3682 <= ((+$signed((reg3681 ?
                          forvar3678 : reg3670))) + reg3681[(3'h7):(3'h6)]);
                    end
                  reg3683 <= $unsigned(forvar3689[(3'h4):(1'h1)]);
                  for (forvar3684 = (1'h0); (forvar3684 < (1'h1)); forvar3684 = (forvar3684 + (1'h1)))
                    begin
                      reg3685 <= reg3646;
                      reg3686 <= reg3675;
                    end
                  if (reg3678[(1'h0):(1'h0)])
                    begin
                      reg3687 <= reg3678;
                      reg3688 <= forvar3636[(2'h3):(2'h2)];
                      reg3689 <= (|$unsigned(wire1156));
                    end
                  else
                    begin
                      reg3687 <= (~^forvar3684[(4'h8):(1'h1)]);
                      reg3688 <= ($unsigned(reg3660) ^ wire1154[(4'h9):(2'h3)]);
                      reg3689 <= $unsigned(($unsigned({reg3674}) << (^wire1159)));
                    end
                end
              for (forvar3692 = (1'h0); (forvar3692 < (1'h0)); forvar3692 = (forvar3692 + (1'h1)))
                begin
                  for (forvar3693 = (1'h0); (forvar3693 < (1'h1)); forvar3693 = (forvar3693 + (1'h1)))
                    begin
                      reg3694 <= $signed((8'haf));
                      reg3695 <= $signed($unsigned($signed((8'ha7))));
                    end
                end
            end
          if (wire2166[(1'h1):(1'h1)])
            begin
              for (forvar3696 = (1'h0); (forvar3696 < (2'h2)); forvar3696 = (forvar3696 + (1'h1)))
                begin
                  if ((~$signed(wire2165)))
                    begin
                      reg3697 <= $signed((reg3690[(2'h2):(2'h2)] ?
                          $signed($signed((8'ha2))) : $unsigned(reg3658)));
                    end
                  else
                    begin
                      reg3697 <= reg3654;
                    end
                end
              if ((&reg3680[(1'h1):(1'h0)]))
                begin
                  reg3698 <= $signed(reg3660[(4'ha):(2'h3)]);
                end
              else
                begin
                  if ($unsigned($signed($unsigned($signed(forvar3663)))))
                    begin
                      reg3698 <= reg3672;
                      reg3699 <= ($unsigned((+(8'h9e))) ?
                          (reg3690 ?
                              (wire1156 >> (reg3654 != wire3631)) : reg3669[(3'h4):(3'h4)]) : $signed((~&(&(8'h9f)))));
                    end
                  else
                    begin
                      reg3698 <= reg3671[(3'h6):(1'h1)];
                      reg3699 <= wire1157[(2'h2):(2'h2)];
                    end
                  if (reg3688[(4'h9):(3'h5)])
                    begin
                      reg3700 <= (^reg3688[(3'h5):(1'h0)]);
                      reg3701 <= forvar3637;
                      reg3702 <= (reg3661 ?
                          forvar3655 : ($unsigned((forvar3638 ?
                                  forvar3644 : reg3667)) ?
                              (wire2165 ?
                                  (reg3701 * forvar3682) : $unsigned(forvar3682)) : $unsigned((!reg3640))));
                      reg3703 <= ($unsigned({(wire3634 + reg3653)}) ?
                          wire1157[(2'h3):(2'h3)] : $unsigned($unsigned($signed((8'ha2)))));
                    end
                  else
                    begin
                      reg3700 <= (wire1155[(1'h0):(1'h0)] ?
                          reg3643[(3'h5):(1'h0)] : reg3668[(3'h4):(1'h1)]);
                      reg3701 <= wire1158;
                      reg3702 <= ($unsigned({(reg3698 ?
                                  forvar3673 : (8'ha3))}) ?
                          $unsigned((reg3646 ?
                              forvar3637[(4'hb):(4'h9)] : (reg3703 ^ forvar3689))) : (((8'hae) <= (reg3669 >= reg3671)) - ({(8'h9d)} || reg3652[(3'h7):(2'h2)])));
                    end
                  if ((reg3687[(4'h9):(4'h8)] ^~ wire1159[(1'h1):(1'h0)]))
                    begin
                      reg3704 <= reg3694;
                      reg3705 <= (({reg3649[(3'h4):(2'h2)]} ?
                              reg3665 : {((8'h9d) ? (8'hac) : forvar3684)}) ?
                          $signed({(~|(8'ha6))}) : (($signed(reg3653) * (reg3697 || forvar3696)) ?
                              $unsigned((reg3643 >>> reg3678)) : forvar3693[(4'hb):(3'h5)]));
                      reg3706 <= (($unsigned(forvar3642) ?
                              (reg3677[(1'h1):(1'h1)] ?
                                  $unsigned(reg3695) : $unsigned(reg3660)) : (~(-reg3701))) ?
                          (8'ha2) : reg3661);
                    end
                  else
                    begin
                      reg3704 <= (8'ha6);
                      reg3705 <= reg3683[(2'h3):(2'h2)];
                      reg3706 <= {$signed($signed((wire3365 >> (8'h9c))))};
                    end
                end
              for (forvar3707 = (1'h0); (forvar3707 < (2'h3)); forvar3707 = (forvar3707 + (1'h1)))
                begin
                  for (forvar3708 = (1'h0); (forvar3708 < (1'h1)); forvar3708 = (forvar3708 + (1'h1)))
                    begin
                      reg3709 <= $unsigned((^(forvar3659[(2'h3):(1'h1)] ?
                          reg3671[(3'h5):(1'h1)] : (reg3704 <= (8'ha7)))));
                    end
                end
              if (forvar3656[(4'ha):(3'h4)])
                begin
                  if ($signed(wire2167[(1'h1):(1'h1)]))
                    begin
                      reg3710 <= (~&(^~reg3681[(1'h1):(1'h0)]));
                      reg3711 <= (reg3710 ? wire2166 : (reg3678 > (^wire3631)));
                      reg3712 <= $unsigned((!(reg3690[(3'h6):(2'h2)] ?
                          (reg3681 ?
                              wire1159 : (8'ha3)) : (reg3680 * reg3700))));
                      reg3713 <= ($signed((&reg3668)) && (~^(reg3652 ?
                          {forvar3638} : (forvar3662 ? reg3647 : reg3711))));
                    end
                  else
                    begin
                      reg3710 <= {(!($unsigned(reg3671) | (reg3703 ~^ wire3634)))};
                      reg3711 <= (&((8'hb6) > reg3660[(1'h0):(1'h0)]));
                      reg3712 <= reg3687;
                    end
                end
              else
                begin
                  if ($unsigned($unsigned($signed($signed(reg3666)))))
                    begin
                      reg3710 <= $signed((8'ha7));
                      reg3711 <= $unsigned($unsigned($unsigned($unsigned(reg3710))));
                      reg3712 <= reg3646[(3'h5):(1'h0)];
                      reg3713 <= wire3634[(4'ha):(1'h1)];
                    end
                  else
                    begin
                      reg3710 <= (&forvar3708[(2'h2):(1'h1)]);
                      reg3711 <= reg3676;
                      reg3712 <= ((^{$signed(wire3631)}) ?
                          (|((~&reg3645) >>> (^~reg3653))) : (~&(~&$signed(reg3668))));
                    end
                end
            end
          else
            begin
              if ((-forvar3637[(4'ha):(3'h6)]))
                begin
                  for (forvar3696 = (1'h0); (forvar3696 < (1'h0)); forvar3696 = (forvar3696 + (1'h1)))
                    begin
                      reg3697 <= $unsigned($unsigned($unsigned((reg3695 ?
                          wire1159 : reg3678))));
                    end
                end
              else
                begin
                  if ($signed($unsigned({$unsigned((8'h9e))})))
                    begin
                      reg3696 <= $unsigned((reg3651[(4'h9):(2'h3)] <<< (|$signed(reg3698))));
                    end
                  else
                    begin
                      reg3696 <= {($signed(reg3704) ?
                              $unsigned(wire3631[(4'h9):(4'h9)]) : $unsigned((reg3647 ?
                                  reg3679 : reg3660)))};
                      reg3697 <= $signed((({wire3633} ?
                              $unsigned(reg3675) : (wire2166 ?
                                  reg3698 : (8'hb6))) ?
                          (((8'hb7) && reg3705) ?
                              $unsigned(wire2162) : (8'ha5)) : $signed($signed((8'ha6)))));
                      reg3698 <= wire3365;
                      reg3699 <= reg3689[(1'h0):(1'h0)];
                    end
                end
              if ((8'hb9))
                begin
                  if (reg3645)
                    begin
                      reg3700 <= (8'hb0);
                      reg3701 <= (((reg3666 & forvar3656) ?
                              reg3675 : wire3631) ?
                          reg3699 : $unsigned(wire2164[(2'h3):(2'h3)]));
                      reg3702 <= reg3695;
                      reg3703 <= reg3712[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3700 <= ((~forvar3696) ?
                          ((~|forvar3682[(1'h0):(1'h0)]) ?
                              (reg3690[(2'h3):(2'h2)] ?
                                  (~|reg3675) : (reg3697 == reg3647)) : {wire1156[(4'ha):(2'h3)]}) : reg3652);
                      reg3701 <= ((8'hac) ?
                          reg3682 : $signed(reg3671[(3'h7):(1'h1)]));
                      reg3702 <= (wire2162 || (+{{forvar3655}}));
                    end
                  if ({($signed((+wire1158)) << $signed((~^reg3676)))})
                    begin
                      reg3704 <= $signed((reg3667[(4'h9):(1'h0)] ?
                          forvar3638 : wire1157));
                      reg3705 <= reg3690;
                      reg3706 <= $unsigned((forvar3655[(3'h7):(3'h7)] ?
                          forvar3696 : ($signed(forvar3673) ?
                              $unsigned(reg3645) : forvar3662[(4'h9):(4'h9)])));
                    end
                  else
                    begin
                      reg3704 <= $signed(forvar3707);
                    end
                end
              else
                begin
                  for (forvar3700 = (1'h0); (forvar3700 < (2'h3)); forvar3700 = (forvar3700 + (1'h1)))
                    begin
                      reg3701 <= {$unsigned($signed({reg3643}))};
                      reg3702 <= (^~$signed(($signed((8'ha3)) <= (&reg3652))));
                      reg3703 <= $signed((8'hb8));
                    end
                  for (forvar3704 = (1'h0); (forvar3704 < (1'h0)); forvar3704 = (forvar3704 + (1'h1)))
                    begin
                      reg3705 <= $unsigned($signed($unsigned((reg3696 ?
                          forvar3689 : reg3676))));
                    end
                end
              reg3707 <= {$signed(wire1156[(3'h5):(3'h5)])};
            end
        end
      else
        begin
          for (forvar3641 = (1'h0); (forvar3641 < (1'h0)); forvar3641 = (forvar3641 + (1'h1)))
            begin
              if ($unsigned($unsigned($signed((~&reg3712)))))
                begin
                  for (forvar3642 = (1'h0); (forvar3642 < (2'h2)); forvar3642 = (forvar3642 + (1'h1)))
                    begin
                      reg3643 <= {(reg3712 && {forvar3684})};
                      reg3644 <= $signed((((8'hb8) ?
                          (reg3699 <= wire3631) : ((8'h9f) ?
                              wire3631 : (8'hb8))) == (~&wire3633)));
                    end
                end
              else
                begin
                  reg3642 <= ({{forvar3692[(3'h4):(2'h3)]}} ?
                      ($unsigned(wire3365) | ({wire1158} ?
                          (reg3705 > reg3689) : $unsigned(reg3677))) : {$signed((-reg3712))});
                  if ((reg3711 != (8'ha4)))
                    begin
                      reg3643 <= (($unsigned({forvar3687}) ?
                          reg3648 : (8'h9e)) >> reg3713[(4'hc):(4'hb)]);
                      reg3644 <= ((~{forvar3693[(2'h2):(1'h0)]}) ?
                          reg3689 : $signed($signed((~&reg3639))));
                      reg3645 <= $signed((((forvar3678 ?
                              reg3709 : (8'ha5)) > (forvar3700 ?
                              reg3649 : reg3694)) ?
                          (&(reg3668 <<< forvar3708)) : reg3652[(4'h9):(2'h3)]));
                    end
                  else
                    begin
                      reg3643 <= $signed(forvar3707[(3'h6):(3'h6)]);
                      reg3644 <= reg3661;
                      reg3645 <= (+$signed((reg3682 ?
                          (forvar3684 ? reg3684 : reg3644) : wire1154)));
                    end
                end
              for (forvar3646 = (1'h0); (forvar3646 < (2'h3)); forvar3646 = (forvar3646 + (1'h1)))
                begin
                  for (forvar3647 = (1'h0); (forvar3647 < (1'h0)); forvar3647 = (forvar3647 + (1'h1)))
                    begin
                      reg3648 <= (8'hb2);
                      reg3649 <= (-(&(~|$unsigned(forvar3657))));
                      reg3650 <= ($unsigned($signed($unsigned(forvar3689))) ?
                          reg3690[(1'h1):(1'h1)] : $signed({reg3646[(3'h5):(2'h3)]}));
                    end
                  if ((8'hae))
                    begin
                      reg3651 <= (($signed($unsigned(reg3643)) ?
                          $signed(reg3702[(4'h8):(3'h7)]) : forvar3682) * ($signed({reg3661}) ?
                          reg3709[(2'h2):(2'h2)] : (reg3684 ^~ (reg3707 ?
                              forvar3704 : reg3689))));
                      reg3652 <= ({((reg3678 ^~ reg3713) ~^ (reg3643 ?
                                  reg3698 : forvar3682))} ?
                          {(((8'hae) ? reg3701 : reg3642) ?
                                  (wire3631 ?
                                      reg3696 : reg3711) : reg3669[(2'h3):(1'h1)])} : $unsigned(($signed((8'hba)) ?
                              (forvar3662 ?
                                  reg3684 : wire2162) : (~^reg3691))));
                      reg3653 <= ({reg3678[(2'h2):(2'h2)]} ?
                          {$signed((reg3658 == reg3688))} : ((8'hb5) ^~ ((-reg3680) ?
                              ((8'hba) >= reg3689) : ((8'hb8) + reg3689))));
                      reg3654 <= $unsigned(reg3691);
                    end
                  else
                    begin
                      reg3651 <= ((~((reg3640 ?
                              reg3660 : forvar3708) << (wire2166 ?
                              reg3658 : reg3667))) ?
                          reg3696[(3'h5):(1'h1)] : $unsigned({$signed((8'h9d))}));
                    end
                end
              if ($signed($unsigned(forvar3642)))
                begin
                  if ({$unsigned($unsigned((!(8'h9f))))})
                    begin
                      reg3655 <= $signed(forvar3707);
                      reg3656 <= ($unsigned(reg3691) ~^ $unsigned(forvar3642));
                      reg3657 <= (~|$signed(($unsigned(reg3688) ?
                          reg3654 : $signed(wire3631))));
                      reg3658 <= (&$signed((~&reg3680[(3'h5):(1'h1)])));
                    end
                  else
                    begin
                      reg3655 <= (reg3695 ?
                          reg3681[(2'h2):(2'h2)] : (&$unsigned($signed(forvar3684))));
                      reg3656 <= forvar3647[(3'h7):(3'h7)];
                      reg3657 <= ($signed((&(&(8'hb9)))) ?
                          ($signed((forvar3689 ? wire3631 : (8'hb4))) ?
                              $unsigned($unsigned(wire2162)) : $signed($signed(reg3640))) : ($signed($signed(wire1158)) * $unsigned($signed(reg3672))));
                      reg3658 <= (((~^$unsigned((8'hb2))) ?
                              (^~$signed(reg3668)) : reg3706) ?
                          reg3689[(1'h0):(1'h0)] : forvar3692);
                    end
                  if ((+$signed((~&(|reg3681)))))
                    begin
                      reg3659 <= (^~$unsigned($unsigned($signed(reg3683))));
                      reg3660 <= (|$signed($unsigned(reg3684)));
                      reg3661 <= (~^(((|reg3650) ?
                          $unsigned(forvar3684) : wire2167[(2'h2):(2'h2)]) && ((~|reg3670) ?
                          $unsigned(forvar3687) : {reg3711})));
                    end
                  else
                    begin
                      reg3659 <= forvar3692[(4'h8):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar3655 = (1'h0); (forvar3655 < (1'h1)); forvar3655 = (forvar3655 + (1'h1)))
                    begin
                      reg3656 <= {(($signed(forvar3638) ?
                                  $signed(reg3667) : forvar3682[(2'h2):(1'h1)]) ?
                              reg3646[(1'h1):(1'h0)] : $signed(forvar3663))};
                      reg3657 <= (!(forvar3684 != (^$unsigned(reg3684))));
                    end
                end
              for (forvar3662 = (1'h0); (forvar3662 < (1'h0)); forvar3662 = (forvar3662 + (1'h1)))
                begin
                  if ($signed(reg3650[(3'h7):(3'h4)]))
                    begin
                      reg3663 <= $unsigned($unsigned($signed($signed(reg3695))));
                      reg3664 <= $signed((8'hae));
                    end
                  else
                    begin
                      reg3663 <= (-reg3703[(4'h9):(4'h8)]);
                      reg3664 <= forvar3684[(1'h0):(1'h0)];
                      reg3665 <= ((forvar3689[(1'h1):(1'h0)] ?
                          $unsigned({reg3652}) : ((reg3683 ?
                              reg3667 : reg3660) ^ (-wire1157))) + {forvar3696});
                    end
                  for (forvar3666 = (1'h0); (forvar3666 < (1'h1)); forvar3666 = (forvar3666 + (1'h1)))
                    begin
                      reg3667 <= $signed(((^~$unsigned(wire1155)) ?
                          reg3696 : (((8'h9f) ? forvar3678 : wire3631) ?
                              (~^reg3699) : ((8'haf) ? reg3704 : (8'hb8)))));
                      reg3668 <= wire3365;
                      reg3669 <= $unsigned($signed((8'hb7)));
                    end
                  for (forvar3670 = (1'h0); (forvar3670 < (1'h1)); forvar3670 = (forvar3670 + (1'h1)))
                    begin
                      reg3671 <= $signed(forvar3663);
                      reg3672 <= ($signed(wire1154[(4'h9):(3'h7)]) < forvar3684);
                      reg3673 <= ($signed((~^((8'ha3) ? wire1158 : wire2166))) ?
                          forvar3644[(2'h3):(2'h2)] : (reg3653[(3'h5):(3'h4)] ?
                              (&$unsigned(forvar3670)) : reg3659));
                    end
                end
            end
        end
      for (forvar3714 = (1'h0); (forvar3714 < (2'h2)); forvar3714 = (forvar3714 + (1'h1)))
        begin
          if ((reg3679[(4'h9):(1'h0)] ?
              forvar3644[(3'h5):(2'h2)] : $unsigned($signed($signed((8'ha6))))))
            begin
              reg3715 <= (&$unsigned(((reg3654 ? forvar3657 : reg3711) ?
                  $unsigned(reg3639) : (reg3657 >>> wire1158))));
              for (forvar3716 = (1'h0); (forvar3716 < (2'h2)); forvar3716 = (forvar3716 + (1'h1)))
                begin
                  for (forvar3717 = (1'h0); (forvar3717 < (2'h2)); forvar3717 = (forvar3717 + (1'h1)))
                    begin
                      reg3718 <= $unsigned((&reg3672[(3'h5):(1'h1)]));
                    end
                  for (forvar3719 = (1'h0); (forvar3719 < (1'h0)); forvar3719 = (forvar3719 + (1'h1)))
                    begin
                      reg3720 <= reg3696[(3'h5):(2'h2)];
                      reg3721 <= forvar3663;
                      reg3722 <= $signed(forvar3659);
                      reg3723 <= (^$unsigned(reg3675));
                    end
                  for (forvar3724 = (1'h0); (forvar3724 < (1'h0)); forvar3724 = (forvar3724 + (1'h1)))
                    begin
                      reg3725 <= (wire2167[(2'h3):(2'h3)] >>> $unsigned(reg3647[(4'he):(4'hc)]));
                      reg3726 <= ((^~(!$signed(reg3654))) ?
                          $unsigned($signed($signed(reg3722))) : (+reg3715));
                      reg3727 <= (~&reg3673[(1'h0):(1'h0)]);
                      reg3728 <= ($signed((forvar3657[(4'he):(3'h6)] ?
                          ((8'ha7) ^~ wire1159) : $unsigned((8'ha1)))) << (($unsigned(reg3644) ?
                          (|reg3691) : $signed((8'ha8))) || reg3648));
                    end
                  if ((|$unsigned(forvar3638[(3'h6):(3'h4)])))
                    begin
                      reg3729 <= $unsigned({forvar3693});
                      reg3730 <= forvar3693;
                    end
                  else
                    begin
                      reg3729 <= reg3713;
                      reg3730 <= $signed($signed(forvar3673));
                      reg3731 <= {((reg3667[(2'h3):(1'h0)] ?
                                  (wire2164 ? reg3695 : (8'ha4)) : forvar3693) ?
                              $signed((forvar3692 ?
                                  reg3712 : reg3695)) : ((reg3674 <= reg3672) ?
                                  $signed(reg3697) : $unsigned(reg3709)))};
                    end
                end
              for (forvar3732 = (1'h0); (forvar3732 < (2'h2)); forvar3732 = (forvar3732 + (1'h1)))
                begin
                  if ({(~|reg3715)})
                    begin
                      reg3733 <= (($signed((reg3676 >>> wire1155)) ?
                          ({reg3677} << reg3639) : {reg3647}) >= reg3657);
                    end
                  else
                    begin
                      reg3733 <= (({{reg3648}} >= ((reg3671 ?
                              reg3640 : reg3696) << reg3713[(4'hb):(1'h0)])) ?
                          reg3688 : $unsigned((|$unsigned(reg3648))));
                    end
                  if (reg3689[(4'hb):(4'h8)])
                    begin
                      reg3734 <= $signed((~|$signed($signed(wire1156))));
                    end
                  else
                    begin
                      reg3734 <= ((^(^$unsigned((8'hb0)))) ?
                          reg3723[(3'h7):(1'h1)] : {(-(&reg3729))});
                      reg3735 <= (-reg3690[(3'h6):(3'h5)]);
                      reg3736 <= {{{$signed(reg3731)}}};
                    end
                  for (forvar3737 = (1'h0); (forvar3737 < (1'h0)); forvar3737 = (forvar3737 + (1'h1)))
                    begin
                      reg3738 <= (!(~&forvar3650[(4'hd):(2'h3)]));
                    end
                  if (forvar3687[(3'h7):(2'h3)])
                    begin
                      reg3739 <= reg3709;
                    end
                  else
                    begin
                      reg3739 <= $unsigned((~((reg3653 ?
                          reg3700 : reg3715) > wire1156)));
                      reg3740 <= ($unsigned(wire1158) >>> {((reg3699 ?
                              forvar3636 : reg3711) - {wire2162})});
                    end
                end
              if (($unsigned(((reg3738 >> reg3676) ?
                      $signed((8'hb9)) : (reg3712 ? wire1154 : reg3672))) ?
                  $unsigned(((wire3365 >>> (8'hb1)) ?
                      reg3683[(3'h4):(3'h4)] : reg3645[(1'h0):(1'h0)])) : $unsigned(reg3687)))
                begin
                  reg3741 <= forvar3641[(3'h5):(3'h4)];
                  for (forvar3742 = (1'h0); (forvar3742 < (1'h0)); forvar3742 = (forvar3742 + (1'h1)))
                    begin
                      reg3743 <= $signed($unsigned($unsigned($signed(forvar3708))));
                      reg3744 <= {$unsigned((^(~^forvar3742)))};
                      reg3745 <= (forvar3636 != (~((^~reg3668) ?
                          reg3647[(4'h9):(1'h1)] : (reg3715 ?
                              reg3743 : forvar3682))));
                    end
                  for (forvar3746 = (1'h0); (forvar3746 < (1'h1)); forvar3746 = (forvar3746 + (1'h1)))
                    begin
                      reg3747 <= forvar3650;
                      reg3748 <= wire3631;
                    end
                  reg3749 <= ((~($signed(reg3738) ?
                      (!wire2165) : (8'hb9))) && forvar3659[(1'h0):(1'h0)]);
                end
              else
                begin
                  reg3741 <= reg3677[(1'h0):(1'h0)];
                end
            end
          else
            begin
              if (($signed((8'hb4)) <= $unsigned($unsigned((reg3718 ?
                  (8'hac) : reg3667)))))
                begin
                  if ($unsigned(((~&(reg3740 ? forvar3704 : reg3691)) ?
                      (-(~|wire1154)) : $signed((-reg3660)))))
                    begin
                      reg3715 <= (($unsigned($unsigned(reg3706)) ?
                          {$signed(wire1157)} : ($signed(wire1158) <<< (~|forvar3717))) << $unsigned(forvar3659[(2'h3):(1'h0)]));
                      reg3716 <= ($signed($signed((wire1154 ?
                              reg3723 : (8'hb5)))) ?
                          ({reg3657[(3'h5):(3'h5)]} < ($unsigned(forvar3650) ?
                              (reg3744 == (8'hba)) : reg3650)) : {$unsigned($unsigned(reg3699))});
                      reg3717 <= ((((~|(8'ha0)) >= $unsigned((8'hb5))) ?
                              (8'ha3) : forvar3650[(3'h4):(1'h1)]) ?
                          $signed((^$signed(reg3741))) : reg3747);
                    end
                  else
                    begin
                      reg3715 <= (reg3734 == (reg3720[(3'h7):(3'h6)] >>> $unsigned((~&wire1157))));
                      reg3716 <= reg3713;
                    end
                  reg3718 <= (-{(~&reg3713)});
                  for (forvar3719 = (1'h0); (forvar3719 < (2'h3)); forvar3719 = (forvar3719 + (1'h1)))
                    begin
                      reg3720 <= $signed($signed((^reg3712)));
                    end
                  if (reg3669)
                    begin
                      reg3721 <= reg3730;
                      reg3722 <= (reg3735[(2'h2):(1'h0)] | (+{reg3712}));
                    end
                  else
                    begin
                      reg3721 <= reg3651[(3'h5):(2'h2)];
                    end
                end
              else
                begin
                  if ({reg3667})
                    begin
                      reg3715 <= ($signed(reg3712) ?
                          {reg3701} : $signed($signed((~(8'hb5)))));
                      reg3716 <= $unsigned((&reg3718[(3'h7):(1'h1)]));
                    end
                  else
                    begin
                      reg3715 <= {{((reg3678 && reg3669) < forvar3638)}};
                      reg3716 <= $unsigned((^{{reg3739}}));
                      reg3717 <= $signed(forvar3700);
                      reg3718 <= (~|$unsigned((&(forvar3708 > reg3661))));
                    end
                end
              reg3723 <= $unsigned(reg3720[(4'ha):(4'ha)]);
            end
        end
      reg3750 <= {(wire2164[(3'h4):(3'h4)] ?
              $unsigned(reg3645[(1'h0):(1'h0)]) : reg3658[(1'h0):(1'h0)])};
    end
  always
    @(posedge clk) begin
      for (forvar3751 = (1'h0); (forvar3751 < (2'h3)); forvar3751 = (forvar3751 + (1'h1)))
        begin
          if ($unsigned($unsigned($signed(reg3749))))
            begin
              if (reg3706[(1'h1):(1'h1)])
                begin
                  for (forvar3752 = (1'h0); (forvar3752 < (2'h2)); forvar3752 = (forvar3752 + (1'h1)))
                    begin
                      reg3753 <= ((^~(reg3750 & (-reg3654))) >= reg3749[(3'h7):(1'h1)]);
                      reg3754 <= $signed(reg3729[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  reg3752 <= (+$signed(forvar3708));
                  for (forvar3753 = (1'h0); (forvar3753 < (1'h1)); forvar3753 = (forvar3753 + (1'h1)))
                    begin
                      reg3754 <= ($unsigned(reg3640) <= $unsigned((+(reg3740 ?
                          reg3726 : reg3727))));
                    end
                end
            end
          else
            begin
              for (forvar3752 = (1'h0); (forvar3752 < (1'h1)); forvar3752 = (forvar3752 + (1'h1)))
                begin
                  for (forvar3753 = (1'h0); (forvar3753 < (2'h2)); forvar3753 = (forvar3753 + (1'h1)))
                    begin
                      reg3754 <= $signed($signed((^$unsigned(reg3748))));
                    end
                  for (forvar3755 = (1'h0); (forvar3755 < (1'h0)); forvar3755 = (forvar3755 + (1'h1)))
                    begin
                      reg3756 <= $unsigned(((reg3695[(3'h6):(1'h1)] ?
                              reg3740[(3'h4):(3'h4)] : $signed(reg3752)) ?
                          (forvar3704 ?
                              $signed(reg3748) : reg3720[(3'h7):(2'h3)]) : ({reg3695} ?
                              $signed(forvar3724) : $signed(forvar3656))));
                      reg3757 <= (~|{({reg3647} ?
                              (~&forvar3662) : (reg3712 ?
                                  reg3727 : forvar3641))});
                      reg3758 <= $signed((|$signed(reg3749)));
                    end
                  if ({(~|(reg3647 + {reg3745}))})
                    begin
                      reg3759 <= (($signed(forvar3657) * $signed({reg3758})) ?
                          reg3640[(3'h6):(2'h3)] : (!((~|forvar3638) + $signed(reg3682))));
                      reg3760 <= reg3694;
                      reg3761 <= $signed($unsigned(reg3668[(3'h4):(1'h0)]));
                      reg3762 <= ($unsigned(wire3633[(3'h6):(2'h2)]) ?
                          (($unsigned(reg3759) >> $signed(reg3657)) == ((^forvar3666) & $signed(reg3658))) : $signed(reg3640[(4'hb):(2'h3)]));
                    end
                  else
                    begin
                      reg3759 <= (|forvar3724[(2'h2):(2'h2)]);
                      reg3760 <= forvar3708;
                      reg3761 <= (($unsigned(reg3669) ?
                              $signed(reg3699[(3'h4):(2'h3)]) : reg3731[(1'h0):(1'h0)]) ?
                          ((reg3681 ? reg3747[(3'h5):(3'h5)] : reg3728) ?
                              $unsigned((8'haf)) : (reg3729[(3'h6):(3'h4)] << {reg3761})) : (~&reg3663));
                      reg3762 <= (($signed(reg3688[(1'h0):(1'h0)]) ^ forvar3644[(1'h1):(1'h1)]) | ($signed($signed(reg3727)) ?
                          reg3749[(1'h1):(1'h0)] : reg3645));
                    end
                end
              for (forvar3763 = (1'h0); (forvar3763 < (2'h3)); forvar3763 = (forvar3763 + (1'h1)))
                begin
                  for (forvar3764 = (1'h0); (forvar3764 < (2'h2)); forvar3764 = (forvar3764 + (1'h1)))
                    begin
                      reg3765 <= {forvar3673};
                      reg3766 <= ($unsigned(reg3727) && reg3734);
                      reg3767 <= reg3697;
                      reg3768 <= (((|{wire1158}) >> reg3739[(3'h4):(1'h1)]) != $unsigned(reg3756));
                    end
                  reg3769 <= reg3666[(4'h9):(4'h9)];
                  for (forvar3770 = (1'h0); (forvar3770 < (2'h2)); forvar3770 = (forvar3770 + (1'h1)))
                    begin
                      reg3771 <= (&wire2166[(4'hd):(3'h7)]);
                      reg3772 <= $signed(reg3744);
                      reg3773 <= $signed((({wire1154} ?
                          $signed((8'hb1)) : forvar3751) & {{forvar3673}}));
                      reg3774 <= forvar3763;
                    end
                  if ((forvar3678 == ((8'ha1) ?
                      forvar3751[(4'h8):(1'h0)] : (~wire1158))))
                    begin
                      reg3775 <= $signed($signed($signed($signed(reg3758))));
                      reg3776 <= (($unsigned($signed(forvar3755)) & ((^forvar3650) ~^ {reg3773})) <= ({forvar3670} < reg3664));
                    end
                  else
                    begin
                      reg3775 <= reg3655;
                      reg3776 <= $signed((forvar3642[(2'h2):(1'h1)] ?
                          (wire1159[(4'h8):(3'h7)] ?
                              (forvar3670 ? forvar3704 : reg3661) : (reg3645 ?
                                  wire1159 : (8'hb5))) : $signed((forvar3742 ~^ reg3727))));
                      reg3777 <= (reg3664[(4'hc):(3'h5)] ?
                          ((~(reg3685 || reg3762)) >= wire3365[(1'h1):(1'h1)]) : {wire1154});
                    end
                end
            end
          for (forvar3778 = (1'h0); (forvar3778 < (2'h3)); forvar3778 = (forvar3778 + (1'h1)))
            begin
              for (forvar3779 = (1'h0); (forvar3779 < (2'h3)); forvar3779 = (forvar3779 + (1'h1)))
                begin
                  for (forvar3780 = (1'h0); (forvar3780 < (1'h1)); forvar3780 = (forvar3780 + (1'h1)))
                    begin
                      reg3781 <= $unsigned($signed(((reg3753 ?
                              reg3758 : forvar3693) ?
                          (reg3639 > forvar3732) : {wire1158})));
                    end
                  for (forvar3782 = (1'h0); (forvar3782 < (2'h2)); forvar3782 = (forvar3782 + (1'h1)))
                    begin
                      reg3783 <= (($unsigned(reg3694) & (~^$unsigned(forvar3684))) ?
                          (8'h9d) : forvar3693);
                    end
                  reg3784 <= (reg3750 ?
                      $unsigned(((reg3727 <= (8'hab)) ?
                          (~|reg3776) : wire1154[(3'h7):(3'h7)])) : $unsigned($signed(reg3669[(1'h1):(1'h0)])));
                  if ((&reg3652))
                    begin
                      reg3785 <= reg3717[(2'h3):(1'h0)];
                      reg3786 <= $unsigned(((^(reg3678 ?
                          reg3679 : reg3769)) & $signed((forvar3692 ?
                          (8'h9f) : reg3726))));
                      reg3787 <= $unsigned((reg3711 || reg3720));
                    end
                  else
                    begin
                      reg3785 <= $unsigned($signed($unsigned((^reg3721))));
                      reg3786 <= ($signed(forvar3644) ?
                          (((forvar3693 * reg3660) ?
                                  $unsigned(reg3736) : reg3697[(1'h0):(1'h0)]) ?
                              ($signed(forvar3782) <<< (~^forvar3737)) : (~(~&forvar3707))) : ((^reg3784[(4'h8):(3'h4)]) != (|{forvar3716})));
                      reg3787 <= reg3700[(1'h0):(1'h0)];
                      reg3788 <= reg3720[(4'hb):(3'h7)];
                    end
                end
              for (forvar3789 = (1'h0); (forvar3789 < (2'h2)); forvar3789 = (forvar3789 + (1'h1)))
                begin
                  reg3790 <= ({{$unsigned(forvar3763)}} + $unsigned(((^~reg3668) != $unsigned(forvar3689))));
                end
              for (forvar3791 = (1'h0); (forvar3791 < (1'h0)); forvar3791 = (forvar3791 + (1'h1)))
                begin
                  if (($signed(reg3711) * $signed((~|$unsigned(reg3661)))))
                    begin
                      reg3792 <= forvar3684[(2'h3):(1'h1)];
                      reg3793 <= $unsigned((((reg3769 ?
                              reg3686 : wire1154) ^ reg3750) ?
                          $signed((forvar3637 ?
                              reg3712 : forvar3636)) : (^$unsigned(reg3753))));
                    end
                  else
                    begin
                      reg3792 <= $signed(reg3672[(4'h8):(3'h5)]);
                      reg3793 <= (8'hac);
                      reg3794 <= (~&(^~($unsigned(wire3633) || (forvar3637 ?
                          reg3694 : forvar3789))));
                      reg3795 <= reg3792[(2'h3):(2'h3)];
                    end
                  if ($unsigned((^~reg3704)))
                    begin
                      reg3796 <= $signed((reg3659 ?
                          (forvar3704 ?
                              $unsigned(reg3786) : forvar3684) : $unsigned(reg3728)));
                      reg3797 <= $signed(($unsigned((reg3781 ?
                              reg3661 : reg3749)) ?
                          ($signed(reg3690) ?
                              (forvar3746 ?
                                  forvar3770 : forvar3673) : reg3715) : ((reg3666 >>> reg3739) ^ (-reg3790))));
                    end
                  else
                    begin
                      reg3796 <= (8'haa);
                      reg3797 <= $signed(($unsigned((8'h9d)) ?
                          reg3698[(1'h1):(1'h0)] : {(reg3750 ?
                                  (8'hb8) : reg3743)}));
                    end
                end
              reg3798 <= {($signed(forvar3662[(4'hd):(3'h5)]) ?
                      ({wire2167} ?
                          reg3689[(4'hb):(4'hb)] : wire1156[(2'h2):(1'h1)]) : {{forvar3752}})};
            end
          reg3799 <= reg3670[(4'h9):(3'h4)];
        end
      for (forvar3800 = (1'h0); (forvar3800 < (2'h3)); forvar3800 = (forvar3800 + (1'h1)))
        begin
          if (($signed((~&$signed(reg3674))) ?
              ($unsigned((^~reg3715)) ?
                  {((8'haf) ?
                          reg3640 : forvar3682)} : reg3651[(2'h2):(1'h1)]) : forvar3764[(1'h1):(1'h1)]))
            begin
              reg3801 <= ($signed(reg3668[(2'h2):(2'h2)]) < ((8'ha6) ?
                  reg3657 : (reg3727[(1'h1):(1'h0)] & forvar3751)));
            end
          else
            begin
              for (forvar3801 = (1'h0); (forvar3801 < (1'h1)); forvar3801 = (forvar3801 + (1'h1)))
                begin
                  for (forvar3802 = (1'h0); (forvar3802 < (1'h1)); forvar3802 = (forvar3802 + (1'h1)))
                    begin
                      reg3803 <= reg3695[(3'h4):(1'h0)];
                      reg3804 <= reg3696;
                      reg3805 <= (reg3689 >> forvar3655[(4'h8):(3'h6)]);
                      reg3806 <= $signed(((wire2167 == reg3717) ?
                          (!(!reg3768)) : $signed({forvar3682})));
                    end
                  reg3807 <= (|(reg3721[(3'h6):(3'h4)] > reg3743));
                  if (($unsigned(reg3667) * (({(8'ha6)} ?
                          (reg3690 ? reg3681 : wire1155) : $unsigned(reg3652)) ?
                      forvar3752 : $signed(((8'ha6) >= reg3761)))))
                    begin
                      reg3808 <= (((forvar3673 ^ (reg3659 ?
                              reg3673 : wire3634)) ?
                          wire2167[(1'h0):(1'h0)] : reg3640[(4'h9):(1'h0)]) >> $unsigned({((8'ha2) >= wire1157)}));
                      reg3809 <= reg3741;
                    end
                  else
                    begin
                      reg3808 <= forvar3657;
                      reg3809 <= (((8'hb4) >> ($unsigned(reg3723) << $signed(reg3677))) ?
                          $unsigned(reg3793[(1'h1):(1'h1)]) : $signed(reg3747));
                      reg3810 <= $signed(reg3677[(1'h0):(1'h0)]);
                    end
                  for (forvar3811 = (1'h0); (forvar3811 < (2'h2)); forvar3811 = (forvar3811 + (1'h1)))
                    begin
                      reg3812 <= $unsigned($unsigned($unsigned((8'h9c))));
                    end
                end
              reg3813 <= $unsigned(($signed(forvar3659[(3'h4):(2'h2)]) ?
                  forvar3678[(4'h9):(1'h0)] : {$unsigned(reg3758)}));
              for (forvar3814 = (1'h0); (forvar3814 < (2'h3)); forvar3814 = (forvar3814 + (1'h1)))
                begin
                  reg3815 <= $signed({(reg3804 <= {reg3807})});
                  reg3816 <= {forvar3719};
                end
            end
          for (forvar3817 = (1'h0); (forvar3817 < (2'h3)); forvar3817 = (forvar3817 + (1'h1)))
            begin
              if (reg3794)
                begin
                  for (forvar3818 = (1'h0); (forvar3818 < (2'h2)); forvar3818 = (forvar3818 + (1'h1)))
                    begin
                      reg3819 <= forvar3636[(2'h2):(2'h2)];
                      reg3820 <= {$unsigned(((~|reg3704) <<< forvar3696))};
                    end
                  for (forvar3821 = (1'h0); (forvar3821 < (1'h1)); forvar3821 = (forvar3821 + (1'h1)))
                    begin
                      reg3822 <= (reg3660[(1'h0):(1'h0)] ?
                          (~&$unsigned((reg3804 < forvar3696))) : ((~^{reg3694}) >> (^~(reg3695 ?
                              reg3653 : reg3643))));
                      reg3823 <= ($signed($unsigned((forvar3770 ?
                          forvar3687 : reg3679))) | $signed(reg3792[(4'h8):(3'h4)]));
                    end
                  if (reg3790)
                    begin
                      reg3824 <= $unsigned($unsigned($unsigned(reg3823)));
                      reg3825 <= (^reg3677);
                    end
                  else
                    begin
                      reg3824 <= wire1157;
                      reg3825 <= ($unsigned((~$unsigned(reg3799))) * ((8'haf) == $signed((forvar3641 ?
                          reg3772 : reg3776))));
                      reg3826 <= forvar3673[(3'h6):(1'h1)];
                    end
                  for (forvar3827 = (1'h0); (forvar3827 < (2'h2)); forvar3827 = (forvar3827 + (1'h1)))
                    begin
                      reg3828 <= $unsigned($unsigned($signed($unsigned(forvar3814))));
                      reg3829 <= reg3741[(3'h5):(2'h3)];
                      reg3830 <= (forvar3814 ?
                          {((reg3684 ?
                                  (8'hb3) : reg3727) * reg3774[(4'h9):(1'h1)])} : reg3799[(3'h6):(2'h3)]);
                      reg3831 <= ((-forvar3716[(2'h2):(2'h2)]) ?
                          (8'h9e) : reg3786);
                    end
                end
              else
                begin
                  reg3818 <= reg3819[(1'h0):(1'h0)];
                  for (forvar3819 = (1'h0); (forvar3819 < (2'h3)); forvar3819 = (forvar3819 + (1'h1)))
                    begin
                      reg3820 <= $signed((((^~reg3820) >> (reg3754 && (8'haa))) <= reg3687[(4'hd):(3'h6)]));
                      reg3821 <= ({(!$signed(wire2165))} ?
                          $signed((~^(forvar3752 ^ reg3711))) : ({$signed((8'haf))} ?
                              (^~reg3762) : $signed((8'hb8))));
                      reg3822 <= $unsigned($unsigned(reg3775[(2'h2):(1'h0)]));
                      reg3823 <= reg3653;
                    end
                  for (forvar3824 = (1'h0); (forvar3824 < (2'h2)); forvar3824 = (forvar3824 + (1'h1)))
                    begin
                      reg3825 <= reg3682;
                      reg3826 <= ({($signed(reg3665) ?
                              (reg3705 ^ forvar3819) : (reg3808 << forvar3687))} == ($signed($signed(forvar3724)) ^ {(~(8'hac))}));
                    end
                end
              reg3832 <= $signed($signed($signed(reg3741[(1'h1):(1'h1)])));
            end
          reg3833 <= (^reg3666);
          reg3834 <= reg3819;
        end
    end
  assign wire3835 = reg3728[(4'hb):(3'h5)];
  always
    @(posedge clk) begin
      if (($unsigned(forvar3656) > (((forvar3657 > reg3640) || (reg3834 ?
              reg3769 : forvar3678)) ?
          {$signed(reg3783)} : $signed((reg3740 && reg3786)))))
        begin
          if (({$signed(reg3743)} ?
              $signed((^(~reg3807))) : (~^{(reg3765 ^~ reg3752)})))
            begin
              if (($unsigned(reg3738[(3'h5):(3'h4)]) ?
                  reg3691[(4'hc):(2'h3)] : reg3664))
                begin
                  reg3836 <= $signed((~&forvar3678));
                  for (forvar3837 = (1'h0); (forvar3837 < (1'h0)); forvar3837 = (forvar3837 + (1'h1)))
                    begin
                      reg3838 <= $signed((^~$unsigned($unsigned(reg3781))));
                    end
                  if (({{(|forvar3801)}} ^ reg3774))
                    begin
                      reg3839 <= {{($unsigned(forvar3719) * forvar3666)}};
                    end
                  else
                    begin
                      reg3839 <= forvar3789[(2'h3):(1'h1)];
                      reg3840 <= (($signed((forvar3764 ? reg3794 : (8'ha0))) ?
                              ((reg3722 ?
                                  reg3639 : reg3676) <<< (^~reg3725)) : (~(forvar3666 ~^ forvar3657))) ?
                          $unsigned((forvar3753 == reg3678)) : (!$signed(reg3663)));
                    end
                  for (forvar3841 = (1'h0); (forvar3841 < (1'h0)); forvar3841 = (forvar3841 + (1'h1)))
                    begin
                      reg3842 <= reg3661[(4'h8):(3'h6)];
                    end
                end
              else
                begin
                  for (forvar3836 = (1'h0); (forvar3836 < (2'h3)); forvar3836 = (forvar3836 + (1'h1)))
                    begin
                      reg3837 <= wire2162[(4'he):(4'he)];
                      reg3838 <= $signed(forvar3841);
                      reg3839 <= $unsigned((8'ha6));
                    end
                  if ($signed((^(reg3803[(2'h3):(2'h2)] ^~ {(8'h9e)}))))
                    begin
                      reg3840 <= (reg3677[(1'h1):(1'h0)] + forvar3670[(4'h9):(3'h5)]);
                      reg3841 <= (wire2166 || (reg3788[(2'h2):(2'h2)] ?
                          ((reg3785 ?
                              reg3775 : forvar3637) ^ (~&reg3769)) : forvar3682[(2'h2):(1'h1)]));
                      reg3842 <= $signed($signed($unsigned({reg3695})));
                      reg3843 <= forvar3687[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3840 <= {reg3733[(3'h5):(2'h3)]};
                      reg3841 <= (reg3760[(2'h2):(1'h1)] == $signed({wire2165[(4'h9):(3'h6)]}));
                      reg3842 <= $unsigned((((reg3715 ?
                              reg3767 : reg3706) + forvar3687[(3'h4):(2'h2)]) ?
                          (^~$signed(reg3838)) : ({reg3794} > $signed(reg3820))));
                      reg3843 <= (8'hb7);
                    end
                  if (($signed(((forvar3801 << forvar3659) ?
                      reg3793 : $unsigned(reg3796))) && $unsigned({(+reg3685)})))
                    begin
                      reg3844 <= ((reg3753[(1'h1):(1'h1)] | reg3707) == reg3716);
                      reg3845 <= (($signed($signed(reg3805)) ?
                              ((forvar3737 > reg3762) >= (reg3793 ^ reg3663)) : {(+forvar3717)}) ?
                          (forvar3778[(3'h6):(3'h5)] ?
                              reg3834[(4'ha):(3'h5)] : ($unsigned(wire1158) ^ $unsigned(forvar3707))) : $unsigned((wire2166[(3'h6):(2'h2)] ~^ reg3841[(4'hf):(4'h9)])));
                      reg3846 <= reg3747;
                    end
                  else
                    begin
                      reg3844 <= wire1156[(4'hc):(4'ha)];
                      reg3845 <= forvar3791[(1'h1):(1'h0)];
                      reg3846 <= ((8'hab) ?
                          (8'ha0) : forvar3811[(4'h8):(4'h8)]);
                      reg3847 <= reg3706[(1'h1):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar3836 = (1'h0); (forvar3836 < (1'h0)); forvar3836 = (forvar3836 + (1'h1)))
                begin
                  for (forvar3837 = (1'h0); (forvar3837 < (1'h1)); forvar3837 = (forvar3837 + (1'h1)))
                    begin
                      reg3838 <= {reg3696[(3'h5):(3'h4)]};
                      reg3839 <= $unsigned((^reg3736));
                      reg3840 <= {{$unsigned((forvar3824 + reg3716))}};
                      reg3841 <= (+(forvar3707 | $unsigned($unsigned(reg3847))));
                    end
                  reg3842 <= {(-$unsigned($unsigned(wire1158)))};
                  for (forvar3843 = (1'h0); (forvar3843 < (2'h2)); forvar3843 = (forvar3843 + (1'h1)))
                    begin
                      reg3844 <= (~((wire1155[(2'h3):(2'h3)] ^ ((8'haa) ?
                          reg3700 : reg3822)) * (reg3795[(3'h4):(1'h0)] ?
                          $signed(reg3767) : $signed(forvar3818))));
                      reg3845 <= $unsigned(((reg3717 ?
                          ((8'hb2) ? reg3756 : reg3707) : (reg3820 ?
                              reg3718 : (8'h9f))) >>> (^$unsigned((8'hb6)))));
                      reg3846 <= (reg3828[(2'h2):(2'h2)] <= ($unsigned((reg3734 ?
                              reg3830 : forvar3824)) ?
                          ((^~reg3820) ~^ reg3701) : {reg3706[(3'h5):(2'h2)]}));
                    end
                end
              for (forvar3847 = (1'h0); (forvar3847 < (1'h0)); forvar3847 = (forvar3847 + (1'h1)))
                begin
                  for (forvar3848 = (1'h0); (forvar3848 < (2'h2)); forvar3848 = (forvar3848 + (1'h1)))
                    begin
                      reg3849 <= ({$signed(forvar3763[(1'h1):(1'h1)])} ?
                          {{(forvar3666 ?
                                      (8'hb4) : (8'had))}} : {$signed(forvar3637[(3'h6):(1'h1)])});
                    end
                  if ($unsigned((~|$signed({reg3656}))))
                    begin
                      reg3850 <= reg3759;
                      reg3851 <= (~^(($unsigned(reg3820) ^~ (8'hb3)) >= $unsigned({reg3716})));
                      reg3852 <= (({reg3710} ^~ (~(8'ha2))) ?
                          (&((|reg3699) ?
                              (reg3650 >= reg3655) : $unsigned((8'hba)))) : reg3807);
                    end
                  else
                    begin
                      reg3850 <= (&forvar3752[(1'h0):(1'h0)]);
                    end
                  for (forvar3853 = (1'h0); (forvar3853 < (1'h1)); forvar3853 = (forvar3853 + (1'h1)))
                    begin
                      reg3854 <= {$unsigned(((-forvar3673) ?
                              (8'hba) : reg3698[(2'h2):(1'h1)]))};
                      reg3855 <= ($signed((~(reg3690 <<< reg3830))) ^~ reg3806);
                      reg3856 <= (reg3670[(1'h0):(1'h0)] ?
                          ((8'hb6) || $signed(wire1158[(1'h0):(1'h0)])) : (+reg3645[(1'h0):(1'h0)]));
                      reg3857 <= $signed((reg3783[(2'h3):(1'h0)] ^~ reg3819[(2'h3):(1'h0)]));
                    end
                  if (($unsigned(((~^forvar3684) ?
                      {(8'ha0)} : (forvar3737 * reg3667))) != $signed((^~(^(8'ha9))))))
                    begin
                      reg3858 <= (8'h9e);
                      reg3859 <= wire2165[(4'hd):(1'h0)];
                    end
                  else
                    begin
                      reg3858 <= (8'ha4);
                      reg3859 <= ({reg3721} >> reg3808[(4'he):(4'ha)]);
                      reg3860 <= forvar3843[(1'h1):(1'h0)];
                    end
                end
            end
        end
      else
        begin
          for (forvar3836 = (1'h0); (forvar3836 < (1'h0)); forvar3836 = (forvar3836 + (1'h1)))
            begin
              for (forvar3837 = (1'h0); (forvar3837 < (1'h1)); forvar3837 = (forvar3837 + (1'h1)))
                begin
                  for (forvar3838 = (1'h0); (forvar3838 < (1'h0)); forvar3838 = (forvar3838 + (1'h1)))
                    begin
                      reg3839 <= {(^~(^~$signed(reg3829)))};
                      reg3840 <= (|((^~((8'haf) ? (8'hb1) : reg3730)) ?
                          reg3701 : reg3680));
                    end
                end
            end
          if ((8'ha2))
            begin
              for (forvar3841 = (1'h0); (forvar3841 < (1'h0)); forvar3841 = (forvar3841 + (1'h1)))
                begin
                  for (forvar3842 = (1'h0); (forvar3842 < (2'h2)); forvar3842 = (forvar3842 + (1'h1)))
                    begin
                      reg3843 <= (((8'hb9) >>> {(reg3842 ?
                                  reg3759 : reg3812)}) ?
                          ($signed(forvar3827) - (~|$unsigned(forvar3764))) : $signed({(forvar3746 ?
                                  reg3665 : reg3698)}));
                      reg3844 <= $unsigned($unsigned(forvar3636[(1'h1):(1'h1)]));
                      reg3845 <= (!$unsigned($signed((^forvar3838))));
                    end
                end
            end
          else
            begin
              for (forvar3841 = (1'h0); (forvar3841 < (2'h2)); forvar3841 = (forvar3841 + (1'h1)))
                begin
                  for (forvar3842 = (1'h0); (forvar3842 < (2'h2)); forvar3842 = (forvar3842 + (1'h1)))
                    begin
                      reg3843 <= $signed(({(reg3818 | reg3754)} != $signed((reg3659 ?
                          reg3825 : reg3855))));
                      reg3844 <= (~&$unsigned(forvar3780[(2'h3):(2'h3)]));
                      reg3845 <= (~|(!$signed($unsigned((8'hb7)))));
                      reg3846 <= $signed($signed(((forvar3824 || (8'h9d)) ?
                          (forvar3737 ?
                              forvar3637 : reg3768) : reg3801[(2'h2):(1'h0)])));
                    end
                  reg3847 <= reg3666[(3'h6):(1'h1)];
                end
            end
          for (forvar3848 = (1'h0); (forvar3848 < (2'h2)); forvar3848 = (forvar3848 + (1'h1)))
            begin
              for (forvar3849 = (1'h0); (forvar3849 < (2'h2)); forvar3849 = (forvar3849 + (1'h1)))
                begin
                  for (forvar3850 = (1'h0); (forvar3850 < (1'h1)); forvar3850 = (forvar3850 + (1'h1)))
                    begin
                      reg3851 <= $unsigned(((8'hb8) ^ $signed((reg3668 ?
                          reg3651 : forvar3779))));
                    end
                  if ($unsigned((reg3851[(2'h3):(2'h2)] & $unsigned((~|forvar3684)))))
                    begin
                      reg3852 <= $signed({{(reg3750 - reg3843)}});
                      reg3853 <= reg3702;
                      reg3854 <= (($signed((reg3674 ? reg3840 : (8'ha8))) ?
                          forvar3670 : forvar3714) <<< forvar3811[(3'h7):(3'h4)]);
                    end
                  else
                    begin
                      reg3852 <= reg3760[(3'h6):(2'h2)];
                    end
                  for (forvar3855 = (1'h0); (forvar3855 < (2'h2)); forvar3855 = (forvar3855 + (1'h1)))
                    begin
                      reg3856 <= reg3823;
                    end
                  reg3857 <= $signed(reg3799[(3'h5):(1'h1)]);
                end
            end
          reg3858 <= (~|(($unsigned(forvar3708) ?
              (^reg3777) : forvar3657[(1'h0):(1'h0)]) == ((~|reg3808) ~^ (reg3678 < forvar3801))));
        end
      if ($signed(reg3793[(4'h8):(2'h2)]))
        begin
          for (forvar3861 = (1'h0); (forvar3861 < (2'h2)); forvar3861 = (forvar3861 + (1'h1)))
            begin
              for (forvar3862 = (1'h0); (forvar3862 < (2'h3)); forvar3862 = (forvar3862 + (1'h1)))
                begin
                  for (forvar3863 = (1'h0); (forvar3863 < (2'h3)); forvar3863 = (forvar3863 + (1'h1)))
                    begin
                      reg3864 <= ((reg3792[(4'h8):(1'h0)] ?
                          $signed((|reg3688)) : ($signed(reg3833) & reg3720[(3'h4):(1'h1)])) | wire2164);
                      reg3865 <= ($unsigned(reg3685) ?
                          (reg3758 ?
                              reg3822 : forvar3746) : $unsigned((~|reg3706[(2'h2):(1'h1)])));
                      reg3866 <= (^~$signed(((^~forvar3853) ?
                          $signed(wire2167) : (reg3787 ~^ wire2166))));
                      reg3867 <= $unsigned(reg3656[(3'h5):(2'h2)]);
                    end
                  for (forvar3868 = (1'h0); (forvar3868 < (2'h2)); forvar3868 = (forvar3868 + (1'h1)))
                    begin
                      reg3869 <= (reg3801 ?
                          (((&reg3839) ? {reg3851} : reg3769[(2'h3):(1'h1)]) ?
                              {(!reg3824)} : reg3734[(1'h0):(1'h0)]) : {reg3783[(1'h0):(1'h0)]});
                    end
                  reg3870 <= ({($unsigned(reg3864) != (^reg3815))} ?
                      reg3776[(3'h5):(1'h0)] : reg3663[(3'h4):(2'h2)]);
                  reg3871 <= ($unsigned(((forvar3850 || reg3781) + (~|forvar3753))) ~^ forvar3678);
                end
              for (forvar3872 = (1'h0); (forvar3872 < (1'h1)); forvar3872 = (forvar3872 + (1'h1)))
                begin
                  for (forvar3873 = (1'h0); (forvar3873 < (2'h2)); forvar3873 = (forvar3873 + (1'h1)))
                    begin
                      reg3874 <= forvar3753[(2'h3):(2'h2)];
                      reg3875 <= ($signed({reg3783}) & (!reg3843));
                      reg3876 <= (~|reg3810);
                    end
                end
              if (reg3667[(4'hb):(4'ha)])
                begin
                  for (forvar3877 = (1'h0); (forvar3877 < (1'h1)); forvar3877 = (forvar3877 + (1'h1)))
                    begin
                      reg3878 <= {forvar3819[(2'h2):(1'h1)]};
                      reg3879 <= $unsigned($unsigned((reg3709 ?
                          ((8'ha5) + reg3870) : reg3831)));
                    end
                  for (forvar3880 = (1'h0); (forvar3880 < (1'h1)); forvar3880 = (forvar3880 + (1'h1)))
                    begin
                      reg3881 <= $unsigned(((+(^~(8'ha0))) ~^ (-$signed(reg3642))));
                      reg3882 <= ($signed((|reg3819[(3'h7):(3'h5)])) ?
                          ((+$signed((8'hba))) || ($signed(reg3740) >>> (^~forvar3753))) : $unsigned((reg3660 & reg3722)));
                      reg3883 <= $signed($unsigned(reg3851));
                      reg3884 <= ((({reg3843} ?
                              forvar3818[(2'h2):(1'h1)] : reg3740) ?
                          (forvar3708 && (|forvar3861)) : (~reg3836)) << $unsigned($signed(reg3858)));
                    end
                end
              else
                begin
                  for (forvar3877 = (1'h0); (forvar3877 < (2'h2)); forvar3877 = (forvar3877 + (1'h1)))
                    begin
                      reg3878 <= $signed($unsigned(reg3669[(2'h3):(1'h0)]));
                    end
                  reg3879 <= (+((+reg3675[(2'h3):(1'h1)]) + $signed($signed(reg3642))));
                  if ($unsigned((~&{(~|reg3744)})))
                    begin
                      reg3880 <= ({$signed(reg3707)} ?
                          (&($unsigned(reg3866) ?
                              $unsigned(reg3679) : forvar3868[(4'hb):(2'h2)])) : (&(~^(forvar3678 + reg3699))));
                      reg3881 <= (8'hb1);
                    end
                  else
                    begin
                      reg3880 <= $unsigned((~^(~&forvar3663)));
                      reg3881 <= ($unsigned($signed($signed(reg3837))) ?
                          (8'ha3) : {(8'h9d)});
                      reg3882 <= $signed($signed((!(+reg3671))));
                    end
                end
            end
          reg3885 <= ($unsigned((|$unsigned(forvar3877))) ?
              forvar3638[(4'hd):(2'h2)] : ({(-(8'hb6))} && $signed($unsigned((8'hab)))));
          for (forvar3886 = (1'h0); (forvar3886 < (2'h2)); forvar3886 = (forvar3886 + (1'h1)))
            begin
              for (forvar3887 = (1'h0); (forvar3887 < (2'h2)); forvar3887 = (forvar3887 + (1'h1)))
                begin
                  for (forvar3888 = (1'h0); (forvar3888 < (2'h2)); forvar3888 = (forvar3888 + (1'h1)))
                    begin
                      reg3889 <= wire2164[(4'hb):(3'h6)];
                      reg3890 <= $unsigned((reg3867[(1'h1):(1'h0)] || ($unsigned(reg3658) ?
                          $unsigned((8'ha4)) : (~^reg3653))));
                      reg3891 <= $signed(($signed(reg3765[(1'h1):(1'h0)]) ?
                          wire3835[(4'hd):(4'hd)] : reg3857));
                    end
                  for (forvar3892 = (1'h0); (forvar3892 < (1'h0)); forvar3892 = (forvar3892 + (1'h1)))
                    begin
                      reg3893 <= $signed(($unsigned((^(8'hac))) ?
                          forvar3892[(1'h1):(1'h1)] : reg3668));
                    end
                  if (((+{(forvar3663 ? (8'haa) : forvar3791)}) ?
                      reg3694 : forvar3689[(2'h2):(2'h2)]))
                    begin
                      reg3894 <= $unsigned((^~(~&((8'hb4) ?
                          forvar3850 : reg3824))));
                    end
                  else
                    begin
                      reg3894 <= $unsigned(reg3750);
                      reg3895 <= $signed(wire1157);
                      reg3896 <= reg3761;
                    end
                  for (forvar3897 = (1'h0); (forvar3897 < (2'h3)); forvar3897 = (forvar3897 + (1'h1)))
                    begin
                      reg3898 <= ((~&reg3823[(1'h1):(1'h1)]) ?
                          reg3845[(1'h1):(1'h0)] : reg3674);
                      reg3899 <= $signed($unsigned({$unsigned(reg3864)}));
                    end
                end
              for (forvar3900 = (1'h0); (forvar3900 < (2'h2)); forvar3900 = (forvar3900 + (1'h1)))
                begin
                  if ((((-reg3783) ?
                      reg3843[(4'h8):(3'h5)] : (reg3698 ?
                          (reg3722 ? reg3651 : forvar3888) : (reg3735 ?
                              (8'ha0) : reg3845))) <<< ((^~reg3768[(2'h3):(2'h2)]) != ($signed(reg3871) < $unsigned(reg3810)))))
                    begin
                      reg3901 <= forvar3873;
                    end
                  else
                    begin
                      reg3901 <= forvar3887;
                      reg3902 <= reg3890[(2'h3):(2'h3)];
                    end
                end
              for (forvar3903 = (1'h0); (forvar3903 < (1'h0)); forvar3903 = (forvar3903 + (1'h1)))
                begin
                  if ({$unsigned($signed(reg3713))})
                    begin
                      reg3904 <= $unsigned(reg3668);
                      reg3905 <= (~reg3843);
                      reg3906 <= forvar3666[(2'h3):(2'h3)];
                      reg3907 <= $signed($signed({$unsigned(reg3905)}));
                    end
                  else
                    begin
                      reg3904 <= forvar3737;
                    end
                  if ($signed(((&$unsigned(wire2167)) ?
                      (~&(forvar3877 < forvar3821)) : forvar3847[(3'h5):(1'h0)])))
                    begin
                      reg3908 <= $unsigned(($signed(forvar3684[(3'h6):(3'h5)]) < {reg3893}));
                      reg3909 <= $signed($unsigned(((forvar3708 <= forvar3693) == forvar3647[(4'h9):(3'h5)])));
                      reg3910 <= {{(-reg3798)}};
                      reg3911 <= reg3851[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3908 <= (reg3796 ?
                          (&($signed(reg3829) ~^ $unsigned(reg3777))) : reg3832);
                      reg3909 <= ((forvar3872[(4'hd):(3'h7)] ?
                          ((8'ha6) | reg3781[(1'h0):(1'h0)]) : reg3712) | $signed(reg3905[(2'h3):(1'h1)]));
                      reg3910 <= reg3690[(1'h1):(1'h1)];
                    end
                  for (forvar3912 = (1'h0); (forvar3912 < (1'h1)); forvar3912 = (forvar3912 + (1'h1)))
                    begin
                      reg3913 <= ((((reg3910 ? reg3696 : forvar3892) ?
                                  reg3758 : {reg3860}) ?
                              $unsigned((~^forvar3853)) : (-(wire3634 >> reg3845))) ?
                          $unsigned((|(reg3899 ?
                              (8'hb4) : reg3658))) : $signed(($signed(reg3667) ?
                              $signed((8'hb5)) : (~forvar3837))));
                      reg3914 <= reg3642;
                      reg3915 <= (reg3819[(1'h1):(1'h0)] ?
                          ((reg3730[(1'h0):(1'h0)] ?
                              (~&(8'hb7)) : (forvar3717 == reg3684)) >>> forvar3888[(3'h5):(1'h0)]) : $unsigned($signed((reg3674 - reg3654))));
                      reg3916 <= $unsigned((8'ha7));
                    end
                  for (forvar3917 = (1'h0); (forvar3917 < (2'h2)); forvar3917 = (forvar3917 + (1'h1)))
                    begin
                      reg3918 <= $signed($signed(reg3781[(3'h7):(2'h3)]));
                      reg3919 <= (|(reg3844 ^ reg3653));
                    end
                end
            end
          for (forvar3920 = (1'h0); (forvar3920 < (1'h0)); forvar3920 = (forvar3920 + (1'h1)))
            begin
              if ($signed($signed(($unsigned(forvar3814) ?
                  $unsigned(reg3907) : (forvar3877 ? (8'ha5) : reg3830)))))
                begin
                  reg3921 <= $unsigned((~^reg3831[(1'h0):(1'h0)]));
                  for (forvar3922 = (1'h0); (forvar3922 < (1'h0)); forvar3922 = (forvar3922 + (1'h1)))
                    begin
                      reg3923 <= ($unsigned(wire3631[(1'h1):(1'h0)]) ?
                          $unsigned(reg3883[(3'h5):(1'h1)]) : (($signed(forvar3827) - $unsigned(forvar3684)) <= (~reg3830)));
                      reg3924 <= $unsigned($unsigned($unsigned((reg3652 << reg3860))));
                      reg3925 <= ($unsigned(reg3760) < $unsigned((-$signed(reg3772))));
                    end
                end
              else
                begin
                  for (forvar3921 = (1'h0); (forvar3921 < (2'h3)); forvar3921 = (forvar3921 + (1'h1)))
                    begin
                      reg3922 <= (((~&$unsigned(reg3808)) <= forvar3779) ?
                          $signed(((reg3722 ? reg3884 : (8'hb9)) ?
                              {reg3743} : (reg3663 - reg3853))) : (+reg3867[(1'h0):(1'h0)]));
                      reg3923 <= $unsigned((reg3792 ?
                          forvar3863 : (((8'hb7) << (8'hab)) * $unsigned(reg3788))));
                      reg3924 <= (wire2165 ?
                          (reg3726[(1'h0):(1'h0)] ?
                              reg3833 : forvar3850[(2'h3):(1'h1)]) : ((|((8'hb2) ?
                              reg3773 : (8'hb1))) | $unsigned(reg3721[(2'h3):(2'h3)])));
                      reg3925 <= reg3667;
                    end
                  for (forvar3926 = (1'h0); (forvar3926 < (2'h3)); forvar3926 = (forvar3926 + (1'h1)))
                    begin
                      reg3927 <= (-{$unsigned(((8'hba) ? reg3658 : reg3740))});
                      reg3928 <= wire3365;
                    end
                end
              for (forvar3929 = (1'h0); (forvar3929 < (1'h1)); forvar3929 = (forvar3929 + (1'h1)))
                begin
                  if (forvar3704[(3'h4):(1'h0)])
                    begin
                      reg3930 <= reg3825;
                      reg3931 <= (($signed((~&(8'ha8))) ^ reg3841[(3'h5):(3'h4)]) ?
                          ((((8'hb8) == wire1155) ?
                              $signed(reg3758) : ((8'ha9) + reg3781)) * ((reg3728 * reg3787) > $unsigned(reg3830))) : {$signed($signed(reg3700))});
                    end
                  else
                    begin
                      reg3930 <= (-reg3865);
                      reg3931 <= (8'ha4);
                      reg3932 <= $signed($unsigned(((~&(8'h9c)) ^~ (+reg3786))));
                    end
                  for (forvar3933 = (1'h0); (forvar3933 < (2'h2)); forvar3933 = (forvar3933 + (1'h1)))
                    begin
                      reg3934 <= reg3816;
                      reg3935 <= (^~reg3806[(3'h6):(3'h4)]);
                      reg3936 <= $signed($signed((~&$unsigned(reg3881))));
                    end
                end
              reg3937 <= ({((reg3750 == reg3907) ?
                          (|(8'ha0)) : $unsigned(forvar3657))} ?
                  reg3828[(4'h9):(3'h7)] : $signed((~^(reg3909 ~^ reg3745))));
              reg3938 <= $signed($signed(($signed(reg3840) ^ $signed(reg3927))));
            end
        end
      else
        begin
          for (forvar3861 = (1'h0); (forvar3861 < (1'h0)); forvar3861 = (forvar3861 + (1'h1)))
            begin
              for (forvar3862 = (1'h0); (forvar3862 < (2'h2)); forvar3862 = (forvar3862 + (1'h1)))
                begin
                  if (reg3830[(4'h8):(2'h2)])
                    begin
                      reg3863 <= $unsigned(forvar3853);
                    end
                  else
                    begin
                      reg3863 <= {$signed(reg3703[(3'h6):(1'h0)])};
                      reg3864 <= forvar3724;
                    end
                  for (forvar3865 = (1'h0); (forvar3865 < (1'h1)); forvar3865 = (forvar3865 + (1'h1)))
                    begin
                      reg3866 <= (forvar3770 ?
                          {((+reg3882) ?
                                  $unsigned(reg3657) : (reg3839 | (8'hb2)))} : reg3870[(4'hd):(3'h4)]);
                      reg3867 <= reg3720[(1'h0):(1'h0)];
                      reg3868 <= reg3703[(3'h6):(2'h3)];
                    end
                  for (forvar3869 = (1'h0); (forvar3869 < (1'h1)); forvar3869 = (forvar3869 + (1'h1)))
                    begin
                      reg3870 <= (8'h9c);
                      reg3871 <= (reg3858[(3'h4):(3'h4)] * (^~forvar3872[(2'h2):(1'h1)]));
                      reg3872 <= $unsigned((({(8'hb2)} ?
                              $unsigned(forvar3644) : (~&forvar3789)) ?
                          $unsigned(reg3870[(4'h9):(2'h3)]) : (reg3881 ^~ forvar3666)));
                      reg3873 <= $unsigned({((~^reg3684) ?
                              (-reg3670) : reg3740[(2'h2):(1'h0)])});
                    end
                end
              if (reg3765)
                begin
                  for (forvar3874 = (1'h0); (forvar3874 < (2'h2)); forvar3874 = (forvar3874 + (1'h1)))
                    begin
                      reg3875 <= ((($unsigned(reg3650) ?
                                  reg3785 : $signed((8'ha3))) ?
                              wire3365 : reg3808[(4'hb):(1'h1)]) ?
                          $unsigned((^~((8'ha7) ?
                              reg3781 : reg3804))) : $signed(reg3674[(2'h3):(2'h2)]));
                      reg3876 <= {forvar3684};
                    end
                  reg3877 <= (~&(~&($unsigned(reg3657) ?
                      (^~reg3918) : reg3890)));
                  if ((!(^{$signed(reg3759)})))
                    begin
                      reg3878 <= {(((forvar3659 == reg3703) ~^ $unsigned(reg3649)) ?
                              (8'hab) : forvar3641)};
                    end
                  else
                    begin
                      reg3878 <= ($unsigned(reg3660) || (+$unsigned((reg3878 >>> reg3656))));
                      reg3879 <= {forvar3814};
                      reg3880 <= {((~^(reg3720 ? forvar3638 : reg3685)) ?
                              forvar3865[(2'h2):(1'h1)] : reg3729[(3'h6):(1'h1)])};
                      reg3881 <= wire1159;
                    end
                  for (forvar3882 = (1'h0); (forvar3882 < (2'h2)); forvar3882 = (forvar3882 + (1'h1)))
                    begin
                      reg3883 <= ((8'hb4) <<< reg3646);
                      reg3884 <= (((-reg3664[(3'h5):(2'h2)]) ?
                              {$unsigned(reg3710)} : forvar3892[(2'h2):(1'h0)]) ?
                          ({(wire1157 ? reg3874 : reg3656)} ?
                              reg3859 : (~^{wire3633})) : (reg3691[(3'h6):(2'h2)] ?
                              $signed((reg3858 || reg3851)) : reg3774));
                      reg3885 <= reg3655;
                    end
                end
              else
                begin
                  for (forvar3874 = (1'h0); (forvar3874 < (1'h1)); forvar3874 = (forvar3874 + (1'h1)))
                    begin
                      reg3875 <= $signed($signed((-$signed((8'hab)))));
                      reg3876 <= reg3727;
                      reg3877 <= {reg3822[(3'h4):(1'h0)]};
                    end
                  reg3878 <= ($signed(((reg3863 ?
                          (8'hb9) : reg3699) || (-reg3882))) ?
                      $signed(((8'had) || (8'hba))) : $signed($signed($unsigned((8'hae)))));
                  for (forvar3879 = (1'h0); (forvar3879 < (2'h3)); forvar3879 = (forvar3879 + (1'h1)))
                    begin
                      reg3880 <= ((((forvar3666 ?
                                  forvar3779 : wire2164) != (^~forvar3707)) ?
                              ($signed(reg3739) ?
                                  ((8'ha8) * wire3835) : (-(8'hb1))) : (forvar3638 | (+wire1155))) ?
                          forvar3861 : $signed(($signed(reg3899) ?
                              (reg3839 > reg3832) : reg3659[(2'h2):(1'h0)])));
                      reg3881 <= ((|$unsigned(reg3844[(1'h1):(1'h0)])) ?
                          (8'ha5) : $unsigned(($unsigned(forvar3656) && (reg3922 ?
                              wire2162 : reg3767))));
                    end
                end
            end
          reg3886 <= ($signed({(+reg3804)}) - forvar3817);
          reg3887 <= ($signed((~$unsigned(reg3757))) << ($unsigned((reg3652 && (8'h9d))) ~^ reg3860));
        end
      for (forvar3939 = (1'h0); (forvar3939 < (2'h3)); forvar3939 = (forvar3939 + (1'h1)))
        begin
          for (forvar3940 = (1'h0); (forvar3940 < (2'h3)); forvar3940 = (forvar3940 + (1'h1)))
            begin
              if ((reg3715[(4'h9):(4'h9)] ?
                  (reg3765 >= $signed(reg3752[(4'h8):(1'h0)])) : ({(reg3691 ?
                          reg3659 : forvar3873)} <= $signed((8'ha3)))))
                begin
                  if ($signed($signed(reg3910)))
                    begin
                      reg3941 <= $signed(($signed($signed(forvar3929)) && (8'hb5)));
                      reg3942 <= (^~{(!((8'hb4) << reg3786))});
                      reg3943 <= reg3682[(1'h0):(1'h0)];
                      reg3944 <= ((forvar3655[(3'h6):(1'h0)] ?
                          reg3669[(1'h0):(1'h0)] : ($signed(reg3713) || $unsigned(forvar3716))) ^ $signed((~&(forvar3646 ?
                          reg3813 : forvar3655))));
                    end
                  else
                    begin
                      reg3941 <= (|forvar3912);
                      reg3942 <= $unsigned(reg3713[(1'h1):(1'h1)]);
                      reg3943 <= {(~^forvar3887[(2'h3):(1'h0)])};
                      reg3944 <= $signed(reg3705);
                    end
                end
              else
                begin
                  if ($unsigned((8'hb0)))
                    begin
                      reg3941 <= (reg3657[(2'h2):(2'h2)] ^ (forvar3861[(3'h5):(1'h0)] ?
                          $unsigned((+(8'hb9))) : $signed((forvar3862 ?
                              reg3793 : (8'ha3)))));
                    end
                  else
                    begin
                      reg3941 <= $signed((~$unsigned((reg3775 ?
                          (8'h9e) : reg3783))));
                      reg3942 <= (reg3884[(3'h5):(3'h5)] ?
                          (reg3729[(4'ha):(4'h9)] ?
                              (~|$signed(reg3887)) : ((reg3752 ~^ wire1159) ?
                                  (forvar3684 ?
                                      reg3726 : (8'ha8)) : $signed(reg3849))) : ($unsigned(reg3921[(2'h3):(2'h3)]) >= (reg3846 ^~ reg3694)));
                      reg3943 <= ((~(8'ha1)) * (|{(~&reg3875)}));
                      reg3944 <= {$unsigned(reg3775)};
                    end
                  for (forvar3945 = (1'h0); (forvar3945 < (2'h2)); forvar3945 = (forvar3945 + (1'h1)))
                    begin
                      reg3946 <= $signed((8'h9e));
                      reg3947 <= ({wire1157} + $unsigned(reg3902[(4'ha):(4'h9)]));
                      reg3948 <= (+(~&($signed(forvar3719) ?
                          reg3695 : $signed(reg3691))));
                    end
                  for (forvar3949 = (1'h0); (forvar3949 < (1'h1)); forvar3949 = (forvar3949 + (1'h1)))
                    begin
                      reg3950 <= ($unsigned($signed((reg3738 >>> reg3777))) & forvar3641[(3'h4):(2'h2)]);
                      reg3951 <= {reg3752};
                      reg3952 <= (~^(reg3776 - $signed((reg3758 - (8'ha4)))));
                    end
                end
            end
          for (forvar3953 = (1'h0); (forvar3953 < (1'h1)); forvar3953 = (forvar3953 + (1'h1)))
            begin
              for (forvar3954 = (1'h0); (forvar3954 < (1'h1)); forvar3954 = (forvar3954 + (1'h1)))
                begin
                  if ($signed((({wire1157} ?
                      {reg3666} : $unsigned(reg3887)) + $signed($unsigned((8'hb8))))))
                    begin
                      reg3955 <= forvar3818[(3'h6):(2'h2)];
                      reg3956 <= $unsigned({({reg3880} ?
                              (|reg3735) : (reg3941 ? wire1157 : reg3786))});
                      reg3957 <= $signed($unsigned((-(reg3739 > reg3868))));
                    end
                  else
                    begin
                      reg3955 <= $signed($unsigned(($unsigned(forvar3861) ?
                          reg3870 : (8'h9c))));
                      reg3956 <= $signed($unsigned(wire2167));
                      reg3957 <= $unsigned(forvar3763[(5'h10):(4'h8)]);
                    end
                  for (forvar3958 = (1'h0); (forvar3958 < (2'h3)); forvar3958 = (forvar3958 + (1'h1)))
                    begin
                      reg3959 <= ({{forvar3802}} <<< (|reg3864));
                      reg3960 <= reg3831;
                      reg3961 <= forvar3650;
                      reg3962 <= (-(reg3934 ?
                          ($unsigned(forvar3872) ?
                              forvar3818 : ((8'hb1) == forvar3689)) : forvar3861[(4'h8):(1'h1)]));
                    end
                end
              reg3963 <= reg3798[(3'h6):(3'h4)];
              for (forvar3964 = (1'h0); (forvar3964 < (1'h0)); forvar3964 = (forvar3964 + (1'h1)))
                begin
                  for (forvar3965 = (1'h0); (forvar3965 < (1'h0)); forvar3965 = (forvar3965 + (1'h1)))
                    begin
                      reg3966 <= $signed($unsigned($unsigned(wire1158)));
                      reg3967 <= (-reg3886);
                      reg3968 <= reg3651;
                      reg3969 <= $unsigned($signed(reg3913[(2'h3):(2'h2)]));
                    end
                end
              reg3970 <= reg3834;
            end
          for (forvar3971 = (1'h0); (forvar3971 < (2'h2)); forvar3971 = (forvar3971 + (1'h1)))
            begin
              reg3972 <= $unsigned(forvar3861);
              reg3973 <= (($unsigned($signed((8'h9d))) >> reg3741) ?
                  (~|$signed(reg3921[(4'hd):(3'h4)])) : $unsigned(reg3673));
              reg3974 <= $signed(({forvar3717[(4'h8):(3'h7)]} ~^ (reg3787 ?
                  $signed(reg3682) : (forvar3647 ^~ reg3915))));
              if ($unsigned(($signed($signed((8'h9d))) + (&forvar3920))))
                begin
                  reg3975 <= reg3715[(3'h7):(3'h6)];
                  if (wire3633[(3'h6):(2'h3)])
                    begin
                      reg3976 <= reg3718;
                    end
                  else
                    begin
                      reg3976 <= ({$signed($signed(reg3844))} ?
                          $signed((|(^~reg3866))) : reg3891[(4'hc):(2'h3)]);
                      reg3977 <= $unsigned(((~&{forvar3646}) ?
                          (forvar3920[(1'h0):(1'h0)] ?
                              (^forvar3912) : reg3809) : (^~$unsigned(forvar3929))));
                      reg3978 <= $signed((forvar3673 ^ $signed((+reg3680))));
                      reg3979 <= reg3845;
                    end
                end
              else
                begin
                  for (forvar3975 = (1'h0); (forvar3975 < (1'h1)); forvar3975 = (forvar3975 + (1'h1)))
                    begin
                      reg3976 <= $unsigned(forvar3971[(2'h2):(2'h2)]);
                      reg3977 <= reg3688[(3'h5):(2'h2)];
                      reg3978 <= (~reg3875);
                    end
                  reg3979 <= ((^(~|reg3806[(1'h0):(1'h0)])) ?
                      {$signed($signed(forvar3929))} : forvar3892);
                end
            end
          for (forvar3980 = (1'h0); (forvar3980 < (1'h1)); forvar3980 = (forvar3980 + (1'h1)))
            begin
              for (forvar3981 = (1'h0); (forvar3981 < (2'h3)); forvar3981 = (forvar3981 + (1'h1)))
                begin
                  for (forvar3982 = (1'h0); (forvar3982 < (2'h2)); forvar3982 = (forvar3982 + (1'h1)))
                    begin
                      reg3983 <= reg3697;
                      reg3984 <= (($signed($unsigned(reg3977)) ?
                          $unsigned(forvar3780[(4'h9):(2'h3)]) : ($unsigned(forvar3922) || (reg3664 > reg3787))) && $signed(((~reg3801) ?
                          forvar3940 : reg3656[(1'h0):(1'h0)])));
                      reg3985 <= reg3901[(1'h0):(1'h0)];
                      reg3986 <= (({reg3768} ^~ reg3783) >>> $signed(reg3749[(1'h0):(1'h0)]));
                    end
                  if (({$unsigned(forvar3662)} ?
                      $signed($unsigned((reg3913 & reg3894))) : reg3985[(3'h4):(2'h3)]))
                    begin
                      reg3987 <= $signed((!$unsigned((reg3871 ~^ reg3680))));
                      reg3988 <= reg3936;
                      reg3989 <= ({$unsigned(reg3935)} - ({(reg3943 ?
                              reg3713 : reg3871)} & reg3932));
                    end
                  else
                    begin
                      reg3987 <= ($signed(reg3651[(1'h0):(1'h0)]) ?
                          forvar3644 : reg3832[(4'h9):(1'h0)]);
                      reg3988 <= $signed(($unsigned(forvar3940) ?
                          ($signed(reg3959) ?
                              (!reg3973) : (reg3653 ?
                                  (8'ha2) : reg3907)) : $unsigned((reg3883 ?
                              (8'ha2) : (8'hae)))));
                    end
                  reg3990 <= $signed((reg3739[(2'h3):(1'h0)] - reg3944));
                end
            end
        end
      reg3991 <= $signed((~^$signed((reg3813 ? (8'hb5) : forvar3861))));
    end
  assign wire3992 = ((($signed(reg3880) ?
                            (reg3801 >>> reg3901) : wire2166[(1'h0):(1'h0)]) ?
                        (8'ha7) : reg3654) ^ ($unsigned({forvar3642}) ?
                        (8'ha1) : reg3768));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module647
#( parameter param1055 = (((~&((8'h9d) ? (8'hab) : (8'hb4))) || ({(8'hb9)} ? ((8'hab) ? (8'ha9) : (8'hb4)) : {(8'hab)})) + (~&(8'hb1))) )
(y, clk, wire652, wire651, wire650, wire649, wire648);
  output wire [(32'h83):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire652;
  input wire [(2'h2):(1'h0)] wire651;
  input wire signed [(3'h5):(1'h0)] wire650;
  input wire signed [(4'he):(1'h0)] wire649;
  input wire [(4'he):(1'h0)] wire648;
  wire [(4'h9):(1'h0)] wire1054;
  wire signed [(4'h9):(1'h0)] wire1053;
  wire signed [(4'h9):(1'h0)] wire1051;
  wire signed [(5'h10):(1'h0)] wire659;
  wire [(4'hf):(1'h0)] wire658;
  wire [(4'he):(1'h0)] wire657;
  reg signed [(4'hf):(1'h0)] reg656 = (1'h0);
  wire [(4'he):(1'h0)] wire655;
  wire [(5'h10):(1'h0)] wire654;
  wire signed [(4'hd):(1'h0)] wire653;
  assign y = {wire1054,
                 wire1053,
                 wire1051,
                 wire659,
                 wire658,
                 wire657,
                 reg656,
                 wire655,
                 wire654,
                 wire653,
                 (1'h0)};
  assign wire653 = {(|(wire650[(3'h5):(2'h3)] ?
                           $signed(wire650) : ((8'h9d) >> wire649)))};
  assign wire654 = $signed($unsigned((^(wire650 ? wire648 : wire648))));
  assign wire655 = (&(wire650 ?
                       (wire654[(3'h4):(2'h3)] >>> wire650[(2'h2):(2'h2)]) : $signed((~&wire649))));
  always
    @(posedge clk) begin
      reg656 <= $signed($unsigned({(wire654 ? wire649 : wire655)}));
    end
  assign wire657 = wire651;
  assign wire658 = wire650;
  assign wire659 = ($unsigned($signed({(8'ha8)})) ?
                       (((wire655 + wire648) ?
                               ((8'haa) - wire651) : $unsigned(wire650)) ?
                           $unsigned(wire653[(3'h6):(2'h2)]) : (!wire651)) : {($unsigned(wire655) ?
                               (wire654 ? wire653 : (8'had)) : wire651)});
  module660 modinst1052 (wire1051, clk, wire648, wire650, wire659, wire649);
  assign wire1053 = $signed($signed({wire649}));
  assign wire1054 = reg656[(2'h3):(2'h3)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module660  (y, clk, wire664, wire663, wire662, wire661);
  output wire [(32'h1111):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire664;
  input wire [(2'h2):(1'h0)] wire663;
  input wire [(5'h10):(1'h0)] wire662;
  input wire signed [(4'he):(1'h0)] wire661;
  wire signed [(4'hf):(1'h0)] wire1050;
  reg [(4'ha):(1'h0)] reg1036 = (1'h0);
  reg [(4'hf):(1'h0)] reg1035 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1034 = (1'h0);
  reg [(4'hc):(1'h0)] reg1033 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1049 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1048 = (1'h0);
  reg [(5'h10):(1'h0)] reg1047 = (1'h0);
  reg [(3'h5):(1'h0)] reg1046 = (1'h0);
  reg [(4'ha):(1'h0)] reg1045 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1044 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1043 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1042 = (1'h0);
  reg [(4'hc):(1'h0)] reg1041 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1040 = (1'h0);
  reg [(4'hf):(1'h0)] reg1039 = (1'h0);
  reg [(4'h9):(1'h0)] reg1038 = (1'h0);
  reg [(5'h10):(1'h0)] reg1037 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1036 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1035 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1034 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1033 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1032 = (1'h0);
  reg [(3'h4):(1'h0)] reg1031 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1030 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1029 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1028 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1027 = (1'h0);
  reg [(4'hb):(1'h0)] reg1026 = (1'h0);
  reg [(4'hd):(1'h0)] reg1025 = (1'h0);
  reg [(4'ha):(1'h0)] reg1024 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1023 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1022 = (1'h0);
  reg [(4'h9):(1'h0)] reg1006 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1002 = (1'h0);
  reg [(4'he):(1'h0)] forvar1001 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg998 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar996 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg993 = (1'h0);
  reg [(3'h4):(1'h0)] reg1021 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1020 = (1'h0);
  reg [(2'h2):(1'h0)] reg1019 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1018 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1016 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1015 = (1'h0);
  reg [(5'h10):(1'h0)] reg1014 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1013 = (1'h0);
  reg [(4'hc):(1'h0)] reg1012 = (1'h0);
  reg [(3'h5):(1'h0)] reg1011 = (1'h0);
  reg [(3'h5):(1'h0)] reg1010 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1009 = (1'h0);
  reg [(4'ha):(1'h0)] reg1008 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1007 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1006 = (1'h0);
  reg [(4'he):(1'h0)] reg1005 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1004 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1003 = (1'h0);
  reg [(5'h10):(1'h0)] reg1002 = (1'h0);
  reg [(3'h7):(1'h0)] reg1001 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1000 = (1'h0);
  reg [(4'h8):(1'h0)] reg999 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar998 = (1'h0);
  reg [(4'hf):(1'h0)] reg997 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg996 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg995 = (1'h0);
  reg [(4'hd):(1'h0)] reg994 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar993 = (1'h0);
  reg signed [(4'he):(1'h0)] reg992 = (1'h0);
  reg [(4'h8):(1'h0)] reg991 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg990 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg989 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg986 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar983 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar982 = (1'h0);
  reg [(2'h3):(1'h0)] reg988 = (1'h0);
  reg [(4'hf):(1'h0)] reg987 = (1'h0);
  reg [(4'hc):(1'h0)] forvar986 = (1'h0);
  reg [(3'h5):(1'h0)] reg985 = (1'h0);
  reg [(4'hf):(1'h0)] reg984 = (1'h0);
  reg [(4'hc):(1'h0)] reg983 = (1'h0);
  reg [(3'h6):(1'h0)] reg982 = (1'h0);
  reg [(2'h3):(1'h0)] forvar978 = (1'h0);
  reg [(4'h8):(1'h0)] reg981 = (1'h0);
  reg [(3'h6):(1'h0)] reg980 = (1'h0);
  reg [(4'hf):(1'h0)] reg979 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg978 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg977 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg970 = (1'h0);
  reg [(4'he):(1'h0)] forvar968 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg976 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg975 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg974 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg973 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg972 = (1'h0);
  reg [(4'h8):(1'h0)] reg971 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar970 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg969 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg968 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg967 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar966 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg965 = (1'h0);
  reg [(3'h7):(1'h0)] reg964 = (1'h0);
  reg [(4'h9):(1'h0)] reg963 = (1'h0);
  reg signed [(4'he):(1'h0)] reg962 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar960 = (1'h0);
  reg signed [(4'he):(1'h0)] reg961 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg960 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg959 = (1'h0);
  reg signed [(4'he):(1'h0)] reg958 = (1'h0);
  reg [(4'hc):(1'h0)] reg957 = (1'h0);
  reg [(3'h4):(1'h0)] forvar956 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar955 = (1'h0);
  reg signed [(4'he):(1'h0)] reg954 = (1'h0);
  reg [(4'ha):(1'h0)] reg953 = (1'h0);
  reg [(4'hc):(1'h0)] reg952 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg951 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg950 = (1'h0);
  reg signed [(4'he):(1'h0)] reg949 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar948 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar947 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg946 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg939 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg945 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg944 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg942 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar941 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg940 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar939 = (1'h0);
  reg [(5'h10):(1'h0)] reg938 = (1'h0);
  reg [(4'he):(1'h0)] forvar937 = (1'h0);
  reg [(4'h9):(1'h0)] forvar936 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire935;
  reg signed [(5'h10):(1'h0)] reg926 = (1'h0);
  reg [(4'ha):(1'h0)] forvar912 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg921 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar919 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg916 = (1'h0);
  reg [(3'h7):(1'h0)] reg915 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar908 = (1'h0);
  reg [(4'hf):(1'h0)] reg934 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg933 = (1'h0);
  reg [(4'hb):(1'h0)] reg932 = (1'h0);
  reg [(2'h2):(1'h0)] reg931 = (1'h0);
  reg [(3'h7):(1'h0)] reg930 = (1'h0);
  reg [(4'hb):(1'h0)] forvar929 = (1'h0);
  reg [(3'h7):(1'h0)] reg928 = (1'h0);
  reg signed [(4'he):(1'h0)] reg927 = (1'h0);
  reg [(4'ha):(1'h0)] forvar926 = (1'h0);
  reg [(4'hf):(1'h0)] reg925 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg924 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar923 = (1'h0);
  reg [(3'h7):(1'h0)] reg922 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar921 = (1'h0);
  reg [(2'h2):(1'h0)] reg920 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg919 = (1'h0);
  reg [(3'h6):(1'h0)] reg918 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg917 = (1'h0);
  reg [(2'h3):(1'h0)] forvar916 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar915 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg911 = (1'h0);
  reg [(4'hd):(1'h0)] forvar909 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar906 = (1'h0);
  reg [(2'h2):(1'h0)] reg914 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg913 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg912 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar911 = (1'h0);
  reg [(3'h6):(1'h0)] reg910 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg909 = (1'h0);
  reg [(4'h9):(1'h0)] reg908 = (1'h0);
  reg [(3'h4):(1'h0)] reg907 = (1'h0);
  reg signed [(4'he):(1'h0)] reg906 = (1'h0);
  reg [(4'h8):(1'h0)] reg905 = (1'h0);
  wire [(4'he):(1'h0)] wire904;
  reg signed [(3'h4):(1'h0)] reg871 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar868 = (1'h0);
  reg [(2'h3):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg902 = (1'h0);
  reg [(2'h2):(1'h0)] reg901 = (1'h0);
  reg [(4'ha):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg899 = (1'h0);
  reg [(4'h9):(1'h0)] reg898 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg897 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg896 = (1'h0);
  reg [(4'hc):(1'h0)] forvar895 = (1'h0);
  reg [(5'h10):(1'h0)] forvar894 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg893 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg892 = (1'h0);
  reg [(4'hc):(1'h0)] reg891 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg890 = (1'h0);
  reg [(2'h2):(1'h0)] reg889 = (1'h0);
  reg [(5'h10):(1'h0)] reg888 = (1'h0);
  reg [(4'hf):(1'h0)] reg887 = (1'h0);
  reg [(3'h6):(1'h0)] reg886 = (1'h0);
  reg [(2'h3):(1'h0)] forvar885 = (1'h0);
  reg [(4'h9):(1'h0)] forvar884 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg883 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg882 = (1'h0);
  reg [(4'hb):(1'h0)] reg881 = (1'h0);
  reg [(3'h5):(1'h0)] reg880 = (1'h0);
  reg [(4'ha):(1'h0)] reg879 = (1'h0);
  reg [(4'h8):(1'h0)] reg878 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg876 = (1'h0);
  reg [(4'he):(1'h0)] forvar875 = (1'h0);
  reg [(4'hc):(1'h0)] reg874 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg873 = (1'h0);
  reg signed [(4'he):(1'h0)] reg872 = (1'h0);
  reg [(4'hc):(1'h0)] forvar871 = (1'h0);
  reg [(4'h8):(1'h0)] reg870 = (1'h0);
  reg [(4'h8):(1'h0)] reg869 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg868 = (1'h0);
  reg [(3'h7):(1'h0)] forvar855 = (1'h0);
  reg [(3'h7):(1'h0)] reg854 = (1'h0);
  reg [(4'h8):(1'h0)] reg853 = (1'h0);
  reg [(3'h5):(1'h0)] forvar851 = (1'h0);
  reg [(2'h3):(1'h0)] forvar845 = (1'h0);
  reg [(4'h9):(1'h0)] reg867 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg866 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg865 = (1'h0);
  reg [(3'h6):(1'h0)] forvar864 = (1'h0);
  reg [(2'h3):(1'h0)] reg863 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg862 = (1'h0);
  reg [(3'h6):(1'h0)] reg861 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg860 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg859 = (1'h0);
  reg [(2'h2):(1'h0)] reg858 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg857 = (1'h0);
  reg [(5'h10):(1'h0)] reg856 = (1'h0);
  reg signed [(4'he):(1'h0)] reg855 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar854 = (1'h0);
  reg [(4'h8):(1'h0)] forvar853 = (1'h0);
  reg [(4'hd):(1'h0)] forvar850 = (1'h0);
  reg [(4'hc):(1'h0)] reg852 = (1'h0);
  reg [(4'hc):(1'h0)] reg851 = (1'h0);
  reg [(4'hb):(1'h0)] reg850 = (1'h0);
  reg [(4'ha):(1'h0)] reg847 = (1'h0);
  reg [(5'h10):(1'h0)] reg846 = (1'h0);
  reg [(4'hd):(1'h0)] forvar844 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar838 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar837 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar834 = (1'h0);
  reg [(3'h4):(1'h0)] reg832 = (1'h0);
  reg [(4'hc):(1'h0)] forvar829 = (1'h0);
  reg [(4'h8):(1'h0)] forvar824 = (1'h0);
  reg [(3'h5):(1'h0)] forvar816 = (1'h0);
  reg [(4'hd):(1'h0)] forvar811 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg849 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg848 = (1'h0);
  reg [(3'h5):(1'h0)] forvar847 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar846 = (1'h0);
  reg [(3'h7):(1'h0)] reg839 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg845 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg844 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg843 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg842 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg841 = (1'h0);
  reg [(2'h3):(1'h0)] reg840 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar839 = (1'h0);
  reg [(3'h4):(1'h0)] forvar836 = (1'h0);
  reg [(3'h7):(1'h0)] reg838 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg837 = (1'h0);
  reg [(3'h5):(1'h0)] reg836 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg834 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg833 = (1'h0);
  reg [(4'he):(1'h0)] forvar832 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg831 = (1'h0);
  reg [(4'hd):(1'h0)] reg830 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg829 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg828 = (1'h0);
  reg [(5'h10):(1'h0)] reg827 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg826 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg825 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg824 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg823 = (1'h0);
  reg [(4'hc):(1'h0)] forvar822 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg821 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg817 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar815 = (1'h0);
  reg [(3'h7):(1'h0)] forvar813 = (1'h0);
  reg [(4'hb):(1'h0)] reg812 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg820 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg819 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg818 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar817 = (1'h0);
  reg [(4'h8):(1'h0)] reg816 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg815 = (1'h0);
  reg signed [(4'he):(1'h0)] reg814 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg813 = (1'h0);
  reg [(3'h4):(1'h0)] forvar812 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg811 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar810 = (1'h0);
  wire [(3'h6):(1'h0)] wire809;
  wire [(2'h2):(1'h0)] wire808;
  reg [(4'hd):(1'h0)] reg784 = (1'h0);
  reg [(4'h8):(1'h0)] reg785 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar778 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar774 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg771 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg807 = (1'h0);
  reg [(3'h5):(1'h0)] forvar806 = (1'h0);
  reg [(3'h5):(1'h0)] reg805 = (1'h0);
  reg [(3'h7):(1'h0)] reg804 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg803 = (1'h0);
  reg [(3'h7):(1'h0)] reg802 = (1'h0);
  reg [(3'h4):(1'h0)] forvar801 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg800 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg799 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg798 = (1'h0);
  reg [(4'hb):(1'h0)] reg797 = (1'h0);
  reg [(4'h9):(1'h0)] reg796 = (1'h0);
  reg [(4'h8):(1'h0)] reg795 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg794 = (1'h0);
  reg [(4'h9):(1'h0)] reg793 = (1'h0);
  reg [(3'h4):(1'h0)] reg792 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg791 = (1'h0);
  reg [(4'ha):(1'h0)] reg790 = (1'h0);
  reg [(5'h10):(1'h0)] forvar789 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg788 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg787 = (1'h0);
  reg [(4'hf):(1'h0)] reg786 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar785 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar784 = (1'h0);
  reg [(2'h3):(1'h0)] reg783 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg782 = (1'h0);
  reg [(3'h4):(1'h0)] reg781 = (1'h0);
  reg [(4'hf):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg779 = (1'h0);
  reg [(5'h10):(1'h0)] reg778 = (1'h0);
  reg [(2'h2):(1'h0)] reg777 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg776 = (1'h0);
  reg [(4'hc):(1'h0)] reg775 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg774 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar773 = (1'h0);
  reg [(5'h10):(1'h0)] forvar772 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar771 = (1'h0);
  reg [(3'h4):(1'h0)] reg770 = (1'h0);
  reg [(3'h7):(1'h0)] reg769 = (1'h0);
  reg signed [(4'he):(1'h0)] reg768 = (1'h0);
  reg [(2'h2):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar763 = (1'h0);
  reg [(3'h4):(1'h0)] reg758 = (1'h0);
  reg [(4'he):(1'h0)] reg754 = (1'h0);
  reg [(4'h8):(1'h0)] forvar753 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar752 = (1'h0);
  reg [(3'h7):(1'h0)] reg751 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg750 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar747 = (1'h0);
  reg [(4'h9):(1'h0)] reg744 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg766 = (1'h0);
  reg [(4'h9):(1'h0)] reg765 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg764 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg763 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg762 = (1'h0);
  reg [(2'h2):(1'h0)] reg761 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg760 = (1'h0);
  reg signed [(4'he):(1'h0)] reg759 = (1'h0);
  reg [(4'h9):(1'h0)] forvar758 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg757 = (1'h0);
  reg [(2'h3):(1'h0)] reg756 = (1'h0);
  reg [(3'h7):(1'h0)] reg755 = (1'h0);
  reg [(3'h7):(1'h0)] forvar754 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg753 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg752 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar751 = (1'h0);
  reg [(3'h5):(1'h0)] forvar750 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg746 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg742 = (1'h0);
  reg [(3'h4):(1'h0)] reg749 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg748 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg747 = (1'h0);
  reg [(3'h7):(1'h0)] forvar746 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg745 = (1'h0);
  reg [(3'h5):(1'h0)] forvar744 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg743 = (1'h0);
  reg [(4'hc):(1'h0)] forvar742 = (1'h0);
  reg [(3'h4):(1'h0)] reg741 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg740 = (1'h0);
  reg [(4'ha):(1'h0)] reg739 = (1'h0);
  reg [(4'he):(1'h0)] forvar738 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar737 = (1'h0);
  reg [(2'h2):(1'h0)] forvar736 = (1'h0);
  reg [(4'ha):(1'h0)] forvar735 = (1'h0);
  reg [(5'h10):(1'h0)] reg734 = (1'h0);
  reg [(4'ha):(1'h0)] reg733 = (1'h0);
  reg [(4'hf):(1'h0)] reg732 = (1'h0);
  reg [(4'hd):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg730 = (1'h0);
  reg [(5'h10):(1'h0)] reg729 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar728 = (1'h0);
  reg [(4'hd):(1'h0)] reg727 = (1'h0);
  reg [(4'hd):(1'h0)] reg726 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg725 = (1'h0);
  reg [(2'h2):(1'h0)] reg724 = (1'h0);
  reg [(4'h9):(1'h0)] reg723 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg722 = (1'h0);
  reg [(4'hf):(1'h0)] reg721 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg720 = (1'h0);
  reg [(4'hb):(1'h0)] forvar719 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar718 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar714 = (1'h0);
  reg [(4'hd):(1'h0)] reg710 = (1'h0);
  reg [(4'h9):(1'h0)] reg708 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar707 = (1'h0);
  reg [(4'hf):(1'h0)] reg704 = (1'h0);
  reg [(4'he):(1'h0)] forvar702 = (1'h0);
  reg [(4'hf):(1'h0)] reg699 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg718 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar717 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg716 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar715 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg714 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg713 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg712 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg711 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar710 = (1'h0);
  reg [(4'hf):(1'h0)] reg709 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar708 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg707 = (1'h0);
  reg [(3'h6):(1'h0)] reg706 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg705 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar704 = (1'h0);
  reg [(2'h2):(1'h0)] reg703 = (1'h0);
  reg [(4'hf):(1'h0)] reg702 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg701 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg700 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar699 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg698 = (1'h0);
  reg [(5'h10):(1'h0)] forvar697 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg696 = (1'h0);
  reg [(4'h9):(1'h0)] reg695 = (1'h0);
  reg [(2'h2):(1'h0)] reg694 = (1'h0);
  reg signed [(4'he):(1'h0)] reg687 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar683 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg682 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar667 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg693 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar692 = (1'h0);
  reg [(4'hb):(1'h0)] reg691 = (1'h0);
  reg [(3'h7):(1'h0)] reg690 = (1'h0);
  reg [(3'h4):(1'h0)] reg689 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg688 = (1'h0);
  reg [(2'h3):(1'h0)] forvar687 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg686 = (1'h0);
  reg [(3'h4):(1'h0)] reg685 = (1'h0);
  reg [(3'h6):(1'h0)] reg684 = (1'h0);
  reg [(4'hb):(1'h0)] reg683 = (1'h0);
  reg [(4'he):(1'h0)] forvar682 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg681 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar680 = (1'h0);
  reg [(3'h6):(1'h0)] forvar679 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg669 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar668 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg678 = (1'h0);
  reg [(3'h6):(1'h0)] reg677 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg676 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg675 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg674 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar673 = (1'h0);
  reg [(4'hb):(1'h0)] reg672 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg671 = (1'h0);
  reg [(3'h7):(1'h0)] reg670 = (1'h0);
  reg [(4'hc):(1'h0)] forvar669 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg668 = (1'h0);
  reg [(4'hc):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar666 = (1'h0);
  wire [(4'hd):(1'h0)] wire665;
  assign y = {wire1050,
                 reg1036,
                 reg1035,
                 forvar1034,
                 reg1033,
                 reg1049,
                 reg1048,
                 reg1047,
                 reg1046,
                 reg1045,
                 forvar1044,
                 reg1043,
                 forvar1042,
                 reg1041,
                 forvar1040,
                 reg1039,
                 reg1038,
                 reg1037,
                 forvar1036,
                 forvar1035,
                 reg1034,
                 forvar1033,
                 reg1032,
                 reg1031,
                 reg1030,
                 forvar1029,
                 forvar1028,
                 reg1027,
                 reg1026,
                 reg1025,
                 reg1024,
                 forvar1023,
                 forvar1022,
                 reg1006,
                 forvar1002,
                 forvar1001,
                 reg998,
                 forvar996,
                 reg993,
                 reg1021,
                 forvar1020,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 reg1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1008,
                 forvar1007,
                 forvar1006,
                 reg1005,
                 reg1004,
                 reg1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 reg999,
                 forvar998,
                 reg997,
                 reg996,
                 reg995,
                 reg994,
                 forvar993,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 reg986,
                 forvar983,
                 forvar982,
                 reg988,
                 reg987,
                 forvar986,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 forvar978,
                 reg981,
                 reg980,
                 reg979,
                 reg978,
                 reg977,
                 reg970,
                 forvar968,
                 reg976,
                 reg975,
                 reg974,
                 reg973,
                 reg972,
                 reg971,
                 forvar970,
                 reg969,
                 reg968,
                 reg967,
                 forvar966,
                 reg965,
                 reg964,
                 reg963,
                 reg962,
                 forvar960,
                 reg961,
                 reg960,
                 reg959,
                 reg958,
                 reg957,
                 forvar956,
                 forvar955,
                 reg954,
                 reg953,
                 reg952,
                 reg951,
                 reg950,
                 reg949,
                 forvar948,
                 forvar947,
                 reg946,
                 reg939,
                 reg945,
                 reg944,
                 reg943,
                 reg942,
                 forvar941,
                 reg940,
                 forvar939,
                 reg938,
                 forvar937,
                 forvar936,
                 wire935,
                 reg926,
                 forvar912,
                 reg921,
                 forvar919,
                 reg916,
                 reg915,
                 forvar908,
                 reg934,
                 reg933,
                 reg932,
                 reg931,
                 reg930,
                 forvar929,
                 reg928,
                 reg927,
                 forvar926,
                 reg925,
                 reg924,
                 forvar923,
                 reg922,
                 forvar921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 forvar916,
                 forvar915,
                 reg911,
                 forvar909,
                 forvar906,
                 reg914,
                 reg913,
                 reg912,
                 forvar911,
                 reg910,
                 reg909,
                 reg908,
                 reg907,
                 reg906,
                 reg905,
                 wire904,
                 reg871,
                 forvar868,
                 reg903,
                 reg902,
                 reg901,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 forvar895,
                 forvar894,
                 reg893,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg886,
                 forvar885,
                 forvar884,
                 reg883,
                 reg882,
                 reg881,
                 reg880,
                 reg879,
                 reg878,
                 reg877,
                 reg876,
                 forvar875,
                 reg874,
                 reg873,
                 reg872,
                 forvar871,
                 reg870,
                 reg869,
                 reg868,
                 forvar855,
                 reg854,
                 reg853,
                 forvar851,
                 forvar845,
                 reg867,
                 reg866,
                 reg865,
                 forvar864,
                 reg863,
                 reg862,
                 reg861,
                 reg860,
                 reg859,
                 reg858,
                 reg857,
                 reg856,
                 reg855,
                 forvar854,
                 forvar853,
                 forvar850,
                 reg852,
                 reg851,
                 reg850,
                 reg847,
                 reg846,
                 forvar844,
                 forvar838,
                 forvar837,
                 forvar834,
                 reg832,
                 forvar829,
                 forvar824,
                 forvar816,
                 forvar811,
                 reg849,
                 reg848,
                 forvar847,
                 forvar846,
                 reg839,
                 reg845,
                 reg844,
                 reg843,
                 reg842,
                 reg841,
                 reg840,
                 forvar839,
                 forvar836,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 reg834,
                 reg833,
                 forvar832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 reg825,
                 reg824,
                 reg823,
                 forvar822,
                 reg821,
                 reg817,
                 forvar815,
                 forvar813,
                 reg812,
                 reg820,
                 reg819,
                 reg818,
                 forvar817,
                 reg816,
                 reg815,
                 reg814,
                 reg813,
                 forvar812,
                 reg811,
                 forvar810,
                 wire809,
                 wire808,
                 reg784,
                 reg785,
                 forvar778,
                 forvar774,
                 reg771,
                 reg807,
                 forvar806,
                 reg805,
                 reg804,
                 reg803,
                 reg802,
                 forvar801,
                 reg800,
                 reg799,
                 reg798,
                 reg797,
                 reg796,
                 reg795,
                 reg794,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 forvar789,
                 reg788,
                 reg787,
                 reg786,
                 forvar785,
                 forvar784,
                 reg783,
                 reg782,
                 reg781,
                 reg780,
                 reg779,
                 reg778,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 forvar773,
                 forvar772,
                 forvar771,
                 reg770,
                 reg769,
                 reg768,
                 reg767,
                 forvar763,
                 reg758,
                 reg754,
                 forvar753,
                 forvar752,
                 reg751,
                 reg750,
                 forvar747,
                 reg744,
                 reg766,
                 reg765,
                 reg764,
                 reg763,
                 reg762,
                 reg761,
                 reg760,
                 reg759,
                 forvar758,
                 reg757,
                 reg756,
                 reg755,
                 forvar754,
                 reg753,
                 reg752,
                 forvar751,
                 forvar750,
                 reg746,
                 reg742,
                 reg749,
                 reg748,
                 reg747,
                 forvar746,
                 reg745,
                 forvar744,
                 reg743,
                 forvar742,
                 reg741,
                 reg740,
                 reg739,
                 forvar738,
                 forvar737,
                 forvar736,
                 forvar735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 forvar728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 reg720,
                 forvar719,
                 forvar718,
                 forvar714,
                 reg710,
                 reg708,
                 forvar707,
                 reg704,
                 forvar702,
                 reg699,
                 reg718,
                 forvar717,
                 reg716,
                 forvar715,
                 reg714,
                 reg713,
                 reg712,
                 reg711,
                 forvar710,
                 reg709,
                 forvar708,
                 reg707,
                 reg706,
                 reg705,
                 forvar704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 forvar699,
                 reg698,
                 forvar697,
                 reg696,
                 reg695,
                 reg694,
                 reg687,
                 forvar683,
                 reg682,
                 forvar667,
                 reg693,
                 forvar692,
                 reg691,
                 reg690,
                 reg689,
                 reg688,
                 forvar687,
                 reg686,
                 reg685,
                 reg684,
                 reg683,
                 forvar682,
                 reg681,
                 forvar680,
                 forvar679,
                 reg669,
                 forvar668,
                 reg678,
                 reg677,
                 reg676,
                 reg675,
                 reg674,
                 forvar673,
                 reg672,
                 reg671,
                 reg670,
                 forvar669,
                 reg668,
                 reg667,
                 forvar666,
                 wire665,
                 (1'h0)};
  assign wire665 = wire663[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar666 = (1'h0); (forvar666 < (2'h3)); forvar666 = (forvar666 + (1'h1)))
        begin
          if (((+wire661[(4'h9):(4'h8)]) ? (!wire665[(1'h1):(1'h1)]) : wire665))
            begin
              reg667 <= ($signed($unsigned((|wire664))) ?
                  $signed(wire662) : wire663);
              if ($signed($unsigned((~^(wire665 ^ wire664)))))
                begin
                  reg668 <= ((wire664[(4'h8):(3'h4)] ?
                      $unsigned((reg667 != wire664)) : (^~(!wire662))) <= reg667);
                  for (forvar669 = (1'h0); (forvar669 < (2'h3)); forvar669 = (forvar669 + (1'h1)))
                    begin
                      reg670 <= {({$unsigned(wire661)} ?
                              $unsigned((!forvar666)) : $unsigned((~|wire663)))};
                      reg671 <= (-{((forvar669 == reg670) && $unsigned(forvar669))});
                      reg672 <= (reg667[(4'hc):(3'h4)] ?
                          $signed(forvar666) : ({((8'hb4) || forvar666)} ?
                              $signed({wire663}) : reg671[(4'h9):(3'h5)]));
                    end
                  for (forvar673 = (1'h0); (forvar673 < (2'h2)); forvar673 = (forvar673 + (1'h1)))
                    begin
                      reg674 <= $unsigned($signed((|$signed(wire661))));
                      reg675 <= {(|{$signed(reg667)})};
                      reg676 <= $unsigned({{(8'h9f)}});
                      reg677 <= $signed($signed($unsigned($unsigned(wire661))));
                    end
                  reg678 <= $unsigned((~^((reg670 ? wire662 : reg676) ?
                      ((8'h9c) ? wire665 : wire661) : reg671)));
                end
              else
                begin
                  for (forvar668 = (1'h0); (forvar668 < (1'h1)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg669 <= $unsigned($signed($signed($unsigned(reg671))));
                      reg670 <= (~^wire664[(4'h9):(2'h3)]);
                    end
                end
              for (forvar679 = (1'h0); (forvar679 < (1'h1)); forvar679 = (forvar679 + (1'h1)))
                begin
                  for (forvar680 = (1'h0); (forvar680 < (2'h3)); forvar680 = (forvar680 + (1'h1)))
                    begin
                      reg681 <= forvar668;
                    end
                  for (forvar682 = (1'h0); (forvar682 < (1'h0)); forvar682 = (forvar682 + (1'h1)))
                    begin
                      reg683 <= ($signed($unsigned((8'ha6))) ?
                          (~&$signed(wire662[(3'h6):(3'h4)])) : (~^reg681));
                      reg684 <= {$unsigned(forvar682)};
                      reg685 <= (($unsigned((+wire664)) ?
                              (^~(^~(8'hb1))) : (~(reg674 & (8'ha8)))) ?
                          {$unsigned(reg670[(1'h1):(1'h0)])} : wire665);
                      reg686 <= ((8'hba) ?
                          reg676[(1'h1):(1'h1)] : $signed((&(^forvar679))));
                    end
                  for (forvar687 = (1'h0); (forvar687 < (2'h3)); forvar687 = (forvar687 + (1'h1)))
                    begin
                      reg688 <= $unsigned((~^wire664[(2'h2):(1'h0)]));
                      reg689 <= ((^~reg676) && ($signed($unsigned(forvar668)) ?
                          (+(wire661 < wire662)) : ((reg674 <<< wire664) ?
                              (~|forvar679) : (8'ha0))));
                      reg690 <= (forvar673 ?
                          reg671 : ($unsigned(forvar668[(2'h2):(1'h1)]) ~^ reg670));
                      reg691 <= (+(reg677 <<< (reg686 ?
                          $unsigned(reg675) : $signed(reg668))));
                    end
                  for (forvar692 = (1'h0); (forvar692 < (2'h3)); forvar692 = (forvar692 + (1'h1)))
                    begin
                      reg693 <= $signed((&reg674[(3'h5):(3'h5)]));
                    end
                end
            end
          else
            begin
              for (forvar667 = (1'h0); (forvar667 < (1'h1)); forvar667 = (forvar667 + (1'h1)))
                begin
                  for (forvar668 = (1'h0); (forvar668 < (1'h0)); forvar668 = (forvar668 + (1'h1)))
                    begin
                      reg669 <= $unsigned($unsigned($signed((forvar667 ?
                          reg691 : forvar692))));
                      reg670 <= reg690[(2'h2):(1'h0)];
                      reg671 <= ($signed($signed($unsigned(wire663))) >= reg672[(3'h4):(1'h1)]);
                      reg672 <= {$signed((-$signed((8'hb1))))};
                    end
                  for (forvar673 = (1'h0); (forvar673 < (2'h3)); forvar673 = (forvar673 + (1'h1)))
                    begin
                      reg674 <= (|(((~^forvar673) ?
                          (wire665 ? reg691 : (8'hb6)) : (reg684 ?
                              forvar673 : forvar687)) <<< {reg671}));
                      reg675 <= {((((8'hb8) + forvar680) >>> (wire664 >> forvar682)) * forvar666[(4'he):(4'he)])};
                      reg676 <= $unsigned({(|(~forvar668))});
                    end
                  if ((~^(reg669[(2'h2):(1'h1)] ?
                      $signed($signed(reg672)) : $signed(reg691[(4'hb):(1'h0)]))))
                    begin
                      reg677 <= {$signed($unsigned((reg668 ?
                              reg683 : wire663)))};
                      reg678 <= ($signed(($signed(reg681) >>> (reg689 == (8'ha3)))) == reg672);
                    end
                  else
                    begin
                      reg677 <= $signed((8'ha1));
                    end
                end
              for (forvar679 = (1'h0); (forvar679 < (1'h0)); forvar679 = (forvar679 + (1'h1)))
                begin
                  for (forvar680 = (1'h0); (forvar680 < (1'h1)); forvar680 = (forvar680 + (1'h1)))
                    begin
                      reg681 <= ((+$unsigned(forvar667)) ^ reg671[(4'h8):(3'h7)]);
                      reg682 <= reg677;
                    end
                end
              for (forvar683 = (1'h0); (forvar683 < (2'h2)); forvar683 = (forvar683 + (1'h1)))
                begin
                  reg684 <= (8'hb6);
                  if ({reg683})
                    begin
                      reg685 <= $signed($unsigned($unsigned((reg681 != (8'haf)))));
                      reg686 <= wire665;
                    end
                  else
                    begin
                      reg685 <= $signed(wire663);
                      reg686 <= $unsigned(reg684);
                      reg687 <= ($unsigned($unsigned(reg691)) ?
                          reg686 : $signed(((reg674 >= (8'h9d)) ?
                              reg683[(3'h4):(2'h2)] : {reg683})));
                      reg688 <= $unsigned($unsigned($signed((reg683 ?
                          forvar669 : reg683))));
                    end
                  if ((~^((+(forvar682 ?
                      reg684 : forvar667)) || (forvar668[(2'h3):(2'h3)] ?
                      (reg685 && reg669) : {reg674}))))
                    begin
                      reg689 <= $unsigned((~$signed(((8'h9c) ?
                          reg683 : reg691))));
                      reg690 <= ($signed(reg682) > forvar667[(4'h8):(2'h3)]);
                      reg691 <= $signed(({wire664[(3'h7):(3'h4)]} ~^ forvar692[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg689 <= $signed((wire662 << ((forvar679 <= wire663) >> (!reg687))));
                    end
                  for (forvar692 = (1'h0); (forvar692 < (1'h1)); forvar692 = (forvar692 + (1'h1)))
                    begin
                      reg693 <= reg687[(2'h3):(2'h2)];
                      reg694 <= ((((~wire664) ^~ (forvar669 & reg672)) ?
                          reg668[(4'hf):(4'he)] : reg678[(2'h2):(1'h1)]) * $unsigned(reg691[(4'h9):(4'h9)]));
                      reg695 <= $signed((^~(8'ha1)));
                      reg696 <= (($unsigned($unsigned(forvar680)) >>> (reg688[(3'h5):(3'h4)] ~^ $signed(reg675))) && ((|reg670) ~^ $unsigned(wire665)));
                    end
                end
            end
        end
      if (reg676[(3'h7):(1'h1)])
        begin
          for (forvar697 = (1'h0); (forvar697 < (1'h0)); forvar697 = (forvar697 + (1'h1)))
            begin
              reg698 <= {(($unsigned(reg687) >> $signed(reg691)) ?
                      wire663[(1'h0):(1'h0)] : $signed({(8'haf)}))};
              for (forvar699 = (1'h0); (forvar699 < (2'h3)); forvar699 = (forvar699 + (1'h1)))
                begin
                  reg700 <= wire663;
                  if ((forvar673 ?
                      $unsigned((8'ha8)) : (^reg678[(3'h4):(2'h3)])))
                    begin
                      reg701 <= reg678;
                      reg702 <= $unsigned((-reg674[(4'hc):(4'h9)]));
                      reg703 <= ({$unsigned((reg701 != (8'haa)))} && (^~((~|reg687) ?
                          $signed(forvar669) : forvar692[(2'h3):(2'h2)])));
                    end
                  else
                    begin
                      reg701 <= forvar683[(1'h1):(1'h1)];
                    end
                  for (forvar704 = (1'h0); (forvar704 < (1'h1)); forvar704 = (forvar704 + (1'h1)))
                    begin
                      reg705 <= ((~^{$unsigned(reg675)}) == ($signed((+(8'hb1))) < (8'hb0)));
                      reg706 <= ($signed((~^(wire661 << reg701))) > $unsigned(reg690));
                      reg707 <= (|($signed((~^reg671)) <<< $unsigned((~^reg689))));
                    end
                end
              for (forvar708 = (1'h0); (forvar708 < (2'h3)); forvar708 = (forvar708 + (1'h1)))
                begin
                  reg709 <= reg675[(4'h9):(1'h0)];
                  for (forvar710 = (1'h0); (forvar710 < (1'h1)); forvar710 = (forvar710 + (1'h1)))
                    begin
                      reg711 <= $unsigned({(!forvar682)});
                      reg712 <= $signed($unsigned($signed((forvar699 ?
                          forvar704 : forvar683))));
                      reg713 <= (~|forvar710[(1'h0):(1'h0)]);
                      reg714 <= (&reg695);
                    end
                end
              for (forvar715 = (1'h0); (forvar715 < (2'h3)); forvar715 = (forvar715 + (1'h1)))
                begin
                  reg716 <= $unsigned(forvar680[(3'h6):(1'h1)]);
                  for (forvar717 = (1'h0); (forvar717 < (1'h0)); forvar717 = (forvar717 + (1'h1)))
                    begin
                      reg718 <= (forvar715 ^ $unsigned((+((8'ha4) <<< reg695))));
                    end
                end
            end
        end
      else
        begin
          if ($unsigned((8'hb0)))
            begin
              if ($unsigned((reg690[(2'h3):(1'h0)] ?
                  (|reg683) : reg691[(3'h5):(1'h0)])))
                begin
                  for (forvar697 = (1'h0); (forvar697 < (1'h0)); forvar697 = (forvar697 + (1'h1)))
                    begin
                      reg698 <= reg671;
                      reg699 <= reg676[(3'h6):(1'h1)];
                      reg700 <= (reg696[(2'h3):(2'h3)] ?
                          reg718 : $unsigned({(~forvar683)}));
                      reg701 <= $unsigned((~^($signed(forvar699) ?
                          $signed(reg691) : (forvar687 == reg678))));
                    end
                  for (forvar702 = (1'h0); (forvar702 < (1'h1)); forvar702 = (forvar702 + (1'h1)))
                    begin
                      reg703 <= $signed(((8'hae) | reg678[(2'h2):(1'h0)]));
                      reg704 <= forvar669[(3'h4):(1'h1)];
                      reg705 <= ((~|(&(forvar682 ? forvar666 : reg675))) ?
                          $unsigned({$signed((8'hb3))}) : {((~|reg687) ?
                                  (+reg686) : reg700)});
                      reg706 <= forvar702;
                    end
                  for (forvar707 = (1'h0); (forvar707 < (1'h0)); forvar707 = (forvar707 + (1'h1)))
                    begin
                      reg708 <= ($unsigned((forvar683[(1'h1):(1'h0)] & (reg714 ?
                          reg695 : (8'hb0)))) >= reg711[(2'h3):(1'h1)]);
                      reg709 <= reg703;
                      reg710 <= reg670[(3'h6):(3'h6)];
                    end
                  if (((~^reg672[(3'h4):(3'h4)]) << reg711))
                    begin
                      reg711 <= (reg678[(3'h6):(2'h3)] && $signed((~$unsigned((8'hab)))));
                    end
                  else
                    begin
                      reg711 <= forvar668[(2'h2):(1'h0)];
                      reg712 <= (8'ha1);
                      reg713 <= ($unsigned(forvar666) * (reg690[(3'h5):(3'h4)] ^~ (&reg695[(4'h9):(3'h6)])));
                    end
                end
              else
                begin
                  for (forvar697 = (1'h0); (forvar697 < (1'h0)); forvar697 = (forvar697 + (1'h1)))
                    begin
                      reg698 <= $signed((reg675[(4'h8):(1'h0)] <= $unsigned((^~forvar702))));
                      reg699 <= ({({forvar707} ?
                              (reg710 ?
                                  (8'ha4) : reg689) : reg718)} <<< $signed((~(~|reg707))));
                      reg700 <= $unsigned((($signed(reg677) ?
                          (reg714 ?
                              forvar667 : reg678) : $signed((8'ha7))) >= (-(~^wire662))));
                    end
                end
              for (forvar714 = (1'h0); (forvar714 < (1'h1)); forvar714 = (forvar714 + (1'h1)))
                begin
                  for (forvar715 = (1'h0); (forvar715 < (2'h2)); forvar715 = (forvar715 + (1'h1)))
                    begin
                      reg716 <= ($unsigned($signed((forvar707 > reg669))) && ((reg702[(4'hf):(2'h3)] * forvar704[(1'h0):(1'h0)]) ?
                          (&$unsigned(forvar668)) : {(-wire664)}));
                    end
                end
            end
          else
            begin
              if (($signed(forvar667) < forvar687[(1'h0):(1'h0)]))
                begin
                  for (forvar697 = (1'h0); (forvar697 < (1'h0)); forvar697 = (forvar697 + (1'h1)))
                    begin
                      reg698 <= $signed($signed({reg710}));
                      reg699 <= ((reg704 * {reg685[(2'h2):(2'h2)]}) ?
                          (((reg684 && forvar692) << (reg695 ?
                                  reg718 : reg672)) ?
                              forvar702 : $signed($unsigned((8'hb7)))) : forvar669);
                      reg700 <= ($unsigned({reg688[(2'h2):(1'h1)]}) ?
                          ((wire661[(3'h6):(2'h2)] ^~ wire665) ?
                              $signed((reg671 > (8'haa))) : (-$signed(wire663))) : reg670[(3'h5):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar697 = (1'h0); (forvar697 < (1'h0)); forvar697 = (forvar697 + (1'h1)))
                    begin
                      reg698 <= $unsigned($signed(reg667[(1'h0):(1'h0)]));
                      reg699 <= forvar666[(4'he):(1'h1)];
                    end
                  if (wire661[(4'h9):(4'h9)])
                    begin
                      reg700 <= (8'hb9);
                      reg701 <= {$unsigned((reg669[(1'h1):(1'h1)] || $signed((8'h9f))))};
                      reg702 <= forvar699;
                      reg703 <= (!reg686[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg700 <= ($unsigned({reg705}) ?
                          $signed($signed($unsigned(reg683))) : reg677);
                      reg701 <= (($unsigned(reg710[(3'h7):(3'h5)]) != $signed({reg681})) ?
                          (reg712 ?
                              $signed(reg675[(4'h8):(1'h0)]) : reg671) : (+($signed(wire661) ?
                              ((8'ha5) ?
                                  forvar714 : (8'ha9)) : $unsigned(reg706))));
                    end
                end
            end
          for (forvar717 = (1'h0); (forvar717 < (2'h3)); forvar717 = (forvar717 + (1'h1)))
            begin
              for (forvar718 = (1'h0); (forvar718 < (1'h0)); forvar718 = (forvar718 + (1'h1)))
                begin
                  for (forvar719 = (1'h0); (forvar719 < (1'h0)); forvar719 = (forvar719 + (1'h1)))
                    begin
                      reg720 <= forvar710[(2'h3):(2'h2)];
                      reg721 <= ($signed($unsigned((reg714 ?
                          reg683 : reg708))) <<< wire665);
                      reg722 <= $unsigned((8'hac));
                      reg723 <= ($signed($signed((^~(8'hb8)))) ^~ (8'hb7));
                    end
                  if ((^~$signed($signed($unsigned(reg669)))))
                    begin
                      reg724 <= (forvar718 & $unsigned({$signed(reg694)}));
                      reg725 <= {reg694};
                      reg726 <= ((+{(forvar715 ? reg695 : reg670)}) | reg674);
                    end
                  else
                    begin
                      reg724 <= $signed(($signed(((8'ha9) ? reg690 : reg668)) ?
                          reg704 : forvar667));
                      reg725 <= $unsigned((({forvar687} ?
                              $unsigned((8'hac)) : (wire662 ~^ forvar719)) ?
                          $unsigned((reg677 ?
                              reg696 : wire664)) : {(reg691 || reg704)}));
                      reg726 <= $signed(reg709);
                      reg727 <= forvar682;
                    end
                end
              if (forvar708[(4'hd):(1'h1)])
                begin
                  for (forvar728 = (1'h0); (forvar728 < (1'h0)); forvar728 = (forvar728 + (1'h1)))
                    begin
                      reg729 <= (~|(~|(((8'ha3) ?
                          reg667 : forvar702) * forvar702[(1'h1):(1'h1)])));
                      reg730 <= ($signed($unsigned((!forvar717))) ?
                          (&forvar717[(3'h6):(1'h0)]) : (8'h9e));
                    end
                  if (reg709[(4'h8):(3'h5)])
                    begin
                      reg731 <= reg707;
                      reg732 <= (^reg681);
                      reg733 <= $unsigned((reg691[(3'h5):(2'h3)] >>> $signed($unsigned(reg703))));
                      reg734 <= {(((reg686 >= reg693) ?
                              $signed(forvar666) : reg682[(1'h0):(1'h0)]) >> $signed($signed((8'ha0))))};
                    end
                  else
                    begin
                      reg731 <= ({(reg701 ? {reg699} : (forvar707 < reg707))} ?
                          ((!$unsigned((8'ha7))) - {$signed((8'hb6))}) : $signed((^$unsigned(reg725))));
                      reg732 <= reg723[(4'h8):(4'h8)];
                      reg733 <= $unsigned($signed((8'h9c)));
                    end
                end
              else
                begin
                  for (forvar728 = (1'h0); (forvar728 < (2'h3)); forvar728 = (forvar728 + (1'h1)))
                    begin
                      reg729 <= (+(-reg694));
                      reg730 <= reg727[(3'h5):(3'h4)];
                      reg731 <= {($unsigned(((8'ha9) < forvar704)) >= (reg691 < ((8'hb2) ?
                              (8'hb3) : reg708)))};
                      reg732 <= reg695;
                    end
                end
            end
        end
      for (forvar735 = (1'h0); (forvar735 < (1'h0)); forvar735 = (forvar735 + (1'h1)))
        begin
          for (forvar736 = (1'h0); (forvar736 < (1'h0)); forvar736 = (forvar736 + (1'h1)))
            begin
              for (forvar737 = (1'h0); (forvar737 < (2'h2)); forvar737 = (forvar737 + (1'h1)))
                begin
                  for (forvar738 = (1'h0); (forvar738 < (1'h0)); forvar738 = (forvar738 + (1'h1)))
                    begin
                      reg739 <= (^(reg670[(1'h0):(1'h0)] ?
                          $unsigned((forvar704 ?
                              reg687 : forvar697)) : {reg731}));
                      reg740 <= (~reg733[(3'h4):(3'h4)]);
                      reg741 <= (~^$signed(((reg709 - wire663) ?
                          $signed(forvar707) : (forvar683 ^ forvar704))));
                    end
                end
            end
          if ($signed(($signed(wire662) | $unsigned($unsigned(reg720)))))
            begin
              if (($unsigned($unsigned((~^reg706))) | $signed({(forvar692 ?
                      wire664 : reg686)})))
                begin
                  for (forvar742 = (1'h0); (forvar742 < (1'h0)); forvar742 = (forvar742 + (1'h1)))
                    begin
                      reg743 <= $unsigned((((^(8'hb4)) & forvar742[(2'h2):(2'h2)]) <<< reg730[(3'h7):(1'h0)]));
                    end
                  for (forvar744 = (1'h0); (forvar744 < (1'h1)); forvar744 = (forvar744 + (1'h1)))
                    begin
                      reg745 <= forvar683;
                    end
                  for (forvar746 = (1'h0); (forvar746 < (1'h0)); forvar746 = (forvar746 + (1'h1)))
                    begin
                      reg747 <= $unsigned((~^(~|$signed((8'ha3)))));
                      reg748 <= $unsigned((~^(+forvar680)));
                      reg749 <= (~^(~&reg740));
                    end
                end
              else
                begin
                  if ($unsigned($signed(($signed(reg733) ^~ (^forvar737)))))
                    begin
                      reg742 <= $signed((forvar673[(1'h1):(1'h0)] ?
                          (((8'hb4) ? (8'ha5) : (8'ha8)) ?
                              $unsigned(reg701) : (~reg709)) : forvar738));
                    end
                  else
                    begin
                      reg742 <= (($signed((reg675 >= reg731)) ?
                              $unsigned(wire663[(1'h1):(1'h1)]) : $unsigned((-forvar673))) ?
                          (+reg743) : (~|(~forvar699)));
                      reg743 <= $unsigned((^forvar718[(4'ha):(1'h1)]));
                    end
                  for (forvar744 = (1'h0); (forvar744 < (2'h3)); forvar744 = (forvar744 + (1'h1)))
                    begin
                      reg745 <= $signed(reg742);
                      reg746 <= (!reg707);
                      reg747 <= {$unsigned($unsigned(reg732[(4'hf):(4'hd)]))};
                      reg748 <= $signed((+((forvar680 ?
                          forvar735 : (8'hb6)) < $unsigned(reg670))));
                    end
                  if (wire662[(4'hb):(3'h7)])
                    begin
                      reg749 <= $signed((^~(^~$unsigned(wire662))));
                    end
                  else
                    begin
                      reg749 <= $unsigned((forvar702[(1'h0):(1'h0)] ?
                          $unsigned((reg682 ?
                              forvar702 : forvar715)) : reg688));
                    end
                end
              for (forvar750 = (1'h0); (forvar750 < (1'h0)); forvar750 = (forvar750 + (1'h1)))
                begin
                  for (forvar751 = (1'h0); (forvar751 < (1'h0)); forvar751 = (forvar751 + (1'h1)))
                    begin
                      reg752 <= forvar744;
                      reg753 <= (($signed((|reg748)) ?
                              $signed($signed(forvar738)) : (^~reg686)) ?
                          $signed((8'haa)) : wire664[(4'ha):(1'h1)]);
                    end
                  for (forvar754 = (1'h0); (forvar754 < (2'h2)); forvar754 = (forvar754 + (1'h1)))
                    begin
                      reg755 <= forvar682[(1'h1):(1'h1)];
                      reg756 <= reg720[(1'h1):(1'h1)];
                      reg757 <= reg718[(2'h3):(2'h2)];
                    end
                end
              if (reg752[(3'h5):(1'h0)])
                begin
                  for (forvar758 = (1'h0); (forvar758 < (1'h1)); forvar758 = (forvar758 + (1'h1)))
                    begin
                      reg759 <= (($signed($signed(reg682)) + (forvar692 ^~ $signed(forvar697))) ?
                          $unsigned((((8'hb2) - (8'haf)) ?
                              $signed(forvar717) : (forvar687 ?
                                  reg676 : forvar758))) : reg724[(1'h1):(1'h1)]);
                      reg760 <= $unsigned({$unsigned({forvar718})});
                    end
                  reg761 <= forvar758[(1'h1):(1'h1)];
                  reg762 <= (~$signed((~&reg732)));
                end
              else
                begin
                  for (forvar758 = (1'h0); (forvar758 < (1'h1)); forvar758 = (forvar758 + (1'h1)))
                    begin
                      reg759 <= $signed(({$unsigned((8'hb9))} ?
                          (8'hab) : (8'haf)));
                      reg760 <= ($signed({reg732[(4'ha):(4'h8)]}) >= (8'ha2));
                      reg761 <= (reg703 ?
                          {forvar758} : $signed(((^(8'hb9)) * (~&forvar718))));
                    end
                  if ((-reg700))
                    begin
                      reg762 <= (-wire665[(4'h8):(3'h4)]);
                      reg763 <= reg668[(3'h7):(1'h0)];
                      reg764 <= $signed(forvar707[(4'hb):(3'h5)]);
                    end
                  else
                    begin
                      reg762 <= ($unsigned({reg682[(1'h1):(1'h1)]}) ?
                          (reg701[(2'h3):(1'h0)] + (reg743[(2'h3):(1'h0)] != $signed(forvar736))) : $signed({$unsigned(reg733)}));
                      reg763 <= $unsigned($signed($signed($signed(reg706))));
                      reg764 <= $signed(($signed(reg707) ?
                          {(^~reg722)} : ($unsigned(forvar714) ?
                              (reg706 | (8'ha4)) : $unsigned(reg731))));
                      reg765 <= {(($signed(reg688) ?
                              {reg678} : $unsigned(forvar750)) ~^ ($unsigned(reg763) != $signed(forvar707)))};
                    end
                end
              reg766 <= reg688;
            end
          else
            begin
              for (forvar742 = (1'h0); (forvar742 < (1'h0)); forvar742 = (forvar742 + (1'h1)))
                begin
                  if ($unsigned((+((reg669 ? forvar704 : (8'ha6)) || (reg705 ?
                      reg700 : reg714)))))
                    begin
                      reg743 <= $unsigned(reg742[(3'h5):(1'h0)]);
                      reg744 <= {(+(8'h9e))};
                      reg745 <= reg681;
                    end
                  else
                    begin
                      reg743 <= reg761[(1'h0):(1'h0)];
                      reg744 <= ($signed(({reg670} | (forvar751 ?
                          reg718 : reg711))) * forvar750);
                      reg745 <= ($unsigned(reg747) == wire663);
                      reg746 <= reg748[(2'h2):(1'h1)];
                    end
                  for (forvar747 = (1'h0); (forvar747 < (2'h3)); forvar747 = (forvar747 + (1'h1)))
                    begin
                      reg748 <= $unsigned($signed(reg714));
                      reg749 <= ((^reg723[(1'h1):(1'h1)]) | (&(+reg677)));
                      reg750 <= (8'ha6);
                      reg751 <= (&($signed(forvar708[(3'h7):(2'h3)]) ?
                          (reg739[(1'h1):(1'h0)] ?
                              (reg746 ?
                                  reg711 : reg746) : $signed(reg698)) : ((reg693 ?
                                  reg734 : reg668) ?
                              (!reg729) : (!(8'hab)))));
                    end
                end
              for (forvar752 = (1'h0); (forvar752 < (1'h1)); forvar752 = (forvar752 + (1'h1)))
                begin
                  for (forvar753 = (1'h0); (forvar753 < (2'h2)); forvar753 = (forvar753 + (1'h1)))
                    begin
                      reg754 <= {($signed(forvar719) ?
                              reg703[(2'h2):(1'h1)] : reg683[(1'h1):(1'h0)])};
                    end
                  reg755 <= ($unsigned((~^(forvar673 && reg689))) ?
                      (($unsigned((8'hb1)) & $unsigned((8'ha6))) >> $signed((!reg743))) : {$signed((reg744 ^ reg756))});
                end
              if ($unsigned($unsigned((reg682[(2'h2):(1'h0)] | (!reg765)))))
                begin
                  reg756 <= $signed((reg703 ?
                      (!(8'hab)) : {forvar704[(1'h0):(1'h0)]}));
                end
              else
                begin
                  if ((~(~|{((8'ha8) << reg765)})))
                    begin
                      reg756 <= ($unsigned({forvar702[(2'h3):(2'h2)]}) ?
                          $signed(reg704[(3'h7):(2'h2)]) : reg695);
                    end
                  else
                    begin
                      reg756 <= reg701[(3'h6):(3'h5)];
                      reg757 <= forvar738;
                      reg758 <= (forvar728[(2'h3):(2'h3)] ?
                          {{(wire661 ? forvar736 : (8'h9f))}} : reg764);
                      reg759 <= reg684[(3'h6):(3'h4)];
                    end
                  if (reg742)
                    begin
                      reg760 <= {reg703[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg760 <= $unsigned(forvar738);
                      reg761 <= ((({reg727} ?
                          reg670[(1'h1):(1'h0)] : ((8'hac) ?
                              reg711 : reg705)) << $unsigned(reg672[(2'h3):(1'h1)])) <= reg764[(2'h2):(1'h1)]);
                      reg762 <= reg676[(4'h8):(3'h6)];
                    end
                  for (forvar763 = (1'h0); (forvar763 < (2'h2)); forvar763 = (forvar763 + (1'h1)))
                    begin
                      reg764 <= forvar673;
                      reg765 <= {((|(reg765 <<< reg682)) ^ ((reg730 ~^ forvar750) ?
                              (forvar758 >> forvar717) : forvar666[(4'hb):(2'h3)]))};
                      reg766 <= (reg685 ? forvar679 : $signed((|(~&reg760))));
                    end
                  if ($unsigned(reg684[(3'h6):(2'h2)]))
                    begin
                      reg767 <= reg698[(4'h8):(4'h8)];
                      reg768 <= reg757;
                    end
                  else
                    begin
                      reg767 <= $unsigned(reg684);
                      reg768 <= $signed((($unsigned(reg684) && $signed(forvar699)) << ((|forvar736) ?
                          $signed(reg742) : $unsigned(reg733))));
                      reg769 <= wire663;
                    end
                end
            end
          reg770 <= ((~|reg740[(4'hb):(1'h0)]) && (^~reg674[(2'h2):(2'h2)]));
        end
      if ((forvar692[(2'h2):(2'h2)] << forvar669[(3'h7):(3'h6)]))
        begin
          for (forvar771 = (1'h0); (forvar771 < (1'h0)); forvar771 = (forvar771 + (1'h1)))
            begin
              for (forvar772 = (1'h0); (forvar772 < (1'h1)); forvar772 = (forvar772 + (1'h1)))
                begin
                  for (forvar773 = (1'h0); (forvar773 < (2'h3)); forvar773 = (forvar773 + (1'h1)))
                    begin
                      reg774 <= ($unsigned(((8'hb1) >> $signed(reg741))) ?
                          $signed((^~reg749[(2'h2):(2'h2)])) : $unsigned(($signed(reg678) <= (reg767 ^ reg709))));
                      reg775 <= reg677;
                    end
                  if (reg716[(2'h3):(1'h1)])
                    begin
                      reg776 <= (~|$signed($signed((reg754 != forvar673))));
                      reg777 <= $signed(((&forvar744) << {(&reg720)}));
                      reg778 <= (~&reg754[(4'hb):(1'h0)]);
                      reg779 <= (8'hab);
                    end
                  else
                    begin
                      reg776 <= $unsigned((~&(~&{reg694})));
                      reg777 <= reg739[(2'h2):(1'h0)];
                      reg778 <= forvar679;
                    end
                  if (((forvar715 << $signed(reg704[(2'h2):(2'h2)])) ?
                      reg699 : (~|$unsigned({reg760}))))
                    begin
                      reg780 <= (reg720 == (8'hb3));
                    end
                  else
                    begin
                      reg780 <= ({$unsigned(reg778)} || (^(^$unsigned(forvar758))));
                      reg781 <= (^($signed($signed(reg778)) ?
                          $signed((reg751 - forvar746)) : $unsigned({reg675})));
                      reg782 <= $unsigned($signed(forvar750[(2'h3):(1'h0)]));
                    end
                  reg783 <= $signed($signed($unsigned($signed(reg703))));
                end
              for (forvar784 = (1'h0); (forvar784 < (2'h2)); forvar784 = (forvar784 + (1'h1)))
                begin
                  for (forvar785 = (1'h0); (forvar785 < (1'h1)); forvar785 = (forvar785 + (1'h1)))
                    begin
                      reg786 <= (((!reg667) ?
                              $signed($unsigned(forvar682)) : {$unsigned(reg686)}) ?
                          (forvar668 ?
                              ((~^(8'ha6)) ?
                                  $unsigned(reg724) : (reg710 ?
                                      forvar682 : reg694)) : ($unsigned(forvar747) ?
                                  $signed(reg753) : (wire662 ?
                                      (8'h9f) : (8'ha2)))) : {$signed((forvar715 << reg764))});
                      reg787 <= ($unsigned(forvar717) ?
                          (!$unsigned((reg745 <= reg725))) : reg723);
                      reg788 <= $unsigned($signed({$signed(reg726)}));
                    end
                end
              for (forvar789 = (1'h0); (forvar789 < (1'h1)); forvar789 = (forvar789 + (1'h1)))
                begin
                  if (forvar710[(2'h3):(1'h0)])
                    begin
                      reg790 <= (-(reg766[(4'h8):(3'h6)] | reg770[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg790 <= (~^($signed(((8'hb4) > reg777)) >>> $unsigned({forvar785})));
                      reg791 <= reg762;
                      reg792 <= (~($unsigned($unsigned(reg696)) ~^ ({reg787} << reg727[(2'h2):(1'h1)])));
                    end
                  if ((reg763[(2'h3):(1'h0)] ^~ $signed($unsigned((forvar687 ?
                      reg672 : forvar742)))))
                    begin
                      reg793 <= $unsigned((8'hac));
                      reg794 <= $signed((reg777[(1'h1):(1'h0)] > forvar704[(3'h5):(3'h4)]));
                      reg795 <= reg675;
                      reg796 <= forvar687;
                    end
                  else
                    begin
                      reg793 <= wire661[(4'h9):(2'h2)];
                      reg794 <= $unsigned($unsigned(({reg676} ?
                          (reg769 + (8'hb5)) : forvar736[(2'h2):(1'h1)])));
                      reg795 <= reg754;
                      reg796 <= (&{(8'ha9)});
                    end
                  if (((!forvar669) | $unsigned($unsigned((reg720 - (8'hb4))))))
                    begin
                      reg797 <= $signed((forvar683 ?
                          {forvar737} : $signed(reg694[(1'h1):(1'h0)])));
                      reg798 <= (reg675 <<< (~$unsigned($signed(forvar772))));
                      reg799 <= reg669[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg797 <= (8'h9f);
                      reg798 <= reg798;
                      reg799 <= (reg760[(3'h5):(2'h2)] < forvar789[(4'hf):(3'h7)]);
                      reg800 <= $signed($unsigned(($unsigned(reg700) ?
                          reg675 : (^(8'ha2)))));
                    end
                end
              for (forvar801 = (1'h0); (forvar801 < (1'h1)); forvar801 = (forvar801 + (1'h1)))
                begin
                  reg802 <= (-(8'hb2));
                  if ((~($unsigned(forvar747[(3'h5):(2'h3)]) ?
                      $unsigned(reg676[(3'h4):(2'h3)]) : reg734[(3'h5):(1'h0)])))
                    begin
                      reg803 <= (8'ha3);
                      reg804 <= {(+{$unsigned(reg677)})};
                      reg805 <= reg754;
                    end
                  else
                    begin
                      reg803 <= ((reg708[(1'h1):(1'h1)] > (~^(reg711 == reg780))) <<< forvar784[(4'hd):(4'hc)]);
                    end
                  for (forvar806 = (1'h0); (forvar806 < (1'h1)); forvar806 = (forvar806 + (1'h1)))
                    begin
                      reg807 <= (reg670[(2'h2):(1'h0)] ?
                          (forvar744 ?
                              {{reg723}} : $unsigned((forvar801 ?
                                  reg793 : reg770))) : $signed($signed($signed(reg707))));
                    end
                end
            end
        end
      else
        begin
          reg771 <= (|forvar751[(2'h2):(2'h2)]);
          for (forvar772 = (1'h0); (forvar772 < (2'h3)); forvar772 = (forvar772 + (1'h1)))
            begin
              for (forvar773 = (1'h0); (forvar773 < (1'h1)); forvar773 = (forvar773 + (1'h1)))
                begin
                  for (forvar774 = (1'h0); (forvar774 < (1'h1)); forvar774 = (forvar774 + (1'h1)))
                    begin
                      reg775 <= reg702[(3'h4):(2'h2)];
                      reg776 <= (8'hb2);
                      reg777 <= ($unsigned({(~^reg671)}) ?
                          $unsigned((forvar773[(4'ha):(2'h2)] <= forvar719)) : {reg690[(3'h6):(3'h5)]});
                    end
                  for (forvar778 = (1'h0); (forvar778 < (1'h1)); forvar778 = (forvar778 + (1'h1)))
                    begin
                      reg779 <= (&((reg754 ? (~^forvar752) : $signed((8'ha4))) ?
                          forvar758 : forvar687[(1'h1):(1'h1)]));
                      reg780 <= (((reg693 && (^forvar699)) >> $unsigned(forvar728[(3'h5):(1'h1)])) ~^ $signed((((8'haf) ?
                          (8'hba) : (8'ha5)) != $signed(reg716))));
                    end
                  if ((((-{reg798}) ?
                      ((reg731 > reg712) ?
                          {forvar687} : (reg781 + (8'hb0))) : reg723) ^ $signed(($signed(forvar668) ?
                      ((8'hb5) || (8'h9e)) : (+reg751)))))
                    begin
                      reg781 <= ((+$unsigned((-reg805))) >= reg724[(2'h2):(2'h2)]);
                      reg782 <= reg792[(3'h4):(3'h4)];
                      reg783 <= $signed(((8'had) ?
                          (reg782[(2'h2):(1'h0)] ~^ $unsigned(reg693)) : reg714));
                    end
                  else
                    begin
                      reg781 <= ($signed({$unsigned(reg707)}) << ((~(forvar758 ?
                          reg776 : forvar763)) & ((+reg677) ?
                          (forvar699 <= reg771) : $signed(reg667))));
                      reg782 <= $unsigned($unsigned(reg769[(3'h7):(3'h5)]));
                      reg783 <= (~&reg709);
                    end
                end
              if (reg747)
                begin
                  for (forvar784 = (1'h0); (forvar784 < (2'h3)); forvar784 = (forvar784 + (1'h1)))
                    begin
                      reg785 <= ({reg767[(2'h2):(1'h1)]} != reg796[(4'h9):(2'h2)]);
                      reg786 <= forvar806;
                      reg787 <= reg674;
                    end
                end
              else
                begin
                  reg784 <= $unsigned((reg705 ?
                      reg777[(1'h0):(1'h0)] : reg718[(2'h3):(1'h0)]));
                  for (forvar785 = (1'h0); (forvar785 < (1'h0)); forvar785 = (forvar785 + (1'h1)))
                    begin
                      reg786 <= {reg729[(4'he):(2'h2)]};
                    end
                end
            end
        end
    end
  assign wire808 = $signed(forvar680);
  assign wire809 = {{{(~|reg701)}}};
  always
    @(posedge clk) begin
      if ((|((reg758 ? (~reg784) : reg722) ?
          reg683 : $signed((reg742 ? reg732 : reg783)))))
        begin
          for (forvar810 = (1'h0); (forvar810 < (2'h2)); forvar810 = (forvar810 + (1'h1)))
            begin
              if (reg705)
                begin
                  reg811 <= ((reg794[(1'h1):(1'h1)] ? (!wire665) : (~reg751)) ?
                      $signed((!reg687[(1'h1):(1'h0)])) : ($signed({forvar714}) || (reg753[(1'h0):(1'h0)] > $signed(reg749))));
                  for (forvar812 = (1'h0); (forvar812 < (2'h2)); forvar812 = (forvar812 + (1'h1)))
                    begin
                      reg813 <= reg723[(1'h0):(1'h0)];
                      reg814 <= (|forvar679[(1'h0):(1'h0)]);
                      reg815 <= forvar738[(3'h7):(3'h5)];
                      reg816 <= forvar718;
                    end
                  for (forvar817 = (1'h0); (forvar817 < (2'h3)); forvar817 = (forvar817 + (1'h1)))
                    begin
                      reg818 <= (reg720 || reg770);
                      reg819 <= ($unsigned(((~^reg785) ?
                              $unsigned(reg694) : reg753[(3'h6):(2'h2)])) ?
                          reg766[(3'h7):(3'h4)] : (reg710[(1'h0):(1'h0)] ?
                              $unsigned($unsigned(forvar679)) : (reg727 > reg694)));
                    end
                  reg820 <= ({reg684[(1'h1):(1'h1)]} ?
                      (~&$unsigned({reg684})) : $unsigned($signed((^reg714))));
                end
              else
                begin
                  if ($unsigned(($unsigned((wire808 - reg786)) ?
                      wire665[(1'h0):(1'h0)] : $unsigned((-(8'ha7))))))
                    begin
                      reg811 <= ((reg686[(3'h5):(2'h2)] ?
                          $unsigned((8'hb5)) : {((8'ha4) << reg695)}) == $signed(({reg669} ^ (forvar784 ^ reg732))));
                      reg812 <= {reg724[(2'h2):(1'h0)]};
                    end
                  else
                    begin
                      reg811 <= ((reg746 != ($signed(reg711) - $signed(reg708))) ?
                          reg732 : (($unsigned(reg820) ? {reg798} : reg713) ?
                              reg703 : $unsigned(((8'ha9) ?
                                  reg778 : forvar812))));
                      reg812 <= (~|$signed(forvar679[(3'h6):(3'h5)]));
                    end
                  for (forvar813 = (1'h0); (forvar813 < (1'h0)); forvar813 = (forvar813 + (1'h1)))
                    begin
                      reg814 <= (({(reg751 || (8'ha4))} > reg705[(2'h3):(1'h1)]) ?
                          $unsigned((8'hb5)) : reg700[(4'hf):(4'he)]);
                    end
                  for (forvar815 = (1'h0); (forvar815 < (2'h3)); forvar815 = (forvar815 + (1'h1)))
                    begin
                      reg816 <= {reg775};
                      reg817 <= ((^~$signed((~^reg731))) ?
                          {($unsigned(forvar812) ?
                                  reg671 : (~wire663))} : (~&reg685));
                    end
                  if ($signed($signed(forvar679[(3'h4):(3'h4)])))
                    begin
                      reg818 <= (!(forvar742 ?
                          ($unsigned(reg756) ?
                              ((8'hb7) >>> (8'ha4)) : $signed(wire663)) : (reg780 ?
                              (reg674 ? reg811 : reg694) : $signed(reg769))));
                      reg819 <= $unsigned($signed((8'ha4)));
                      reg820 <= (~{reg793});
                      reg821 <= $unsigned($unsigned(($signed(reg788) ^ {reg704})));
                    end
                  else
                    begin
                      reg818 <= (reg714[(3'h4):(1'h0)] << ($signed($unsigned(reg743)) ?
                          (reg763 ?
                              reg775 : (8'hb9)) : forvar778[(4'hd):(3'h5)]));
                      reg819 <= reg784[(4'ha):(4'h8)];
                    end
                end
              for (forvar822 = (1'h0); (forvar822 < (2'h3)); forvar822 = (forvar822 + (1'h1)))
                begin
                  if ((8'ha5))
                    begin
                      reg823 <= (!$unsigned(reg734));
                      reg824 <= reg669[(3'h4):(1'h1)];
                      reg825 <= forvar817[(3'h5):(2'h2)];
                      reg826 <= ($unsigned(((!forvar815) & reg778)) ?
                          ($unsigned((~reg825)) >> reg765[(3'h7):(1'h1)]) : (~(+((8'hb9) >= reg729))));
                    end
                  else
                    begin
                      reg823 <= ($signed((~|reg800[(2'h2):(1'h1)])) > reg751);
                      reg824 <= reg782[(2'h2):(1'h1)];
                    end
                  if ($unsigned(reg691[(2'h2):(1'h1)]))
                    begin
                      reg827 <= (~^$signed(((reg745 << forvar778) + (reg699 ?
                          (8'hb7) : reg816))));
                    end
                  else
                    begin
                      reg827 <= $unsigned((reg762[(2'h3):(2'h2)] ?
                          forvar679[(1'h1):(1'h1)] : (+(forvar789 >> (8'hb6)))));
                    end
                  if (forvar667)
                    begin
                      reg828 <= ((forvar736 > $signed(reg805[(3'h4):(1'h0)])) <= (~^forvar702));
                      reg829 <= reg745;
                      reg830 <= {($unsigned($unsigned((8'hb2))) ^ reg828)};
                    end
                  else
                    begin
                      reg828 <= reg696;
                      reg829 <= $unsigned((8'hb2));
                      reg830 <= ({{(forvar702 & forvar753)}} && (~reg727[(4'ha):(2'h2)]));
                      reg831 <= (((^~(forvar714 * (8'ha7))) < (8'hac)) <<< $unsigned((+(+reg762))));
                    end
                  for (forvar832 = (1'h0); (forvar832 < (2'h3)); forvar832 = (forvar832 + (1'h1)))
                    begin
                      reg833 <= reg681[(4'h9):(3'h5)];
                      reg834 <= $signed(($unsigned(wire662[(4'hd):(3'h6)]) ?
                          ($unsigned(reg678) ?
                              $signed(reg830) : $signed((8'ha0))) : ((~reg714) <<< wire808)));
                      reg835 <= (-$unsigned($signed(((8'hb8) == reg726))));
                    end
                end
            end
          if ($unsigned((((reg741 | reg759) > (+(8'hb5))) ?
              reg691 : (~|(reg784 <= (8'ha2))))))
            begin
              if ($signed((($unsigned(reg716) - {reg706}) ?
                  ((&forvar666) + reg687[(1'h1):(1'h0)]) : reg745)))
                begin
                  if (reg716)
                    begin
                      reg836 <= reg687;
                      reg837 <= (8'ha8);
                      reg838 <= (+($signed((^reg762)) ?
                          reg700 : $unsigned(reg696)));
                    end
                  else
                    begin
                      reg836 <= reg838;
                    end
                end
              else
                begin
                  for (forvar836 = (1'h0); (forvar836 < (1'h0)); forvar836 = (forvar836 + (1'h1)))
                    begin
                      reg837 <= reg812;
                    end
                end
              if ((~|$unsigned((+(reg803 ? reg742 : reg758)))))
                begin
                  for (forvar839 = (1'h0); (forvar839 < (1'h1)); forvar839 = (forvar839 + (1'h1)))
                    begin
                      reg840 <= $signed(({(reg837 << forvar673)} ?
                          $unsigned((~^(8'ha8))) : reg747[(3'h7):(1'h0)]));
                      reg841 <= reg729;
                      reg842 <= forvar763;
                    end
                  if (reg774)
                    begin
                      reg843 <= $unsigned((8'hb3));
                      reg844 <= forvar680;
                      reg845 <= (-reg724[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg843 <= $unsigned((8'hb9));
                      reg844 <= (forvar718[(3'h4):(2'h2)] ?
                          {{(~(8'ha7))}} : (~&((&forvar746) ?
                              reg812[(3'h5):(3'h5)] : (~&reg716))));
                      reg845 <= (reg731 ?
                          $signed((reg746 ?
                              reg778 : (reg834 ^~ forvar673))) : $unsigned(reg685));
                    end
                end
              else
                begin
                  if ((^~(~&$unsigned(forvar812[(3'h4):(1'h0)]))))
                    begin
                      reg839 <= $signed((reg703 ?
                          $signed(reg705[(1'h0):(1'h0)]) : forvar753));
                      reg840 <= wire808[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg839 <= $unsigned($signed(((forvar718 && wire661) ?
                          $signed(forvar758) : (forvar719 ? reg815 : reg816))));
                      reg840 <= (~{($signed(forvar702) <= (8'hb3))});
                      reg841 <= $signed((forvar758 <= (~^(reg783 != reg743))));
                    end
                end
              for (forvar846 = (1'h0); (forvar846 < (2'h2)); forvar846 = (forvar846 + (1'h1)))
                begin
                  for (forvar847 = (1'h0); (forvar847 < (2'h2)); forvar847 = (forvar847 + (1'h1)))
                    begin
                      reg848 <= (reg767[(2'h2):(1'h1)] > $unsigned({(reg751 ?
                              wire663 : reg721)}));
                      reg849 <= (((~&{reg729}) ?
                              $unsigned(forvar736[(1'h0):(1'h0)]) : ($unsigned(forvar815) >= $signed(forvar714))) ?
                          (({(8'ha2)} ? {forvar784} : $unsigned(reg743)) ?
                              (forvar832[(3'h5):(1'h0)] ^~ (reg760 ?
                                  reg688 : (8'ha2))) : ((reg681 ?
                                      reg799 : forvar669) ?
                                  (~&reg819) : reg836)) : (forvar773 ^~ reg684[(2'h2):(2'h2)]));
                    end
                end
            end
          else
            begin
              reg836 <= ({$unsigned((^reg749))} | reg837[(2'h3):(2'h3)]);
            end
        end
      else
        begin
          for (forvar810 = (1'h0); (forvar810 < (1'h0)); forvar810 = (forvar810 + (1'h1)))
            begin
              for (forvar811 = (1'h0); (forvar811 < (1'h0)); forvar811 = (forvar811 + (1'h1)))
                begin
                  reg812 <= reg712;
                  if (reg671)
                    begin
                      reg813 <= (reg817[(3'h7):(2'h3)] << $unsigned($signed((reg741 ?
                          wire808 : reg774))));
                      reg814 <= {{forvar714}};
                      reg815 <= $signed(($unsigned((^~reg683)) ?
                          reg779 : (~^$unsigned(wire663))));
                    end
                  else
                    begin
                      reg813 <= $signed($signed(reg694));
                      reg814 <= $signed(($signed((reg695 ?
                              reg700 : forvar666)) ?
                          $signed((reg686 ? reg746 : forvar774)) : reg683));
                    end
                end
              if ((^~(((-reg675) != forvar812) | ((reg838 & forvar822) ?
                  (reg844 ? reg849 : reg828) : (!(8'ha1))))))
                begin
                  reg816 <= $signed($unsigned(($signed(reg785) | (~|reg678))));
                end
              else
                begin
                  for (forvar816 = (1'h0); (forvar816 < (1'h1)); forvar816 = (forvar816 + (1'h1)))
                    begin
                      reg817 <= reg791[(3'h6):(1'h1)];
                    end
                  if ({$unsigned($unsigned($unsigned(wire665)))})
                    begin
                      reg818 <= $signed(($signed(forvar697[(1'h1):(1'h1)]) ?
                          forvar687[(1'h0):(1'h0)] : {$unsigned(reg838)}));
                      reg819 <= reg833[(3'h6):(3'h5)];
                      reg820 <= ((~forvar742[(4'h9):(3'h4)]) <<< reg849[(3'h7):(1'h0)]);
                      reg821 <= $signed(($signed($unsigned(reg829)) ~^ $signed((reg829 ?
                          reg842 : forvar668))));
                    end
                  else
                    begin
                      reg818 <= (8'ha8);
                      reg819 <= {forvar785};
                      reg820 <= ($signed({reg686}) != (((forvar812 ?
                                  (8'h9f) : reg790) ?
                              ((8'ha8) >= forvar846) : {reg790}) ?
                          ($signed(reg749) < reg716[(1'h0):(1'h0)]) : wire664));
                      reg821 <= $signed($unsigned((!$signed(reg849))));
                    end
                  for (forvar822 = (1'h0); (forvar822 < (2'h3)); forvar822 = (forvar822 + (1'h1)))
                    begin
                      reg823 <= reg807;
                    end
                end
              for (forvar824 = (1'h0); (forvar824 < (1'h1)); forvar824 = (forvar824 + (1'h1)))
                begin
                  if ((|{((forvar772 ? reg768 : (8'had)) ?
                          {reg743} : (8'hb0))}))
                    begin
                      reg825 <= $unsigned((((~forvar673) ~^ (reg756 ?
                              reg753 : forvar773)) ?
                          (&$signed(reg763)) : ((reg667 ?
                              reg712 : (8'hb4)) <<< $unsigned(forvar832))));
                      reg826 <= forvar744;
                    end
                  else
                    begin
                      reg825 <= $unsigned((((reg825 ? forvar813 : reg844) ?
                          (reg848 ?
                              reg828 : reg676) : ((8'hb2) >> reg688)) || $unsigned(((8'hb0) ^~ (8'ha2)))));
                      reg826 <= ((~&(forvar718 - $unsigned((8'ha3)))) ?
                          $unsigned((reg766[(1'h1):(1'h1)] < (reg748 ?
                              forvar753 : forvar836))) : reg784);
                      reg827 <= ($unsigned((~reg744)) ?
                          reg770[(3'h4):(3'h4)] : $unsigned(((+reg841) ?
                              {reg760} : reg762)));
                      reg828 <= $signed(reg842[(3'h5):(2'h2)]);
                    end
                  for (forvar829 = (1'h0); (forvar829 < (1'h1)); forvar829 = (forvar829 + (1'h1)))
                    begin
                      reg830 <= forvar773;
                      reg831 <= (reg770 ?
                          (~&(~&(8'haa))) : (($signed((8'hac)) ?
                                  $unsigned(reg685) : reg734) ?
                              (^~$signed(forvar697)) : reg823));
                      reg832 <= $unsigned((^$unsigned(reg763)));
                      reg833 <= ($signed($unsigned((reg816 ?
                          reg798 : reg819))) - (($signed(reg797) <= ((8'h9f) ~^ reg672)) ?
                          reg838[(1'h0):(1'h0)] : forvar824));
                    end
                  for (forvar834 = (1'h0); (forvar834 < (2'h3)); forvar834 = (forvar834 + (1'h1)))
                    begin
                      reg835 <= $unsigned({{reg836[(1'h1):(1'h0)]}});
                      reg836 <= $signed((~&{(reg807 ^~ reg830)}));
                    end
                end
              if (((^~($unsigned(reg767) ?
                  {(8'h9f)} : $unsigned(reg708))) >= reg814))
                begin
                  for (forvar837 = (1'h0); (forvar837 < (1'h1)); forvar837 = (forvar837 + (1'h1)))
                    begin
                      reg838 <= $signed(($unsigned((reg764 ?
                          reg672 : reg761)) <<< $unsigned($unsigned(reg766))));
                    end
                  for (forvar839 = (1'h0); (forvar839 < (1'h0)); forvar839 = (forvar839 + (1'h1)))
                    begin
                      reg840 <= reg812[(4'ha):(1'h1)];
                      reg841 <= {forvar735};
                      reg842 <= reg842[(3'h6):(2'h3)];
                    end
                end
              else
                begin
                  reg837 <= $unsigned(wire665[(4'hc):(2'h3)]);
                  for (forvar838 = (1'h0); (forvar838 < (1'h1)); forvar838 = (forvar838 + (1'h1)))
                    begin
                      reg839 <= $signed(forvar707);
                      reg840 <= {$unsigned(((forvar669 - (8'hb4)) ~^ reg705))};
                      reg841 <= ({((forvar669 ? reg751 : (8'hb7)) ?
                                  $unsigned(reg732) : ((8'h9c) ?
                                      reg825 : reg848))} ?
                          reg757 : $signed(reg721));
                      reg842 <= (({(~&forvar751)} ?
                              (reg718[(3'h6):(3'h5)] ?
                                  (reg779 << reg671) : (!(8'hb0))) : $signed($signed(reg826))) ?
                          ((-(reg784 ? reg787 : forvar718)) <<< (+(reg742 ?
                              reg821 : reg710))) : $signed(reg757));
                    end
                end
            end
          reg843 <= reg733[(2'h2):(1'h0)];
          if (((!{(reg792 ^~ reg726)}) <= (~^{wire809})))
            begin
              if ($signed({reg684[(3'h5):(1'h0)]}))
                begin
                  for (forvar844 = (1'h0); (forvar844 < (2'h3)); forvar844 = (forvar844 + (1'h1)))
                    begin
                      reg845 <= (reg713 ?
                          reg757 : ({$unsigned(reg843)} ?
                              $unsigned(forvar667[(4'ha):(4'h8)]) : $signed(wire662)));
                      reg846 <= $unsigned(forvar717);
                      reg847 <= ((+reg794) ~^ (!reg833[(3'h6):(1'h1)]));
                    end
                  if ((^(^$signed($unsigned(reg746)))))
                    begin
                      reg848 <= ($signed({(reg741 >>> wire664)}) ?
                          (8'ha5) : $signed(({reg831} ~^ reg766)));
                      reg849 <= $signed($unsigned(({reg779} >>> (reg834 ?
                          reg726 : reg754))));
                      reg850 <= (reg775[(2'h3):(2'h2)] + (8'hab));
                      reg851 <= {(^~(~^$signed(reg750)))};
                    end
                  else
                    begin
                      reg848 <= ($unsigned(((reg819 ? reg750 : forvar707) ?
                              forvar810[(2'h2):(1'h0)] : (reg818 + reg797))) ?
                          (((forvar669 * forvar784) ?
                                  forvar737 : $signed(forvar785)) ?
                              $unsigned((reg798 || reg848)) : ($unsigned(reg677) ?
                                  $signed(reg763) : ((8'hac) ?
                                      reg776 : forvar750))) : (8'ha6));
                    end
                  reg852 <= {{$signed(reg832[(1'h0):(1'h0)])}};
                end
              else
                begin
                  for (forvar844 = (1'h0); (forvar844 < (2'h3)); forvar844 = (forvar844 + (1'h1)))
                    begin
                      reg845 <= $unsigned(reg774[(2'h2):(1'h0)]);
                    end
                  if (reg677)
                    begin
                      reg846 <= $signed((((reg677 ? reg823 : forvar810) ?
                          forvar817[(2'h2):(1'h1)] : (|(8'hb1))) && $signed($signed(forvar758))));
                      reg847 <= (~|(~|((~|reg748) ?
                          $unsigned(reg675) : reg835[(4'h8):(3'h7)])));
                      reg848 <= reg805[(3'h5):(2'h3)];
                      reg849 <= ({$signed(reg704)} ?
                          (((reg676 <<< reg852) >> $signed(reg726)) * ((~|reg749) ?
                              (&forvar683) : forvar834)) : {$unsigned($signed(reg780))});
                    end
                  else
                    begin
                      reg846 <= reg674[(1'h0):(1'h0)];
                      reg847 <= reg782[(1'h0):(1'h0)];
                    end
                  for (forvar850 = (1'h0); (forvar850 < (1'h0)); forvar850 = (forvar850 + (1'h1)))
                    begin
                      reg851 <= $unsigned($signed($signed(reg821)));
                    end
                end
              for (forvar853 = (1'h0); (forvar853 < (1'h1)); forvar853 = (forvar853 + (1'h1)))
                begin
                  for (forvar854 = (1'h0); (forvar854 < (1'h1)); forvar854 = (forvar854 + (1'h1)))
                    begin
                      reg855 <= reg784[(2'h3):(2'h2)];
                      reg856 <= $signed($unsigned(reg802));
                      reg857 <= $signed(($unsigned($signed(reg690)) ?
                          reg705[(2'h3):(1'h0)] : {$unsigned(reg813)}));
                    end
                  if (({$signed((!forvar710))} ?
                      reg713[(3'h4):(2'h3)] : (({reg721} << forvar850[(4'h9):(3'h4)]) == ($signed(reg802) - (forvar836 ?
                          reg783 : (8'hb4))))))
                    begin
                      reg858 <= $signed(forvar811[(2'h2):(1'h1)]);
                      reg859 <= (~($signed({reg755}) ?
                          $signed($signed(reg743)) : (reg725[(4'h8):(4'h8)] >> (&(8'ha7)))));
                    end
                  else
                    begin
                      reg858 <= reg704[(4'h9):(1'h0)];
                      reg859 <= $signed((!(forvar771[(2'h3):(1'h0)] & {reg668})));
                      reg860 <= ((-($unsigned(forvar673) ?
                              (reg741 ^~ reg829) : (~reg769))) ?
                          ((reg785[(3'h6):(3'h4)] ?
                                  (8'hac) : $unsigned(reg721)) ?
                              $unsigned({forvar763}) : (|{reg688})) : (^$unsigned((reg709 ?
                              forvar824 : reg694))));
                      reg861 <= $unsigned((^~(reg693 ?
                          (forvar784 ? reg729 : (8'h9e)) : {reg684})));
                    end
                  reg862 <= (~^(|reg848[(1'h0):(1'h0)]));
                end
              reg863 <= forvar666[(4'he):(3'h4)];
              for (forvar864 = (1'h0); (forvar864 < (2'h2)); forvar864 = (forvar864 + (1'h1)))
                begin
                  if ((^reg768))
                    begin
                      reg865 <= forvar704[(2'h3):(2'h3)];
                      reg866 <= reg831[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg865 <= $unsigned(($signed({(8'h9d)}) ?
                          (^~(~|forvar669)) : $signed(forvar736)));
                      reg866 <= (reg837 ?
                          reg746[(4'hd):(4'hc)] : reg845[(1'h1):(1'h0)]);
                      reg867 <= forvar753[(3'h7):(3'h5)];
                    end
                end
            end
          else
            begin
              reg844 <= $unsigned($signed((reg747[(3'h4):(2'h2)] ?
                  forvar735 : $unsigned(reg675))));
              for (forvar845 = (1'h0); (forvar845 < (2'h3)); forvar845 = (forvar845 + (1'h1)))
                begin
                  for (forvar846 = (1'h0); (forvar846 < (1'h1)); forvar846 = (forvar846 + (1'h1)))
                    begin
                      reg847 <= ((~&forvar811[(4'h9):(2'h3)]) ?
                          reg799 : (reg782[(1'h0):(1'h0)] >> {$signed(forvar854)}));
                      reg848 <= (+{(reg825 < reg785)});
                      reg849 <= (8'hae);
                      reg850 <= {(~|forvar697)};
                    end
                  for (forvar851 = (1'h0); (forvar851 < (2'h2)); forvar851 = (forvar851 + (1'h1)))
                    begin
                      reg852 <= reg672[(4'h8):(3'h6)];
                      reg853 <= $signed(reg841[(1'h0):(1'h0)]);
                      reg854 <= forvar666;
                    end
                  for (forvar855 = (1'h0); (forvar855 < (2'h3)); forvar855 = (forvar855 + (1'h1)))
                    begin
                      reg856 <= (forvar844[(3'h5):(1'h1)] != (&(~&(forvar692 ?
                          reg783 : forvar680))));
                    end
                end
            end
          if ({{((forvar813 ? (8'ha5) : (8'h9c)) ?
                      forvar697[(4'hf):(1'h1)] : ((8'ha5) || forvar789))}})
            begin
              if ($signed((8'hb1)))
                begin
                  reg868 <= reg807;
                end
              else
                begin
                  if ((reg686 ? $unsigned(reg760) : reg857))
                    begin
                      reg868 <= forvar822;
                      reg869 <= ($unsigned($signed((~(8'had)))) ?
                          $signed(forvar707) : (forvar832[(2'h2):(1'h1)] + (reg713 ?
                              $signed(reg766) : (forvar851 ~^ reg820))));
                    end
                  else
                    begin
                      reg868 <= (+{{(&(8'h9d))}});
                    end
                  reg870 <= {forvar816[(3'h5):(1'h0)]};
                end
              for (forvar871 = (1'h0); (forvar871 < (1'h1)); forvar871 = (forvar871 + (1'h1)))
                begin
                  if ((($signed($signed(reg766)) >>> reg672) && {forvar822[(1'h0):(1'h0)]}))
                    begin
                      reg872 <= ((-(8'ha3)) == ((&(~^reg795)) + ((forvar850 || (8'hb1)) != $signed(forvar744))));
                      reg873 <= forvar871[(3'h6):(2'h3)];
                      reg874 <= $unsigned($signed(((^~reg763) ?
                          (forvar838 | forvar838) : (|reg792))));
                    end
                  else
                    begin
                      reg872 <= ($unsigned((!$unsigned(reg790))) == ((+(~&reg755)) >>> reg796));
                      reg873 <= (~^{{{reg858}}});
                    end
                  for (forvar875 = (1'h0); (forvar875 < (1'h0)); forvar875 = (forvar875 + (1'h1)))
                    begin
                      reg876 <= ((reg771[(4'he):(4'he)] ?
                          ($signed(reg725) & (~reg752)) : ($signed(forvar750) ?
                              reg800 : {reg727})) >= ($unsigned({(8'ha8)}) && reg798[(1'h0):(1'h0)]));
                      reg877 <= (($unsigned((^~(8'hb2))) >> reg683) < ({$unsigned(reg838)} >> forvar864[(1'h0):(1'h0)]));
                    end
                  if ($unsigned(reg854))
                    begin
                      reg878 <= ($signed({reg716[(3'h6):(1'h0)]}) ?
                          (~|(((8'hba) ? reg727 : reg749) & (reg751 ?
                              forvar824 : reg820))) : {reg720});
                      reg879 <= ({($signed(reg857) ?
                                  $signed(forvar822) : (forvar875 ?
                                      reg794 : reg726))} ?
                          ((!{forvar708}) == reg836[(1'h1):(1'h0)]) : {reg774});
                    end
                  else
                    begin
                      reg878 <= ($signed(reg730) + ($signed((+forvar812)) <<< $unsigned(reg820)));
                      reg879 <= ((reg670[(1'h0):(1'h0)] ?
                              ((reg863 ? (8'haa) : reg769) ?
                                  reg861 : $unsigned(forvar839)) : (forvar718[(4'hf):(1'h1)] && (reg691 ?
                                  forvar673 : (8'hb3)))) ?
                          $signed(reg675) : $unsigned((-{reg750})));
                    end
                  if (reg828[(3'h4):(3'h4)])
                    begin
                      reg880 <= {$unsigned($unsigned({reg733}))};
                    end
                  else
                    begin
                      reg880 <= (({$signed(reg855)} ?
                              reg705 : reg765[(3'h4):(1'h0)]) ?
                          $unsigned(forvar715[(3'h4):(1'h1)]) : $signed(((8'haf) >> $signed((8'had)))));
                      reg881 <= $unsigned(reg865[(2'h2):(1'h0)]);
                      reg882 <= $unsigned(reg748[(1'h0):(1'h0)]);
                      reg883 <= $unsigned(((^~(reg855 ? forvar708 : reg757)) ?
                          (8'ha3) : $signed(reg783[(1'h1):(1'h1)])));
                    end
                end
              for (forvar884 = (1'h0); (forvar884 < (1'h1)); forvar884 = (forvar884 + (1'h1)))
                begin
                  for (forvar885 = (1'h0); (forvar885 < (1'h1)); forvar885 = (forvar885 + (1'h1)))
                    begin
                      reg886 <= reg763[(2'h3):(1'h1)];
                      reg887 <= {reg749};
                      reg888 <= (+(~&reg716));
                      reg889 <= reg803;
                    end
                  if (({reg691[(3'h6):(3'h5)]} ?
                      {((~|reg678) == reg703)} : (-$unsigned($signed(forvar785)))))
                    begin
                      reg890 <= (!((8'ha7) <<< reg756));
                      reg891 <= {reg730};
                      reg892 <= ({$signed((forvar702 ?
                              reg849 : reg776))} >= $signed({reg832}));
                      reg893 <= $signed({((reg891 ? reg781 : reg722) ?
                              $unsigned(reg713) : $unsigned(reg852))});
                    end
                  else
                    begin
                      reg890 <= $unsigned(({reg739[(1'h1):(1'h1)]} ?
                          forvar752[(4'h8):(3'h7)] : $unsigned((|forvar738))));
                      reg891 <= reg688;
                    end
                end
              for (forvar894 = (1'h0); (forvar894 < (1'h0)); forvar894 = (forvar894 + (1'h1)))
                begin
                  for (forvar895 = (1'h0); (forvar895 < (2'h3)); forvar895 = (forvar895 + (1'h1)))
                    begin
                      reg896 <= (((-forvar875) ?
                          ($signed(forvar710) ?
                              {(8'ha3)} : reg881[(3'h7):(1'h1)]) : reg869[(1'h0):(1'h0)]) * (($unsigned(reg672) & (reg694 ?
                          (8'hba) : (8'ha2))) >> ((+(8'ha8)) >> reg815[(3'h6):(3'h6)])));
                      reg897 <= {forvar679};
                      reg898 <= (^(~|reg878[(3'h5):(3'h4)]));
                    end
                  reg899 <= (reg691 * reg769[(3'h7):(2'h3)]);
                  if ((|(^reg805)))
                    begin
                      reg900 <= $signed({($signed(reg761) ?
                              (reg816 != reg747) : (8'hb4))});
                      reg901 <= $signed(reg710[(4'hd):(4'h8)]);
                      reg902 <= (~|(reg707 ? reg724 : forvar710));
                    end
                  else
                    begin
                      reg900 <= reg726[(4'hb):(3'h4)];
                      reg901 <= $signed(((reg711[(2'h2):(1'h0)] ?
                              (reg883 ? reg755 : reg889) : ((8'ha9) ?
                                  reg704 : forvar811)) ?
                          reg674 : $unsigned((reg734 >>> (8'ha6)))));
                      reg902 <= reg757[(2'h3):(1'h0)];
                    end
                  reg903 <= {reg843[(2'h3):(1'h0)]};
                end
            end
          else
            begin
              if ((|$unsigned($unsigned((reg869 ? (8'hb2) : reg710)))))
                begin
                  for (forvar868 = (1'h0); (forvar868 < (1'h0)); forvar868 = (forvar868 + (1'h1)))
                    begin
                      reg869 <= $signed((~&$unsigned((reg676 ?
                          reg748 : forvar806))));
                      reg870 <= reg892[(2'h3):(1'h1)];
                      reg871 <= ($signed(({forvar702} ?
                              $signed(wire808) : (reg759 ^ (8'ha2)))) ?
                          $signed($unsigned($unsigned(reg874))) : ($signed(((8'haa) != reg799)) + ((~&reg845) ?
                              $unsigned(reg857) : reg856)));
                      reg872 <= $unsigned($signed($signed({reg898})));
                    end
                end
              else
                begin
                  reg868 <= (~|((~&reg757) ?
                      $unsigned((reg675 ?
                          forvar771 : reg826)) : ($unsigned((8'hab)) != (reg833 ?
                          reg727 : forvar673))));
                  reg869 <= reg687[(3'h4):(3'h4)];
                end
            end
        end
    end
  assign wire904 = ((^~(!(reg689 * reg857))) < ((^~$unsigned(reg694)) ?
                       $unsigned(reg766[(1'h0):(1'h0)]) : $signed(reg765[(3'h5):(2'h3)])));
  always
    @(posedge clk) begin
      reg905 <= ((($signed(reg730) && (8'hb2)) << ({forvar735} ?
              $unsigned((8'ha3)) : forvar710[(1'h0):(1'h0)])) ?
          ({reg903} ^ ($signed(reg734) ?
              $unsigned(reg879) : ((8'hb4) <= reg703))) : forvar667);
      if (forvar682)
        begin
          if (reg683)
            begin
              if ({reg866[(2'h2):(2'h2)]})
                begin
                  reg906 <= {(~&$unsigned((~|reg848)))};
                  if ($unsigned(reg695))
                    begin
                      reg907 <= wire808[(2'h2):(1'h1)];
                      reg908 <= ($unsigned(reg703[(1'h0):(1'h0)]) ?
                          $unsigned(reg838) : reg724);
                      reg909 <= {forvar772};
                    end
                  else
                    begin
                      reg907 <= reg848;
                      reg908 <= wire664[(4'hb):(2'h2)];
                      reg909 <= wire904[(3'h4):(3'h4)];
                      reg910 <= reg813[(1'h1):(1'h0)];
                    end
                  for (forvar911 = (1'h0); (forvar911 < (2'h3)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= {forvar847};
                      reg913 <= (reg726 <= $unsigned((^{(8'hba)})));
                      reg914 <= $unsigned($signed($unsigned((|reg815))));
                    end
                end
              else
                begin
                  for (forvar906 = (1'h0); (forvar906 < (1'h1)); forvar906 = (forvar906 + (1'h1)))
                    begin
                      reg907 <= (~forvar758[(2'h3):(2'h2)]);
                      reg908 <= $unsigned({(^reg724[(1'h1):(1'h0)])});
                      reg909 <= forvar742;
                      reg910 <= ({((reg675 ?
                              reg827 : reg703) < (8'hb0))} ~^ wire904);
                    end
                  for (forvar911 = (1'h0); (forvar911 < (1'h0)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= reg840;
                      reg913 <= reg900[(2'h2):(1'h0)];
                    end
                end
            end
          else
            begin
              if ({reg713})
                begin
                  if ($signed(reg896[(3'h7):(3'h6)]))
                    begin
                      reg906 <= ((^reg909) ? (8'ha5) : reg834);
                    end
                  else
                    begin
                      reg906 <= (wire662[(4'h9):(3'h4)] ?
                          $unsigned(reg888[(4'hb):(2'h3)]) : reg890);
                      reg907 <= $signed($unsigned(reg811));
                      reg908 <= ($unsigned((8'hb1)) ?
                          ($signed($signed((8'hb8))) >> (~&(&reg677))) : $unsigned(($signed(reg790) > (reg731 - (8'hac)))));
                      reg909 <= (reg896[(3'h5):(3'h5)] ?
                          (^~$unsigned({(8'hb7)})) : $unsigned({(forvar753 ?
                                  reg743 : reg857)}));
                    end
                  reg910 <= {wire665[(3'h5):(2'h3)]};
                  for (forvar911 = (1'h0); (forvar911 < (1'h0)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= forvar753[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar906 = (1'h0); (forvar906 < (2'h2)); forvar906 = (forvar906 + (1'h1)))
                    begin
                      reg907 <= $unsigned(($signed((^reg892)) >> $unsigned(forvar758[(3'h5):(2'h3)])));
                    end
                  reg908 <= $unsigned(reg872);
                  for (forvar909 = (1'h0); (forvar909 < (2'h2)); forvar909 = (forvar909 + (1'h1)))
                    begin
                      reg910 <= $unsigned(reg723[(1'h0):(1'h0)]);
                      reg911 <= (reg837[(1'h0):(1'h0)] ?
                          ($signed($unsigned(forvar744)) <= ((^~reg889) ?
                              $signed((8'ha4)) : (-reg866))) : (forvar699 && $signed($signed((8'hae)))));
                      reg912 <= ((reg805 < ($unsigned(forvar894) > reg690[(1'h0):(1'h0)])) + (^reg855));
                    end
                  if ($unsigned(((~&(^reg862)) ~^ (~&$unsigned(forvar666)))))
                    begin
                      reg913 <= reg907[(3'h4):(2'h2)];
                      reg914 <= $unsigned($unsigned(reg751[(2'h3):(1'h1)]));
                    end
                  else
                    begin
                      reg913 <= (forvar834[(2'h3):(1'h0)] <= (forvar666[(4'hb):(1'h1)] >>> ($unsigned((8'hb5)) ?
                          $signed(reg846) : reg883)));
                    end
                end
              for (forvar915 = (1'h0); (forvar915 < (2'h3)); forvar915 = (forvar915 + (1'h1)))
                begin
                  for (forvar916 = (1'h0); (forvar916 < (2'h3)); forvar916 = (forvar916 + (1'h1)))
                    begin
                      reg917 <= ($signed((~|$signed(forvar746))) ?
                          reg881[(2'h2):(1'h0)] : forvar906);
                    end
                  if ($unsigned((reg859 >= reg907)))
                    begin
                      reg918 <= (((reg825[(3'h4):(3'h4)] ^~ reg693[(1'h1):(1'h1)]) ?
                          (reg798[(2'h2):(2'h2)] ^ (reg729 ?
                              forvar772 : reg862)) : {{reg882}}) | reg798);
                      reg919 <= $unsigned(reg812[(3'h4):(1'h0)]);
                      reg920 <= ($unsigned(($unsigned(forvar812) && ((8'ha5) <<< reg770))) ?
                          forvar666[(4'h8):(2'h2)] : ({reg909[(1'h1):(1'h1)]} ?
                              (^(~|reg760)) : reg690[(3'h6):(3'h5)]));
                    end
                  else
                    begin
                      reg918 <= $unsigned($signed(forvar817[(3'h5):(2'h2)]));
                      reg919 <= forvar751;
                      reg920 <= $signed((^~(reg863[(1'h1):(1'h0)] - (forvar667 & reg677))));
                    end
                  for (forvar921 = (1'h0); (forvar921 < (2'h3)); forvar921 = (forvar921 + (1'h1)))
                    begin
                      reg922 <= (^wire661);
                    end
                  for (forvar923 = (1'h0); (forvar923 < (2'h2)); forvar923 = (forvar923 + (1'h1)))
                    begin
                      reg924 <= {(!reg896)};
                      reg925 <= (8'hb6);
                    end
                end
              for (forvar926 = (1'h0); (forvar926 < (1'h0)); forvar926 = (forvar926 + (1'h1)))
                begin
                  if (((8'h9d) ?
                      ((8'ha6) ?
                          $unsigned($signed(forvar692)) : ((forvar717 >> reg868) ?
                              $signed(forvar751) : $unsigned(forvar680))) : {$signed((~|reg725))}))
                    begin
                      reg927 <= {{forvar718[(4'hf):(3'h6)]}};
                      reg928 <= ($unsigned(reg831[(2'h2):(2'h2)]) & (8'hae));
                    end
                  else
                    begin
                      reg927 <= {$signed(reg782)};
                    end
                  for (forvar929 = (1'h0); (forvar929 < (2'h3)); forvar929 = (forvar929 + (1'h1)))
                    begin
                      reg930 <= forvar747[(2'h2):(2'h2)];
                    end
                  if ((^reg681))
                    begin
                      reg931 <= reg729;
                      reg932 <= $unsigned(($signed($unsigned(reg920)) ~^ reg928));
                    end
                  else
                    begin
                      reg931 <= {forvar710[(1'h1):(1'h0)]};
                      reg932 <= ($signed((-(forvar801 >= reg788))) ?
                          ($unsigned((forvar714 ?
                              (8'hb6) : reg912)) ^ (forvar926 == $unsigned(reg785))) : {reg928});
                      reg933 <= (reg927 & ($unsigned($signed(reg910)) ?
                          $signed(reg759[(3'h7):(1'h0)]) : (forvar692[(1'h1):(1'h0)] <<< {reg906})));
                    end
                  reg934 <= {$unsigned($unsigned((forvar754 * forvar771)))};
                end
            end
        end
      else
        begin
          reg906 <= $signed({$signed($unsigned(reg799))});
          reg907 <= (($unsigned({forvar753}) ?
              ((-reg817) ?
                  $unsigned(reg695) : reg671) : $signed(reg732[(4'h9):(1'h0)])) != (|{(reg862 ^ reg876)}));
          for (forvar908 = (1'h0); (forvar908 < (2'h3)); forvar908 = (forvar908 + (1'h1)))
            begin
              for (forvar909 = (1'h0); (forvar909 < (2'h2)); forvar909 = (forvar909 + (1'h1)))
                begin
                  if (($unsigned(forvar753) ?
                      (8'ha7) : ((8'hae) ? {(~&reg901)} : (^$signed(reg706)))))
                    begin
                      reg910 <= $unsigned((reg888 ?
                          $signed((reg851 ?
                              reg824 : reg859)) : ($unsigned(reg914) - (reg674 ?
                              forvar846 : forvar853))));
                      reg911 <= $signed((-((reg792 ? reg865 : (8'ha7)) ?
                          reg699 : (reg743 ? reg825 : reg932))));
                    end
                  else
                    begin
                      reg910 <= {reg787[(3'h6):(2'h2)]};
                      reg911 <= ((+($signed(reg847) || ((8'hb6) ?
                          forvar735 : reg839))) ^ (~|(forvar921[(1'h1):(1'h1)] == $signed(reg837))));
                    end
                end
              if ((|$signed($signed({reg826}))))
                begin
                  if (reg909)
                    begin
                      reg912 <= {$signed(($unsigned(reg733) ?
                              (^~reg701) : $unsigned(wire661)))};
                      reg913 <= ($unsigned(((reg674 ? reg880 : (8'hb2)) ?
                              reg870[(1'h1):(1'h1)] : reg748)) ?
                          reg774 : reg845);
                      reg914 <= (|$signed(reg759[(4'h8):(3'h5)]));
                    end
                  else
                    begin
                      reg912 <= reg741;
                      reg913 <= (~&{{(reg814 ? reg763 : reg752)}});
                    end
                  reg915 <= ((reg780 ?
                          (reg702[(3'h5):(2'h2)] >> forvar871) : $signed((^~reg882))) ?
                      (+$signed($unsigned(reg857))) : (reg840[(1'h1):(1'h0)] << {$unsigned(reg917)}));
                  if ((forvar702 < $unsigned(((8'ha4) ?
                      $unsigned(reg754) : (reg767 || reg832)))))
                    begin
                      reg916 <= ($unsigned(reg777[(1'h1):(1'h1)]) ?
                          $unsigned(reg877) : {(8'ha0)});
                      reg917 <= ({$unsigned($unsigned((8'hb8)))} ?
                          $unsigned(((reg764 ? forvar847 : reg868) ?
                              (reg702 ?
                                  reg880 : reg687) : {reg677})) : (|$signed($signed(reg790))));
                      reg918 <= reg675;
                    end
                  else
                    begin
                      reg916 <= {forvar702};
                    end
                  for (forvar919 = (1'h0); (forvar919 < (2'h3)); forvar919 = (forvar919 + (1'h1)))
                    begin
                      reg920 <= $unsigned((reg748 - (|$signed(reg785))));
                      reg921 <= ({($signed(reg787) ?
                              reg716[(2'h2):(1'h1)] : (~&forvar763))} <<< forvar850[(4'h9):(4'h9)]);
                      reg922 <= reg683;
                    end
                end
              else
                begin
                  for (forvar912 = (1'h0); (forvar912 < (2'h2)); forvar912 = (forvar912 + (1'h1)))
                    begin
                      reg913 <= $signed(($unsigned((reg934 ?
                              forvar923 : reg796)) ?
                          {$signed(forvar667)} : reg686));
                      reg914 <= $unsigned($signed((8'h9c)));
                    end
                  for (forvar915 = (1'h0); (forvar915 < (2'h3)); forvar915 = (forvar915 + (1'h1)))
                    begin
                      reg916 <= {reg670};
                      reg917 <= forvar679;
                    end
                end
              for (forvar923 = (1'h0); (forvar923 < (1'h0)); forvar923 = (forvar923 + (1'h1)))
                begin
                  reg924 <= reg788;
                  if (forvar704[(1'h0):(1'h0)])
                    begin
                      reg925 <= $unsigned(($unsigned({(8'hae)}) ?
                          (^~(|reg922)) : forvar717[(3'h5):(3'h4)]));
                      reg926 <= {(+$unsigned((-reg858)))};
                      reg927 <= ($signed($unsigned((reg814 ?
                          forvar915 : reg874))) ^ (8'ha7));
                      reg928 <= $unsigned($unsigned((8'ha8)));
                    end
                  else
                    begin
                      reg925 <= $unsigned(reg712);
                      reg926 <= ((8'hab) != reg816);
                      reg927 <= (|((^{forvar906}) <= $unsigned((~reg826))));
                      reg928 <= reg686;
                    end
                  for (forvar929 = (1'h0); (forvar929 < (2'h2)); forvar929 = (forvar929 + (1'h1)))
                    begin
                      reg930 <= (((&(reg831 <<< (8'hb2))) ?
                              (reg838 ?
                                  reg797[(1'h1):(1'h1)] : $signed((8'hb0))) : {$unsigned(reg749)}) ?
                          (&($signed(forvar772) ?
                              $signed(forvar778) : $signed(reg882))) : (|$signed({reg764})));
                      reg931 <= forvar752;
                    end
                end
            end
        end
    end
  assign wire935 = $unsigned(wire662[(3'h5):(3'h5)]);
  always
    @(posedge clk) begin
      for (forvar936 = (1'h0); (forvar936 < (2'h2)); forvar936 = (forvar936 + (1'h1)))
        begin
          for (forvar937 = (1'h0); (forvar937 < (1'h0)); forvar937 = (forvar937 + (1'h1)))
            begin
              if ($signed(reg817[(1'h1):(1'h0)]))
                begin
                  reg938 <= (8'hb2);
                  for (forvar939 = (1'h0); (forvar939 < (1'h1)); forvar939 = (forvar939 + (1'h1)))
                    begin
                      reg940 <= (reg866 ~^ reg826[(4'hc):(3'h4)]);
                    end
                  for (forvar941 = (1'h0); (forvar941 < (2'h3)); forvar941 = (forvar941 + (1'h1)))
                    begin
                      reg942 <= {({(~&reg707)} ?
                              reg766 : (reg890 ?
                                  reg751[(3'h6):(1'h0)] : (reg853 ?
                                      reg731 : reg688)))};
                      reg943 <= (^~(|(((8'hba) ~^ (8'ha9)) - reg694[(2'h2):(1'h1)])));
                      reg944 <= (8'ha9);
                      reg945 <= $unsigned(reg816[(3'h7):(3'h7)]);
                    end
                end
              else
                begin
                  if (forvar812[(1'h1):(1'h0)])
                    begin
                      reg938 <= (forvar850[(1'h0):(1'h0)] ^ (forvar855 < {(reg686 ?
                              (8'hb9) : forvar885)}));
                      reg939 <= (($unsigned(((8'hac) ? reg786 : reg684)) ?
                              $unsigned((8'ha0)) : ((reg928 | forvar929) | $unsigned(reg845))) ?
                          ({{forvar747}} <= {reg860[(1'h1):(1'h1)]}) : ($signed($signed(reg762)) ?
                              (reg740 ?
                                  reg695[(3'h7):(3'h7)] : {wire663}) : (^~(wire662 & reg814))));
                    end
                  else
                    begin
                      reg938 <= (~($signed((forvar834 <= reg720)) ?
                          (reg820 >> (forvar845 ?
                              forvar785 : reg785)) : $unsigned((reg708 ?
                              reg854 : (8'haf)))));
                      reg939 <= ($unsigned(reg741[(2'h3):(2'h3)]) ?
                          $unsigned(((forvar752 ? reg749 : reg945) ?
                              (+reg766) : $unsigned(reg775))) : reg807);
                      reg940 <= $signed(((&{reg748}) ?
                          $unsigned((reg862 < reg707)) : (~&reg943[(3'h7):(3'h7)])));
                    end
                  for (forvar941 = (1'h0); (forvar941 < (1'h0)); forvar941 = (forvar941 + (1'h1)))
                    begin
                      reg942 <= $signed({((reg840 ~^ reg800) ?
                              (&reg872) : wire662[(4'h9):(3'h5)])});
                      reg943 <= (&(reg795 ?
                          {forvar850[(3'h4):(1'h0)]} : reg671[(4'ha):(3'h4)]));
                      reg944 <= reg752[(2'h2):(1'h0)];
                      reg945 <= $unsigned(($signed($signed(reg931)) * (reg750[(3'h6):(1'h1)] ?
                          (reg766 >>> (8'hb0)) : (forvar929 ?
                              reg907 : reg874))));
                    end
                end
              reg946 <= (reg899[(1'h0):(1'h0)] && {{reg706}});
              for (forvar947 = (1'h0); (forvar947 < (1'h1)); forvar947 = (forvar947 + (1'h1)))
                begin
                  for (forvar948 = (1'h0); (forvar948 < (2'h2)); forvar948 = (forvar948 + (1'h1)))
                    begin
                      reg949 <= (reg696 * $unsigned(($signed(forvar752) ?
                          (reg707 ? reg896 : (8'h9d)) : reg871)));
                      reg950 <= $signed(reg709);
                    end
                  reg951 <= ((+$signed($unsigned(reg677))) ?
                      $signed(($signed(reg770) << (forvar923 ?
                          forvar838 : reg761))) : forvar772);
                  if ({$unsigned(reg796[(4'h8):(2'h3)])})
                    begin
                      reg952 <= forvar679[(1'h1):(1'h0)];
                      reg953 <= ((8'ha2) ~^ $unsigned((reg722[(3'h5):(3'h5)] ?
                          forvar707 : $signed(forvar773))));
                      reg954 <= ((($unsigned(forvar868) ?
                          (reg749 ?
                              reg892 : (8'hb3)) : $signed(reg741)) || forvar948[(2'h2):(1'h0)]) > reg891);
                    end
                  else
                    begin
                      reg952 <= ((!(forvar699[(1'h1):(1'h1)] ?
                          (-reg691) : reg892[(3'h6):(1'h1)])) ^~ (&$unsigned({reg914})));
                      reg953 <= ($signed((|$signed(forvar939))) < reg819[(2'h3):(1'h0)]);
                      reg954 <= reg694[(1'h0):(1'h0)];
                    end
                end
            end
          if ((~&reg903[(2'h2):(1'h0)]))
            begin
              for (forvar955 = (1'h0); (forvar955 < (2'h3)); forvar955 = (forvar955 + (1'h1)))
                begin
                  for (forvar956 = (1'h0); (forvar956 < (1'h1)); forvar956 = (forvar956 + (1'h1)))
                    begin
                      reg957 <= $unsigned(reg698[(1'h1):(1'h0)]);
                      reg958 <= (+$unsigned((|$unsigned(forvar714))));
                    end
                  if ($unsigned(reg760))
                    begin
                      reg959 <= ($unsigned(($unsigned(reg887) ?
                          $signed(reg934) : $unsigned(reg684))) == (reg920[(1'h1):(1'h0)] != reg681[(3'h7):(3'h5)]));
                      reg960 <= ($signed($unsigned(reg732)) ?
                          (reg674 | forvar668[(2'h2):(1'h1)]) : reg766[(3'h6):(3'h4)]);
                      reg961 <= (8'h9d);
                    end
                  else
                    begin
                      reg959 <= reg730;
                    end
                end
            end
          else
            begin
              for (forvar955 = (1'h0); (forvar955 < (2'h2)); forvar955 = (forvar955 + (1'h1)))
                begin
                  for (forvar956 = (1'h0); (forvar956 < (1'h1)); forvar956 = (forvar956 + (1'h1)))
                    begin
                      reg957 <= reg852[(4'h9):(3'h5)];
                      reg958 <= $signed(forvar785[(2'h2):(1'h0)]);
                      reg959 <= $unsigned(($signed((reg841 ? reg758 : reg695)) ?
                          (+$unsigned(reg838)) : ($signed(wire935) ?
                              (|reg828) : (~&reg831))));
                    end
                  for (forvar960 = (1'h0); (forvar960 < (1'h1)); forvar960 = (forvar960 + (1'h1)))
                    begin
                      reg961 <= forvar916;
                      reg962 <= (forvar687 ?
                          (^~$unsigned((~&forvar948))) : $unsigned((~&(forvar850 ?
                              wire665 : reg677))));
                      reg963 <= forvar832[(3'h7):(1'h0)];
                      reg964 <= {(reg907[(2'h2):(1'h1)] ?
                              reg945[(2'h2):(1'h1)] : ({forvar744} ?
                                  reg918 : forvar687[(1'h1):(1'h1)]))};
                    end
                  reg965 <= ((($unsigned(forvar937) > forvar692) ^ reg678[(3'h6):(1'h0)]) >>> $unsigned(forvar719));
                end
            end
          for (forvar966 = (1'h0); (forvar966 < (2'h3)); forvar966 = (forvar966 + (1'h1)))
            begin
              reg967 <= {$unsigned(($unsigned(reg741) ? reg745 : {reg883}))};
              if ((^(^(^{reg813}))))
                begin
                  if (($signed(((~reg760) - (reg696 ?
                      reg771 : forvar708))) ~^ ($signed(reg920[(1'h0):(1'h0)]) ?
                      {forvar845[(1'h1):(1'h1)]} : $signed(((8'had) & reg930)))))
                    begin
                      reg968 <= reg850[(4'hb):(3'h4)];
                      reg969 <= (~$signed((reg774 > $unsigned(forvar854))));
                    end
                  else
                    begin
                      reg968 <= $signed((8'hae));
                      reg969 <= $signed($unsigned((8'ha3)));
                    end
                  for (forvar970 = (1'h0); (forvar970 < (1'h0)); forvar970 = (forvar970 + (1'h1)))
                    begin
                      reg971 <= $unsigned($unsigned($unsigned({forvar844})));
                      reg972 <= $signed($unsigned($signed({reg685})));
                    end
                  if ($signed($unsigned(reg675)))
                    begin
                      reg973 <= (reg790[(3'h6):(1'h1)] > (~|$signed((reg879 <= forvar801))));
                      reg974 <= $unsigned(($signed((reg891 ?
                          (8'haa) : reg710)) < {$signed(forvar884)}));
                      reg975 <= $unsigned({reg828[(3'h5):(3'h4)]});
                      reg976 <= (forvar714[(3'h7):(1'h0)] ?
                          reg794[(4'hb):(3'h7)] : reg774);
                    end
                  else
                    begin
                      reg973 <= ((($signed(reg790) <<< $unsigned(forvar742)) ?
                              forvar806[(2'h3):(1'h0)] : reg668[(4'ha):(3'h5)]) ?
                          (reg938 ?
                              {reg957[(3'h5):(1'h1)]} : $signed((+reg724))) : {$unsigned(reg676[(3'h7):(3'h5)])});
                      reg974 <= ($signed(($signed(reg780) ?
                          (reg681 ?
                              reg854 : wire663) : wire661[(3'h6):(2'h3)])) ^~ ($unsigned(((8'hb5) ?
                              reg795 : reg793)) ?
                          {reg893[(3'h4):(2'h3)]} : ($unsigned((8'ha9)) ?
                              (^reg921) : (forvar909 >> (8'hb1)))));
                      reg975 <= {forvar747[(2'h3):(2'h2)]};
                    end
                end
              else
                begin
                  for (forvar968 = (1'h0); (forvar968 < (1'h0)); forvar968 = (forvar968 + (1'h1)))
                    begin
                      reg969 <= {(($signed(forvar936) <= (~|forvar847)) >> ($unsigned(forvar845) ?
                              reg957[(3'h4):(3'h4)] : forvar836))};
                      reg970 <= $signed(reg785);
                      reg971 <= reg790;
                      reg972 <= $signed($unsigned($signed((~&reg896))));
                    end
                end
            end
          reg977 <= $unsigned((~^((reg920 ? (8'hb5) : wire935) != {reg832})));
        end
      if ($signed((~^reg916[(3'h6):(3'h6)])))
        begin
          reg978 <= ($unsigned(((forvar708 ^~ reg951) ?
              reg701[(3'h5):(2'h2)] : $signed(forvar822))) && (~|$signed(reg756)));
        end
      else
        begin
          if (reg868)
            begin
              if ((~reg827[(4'hf):(3'h7)]))
                begin
                  if ($unsigned(((reg933[(2'h2):(2'h2)] ^ (forvar707 ?
                      reg838 : reg669)) < (~$unsigned(forvar699)))))
                    begin
                      reg978 <= (8'hac);
                    end
                  else
                    begin
                      reg978 <= reg859[(3'h5):(3'h5)];
                      reg979 <= $unsigned(forvar936[(4'h8):(2'h2)]);
                    end
                  if ((8'hb1))
                    begin
                      reg980 <= {reg835[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg980 <= {forvar669[(4'h9):(1'h1)]};
                    end
                  reg981 <= (reg832[(2'h2):(2'h2)] ?
                      reg918 : $unsigned($signed(forvar784)));
                end
              else
                begin
                  for (forvar978 = (1'h0); (forvar978 < (2'h2)); forvar978 = (forvar978 + (1'h1)))
                    begin
                      reg979 <= (reg916[(3'h4):(3'h4)] ?
                          (~^(8'h9c)) : {{$signed(reg716)}});
                      reg980 <= (+(((~&(8'ha3)) ?
                              (forvar855 ? forvar778 : reg963) : {reg814}) ?
                          reg903[(1'h1):(1'h0)] : ($unsigned(forvar968) >>> (!(8'h9f)))));
                      reg981 <= forvar742;
                    end
                  if (reg722)
                    begin
                      reg982 <= ((((forvar704 >> reg793) <= {reg672}) <= {{forvar847}}) || reg963[(1'h1):(1'h0)]);
                      reg983 <= $signed(forvar839[(4'he):(4'hc)]);
                      reg984 <= ($unsigned($signed(reg765)) ?
                          reg968 : $unsigned({(reg783 ? reg953 : reg916)}));
                      reg985 <= ($signed(((forvar680 == reg862) ?
                              $unsigned(forvar839) : $unsigned(reg983))) ?
                          $signed($signed({forvar683})) : (forvar666[(3'h7):(3'h5)] | reg747[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg982 <= {{((!reg725) ?
                                  (forvar912 | reg708) : reg897[(2'h3):(1'h0)])}};
                      reg983 <= $unsigned((($unsigned(reg972) ?
                              (8'hb3) : $unsigned(forvar746)) ?
                          {(reg893 || (8'ha8))} : ((~|reg879) ?
                              {reg784} : (|reg852))));
                      reg984 <= ({(reg826 ?
                              $signed(reg886) : (reg688 ?
                                  (8'h9c) : forvar824))} || reg982[(3'h6):(3'h6)]);
                      reg985 <= ({reg693} ?
                          ($signed(forvar894[(4'h8):(3'h6)]) ?
                              reg781 : {(reg848 ?
                                      forvar864 : reg867)}) : ({$unsigned(reg709)} ?
                              forvar817 : {(wire661 ? reg976 : reg905)}));
                    end
                  for (forvar986 = (1'h0); (forvar986 < (1'h1)); forvar986 = (forvar986 + (1'h1)))
                    begin
                      reg987 <= ((^$signed((-reg746))) - $signed(({reg950} & (forvar911 ?
                          (8'hb7) : reg827))));
                      reg988 <= ($unsigned((&(reg788 < reg693))) >>> forvar960[(4'ha):(3'h5)]);
                    end
                end
            end
          else
            begin
              for (forvar978 = (1'h0); (forvar978 < (1'h1)); forvar978 = (forvar978 + (1'h1)))
                begin
                  reg979 <= $unsigned(forvar919[(3'h5):(3'h5)]);
                end
              reg980 <= (~^$signed((~^(^reg766))));
              reg981 <= (reg865 ? $signed(reg823) : {$signed({reg938})});
              for (forvar982 = (1'h0); (forvar982 < (2'h2)); forvar982 = (forvar982 + (1'h1)))
                begin
                  for (forvar983 = (1'h0); (forvar983 < (1'h0)); forvar983 = (forvar983 + (1'h1)))
                    begin
                      reg984 <= (~&(&$signed((forvar875 != reg775))));
                      reg985 <= (~|(reg855 + {{reg959}}));
                      reg986 <= (!$signed($signed((reg711 && forvar692))));
                    end
                  if (({$unsigned(reg776)} ?
                      reg774 : ({$unsigned((8'had))} ?
                          (reg747[(2'h2):(1'h1)] << forvar737[(2'h2):(1'h1)]) : (8'ha4))))
                    begin
                      reg987 <= (forvar750[(1'h1):(1'h1)] && reg691[(2'h3):(1'h1)]);
                      reg988 <= ($signed(forvar919) ?
                          (reg891 << $unsigned(forvar966[(1'h1):(1'h1)])) : ($unsigned(wire664[(4'hb):(3'h7)]) ?
                              $signed(reg938[(3'h6):(1'h0)]) : $signed(reg713[(3'h4):(1'h0)])));
                      reg989 <= (|{reg919[(1'h0):(1'h0)]});
                    end
                  else
                    begin
                      reg987 <= (|({$signed(forvar906)} != {(~|reg881)}));
                      reg988 <= $unsigned($signed($unsigned(forvar921)));
                      reg989 <= reg677[(1'h0):(1'h0)];
                      reg990 <= ({{(forvar824 > reg828)}} ?
                          {(+$signed(reg918))} : $signed(reg984[(3'h5):(3'h5)]));
                    end
                  reg991 <= (forvar699[(1'h0):(1'h0)] > reg745);
                  reg992 <= wire664;
                end
            end
          if ($signed((reg756[(2'h2):(1'h1)] ^ $unsigned((+reg694)))))
            begin
              if (($unsigned(reg677[(1'h1):(1'h0)]) | {$signed($unsigned(reg765))}))
                begin
                  for (forvar993 = (1'h0); (forvar993 < (1'h1)); forvar993 = (forvar993 + (1'h1)))
                    begin
                      reg994 <= {forvar753[(4'h8):(2'h2)]};
                      reg995 <= ($signed((8'ha8)) - $unsigned({(&reg770)}));
                      reg996 <= $unsigned({(8'ha0)});
                      reg997 <= (|$signed((-{reg819})));
                    end
                  for (forvar998 = (1'h0); (forvar998 < (1'h0)); forvar998 = (forvar998 + (1'h1)))
                    begin
                      reg999 <= $unsigned((8'ha7));
                      reg1000 <= $signed($unsigned($unsigned((~forvar763))));
                      reg1001 <= ($unsigned($unsigned({forvar919})) == ($unsigned((8'hae)) ?
                          $unsigned(reg881[(4'h8):(2'h3)]) : $unsigned($unsigned(reg769))));
                      reg1002 <= (&$signed($unsigned((^~reg886))));
                    end
                  reg1003 <= $unsigned((~|$signed($signed(reg670))));
                  if ((reg669 >= {((8'hb1) >> (reg870 ? reg712 : reg932))}))
                    begin
                      reg1004 <= ((-$signed((~&reg668))) ^ $signed(forvar746));
                      reg1005 <= (($unsigned({reg776}) << reg739) ?
                          reg786 : ((((8'h9d) ?
                              reg926 : reg759) * $signed(reg836)) <= ((8'h9f) >= (reg865 ?
                              reg721 : reg967))));
                    end
                  else
                    begin
                      reg1004 <= $signed($unsigned(($signed(forvar707) <<< $unsigned((8'had)))));
                    end
                end
              else
                begin
                  for (forvar993 = (1'h0); (forvar993 < (2'h2)); forvar993 = (forvar993 + (1'h1)))
                    begin
                      reg994 <= ((8'h9d) | ((8'h9c) ~^ ((reg741 ^~ reg959) ?
                          (forvar774 <<< (8'had)) : (-reg732))));
                      reg995 <= $unsigned({($unsigned(reg838) << $unsigned((8'hb2)))});
                      reg996 <= ($unsigned((forvar895[(2'h3):(2'h3)] ?
                          (reg802 << reg762) : (reg724 || (8'hb4)))) <= $signed(($unsigned((8'h9d)) >>> (|reg731))));
                      reg997 <= (reg716 ? forvar806[(3'h4):(3'h4)] : reg965);
                    end
                end
              for (forvar1006 = (1'h0); (forvar1006 < (2'h2)); forvar1006 = (forvar1006 + (1'h1)))
                begin
                  for (forvar1007 = (1'h0); (forvar1007 < (1'h1)); forvar1007 = (forvar1007 + (1'h1)))
                    begin
                      reg1008 <= $unsigned((($unsigned(reg987) ?
                              $signed(reg981) : (~|reg770)) ?
                          $unsigned({forvar679}) : forvar845[(2'h2):(1'h0)]));
                      reg1009 <= forvar719;
                      reg1010 <= (($signed(((8'hb2) & reg707)) >>> (|(reg940 ?
                          reg1005 : reg743))) << reg757[(3'h4):(2'h2)]);
                      reg1011 <= (~^(forvar926 ?
                          (reg798 << (^reg882)) : reg672[(3'h6):(3'h4)]));
                    end
                  if (reg1003)
                    begin
                      reg1012 <= $signed({($unsigned(forvar806) ?
                              (reg767 ? forvar846 : forvar772) : reg833)});
                      reg1013 <= $signed((((~|reg897) ?
                              (forvar778 ?
                                  reg816 : reg982) : (reg718 ~^ reg722)) ?
                          reg811[(4'ha):(3'h5)] : ($signed(forvar855) <= (reg739 >>> reg860))));
                      reg1014 <= (^($signed({reg860}) + reg913));
                    end
                  else
                    begin
                      reg1012 <= $signed(($unsigned({reg683}) >> (reg741[(1'h1):(1'h1)] > (^~reg836))));
                      reg1013 <= forvar906;
                      reg1014 <= $unsigned($signed(forvar789[(4'he):(4'ha)]));
                      reg1015 <= reg714[(3'h4):(3'h4)];
                    end
                  if ((!$signed($unsigned((~forvar921)))))
                    begin
                      reg1016 <= $signed(forvar736);
                      reg1017 <= $signed($unsigned((reg687[(1'h0):(1'h0)] ?
                          (~^reg930) : (reg786 ? reg742 : reg1003))));
                      reg1018 <= $unsigned(reg866);
                    end
                  else
                    begin
                      reg1016 <= {((((8'hb3) ?
                                  reg792 : reg970) >> $signed(reg685)) ?
                              ((reg867 << reg1011) - (forvar911 ?
                                  forvar687 : reg690)) : $signed({forvar884}))};
                      reg1017 <= reg676[(3'h7):(2'h3)];
                      reg1018 <= (forvar909[(4'hc):(3'h5)] ?
                          {reg857[(2'h3):(2'h3)]} : reg827[(3'h5):(3'h4)]);
                      reg1019 <= {$signed((+$signed(forvar839)))};
                    end
                  for (forvar1020 = (1'h0); (forvar1020 < (1'h0)); forvar1020 = (forvar1020 + (1'h1)))
                    begin
                      reg1021 <= $signed($signed($signed($unsigned(reg826))));
                    end
                end
            end
          else
            begin
              if ($unsigned(($signed((reg757 ? reg897 : reg760)) ?
                  (~|(-reg922)) : ($signed(reg865) ? (8'ha8) : forvar673))))
                begin
                  reg993 <= $signed((-{(&reg709)}));
                  if ((reg973 ?
                      forvar773 : $unsigned((reg711 ?
                          ((8'hb3) ? reg794 : forvar923) : reg814))))
                    begin
                      reg994 <= forvar839[(4'hd):(2'h2)];
                    end
                  else
                    begin
                      reg994 <= forvar710[(2'h2):(1'h0)];
                      reg995 <= $signed($unsigned(($signed(reg967) + (-reg977))));
                    end
                  for (forvar996 = (1'h0); (forvar996 < (2'h3)); forvar996 = (forvar996 + (1'h1)))
                    begin
                      reg997 <= ({(reg731[(4'h8):(1'h1)] ?
                                  $signed(reg826) : $signed(reg732))} ?
                          ((8'hb3) ?
                              ({reg933} ?
                                  (forvar847 ?
                                      forvar1006 : reg802) : reg814) : {$signed(forvar746)}) : $unsigned((|$signed(reg781))));
                      reg998 <= (reg850[(2'h2):(1'h1)] ?
                          (~|((~|reg882) ?
                              $unsigned(reg925) : {reg816})) : (&forvar871));
                      reg999 <= $unsigned($signed(forvar668));
                      reg1000 <= forvar998;
                    end
                end
              else
                begin
                  for (forvar993 = (1'h0); (forvar993 < (1'h0)); forvar993 = (forvar993 + (1'h1)))
                    begin
                      reg994 <= forvar923;
                    end
                  if ($signed(((+reg868[(2'h3):(1'h0)]) <<< (-$signed(forvar785)))))
                    begin
                      reg995 <= wire665[(3'h6):(2'h2)];
                      reg996 <= reg813[(3'h4):(1'h1)];
                      reg997 <= reg847;
                    end
                  else
                    begin
                      reg995 <= reg749;
                      reg996 <= reg998[(2'h3):(2'h3)];
                      reg997 <= $unsigned((|forvar699[(1'h0):(1'h0)]));
                    end
                end
              for (forvar1001 = (1'h0); (forvar1001 < (2'h3)); forvar1001 = (forvar1001 + (1'h1)))
                begin
                  for (forvar1002 = (1'h0); (forvar1002 < (2'h2)); forvar1002 = (forvar1002 + (1'h1)))
                    begin
                      reg1003 <= $unsigned(reg869[(3'h7):(3'h6)]);
                      reg1004 <= (~$signed(reg766));
                      reg1005 <= reg891[(1'h0):(1'h0)];
                      reg1006 <= (($signed((-(8'ha5))) || {forvar680}) ^~ forvar742);
                    end
                  for (forvar1007 = (1'h0); (forvar1007 < (1'h0)); forvar1007 = (forvar1007 + (1'h1)))
                    begin
                      reg1008 <= (forvar837 ?
                          (~|($unsigned(forvar993) ?
                              (8'ha9) : $unsigned(reg704))) : ({((8'ha4) ^~ reg897)} * (&{reg1010})));
                      reg1009 <= {reg872[(1'h0):(1'h0)]};
                    end
                end
              reg1010 <= $signed($signed($unsigned(reg708)));
              reg1011 <= forvar923[(4'h9):(3'h4)];
            end
          for (forvar1022 = (1'h0); (forvar1022 < (2'h3)); forvar1022 = (forvar1022 + (1'h1)))
            begin
              for (forvar1023 = (1'h0); (forvar1023 < (1'h1)); forvar1023 = (forvar1023 + (1'h1)))
                begin
                  if (wire663[(1'h0):(1'h0)])
                    begin
                      reg1024 <= $signed({(((8'ha0) ^~ forvar774) ?
                              reg845[(3'h6):(3'h5)] : forvar707[(4'h9):(4'h8)])});
                    end
                  else
                    begin
                      reg1024 <= $unsigned($signed(($unsigned((8'ha2)) ^ (reg775 ?
                          reg994 : reg807))));
                      reg1025 <= ((~^reg828[(2'h3):(2'h2)]) ?
                          forvar763[(3'h5):(3'h5)] : (!$signed((&reg868))));
                      reg1026 <= $unsigned(forvar817);
                      reg1027 <= (+({(8'h9e)} ?
                          $signed($unsigned(reg968)) : reg961));
                    end
                end
            end
          if ($unsigned($unsigned((~^(reg768 << reg870)))))
            begin
              for (forvar1028 = (1'h0); (forvar1028 < (2'h2)); forvar1028 = (forvar1028 + (1'h1)))
                begin
                  for (forvar1029 = (1'h0); (forvar1029 < (1'h1)); forvar1029 = (forvar1029 + (1'h1)))
                    begin
                      reg1030 <= (forvar853 > reg757);
                      reg1031 <= (forvar763 ?
                          ($signed($signed(forvar708)) | ((reg888 == reg775) < (wire935 ?
                              forvar810 : reg1027))) : (-((8'hb9) | (reg779 ?
                              reg815 : reg759))));
                      reg1032 <= ((forvar735[(4'ha):(1'h1)] << (^~(forvar744 ?
                              reg714 : reg984))) ?
                          $unsigned(reg836[(1'h1):(1'h0)]) : $unsigned((~|$unsigned(reg730))));
                    end
                end
              for (forvar1033 = (1'h0); (forvar1033 < (1'h1)); forvar1033 = (forvar1033 + (1'h1)))
                begin
                  reg1034 <= reg683;
                end
              for (forvar1035 = (1'h0); (forvar1035 < (2'h3)); forvar1035 = (forvar1035 + (1'h1)))
                begin
                  for (forvar1036 = (1'h0); (forvar1036 < (2'h2)); forvar1036 = (forvar1036 + (1'h1)))
                    begin
                      reg1037 <= reg797;
                      reg1038 <= ((^$unsigned({reg903})) ?
                          (((reg781 | forvar710) & (reg845 ^~ reg930)) << ((^forvar1022) ?
                              (reg800 - reg788) : (reg893 >>> reg734))) : reg981[(3'h4):(3'h4)]);
                      reg1039 <= forvar909;
                    end
                  for (forvar1040 = (1'h0); (forvar1040 < (1'h1)); forvar1040 = (forvar1040 + (1'h1)))
                    begin
                      reg1041 <= ((-(reg901[(2'h2):(1'h0)] ?
                              reg908[(1'h1):(1'h0)] : reg861[(1'h1):(1'h0)])) ?
                          (reg1016[(4'h9):(4'h9)] ~^ ((reg850 ?
                              forvar812 : forvar955) + (reg865 && (8'ha0)))) : {{forvar744}});
                    end
                end
              for (forvar1042 = (1'h0); (forvar1042 < (2'h2)); forvar1042 = (forvar1042 + (1'h1)))
                begin
                  reg1043 <= (-({((8'hba) ^~ reg930)} ?
                      $unsigned($unsigned(forvar812)) : (~(reg825 ?
                          (8'hac) : reg851))));
                  for (forvar1044 = (1'h0); (forvar1044 < (1'h1)); forvar1044 = (forvar1044 + (1'h1)))
                    begin
                      reg1045 <= (~&reg890[(1'h1):(1'h1)]);
                    end
                  if ((^(((|(8'ha9)) ? (&forvar923) : forvar916) ?
                      reg727[(4'hd):(3'h5)] : (-(~&reg1019)))))
                    begin
                      reg1046 <= (~((!(reg803 ^~ reg739)) <<< ($signed(reg761) == {forvar810})));
                      reg1047 <= $unsigned((reg705 * (8'had)));
                      reg1048 <= $signed($signed($unsigned({(8'h9c)})));
                      reg1049 <= reg1039[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg1046 <= reg826;
                      reg1047 <= (+$unsigned($signed(forvar936[(3'h6):(3'h5)])));
                      reg1048 <= reg918;
                    end
                end
            end
          else
            begin
              for (forvar1028 = (1'h0); (forvar1028 < (2'h2)); forvar1028 = (forvar1028 + (1'h1)))
                begin
                  for (forvar1029 = (1'h0); (forvar1029 < (1'h0)); forvar1029 = (forvar1029 + (1'h1)))
                    begin
                      reg1030 <= reg919;
                    end
                  reg1031 <= ((forvar753 < (forvar829 < forvar871)) & forvar960[(3'h6):(2'h3)]);
                  if ((reg669[(2'h2):(2'h2)] >> ((-(reg765 ?
                      (8'hb7) : reg1015)) <= reg800)))
                    begin
                      reg1032 <= $unsigned(($unsigned((~^reg833)) ?
                          $unsigned((~&reg699)) : $signed((~reg990))));
                      reg1033 <= {(|(~^$signed(forvar850)))};
                    end
                  else
                    begin
                      reg1032 <= ($signed($unsigned((reg704 ?
                              reg1027 : reg807))) ?
                          forvar941 : reg795[(1'h0):(1'h0)]);
                      reg1033 <= (reg901[(2'h2):(1'h0)] > reg882[(2'h2):(2'h2)]);
                    end
                  for (forvar1034 = (1'h0); (forvar1034 < (1'h1)); forvar1034 = (forvar1034 + (1'h1)))
                    begin
                      reg1035 <= reg829[(1'h1):(1'h0)];
                      reg1036 <= {forvar885[(1'h0):(1'h0)]};
                    end
                end
            end
        end
    end
  assign wire1050 = (reg856[(5'h10):(3'h6)] ?
                        ($signed((reg755 ? reg828 : forvar853)) ?
                            $unsigned(reg959) : ((reg830 ? (8'hb1) : reg695) ?
                                (reg725 < forvar816) : (~reg846))) : ($signed((reg949 - reg868)) >>> ((~^(8'ha2)) ?
                            reg845 : (&forvar1020))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3367
#( parameter param3630 = ((+(((8'ha8) >= (8'ha4)) ? (+(8'h9e)) : ((8'hb8) | (8'ha7)))) * ((&((8'ha6) >> (8'hac))) ^ (-((8'hb0) > (8'h9f))))) )
(y, clk, wire3368, wire3369, wire3370, wire3371, wire3372);
  output wire [(32'haa9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire3368;
  input wire signed [(4'hb):(1'h0)] wire3369;
  input wire [(3'h4):(1'h0)] wire3370;
  input wire [(3'h4):(1'h0)] wire3371;
  input wire signed [(3'h6):(1'h0)] wire3372;
  wire signed [(4'hb):(1'h0)] wire3629;
  wire [(4'hd):(1'h0)] wire3628;
  reg signed [(2'h2):(1'h0)] reg3627 = (1'h0);
  reg [(3'h7):(1'h0)] reg3626 = (1'h0);
  reg [(3'h6):(1'h0)] reg3625 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3624 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3623 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3622 = (1'h0);
  reg [(4'hd):(1'h0)] reg3621 = (1'h0);
  reg [(4'hd):(1'h0)] reg3620 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3619 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3618 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3617 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3616 = (1'h0);
  wire [(3'h5):(1'h0)] wire3615;
  wire [(3'h6):(1'h0)] wire3614;
  wire signed [(4'hf):(1'h0)] wire3613;
  reg [(2'h3):(1'h0)] reg3612 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3611 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3610 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3609 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3608 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3598 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3590 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3585 = (1'h0);
  reg [(5'h10):(1'h0)] reg3576 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3604 = (1'h0);
  reg [(3'h6):(1'h0)] reg3603 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3595 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3592 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3587 = (1'h0);
  reg [(3'h6):(1'h0)] reg3584 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3583 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3582 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3580 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3577 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3574 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3569 = (1'h0);
  reg [(3'h5):(1'h0)] reg3567 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3566 = (1'h0);
  reg [(4'h8):(1'h0)] reg3563 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3562 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3560 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3556 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3555 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3608 = (1'h0);
  reg [(3'h7):(1'h0)] reg3607 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3606 = (1'h0);
  reg [(3'h6):(1'h0)] reg3605 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3604 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3603 = (1'h0);
  reg [(4'he):(1'h0)] forvar3600 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3597 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3596 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3602 = (1'h0);
  reg [(4'he):(1'h0)] reg3601 = (1'h0);
  reg [(4'ha):(1'h0)] reg3600 = (1'h0);
  reg [(4'hd):(1'h0)] reg3599 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3598 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3597 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3596 = (1'h0);
  reg [(4'he):(1'h0)] forvar3595 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3594 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3593 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3592 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3591 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3590 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3589 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3588 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3587 = (1'h0);
  reg [(4'h8):(1'h0)] reg3586 = (1'h0);
  reg [(4'hb):(1'h0)] reg3585 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3584 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3583 = (1'h0);
  reg [(4'hd):(1'h0)] reg3582 = (1'h0);
  reg [(4'hd):(1'h0)] reg3581 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3580 = (1'h0);
  reg [(3'h7):(1'h0)] reg3579 = (1'h0);
  reg [(2'h2):(1'h0)] reg3578 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3577 = (1'h0);
  reg [(4'he):(1'h0)] forvar3576 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3572 = (1'h0);
  reg [(4'hc):(1'h0)] reg3568 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3575 = (1'h0);
  reg [(4'h9):(1'h0)] reg3574 = (1'h0);
  reg [(4'hf):(1'h0)] reg3573 = (1'h0);
  reg [(3'h4):(1'h0)] reg3572 = (1'h0);
  reg [(3'h5):(1'h0)] reg3571 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3570 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3569 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3568 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3567 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3559 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3558 = (1'h0);
  reg [(4'hb):(1'h0)] reg3566 = (1'h0);
  reg [(3'h7):(1'h0)] reg3565 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3564 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3563 = (1'h0);
  reg [(3'h5):(1'h0)] reg3562 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3561 = (1'h0);
  reg [(4'h9):(1'h0)] reg3560 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3559 = (1'h0);
  reg [(3'h6):(1'h0)] reg3552 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3551 = (1'h0);
  reg [(4'ha):(1'h0)] reg3550 = (1'h0);
  reg [(3'h4):(1'h0)] reg3548 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3547 = (1'h0);
  reg [(3'h5):(1'h0)] reg3558 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3557 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3556 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3555 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3554 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3553 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3552 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3551 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3550 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3549 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3548 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3547 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3546 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3545 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3544 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3543 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3542 = (1'h0);
  reg [(2'h2):(1'h0)] reg3541 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3540 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3539 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3538 = (1'h0);
  reg [(4'hd):(1'h0)] reg3537 = (1'h0);
  reg [(4'hd):(1'h0)] reg3536 = (1'h0);
  reg [(4'h9):(1'h0)] reg3535 = (1'h0);
  reg [(3'h7):(1'h0)] reg3534 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3533 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3532 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3531 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3530 = (1'h0);
  reg [(3'h6):(1'h0)] reg3529 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3528 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3527 = (1'h0);
  reg [(3'h4):(1'h0)] reg3526 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3525 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3524 = (1'h0);
  reg [(3'h6):(1'h0)] reg3523 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3522 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3521 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3520 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3519 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3518 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3517 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3516 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3515 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3514 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3513 = (1'h0);
  reg [(4'ha):(1'h0)] reg3511 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3512 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3511 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3510 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3509 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3508 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3496 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3500 = (1'h0);
  reg [(3'h4):(1'h0)] reg3499 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3498 = (1'h0);
  reg [(4'ha):(1'h0)] reg3495 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3491 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3490 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3488 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3507 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3506 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3503 = (1'h0);
  reg [(4'he):(1'h0)] reg3506 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3505 = (1'h0);
  reg [(4'hc):(1'h0)] reg3504 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3503 = (1'h0);
  reg [(3'h6):(1'h0)] reg3502 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3501 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3500 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3499 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3498 = (1'h0);
  reg [(3'h5):(1'h0)] reg3497 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3496 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3495 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3494 = (1'h0);
  reg [(4'h8):(1'h0)] reg3493 = (1'h0);
  reg [(4'hc):(1'h0)] reg3492 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3491 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3490 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3489 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3488 = (1'h0);
  reg [(4'he):(1'h0)] reg3485 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3478 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3474 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3487 = (1'h0);
  reg [(4'h8):(1'h0)] reg3486 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3485 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3484 = (1'h0);
  reg [(4'hc):(1'h0)] reg3483 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3482 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3481 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3480 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3469 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3464 = (1'h0);
  reg [(3'h7):(1'h0)] reg3458 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3456 = (1'h0);
  reg [(4'hc):(1'h0)] reg3481 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3480 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3476 = (1'h0);
  reg [(3'h6):(1'h0)] reg3479 = (1'h0);
  reg [(3'h6):(1'h0)] reg3478 = (1'h0);
  reg [(3'h7):(1'h0)] reg3477 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3476 = (1'h0);
  reg [(4'h8):(1'h0)] reg3475 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3474 = (1'h0);
  reg [(4'hd):(1'h0)] reg3473 = (1'h0);
  reg [(2'h2):(1'h0)] reg3472 = (1'h0);
  reg [(3'h4):(1'h0)] reg3471 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3470 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3469 = (1'h0);
  reg [(4'hb):(1'h0)] reg3468 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3465 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3467 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3466 = (1'h0);
  reg [(4'h9):(1'h0)] reg3465 = (1'h0);
  reg [(2'h2):(1'h0)] reg3464 = (1'h0);
  reg [(3'h6):(1'h0)] reg3463 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3462 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3461 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3460 = (1'h0);
  reg [(4'he):(1'h0)] reg3459 = (1'h0);
  reg [(4'he):(1'h0)] forvar3458 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3457 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3456 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3455 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3454 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3453 = (1'h0);
  reg [(4'hd):(1'h0)] reg3452 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3451 = (1'h0);
  reg [(4'ha):(1'h0)] reg3450 = (1'h0);
  reg [(4'he):(1'h0)] reg3449 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3448 = (1'h0);
  reg [(4'hd):(1'h0)] reg3447 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3446 = (1'h0);
  reg [(4'hd):(1'h0)] reg3445 = (1'h0);
  reg [(3'h5):(1'h0)] reg3444 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3443 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3442 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3441 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3440 = (1'h0);
  reg [(4'hf):(1'h0)] reg3439 = (1'h0);
  wire [(2'h2):(1'h0)] wire3373;
  wire signed [(3'h6):(1'h0)] wire3374;
  wire signed [(4'hf):(1'h0)] wire3375;
  reg [(5'h10):(1'h0)] forvar3376 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3377 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3378 = (1'h0);
  reg [(4'hf):(1'h0)] reg3379 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3380 = (1'h0);
  reg [(4'hc):(1'h0)] reg3381 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3382 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3383 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3384 = (1'h0);
  reg [(2'h3):(1'h0)] reg3385 = (1'h0);
  reg [(5'h10):(1'h0)] reg3377 = (1'h0);
  reg [(4'ha):(1'h0)] reg3386 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3387 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3388 = (1'h0);
  reg [(3'h5):(1'h0)] reg3389 = (1'h0);
  reg [(2'h2):(1'h0)] reg3390 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3391 = (1'h0);
  reg [(3'h5):(1'h0)] reg3392 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3393 = (1'h0);
  reg [(5'h10):(1'h0)] reg3394 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3395 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3396 = (1'h0);
  reg [(4'hc):(1'h0)] reg3397 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3398 = (1'h0);
  reg [(4'he):(1'h0)] reg3399 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3400 = (1'h0);
  reg [(3'h4):(1'h0)] reg3401 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3402 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3403 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3404 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3405 = (1'h0);
  reg [(3'h6):(1'h0)] reg3406 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3407 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3408 = (1'h0);
  reg [(4'ha):(1'h0)] reg3409 = (1'h0);
  reg [(3'h5):(1'h0)] reg3410 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3411 = (1'h0);
  reg [(3'h4):(1'h0)] reg3387 = (1'h0);
  reg [(4'he):(1'h0)] reg3388 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3386 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3393 = (1'h0);
  reg [(4'h9):(1'h0)] reg3395 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3396 = (1'h0);
  reg [(4'ha):(1'h0)] reg3398 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3399 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3412 = (1'h0);
  reg [(3'h4):(1'h0)] reg3413 = (1'h0);
  wire [(5'h10):(1'h0)] wire3414;
  wire signed [(4'hf):(1'h0)] wire3415;
  wire signed [(2'h2):(1'h0)] wire3437;
  assign y = {wire3629,
                 wire3628,
                 reg3627,
                 reg3626,
                 reg3625,
                 forvar3624,
                 reg3623,
                 forvar3622,
                 reg3621,
                 reg3620,
                 forvar3619,
                 forvar3618,
                 forvar3617,
                 forvar3616,
                 wire3615,
                 wire3614,
                 wire3613,
                 reg3612,
                 reg3611,
                 reg3610,
                 reg3609,
                 forvar3608,
                 forvar3598,
                 forvar3590,
                 forvar3585,
                 reg3576,
                 reg3604,
                 reg3603,
                 reg3595,
                 forvar3592,
                 reg3587,
                 reg3584,
                 reg3583,
                 forvar3582,
                 forvar3580,
                 reg3577,
                 forvar3574,
                 forvar3569,
                 reg3567,
                 forvar3566,
                 reg3563,
                 forvar3562,
                 forvar3560,
                 forvar3556,
                 forvar3555,
                 reg3608,
                 reg3607,
                 reg3606,
                 reg3605,
                 forvar3604,
                 forvar3603,
                 forvar3600,
                 forvar3597,
                 reg3596,
                 reg3602,
                 reg3601,
                 reg3600,
                 reg3599,
                 reg3598,
                 reg3597,
                 forvar3596,
                 forvar3595,
                 reg3594,
                 reg3593,
                 reg3592,
                 reg3591,
                 reg3590,
                 reg3589,
                 reg3588,
                 forvar3587,
                 reg3586,
                 reg3585,
                 forvar3584,
                 forvar3583,
                 reg3582,
                 reg3581,
                 reg3580,
                 reg3579,
                 reg3578,
                 forvar3577,
                 forvar3576,
                 forvar3572,
                 reg3568,
                 reg3575,
                 reg3574,
                 reg3573,
                 reg3572,
                 reg3571,
                 reg3570,
                 reg3569,
                 forvar3568,
                 forvar3567,
                 reg3559,
                 forvar3558,
                 reg3566,
                 reg3565,
                 reg3564,
                 forvar3563,
                 reg3562,
                 reg3561,
                 reg3560,
                 forvar3559,
                 reg3552,
                 forvar3551,
                 reg3550,
                 reg3548,
                 forvar3547,
                 reg3558,
                 reg3557,
                 reg3556,
                 reg3555,
                 reg3554,
                 reg3553,
                 forvar3552,
                 reg3551,
                 forvar3550,
                 reg3549,
                 forvar3548,
                 reg3547,
                 reg3546,
                 forvar3545,
                 reg3544,
                 reg3543,
                 reg3542,
                 reg3541,
                 reg3540,
                 reg3539,
                 reg3538,
                 reg3537,
                 reg3536,
                 reg3535,
                 reg3534,
                 forvar3533,
                 reg3532,
                 reg3531,
                 forvar3530,
                 reg3529,
                 reg3528,
                 reg3527,
                 reg3526,
                 reg3525,
                 forvar3524,
                 reg3523,
                 forvar3522,
                 forvar3521,
                 reg3520,
                 reg3519,
                 forvar3518,
                 reg3517,
                 reg3516,
                 forvar3515,
                 reg3514,
                 reg3513,
                 reg3511,
                 reg3512,
                 forvar3511,
                 forvar3510,
                 reg3509,
                 forvar3508,
                 forvar3496,
                 forvar3500,
                 reg3499,
                 reg3498,
                 reg3495,
                 forvar3491,
                 reg3490,
                 reg3488,
                 reg3507,
                 forvar3506,
                 reg3503,
                 reg3506,
                 reg3505,
                 reg3504,
                 forvar3503,
                 reg3502,
                 reg3501,
                 reg3500,
                 forvar3499,
                 forvar3498,
                 reg3497,
                 reg3496,
                 forvar3495,
                 reg3494,
                 reg3493,
                 reg3492,
                 reg3491,
                 forvar3490,
                 reg3489,
                 forvar3488,
                 reg3485,
                 forvar3478,
                 forvar3474,
                 reg3487,
                 reg3486,
                 forvar3485,
                 reg3484,
                 reg3483,
                 reg3482,
                 forvar3481,
                 reg3480,
                 forvar3469,
                 forvar3464,
                 reg3458,
                 reg3456,
                 reg3481,
                 forvar3480,
                 reg3476,
                 reg3479,
                 reg3478,
                 reg3477,
                 forvar3476,
                 reg3475,
                 reg3474,
                 reg3473,
                 reg3472,
                 reg3471,
                 reg3470,
                 reg3469,
                 reg3468,
                 forvar3465,
                 reg3467,
                 reg3466,
                 reg3465,
                 reg3464,
                 reg3463,
                 reg3462,
                 reg3461,
                 reg3460,
                 reg3459,
                 forvar3458,
                 reg3457,
                 forvar3456,
                 forvar3455,
                 forvar3454,
                 reg3453,
                 reg3452,
                 reg3451,
                 reg3450,
                 reg3449,
                 forvar3448,
                 reg3447,
                 forvar3446,
                 reg3445,
                 reg3444,
                 forvar3443,
                 forvar3442,
                 forvar3441,
                 forvar3440,
                 reg3439,
                 wire3373,
                 wire3374,
                 wire3375,
                 forvar3376,
                 forvar3377,
                 forvar3378,
                 reg3379,
                 reg3380,
                 reg3381,
                 reg3382,
                 forvar3383,
                 reg3384,
                 reg3385,
                 reg3377,
                 reg3386,
                 forvar3387,
                 forvar3388,
                 reg3389,
                 reg3390,
                 reg3391,
                 reg3392,
                 forvar3393,
                 reg3394,
                 forvar3395,
                 forvar3396,
                 reg3397,
                 forvar3398,
                 reg3399,
                 reg3400,
                 reg3401,
                 forvar3402,
                 reg3403,
                 reg3404,
                 forvar3405,
                 reg3406,
                 reg3407,
                 reg3408,
                 reg3409,
                 reg3410,
                 reg3411,
                 reg3387,
                 reg3388,
                 forvar3386,
                 reg3393,
                 reg3395,
                 reg3396,
                 reg3398,
                 forvar3399,
                 reg3412,
                 reg3413,
                 wire3414,
                 wire3415,
                 wire3437,
                 (1'h0)};
  assign wire3373 = (~&($signed($unsigned(wire3369)) * wire3370[(2'h3):(2'h2)]));
  assign wire3374 = $unsigned(wire3373);
  assign wire3375 = $unsigned((~$unsigned($unsigned(wire3373))));
  always
    @(posedge clk) begin
      for (forvar3376 = (1'h0); (forvar3376 < (1'h0)); forvar3376 = (forvar3376 + (1'h1)))
        begin
          if ($signed($signed((forvar3376[(4'hc):(4'h9)] ^~ {wire3370}))))
            begin
              for (forvar3377 = (1'h0); (forvar3377 < (2'h3)); forvar3377 = (forvar3377 + (1'h1)))
                begin
                  for (forvar3378 = (1'h0); (forvar3378 < (1'h1)); forvar3378 = (forvar3378 + (1'h1)))
                    begin
                      reg3379 <= (&$unsigned($signed((^~wire3373))));
                      reg3380 <= forvar3377;
                      reg3381 <= $unsigned(((^wire3371[(1'h0):(1'h0)]) ?
                          {(-reg3380)} : ({wire3372} - ((8'ha9) + forvar3378))));
                      reg3382 <= ({($signed(forvar3376) ?
                                  (wire3369 ~^ forvar3377) : (~|wire3374))} ?
                          ({(reg3381 ? (8'ha4) : forvar3376)} ?
                              (wire3372 < (8'h9c)) : wire3375) : (-wire3373[(2'h2):(2'h2)]));
                    end
                  for (forvar3383 = (1'h0); (forvar3383 < (2'h3)); forvar3383 = (forvar3383 + (1'h1)))
                    begin
                      reg3384 <= $signed($signed((wire3369[(3'h7):(3'h7)] < (-reg3381))));
                      reg3385 <= forvar3378[(3'h4):(1'h0)];
                    end
                end
            end
          else
            begin
              reg3377 <= (8'h9f);
            end
          if ($signed(wire3368))
            begin
              reg3386 <= {($unsigned(wire3371[(1'h1):(1'h0)]) ~^ (+$unsigned(wire3374)))};
              for (forvar3387 = (1'h0); (forvar3387 < (1'h0)); forvar3387 = (forvar3387 + (1'h1)))
                begin
                  for (forvar3388 = (1'h0); (forvar3388 < (2'h3)); forvar3388 = (forvar3388 + (1'h1)))
                    begin
                      reg3389 <= $signed($signed((~reg3386[(3'h4):(1'h1)])));
                      reg3390 <= ($unsigned({(reg3386 ?
                              wire3374 : forvar3376)}) ~^ $unsigned(forvar3387));
                      reg3391 <= {(^$signed(reg3386[(1'h1):(1'h1)]))};
                      reg3392 <= reg3389[(1'h0):(1'h0)];
                    end
                  for (forvar3393 = (1'h0); (forvar3393 < (1'h0)); forvar3393 = (forvar3393 + (1'h1)))
                    begin
                      reg3394 <= forvar3378;
                    end
                end
              for (forvar3395 = (1'h0); (forvar3395 < (1'h1)); forvar3395 = (forvar3395 + (1'h1)))
                begin
                  for (forvar3396 = (1'h0); (forvar3396 < (1'h1)); forvar3396 = (forvar3396 + (1'h1)))
                    begin
                      reg3397 <= ((^~forvar3383) ^~ reg3381[(3'h6):(1'h1)]);
                    end
                  for (forvar3398 = (1'h0); (forvar3398 < (1'h0)); forvar3398 = (forvar3398 + (1'h1)))
                    begin
                      reg3399 <= (reg3392 ^~ (!reg3381));
                      reg3400 <= (~|forvar3395);
                      reg3401 <= (&(~&$unsigned({(8'h9f)})));
                    end
                  for (forvar3402 = (1'h0); (forvar3402 < (2'h2)); forvar3402 = (forvar3402 + (1'h1)))
                    begin
                      reg3403 <= $unsigned(((reg3401 ?
                          $signed((8'haa)) : (-wire3368)) >= reg3380));
                      reg3404 <= $unsigned($unsigned(reg3386));
                    end
                end
              for (forvar3405 = (1'h0); (forvar3405 < (1'h0)); forvar3405 = (forvar3405 + (1'h1)))
                begin
                  if (reg3399)
                    begin
                      reg3406 <= $unsigned(($unsigned((reg3379 ~^ forvar3395)) ?
                          ((8'hae) ?
                              wire3368 : reg3403[(2'h2):(1'h0)]) : reg3389[(3'h5):(2'h3)]));
                    end
                  else
                    begin
                      reg3406 <= $signed((forvar3388[(4'h9):(1'h0)] ?
                          (^$unsigned(forvar3377)) : reg3400[(3'h7):(3'h6)]));
                      reg3407 <= ((^{forvar3396[(1'h1):(1'h1)]}) == {reg3390[(1'h0):(1'h0)]});
                    end
                  if ($signed(($unsigned((&forvar3396)) ^~ $signed($signed(reg3382)))))
                    begin
                      reg3408 <= forvar3395[(2'h3):(2'h2)];
                      reg3409 <= (|(({reg3404} + forvar3402) ?
                          {reg3386} : ((reg3381 + forvar3395) << $signed(forvar3402))));
                    end
                  else
                    begin
                      reg3408 <= (reg3408 ?
                          (~&$unsigned(reg3377)) : (^~$signed((reg3379 ?
                              reg3385 : reg3379))));
                      reg3409 <= (&$signed(($unsigned(reg3407) <= forvar3393)));
                      reg3410 <= $unsigned({reg3397});
                      reg3411 <= {$signed(wire3373)};
                    end
                end
            end
          else
            begin
              if ((+({forvar3395} ?
                  $unsigned($unsigned((8'hb9))) : (-(~reg3409)))))
                begin
                  if ((((-$unsigned(forvar3398)) ?
                      reg3397[(3'h6):(3'h6)] : $signed(wire3372)) | $signed(reg3386)))
                    begin
                      reg3386 <= $unsigned(reg3409);
                    end
                  else
                    begin
                      reg3386 <= ({$signed((~|reg3401))} ?
                          $signed((^(forvar3376 * (8'h9d)))) : (^~(8'ha4)));
                      reg3387 <= (reg3389 ? wire3369 : (!$signed(reg3391)));
                      reg3388 <= reg3409;
                    end
                end
              else
                begin
                  for (forvar3386 = (1'h0); (forvar3386 < (2'h2)); forvar3386 = (forvar3386 + (1'h1)))
                    begin
                      reg3387 <= reg3388;
                    end
                  if ({wire3373[(2'h2):(1'h1)]})
                    begin
                      reg3388 <= (~^(wire3375 ?
                          {(reg3386 && reg3380)} : $signed((!forvar3395))));
                      reg3389 <= $signed($unsigned($signed((reg3386 ?
                          reg3390 : reg3400))));
                    end
                  else
                    begin
                      reg3388 <= ((($unsigned(reg3391) ?
                                  $signed(forvar3383) : (^wire3374)) ?
                              $signed((reg3404 && reg3385)) : reg3408) ?
                          (~^$signed(((8'h9e) ^~ wire3371))) : (forvar3393[(2'h2):(1'h1)] ?
                              ((reg3409 || (8'hb4)) >> (forvar3378 ?
                                  reg3379 : reg3391)) : $unsigned(((8'ha7) * wire3370))));
                    end
                  reg3390 <= $unsigned((~((reg3390 & reg3387) && (^reg3411))));
                  if ((({$signed((8'ha0))} ^~ reg3409[(3'h7):(1'h0)]) ?
                      reg3382[(1'h0):(1'h0)] : (((wire3371 - (8'hb0)) ?
                          (reg3409 * reg3379) : (reg3404 ?
                              reg3399 : reg3407)) <<< $unsigned(reg3380[(1'h0):(1'h0)]))))
                    begin
                      reg3391 <= ((((reg3377 ? reg3385 : (8'h9c)) ?
                              (reg3382 ?
                                  reg3410 : (8'hb5)) : $signed((8'hb0))) ?
                          wire3374[(2'h2):(1'h0)] : $unsigned(forvar3377[(2'h2):(1'h0)])) >= $unsigned($unsigned(reg3401[(1'h1):(1'h1)])));
                      reg3392 <= $signed(((((8'hb0) ?
                          (8'hb7) : reg3404) || {reg3399}) | $unsigned($unsigned((8'haf)))));
                      reg3393 <= $signed((&$unsigned($unsigned(reg3377))));
                      reg3394 <= ((forvar3378 ?
                          {forvar3376[(1'h0):(1'h0)]} : forvar3395) >>> $unsigned(reg3404[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg3391 <= ({($unsigned(reg3391) - $unsigned(forvar3386))} * (forvar3388 ?
                          (reg3397[(4'h8):(3'h4)] >> (wire3370 ^~ (8'h9c))) : (wire3374 > $unsigned(reg3397))));
                      reg3392 <= forvar3387;
                    end
                end
              if (($signed((^~$unsigned(reg3377))) >> $unsigned(reg3388)))
                begin
                  if ((8'ha0))
                    begin
                      reg3395 <= $signed(forvar3398[(2'h3):(1'h0)]);
                      reg3396 <= {$signed(reg3391)};
                      reg3397 <= (~&{reg3391[(2'h2):(1'h1)]});
                    end
                  else
                    begin
                      reg3395 <= $unsigned(reg3403);
                      reg3396 <= (~^((~&(reg3400 ~^ wire3375)) ?
                          forvar3386 : {(reg3410 | reg3388)}));
                      reg3397 <= forvar3383;
                      reg3398 <= $signed((-($signed(reg3411) * (|reg3393))));
                    end
                end
              else
                begin
                  if (reg3382)
                    begin
                      reg3395 <= forvar3386;
                      reg3396 <= (+$unsigned(forvar3378[(4'hc):(2'h2)]));
                    end
                  else
                    begin
                      reg3395 <= (reg3377[(2'h3):(1'h1)] ?
                          $unsigned((&reg3381[(3'h4):(1'h1)])) : $unsigned((reg3379 ?
                              (reg3398 | (8'hb1)) : reg3396[(1'h0):(1'h0)])));
                      reg3396 <= $unsigned({$unsigned(forvar3402[(2'h3):(2'h2)])});
                      reg3397 <= (^~$signed($unsigned((&(8'hb6)))));
                      reg3398 <= $unsigned((reg3390[(1'h1):(1'h0)] ?
                          ((reg3390 ?
                              reg3382 : forvar3387) != {reg3409}) : (forvar3378[(4'hc):(2'h2)] ?
                              $signed(reg3408) : (!forvar3387))));
                    end
                  for (forvar3399 = (1'h0); (forvar3399 < (1'h0)); forvar3399 = (forvar3399 + (1'h1)))
                    begin
                      reg3400 <= reg3394[(4'hd):(4'hd)];
                    end
                end
            end
        end
      reg3412 <= ($unsigned((|((8'h9f) >> reg3399))) ?
          wire3374 : {$signed((reg3386 ? wire3375 : (8'hb8)))});
      reg3413 <= $unsigned(({reg3386} ?
          $signed((forvar3377 ? (8'hb8) : reg3394)) : (wire3371 < reg3406)));
    end
  assign wire3414 = (8'h9f);
  assign wire3415 = (~^reg3403);
  module3416 modinst3438 (wire3437, clk, forvar3398, reg3398, wire3375, reg3399, wire3370);
  always
    @(posedge clk) begin
      reg3439 <= $unsigned(($unsigned($unsigned(forvar3395)) ?
          $unsigned($signed(reg3388)) : reg3407));
      for (forvar3440 = (1'h0); (forvar3440 < (2'h3)); forvar3440 = (forvar3440 + (1'h1)))
        begin
          for (forvar3441 = (1'h0); (forvar3441 < (2'h2)); forvar3441 = (forvar3441 + (1'h1)))
            begin
              for (forvar3442 = (1'h0); (forvar3442 < (1'h1)); forvar3442 = (forvar3442 + (1'h1)))
                begin
                  for (forvar3443 = (1'h0); (forvar3443 < (2'h2)); forvar3443 = (forvar3443 + (1'h1)))
                    begin
                      reg3444 <= (reg3395 <<< forvar3396);
                      reg3445 <= wire3415[(4'hd):(1'h0)];
                    end
                  for (forvar3446 = (1'h0); (forvar3446 < (2'h3)); forvar3446 = (forvar3446 + (1'h1)))
                    begin
                      reg3447 <= {forvar3405};
                    end
                  for (forvar3448 = (1'h0); (forvar3448 < (2'h3)); forvar3448 = (forvar3448 + (1'h1)))
                    begin
                      reg3449 <= reg3390;
                      reg3450 <= $signed($unsigned($signed((reg3445 <= forvar3440))));
                      reg3451 <= $unsigned(reg3391[(1'h0):(1'h0)]);
                      reg3452 <= ((reg3386 ?
                          $signed((reg3398 && forvar3386)) : $unsigned(forvar3393)) << forvar3378);
                    end
                end
            end
          reg3453 <= reg3399;
        end
      if ((8'h9d))
        begin
          for (forvar3454 = (1'h0); (forvar3454 < (2'h3)); forvar3454 = (forvar3454 + (1'h1)))
            begin
              for (forvar3455 = (1'h0); (forvar3455 < (2'h2)); forvar3455 = (forvar3455 + (1'h1)))
                begin
                  for (forvar3456 = (1'h0); (forvar3456 < (2'h3)); forvar3456 = (forvar3456 + (1'h1)))
                    begin
                      reg3457 <= (&reg3394);
                    end
                  for (forvar3458 = (1'h0); (forvar3458 < (1'h0)); forvar3458 = (forvar3458 + (1'h1)))
                    begin
                      reg3459 <= reg3408;
                    end
                end
              if ($signed(forvar3387[(1'h0):(1'h0)]))
                begin
                  reg3460 <= reg3389[(1'h1):(1'h0)];
                  if (reg3450[(1'h1):(1'h1)])
                    begin
                      reg3461 <= {reg3407[(4'ha):(3'h7)]};
                      reg3462 <= $signed((!$unsigned((~(8'hb8)))));
                      reg3463 <= $signed(wire3369[(4'h9):(3'h7)]);
                    end
                  else
                    begin
                      reg3461 <= reg3403;
                    end
                  if (reg3393)
                    begin
                      reg3464 <= reg3447[(4'h8):(1'h1)];
                      reg3465 <= $signed((($unsigned(reg3397) ?
                          reg3464[(1'h1):(1'h0)] : $signed(reg3444)) ^~ $unsigned((reg3404 | reg3452))));
                      reg3466 <= ($unsigned(($signed(forvar3386) ?
                              (reg3409 >>> forvar3402) : reg3380[(2'h3):(1'h0)])) ?
                          (~|((forvar3378 ^ (8'hb9)) > reg3450[(2'h2):(1'h0)])) : (reg3410[(2'h3):(2'h2)] ?
                              ($signed(reg3445) - (+forvar3396)) : reg3465[(3'h4):(1'h0)]));
                      reg3467 <= reg3395[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3464 <= reg3408[(3'h4):(2'h3)];
                      reg3465 <= ({($signed(forvar3455) >>> $unsigned(reg3462))} ?
                          ((~|(reg3399 ? reg3395 : wire3369)) ?
                              reg3388 : $signed($unsigned(reg3466))) : forvar3402);
                      reg3466 <= reg3451;
                      reg3467 <= $signed((-((reg3463 ?
                          reg3391 : forvar3386) ~^ $unsigned(forvar3456))));
                    end
                end
              else
                begin
                  reg3460 <= {wire3370};
                  if ({({{reg3387}} ?
                          ((8'ha2) == (forvar3440 * reg3394)) : reg3461)})
                    begin
                      reg3461 <= (forvar3456 | ($unsigned((reg3451 ?
                          wire3370 : reg3390)) ~^ ((reg3384 | forvar3377) << (reg3447 ?
                          forvar3454 : reg3412))));
                      reg3462 <= reg3377;
                      reg3463 <= reg3467;
                      reg3464 <= reg3459;
                    end
                  else
                    begin
                      reg3461 <= (({forvar3442} ?
                              forvar3386[(4'hd):(4'hb)] : {(reg3449 < forvar3398)}) ?
                          ({{forvar3458}} ?
                              $signed($unsigned(reg3450)) : {(forvar3378 >>> reg3464)}) : forvar3441);
                      reg3462 <= $unsigned((~{forvar3399}));
                    end
                  for (forvar3465 = (1'h0); (forvar3465 < (2'h2)); forvar3465 = (forvar3465 + (1'h1)))
                    begin
                      reg3466 <= (!reg3385);
                      reg3467 <= (reg3403 != {$unsigned({(8'ha4)})});
                      reg3468 <= reg3408[(1'h1):(1'h1)];
                    end
                  reg3469 <= (~($signed($unsigned(reg3465)) ?
                      (reg3381[(3'h7):(3'h4)] <= $unsigned(forvar3393)) : reg3410));
                end
              if ((reg3449 ? (^~$unsigned(forvar3454)) : wire3373))
                begin
                  if ($unsigned((forvar3377[(3'h5):(1'h1)] ?
                      forvar3441[(3'h7):(1'h0)] : $signed((wire3368 ?
                          (8'ha3) : forvar3388)))))
                    begin
                      reg3470 <= (8'ha5);
                      reg3471 <= {{reg3404[(3'h4):(2'h2)]}};
                      reg3472 <= $signed((!{(^~wire3368)}));
                      reg3473 <= $unsigned(($signed((reg3464 | wire3437)) ?
                          {{forvar3465}} : reg3453));
                    end
                  else
                    begin
                      reg3470 <= forvar3376;
                      reg3471 <= (8'ha8);
                      reg3472 <= $signed($unsigned($unsigned({reg3412})));
                    end
                  if (reg3463)
                    begin
                      reg3474 <= (8'hb0);
                      reg3475 <= $signed(reg3445);
                    end
                  else
                    begin
                      reg3474 <= {forvar3442[(2'h2):(1'h0)]};
                    end
                  for (forvar3476 = (1'h0); (forvar3476 < (2'h2)); forvar3476 = (forvar3476 + (1'h1)))
                    begin
                      reg3477 <= {$unsigned($unsigned(wire3373[(1'h0):(1'h0)]))};
                      reg3478 <= (8'ha8);
                      reg3479 <= ((($signed(wire3414) == (forvar3395 < forvar3388)) << $signed((~&reg3400))) && wire3370);
                    end
                end
              else
                begin
                  if (reg3462[(1'h1):(1'h0)])
                    begin
                      reg3470 <= reg3467;
                      reg3471 <= (|reg3475);
                    end
                  else
                    begin
                      reg3470 <= reg3471;
                      reg3471 <= (^~reg3399);
                      reg3472 <= forvar3476[(2'h3):(2'h3)];
                      reg3473 <= (reg3479[(3'h4):(1'h0)] ^ forvar3393);
                    end
                  if (reg3404[(1'h1):(1'h0)])
                    begin
                      reg3474 <= reg3471[(3'h4):(2'h2)];
                      reg3475 <= (forvar3442[(1'h1):(1'h0)] << $signed($signed($unsigned(reg3450))));
                      reg3476 <= (reg3394[(4'hc):(4'ha)] != $signed(reg3398));
                    end
                  else
                    begin
                      reg3474 <= (~|reg3382);
                      reg3475 <= ({($signed((8'had)) ?
                                  reg3471 : $unsigned(forvar3458))} ?
                          reg3476[(4'ha):(4'ha)] : reg3457);
                      reg3476 <= reg3468[(4'ha):(3'h5)];
                    end
                end
              for (forvar3480 = (1'h0); (forvar3480 < (1'h0)); forvar3480 = (forvar3480 + (1'h1)))
                begin
                  reg3481 <= ($unsigned((&(reg3397 ? reg3473 : (8'hb6)))) ?
                      ((reg3462[(1'h1):(1'h0)] == {reg3445}) ?
                          {(^~(8'h9c))} : $signed((forvar3440 + forvar3402))) : ($signed($signed(reg3407)) <= ($unsigned(wire3415) >= $signed(reg3464))));
                end
            end
        end
      else
        begin
          for (forvar3454 = (1'h0); (forvar3454 < (1'h1)); forvar3454 = (forvar3454 + (1'h1)))
            begin
              for (forvar3455 = (1'h0); (forvar3455 < (1'h1)); forvar3455 = (forvar3455 + (1'h1)))
                begin
                  if (reg3478[(1'h0):(1'h0)])
                    begin
                      reg3456 <= ({((reg3399 ~^ forvar3376) ?
                              ((8'h9e) >= wire3437) : $unsigned((8'ha2)))} >> $unsigned((!$unsigned((8'h9c)))));
                      reg3457 <= reg3453;
                      reg3458 <= reg3481[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3456 <= (~&(~^{wire3368}));
                    end
                  reg3459 <= $unsigned($unsigned($signed((reg3410 > forvar3398))));
                  if (reg3400)
                    begin
                      reg3460 <= ((8'hab) ^ (((wire3371 != (8'hac)) ?
                          (+(8'h9c)) : reg3395[(4'h8):(3'h4)]) ^ (~^wire3368[(4'h8):(3'h4)])));
                      reg3461 <= $unsigned((&(reg3379 <<< (reg3379 ?
                          reg3389 : reg3475))));
                      reg3462 <= $unsigned(reg3386[(2'h3):(2'h2)]);
                      reg3463 <= forvar3476;
                    end
                  else
                    begin
                      reg3460 <= $unsigned((~&($signed(reg3456) ?
                          (wire3368 ? forvar3376 : (8'h9e)) : (^forvar3442))));
                      reg3461 <= $unsigned(forvar3476[(1'h1):(1'h1)]);
                      reg3462 <= {($unsigned((~&reg3444)) == (((8'hb4) > (8'haa)) ~^ $signed(wire3414)))};
                      reg3463 <= $unsigned(($signed(reg3462[(1'h0):(1'h0)]) > ($signed(reg3477) ?
                          wire3368[(1'h0):(1'h0)] : wire3368)));
                    end
                end
              for (forvar3464 = (1'h0); (forvar3464 < (1'h0)); forvar3464 = (forvar3464 + (1'h1)))
                begin
                  if ($signed(($signed($unsigned(reg3389)) < ((&(8'ha4)) ?
                      (forvar3378 ? reg3400 : reg3384) : reg3479))))
                    begin
                      reg3465 <= (8'h9d);
                      reg3466 <= $signed((((reg3409 == (8'h9f)) ?
                          {reg3468} : $signed((8'ha0))) >= wire3370));
                      reg3467 <= reg3388;
                      reg3468 <= $unsigned((reg3386 >= $signed({reg3453})));
                    end
                  else
                    begin
                      reg3465 <= wire3415;
                      reg3466 <= $unsigned(reg3397);
                      reg3467 <= ((~&(+(reg3456 ?
                          (8'ha8) : reg3409))) << {(-(reg3393 << reg3410))});
                    end
                  for (forvar3469 = (1'h0); (forvar3469 < (2'h2)); forvar3469 = (forvar3469 + (1'h1)))
                    begin
                      reg3470 <= reg3476[(3'h6):(3'h6)];
                    end
                  if ((&$unsigned(reg3388[(4'he):(3'h7)])))
                    begin
                      reg3471 <= {(((forvar3405 || forvar3465) ?
                                  (reg3481 + reg3469) : $unsigned((8'haf))) ?
                              ($signed(reg3456) & $unsigned(reg3466)) : forvar3464[(2'h2):(1'h0)])};
                      reg3472 <= forvar3386[(4'ha):(4'h9)];
                    end
                  else
                    begin
                      reg3471 <= $signed($unsigned($unsigned((&(8'h9e)))));
                      reg3472 <= (($signed($unsigned(wire3370)) == {(~^(8'ha4))}) ?
                          (8'hb1) : $unsigned(reg3450[(2'h2):(1'h1)]));
                      reg3473 <= reg3451[(2'h2):(1'h1)];
                    end
                end
              if ($signed($unsigned(((reg3468 & forvar3387) ?
                  $signed(reg3466) : $unsigned(forvar3393)))))
                begin
                  if (reg3391[(1'h1):(1'h0)])
                    begin
                      reg3474 <= reg3396[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg3474 <= reg3399;
                      reg3475 <= reg3467[(1'h1):(1'h0)];
                      reg3476 <= reg3395[(3'h7):(3'h6)];
                    end
                  if (wire3415[(3'h6):(1'h0)])
                    begin
                      reg3477 <= {(8'ha9)};
                    end
                  else
                    begin
                      reg3477 <= {$signed((reg3457[(2'h3):(2'h3)] ~^ reg3459))};
                      reg3478 <= $signed(((-$unsigned((8'h9c))) ?
                          (reg3408 << (forvar3454 ?
                              reg3385 : reg3478)) : $signed(reg3413[(1'h0):(1'h0)])));
                      reg3479 <= $unsigned((~^$signed({reg3386})));
                      reg3480 <= $signed($unsigned(reg3450[(1'h0):(1'h0)]));
                    end
                  for (forvar3481 = (1'h0); (forvar3481 < (2'h2)); forvar3481 = (forvar3481 + (1'h1)))
                    begin
                      reg3482 <= (-$unsigned($unsigned($signed(wire3415))));
                      reg3483 <= wire3370[(1'h0):(1'h0)];
                      reg3484 <= (forvar3448 ?
                          (reg3380 ?
                              $signed((8'hba)) : (~&{forvar3454})) : $unsigned(forvar3402));
                    end
                  for (forvar3485 = (1'h0); (forvar3485 < (1'h0)); forvar3485 = (forvar3485 + (1'h1)))
                    begin
                      reg3486 <= ({$signed(wire3375)} ?
                          (forvar3464[(3'h4):(2'h2)] ?
                              (8'hb6) : reg3410[(2'h2):(1'h1)]) : ($unsigned($signed(reg3470)) ^~ ((+forvar3396) & (reg3476 ?
                              reg3460 : forvar3476))));
                      reg3487 <= (8'hb6);
                    end
                end
              else
                begin
                  for (forvar3474 = (1'h0); (forvar3474 < (2'h2)); forvar3474 = (forvar3474 + (1'h1)))
                    begin
                      reg3475 <= forvar3441;
                      reg3476 <= (-(8'hb4));
                      reg3477 <= ($signed((!(^reg3439))) == forvar3458[(4'hd):(3'h5)]);
                    end
                  for (forvar3478 = (1'h0); (forvar3478 < (1'h1)); forvar3478 = (forvar3478 + (1'h1)))
                    begin
                      reg3479 <= $signed(forvar3448[(1'h1):(1'h1)]);
                    end
                  for (forvar3480 = (1'h0); (forvar3480 < (1'h0)); forvar3480 = (forvar3480 + (1'h1)))
                    begin
                      reg3481 <= (|$unsigned($unsigned($signed(reg3453))));
                    end
                  if ($unsigned((+$unsigned((~|reg3472)))))
                    begin
                      reg3482 <= $unsigned(reg3477);
                      reg3483 <= reg3377[(4'hc):(4'h8)];
                      reg3484 <= reg3382[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg3482 <= forvar3485;
                      reg3483 <= ((((&reg3404) && $signed((8'hb1))) ?
                              reg3470 : ((^wire3371) ?
                                  reg3475[(4'h8):(3'h6)] : (forvar3393 == reg3379))) ?
                          wire3372[(2'h2):(1'h1)] : (reg3457 ?
                              $unsigned(reg3458) : reg3482));
                      reg3484 <= ({(&reg3393)} >>> wire3375[(4'hb):(4'hb)]);
                      reg3485 <= $signed($unsigned(($signed(reg3477) ^ $unsigned(forvar3399))));
                    end
                end
            end
          if ({(!(^(^~reg3473)))})
            begin
              for (forvar3488 = (1'h0); (forvar3488 < (2'h2)); forvar3488 = (forvar3488 + (1'h1)))
                begin
                  reg3489 <= {(reg3404[(2'h3):(1'h1)] <= $unsigned(reg3469[(1'h0):(1'h0)]))};
                  for (forvar3490 = (1'h0); (forvar3490 < (1'h1)); forvar3490 = (forvar3490 + (1'h1)))
                    begin
                      reg3491 <= (($unsigned($unsigned(reg3445)) >> reg3384) <<< ((^$signed(reg3407)) & (^~((8'had) + reg3407))));
                      reg3492 <= $signed({((forvar3399 ? reg3384 : forvar3490) ?
                              (^~reg3400) : (forvar3387 && forvar3480))});
                      reg3493 <= {(((reg3411 || reg3466) ?
                              (forvar3377 >= reg3483) : (8'h9f)) <= (~|((8'hb4) ?
                              reg3449 : reg3404)))};
                    end
                  reg3494 <= (reg3404[(1'h1):(1'h0)] == (&({forvar3481} << $unsigned(forvar3481))));
                  for (forvar3495 = (1'h0); (forvar3495 < (1'h1)); forvar3495 = (forvar3495 + (1'h1)))
                    begin
                      reg3496 <= (8'hac);
                      reg3497 <= forvar3485[(3'h4):(1'h0)];
                    end
                end
              for (forvar3498 = (1'h0); (forvar3498 < (2'h2)); forvar3498 = (forvar3498 + (1'h1)))
                begin
                  for (forvar3499 = (1'h0); (forvar3499 < (2'h2)); forvar3499 = (forvar3499 + (1'h1)))
                    begin
                      reg3500 <= (({((8'ha4) ? (8'hba) : wire3371)} ?
                              {(8'had)} : reg3461[(1'h0):(1'h0)]) ?
                          (!reg3404[(1'h1):(1'h1)]) : ($unsigned({reg3452}) ?
                              forvar3377 : reg3493[(1'h1):(1'h1)]));
                      reg3501 <= reg3465[(1'h1):(1'h0)];
                    end
                  reg3502 <= $unsigned($unsigned($signed($unsigned(wire3371))));
                end
              if ((&(~^(~^$unsigned(reg3462)))))
                begin
                  for (forvar3503 = (1'h0); (forvar3503 < (2'h3)); forvar3503 = (forvar3503 + (1'h1)))
                    begin
                      reg3504 <= $unsigned(((^((8'h9d) <= reg3496)) ?
                          $unsigned($signed(wire3374)) : $unsigned($signed(reg3493))));
                      reg3505 <= (forvar3478 ?
                          ((forvar3485 ?
                              $signed((8'haf)) : $signed(reg3388)) + forvar3443[(4'h8):(1'h1)]) : (^~(|$signed(reg3485))));
                    end
                  reg3506 <= ((~^$unsigned(wire3437)) ?
                      (-(~$signed((8'hb1)))) : (8'ha6));
                end
              else
                begin
                  if ((reg3385[(1'h1):(1'h0)] == wire3374[(3'h5):(1'h1)]))
                    begin
                      reg3503 <= {(reg3506 && (8'ha6))};
                      reg3504 <= reg3469;
                      reg3505 <= forvar3387[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg3503 <= (wire3369 ? reg3394[(1'h0):(1'h0)] : (8'h9e));
                      reg3504 <= {forvar3395[(4'h8):(1'h1)]};
                      reg3505 <= (8'hb3);
                    end
                  for (forvar3506 = (1'h0); (forvar3506 < (1'h1)); forvar3506 = (forvar3506 + (1'h1)))
                    begin
                      reg3507 <= $unsigned((+reg3439));
                    end
                end
            end
          else
            begin
              if (forvar3386)
                begin
                  reg3488 <= (8'ha2);
                end
              else
                begin
                  for (forvar3488 = (1'h0); (forvar3488 < (1'h0)); forvar3488 = (forvar3488 + (1'h1)))
                    begin
                      reg3489 <= reg3450[(2'h2):(1'h1)];
                      reg3490 <= ($unsigned(($signed(forvar3469) ?
                              ((8'h9c) ? reg3388 : (8'ha5)) : (!forvar3399))) ?
                          reg3386[(2'h2):(1'h0)] : (reg3467 <= ((8'ha5) ?
                              $signed((8'ha6)) : $unsigned(reg3487))));
                    end
                end
              if ((~&($signed($unsigned(reg3467)) ?
                  (8'h9f) : {$signed(forvar3485)})))
                begin
                  for (forvar3491 = (1'h0); (forvar3491 < (2'h2)); forvar3491 = (forvar3491 + (1'h1)))
                    begin
                      reg3492 <= $signed((reg3377 ?
                          ((~|reg3457) - $signed(reg3480)) : ((reg3388 << forvar3499) ?
                              forvar3396 : {reg3384})));
                      reg3493 <= $unsigned(reg3483);
                      reg3494 <= reg3475;
                    end
                  reg3495 <= reg3382[(3'h5):(3'h5)];
                  if (((({forvar3440} ? $signed((8'haf)) : $signed((8'hb0))) ?
                      wire3375[(4'h9):(3'h4)] : (8'ha9)) ^~ reg3465))
                    begin
                      reg3496 <= $signed($unsigned($signed(reg3379[(4'hb):(3'h4)])));
                      reg3497 <= $signed(reg3480);
                      reg3498 <= reg3407;
                      reg3499 <= reg3380[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg3496 <= {$unsigned(reg3445)};
                      reg3497 <= $signed((~&forvar3481[(3'h4):(2'h2)]));
                      reg3498 <= reg3401;
                      reg3499 <= (!reg3490[(1'h0):(1'h0)]);
                    end
                  for (forvar3500 = (1'h0); (forvar3500 < (2'h3)); forvar3500 = (forvar3500 + (1'h1)))
                    begin
                      reg3501 <= reg3476[(2'h2):(1'h1)];
                      reg3502 <= (reg3396[(3'h5):(3'h4)] <= (reg3385 ?
                          ((8'ha4) ?
                              reg3382 : (reg3384 ?
                                  reg3458 : (8'hb8))) : (|forvar3485)));
                    end
                end
              else
                begin
                  for (forvar3491 = (1'h0); (forvar3491 < (1'h1)); forvar3491 = (forvar3491 + (1'h1)))
                    begin
                      reg3492 <= $signed({reg3495[(3'h4):(1'h0)]});
                      reg3493 <= $signed(reg3461);
                      reg3494 <= ($unsigned(reg3481[(1'h1):(1'h1)]) ?
                          $unsigned($unsigned((8'hb0))) : ((8'hab) >>> {$signed(forvar3469)}));
                      reg3495 <= reg3459[(4'he):(3'h5)];
                    end
                  for (forvar3496 = (1'h0); (forvar3496 < (2'h2)); forvar3496 = (forvar3496 + (1'h1)))
                    begin
                      reg3497 <= reg3479;
                      reg3498 <= $signed($unsigned((~(reg3493 ?
                          reg3396 : forvar3448))));
                      reg3499 <= $unsigned(($unsigned(reg3495[(2'h2):(2'h2)]) && reg3473));
                    end
                end
              for (forvar3503 = (1'h0); (forvar3503 < (1'h1)); forvar3503 = (forvar3503 + (1'h1)))
                begin
                  if ((8'hb9))
                    begin
                      reg3504 <= (+(^~$signed((reg3399 ?
                          reg3452 : forvar3503))));
                    end
                  else
                    begin
                      reg3504 <= forvar3464[(2'h2):(1'h1)];
                      reg3505 <= $unsigned((8'hb2));
                      reg3506 <= (-((~|(8'h9d)) <<< $unsigned((reg3452 ?
                          reg3391 : forvar3500))));
                      reg3507 <= (($signed($signed(reg3445)) ?
                              ((reg3394 ? reg3483 : reg3445) ?
                                  $unsigned(reg3447) : forvar3386[(4'hb):(4'h8)]) : forvar3378) ?
                          ($unsigned($signed(forvar3441)) ~^ (8'hb6)) : (&reg3482[(1'h0):(1'h0)]));
                    end
                  for (forvar3508 = (1'h0); (forvar3508 < (1'h0)); forvar3508 = (forvar3508 + (1'h1)))
                    begin
                      reg3509 <= reg3506[(4'hb):(1'h0)];
                    end
                end
            end
          for (forvar3510 = (1'h0); (forvar3510 < (1'h1)); forvar3510 = (forvar3510 + (1'h1)))
            begin
              if ((~|({(reg3495 ? reg3451 : forvar3402)} ?
                  {reg3497} : $unsigned((-reg3480)))))
                begin
                  for (forvar3511 = (1'h0); (forvar3511 < (1'h1)); forvar3511 = (forvar3511 + (1'h1)))
                    begin
                      reg3512 <= (~^(~(^forvar3441)));
                    end
                end
              else
                begin
                  if (reg3399)
                    begin
                      reg3511 <= ($signed(((reg3507 + forvar3405) + (~&reg3494))) == forvar3478);
                      reg3512 <= reg3491[(2'h3):(2'h2)];
                      reg3513 <= wire3369[(3'h7):(3'h5)];
                      reg3514 <= reg3380;
                    end
                  else
                    begin
                      reg3511 <= (^reg3408[(3'h5):(2'h2)]);
                      reg3512 <= (8'hb4);
                    end
                  for (forvar3515 = (1'h0); (forvar3515 < (1'h1)); forvar3515 = (forvar3515 + (1'h1)))
                    begin
                      reg3516 <= forvar3440;
                    end
                  if ((+$unsigned(reg3494)))
                    begin
                      reg3517 <= (reg3468 << (-{(reg3452 ?
                              reg3468 : reg3394)}));
                    end
                  else
                    begin
                      reg3517 <= reg3502;
                    end
                  for (forvar3518 = (1'h0); (forvar3518 < (1'h0)); forvar3518 = (forvar3518 + (1'h1)))
                    begin
                      reg3519 <= ((forvar3496[(4'ha):(2'h3)] ^~ (!reg3401[(1'h1):(1'h1)])) ?
                          (((reg3497 ? reg3390 : forvar3500) || (reg3386 ?
                              reg3397 : (8'haa))) + ((~^reg3380) || $unsigned(wire3374))) : ((~^(reg3400 ~^ reg3479)) <<< reg3502));
                      reg3520 <= ($unsigned(reg3381[(4'h8):(3'h6)]) - ({{forvar3511}} ?
                          (~reg3499[(2'h3):(2'h2)]) : $signed((forvar3388 ?
                              reg3400 : reg3487))));
                    end
                end
              for (forvar3521 = (1'h0); (forvar3521 < (2'h3)); forvar3521 = (forvar3521 + (1'h1)))
                begin
                  for (forvar3522 = (1'h0); (forvar3522 < (2'h2)); forvar3522 = (forvar3522 + (1'h1)))
                    begin
                      reg3523 <= ($unsigned(forvar3508) <<< (|reg3411));
                    end
                  for (forvar3524 = (1'h0); (forvar3524 < (1'h0)); forvar3524 = (forvar3524 + (1'h1)))
                    begin
                      reg3525 <= forvar3465[(4'h8):(2'h3)];
                      reg3526 <= {(reg3458 | $signed((^~reg3507)))};
                      reg3527 <= (($signed((8'ha7)) << $unsigned($unsigned(reg3466))) >> ({((8'hba) << forvar3454)} <<< (reg3445[(4'hd):(2'h3)] * $unsigned((8'hba)))));
                      reg3528 <= {forvar3488[(2'h3):(2'h3)]};
                    end
                  reg3529 <= $unsigned($signed(reg3494));
                end
              for (forvar3530 = (1'h0); (forvar3530 < (2'h2)); forvar3530 = (forvar3530 + (1'h1)))
                begin
                  if ((-((~^$unsigned(forvar3530)) ?
                      ((reg3457 ? (8'hb3) : forvar3443) ?
                          $signed(reg3382) : {reg3474}) : forvar3498)))
                    begin
                      reg3531 <= {{forvar3443}};
                      reg3532 <= (((forvar3442[(2'h2):(2'h2)] ?
                          $unsigned(reg3493) : (+(8'hb4))) || $signed((!(8'h9e)))) * forvar3498[(4'hc):(3'h5)]);
                    end
                  else
                    begin
                      reg3531 <= reg3527[(2'h2):(1'h0)];
                    end
                end
              for (forvar3533 = (1'h0); (forvar3533 < (2'h3)); forvar3533 = (forvar3533 + (1'h1)))
                begin
                  reg3534 <= $unsigned(($signed({reg3469}) ?
                      ((8'hb0) ?
                          wire3437 : (reg3464 ?
                              reg3465 : reg3465)) : (forvar3398[(4'hd):(4'h9)] || reg3439[(2'h2):(2'h2)])));
                  if ((!$unsigned($signed($signed(reg3472)))))
                    begin
                      reg3535 <= (^(forvar3476 ~^ $unsigned(wire3371)));
                      reg3536 <= (forvar3443[(1'h0):(1'h0)] ?
                          $signed($unsigned(reg3489[(2'h3):(2'h3)])) : $unsigned($unsigned((reg3452 ?
                              reg3382 : reg3452))));
                      reg3537 <= (($signed(forvar3395) - $unsigned((8'hb1))) ?
                          (((reg3397 > forvar3399) ?
                                  (reg3532 <= forvar3500) : {reg3461}) ?
                              {$unsigned((8'ha2))} : reg3488) : reg3393);
                      reg3538 <= $signed(reg3534);
                    end
                  else
                    begin
                      reg3535 <= reg3516[(1'h1):(1'h1)];
                      reg3536 <= reg3496;
                    end
                  reg3539 <= reg3465;
                  if (({(reg3511[(3'h7):(3'h4)] <<< (reg3381 | reg3470))} ?
                      reg3395 : (forvar3377[(1'h0):(1'h0)] >>> reg3472[(2'h2):(1'h0)])))
                    begin
                      reg3540 <= $signed($signed((8'hba)));
                    end
                  else
                    begin
                      reg3540 <= (($signed($unsigned(reg3461)) & wire3371[(2'h2):(1'h1)]) && $unsigned(($unsigned(reg3377) ?
                          forvar3488 : $unsigned(wire3371))));
                      reg3541 <= ((~^$signed((forvar3476 * (8'ha3)))) ?
                          reg3517 : (forvar3395 << {((8'hb4) ?
                                  forvar3469 : wire3368)}));
                      reg3542 <= reg3470[(2'h3):(1'h1)];
                      reg3543 <= reg3501;
                    end
                end
            end
          reg3544 <= {$signed(((8'ha2) ?
                  (forvar3490 ? reg3456 : reg3529) : $unsigned((8'hb8))))};
        end
      for (forvar3545 = (1'h0); (forvar3545 < (1'h1)); forvar3545 = (forvar3545 + (1'h1)))
        begin
          reg3546 <= forvar3393;
        end
    end
  always
    @(posedge clk) begin
      if ($signed((~&$unsigned($signed(reg3490)))))
        begin
          if ($signed(reg3469))
            begin
              reg3547 <= (-{($signed((8'hac)) ?
                      reg3462[(1'h0):(1'h0)] : (!reg3507))});
              for (forvar3548 = (1'h0); (forvar3548 < (2'h3)); forvar3548 = (forvar3548 + (1'h1)))
                begin
                  reg3549 <= forvar3454;
                  for (forvar3550 = (1'h0); (forvar3550 < (1'h1)); forvar3550 = (forvar3550 + (1'h1)))
                    begin
                      reg3551 <= (((reg3480[(3'h4):(1'h1)] < reg3473) ^ (forvar3498 ?
                          $signed(reg3403) : (&reg3491))) <<< forvar3377[(3'h7):(2'h2)]);
                    end
                  for (forvar3552 = (1'h0); (forvar3552 < (1'h0)); forvar3552 = (forvar3552 + (1'h1)))
                    begin
                      reg3553 <= $unsigned({(!(-reg3449))});
                      reg3554 <= ((~$signed($signed((8'hac)))) >= forvar3548);
                      reg3555 <= $signed(forvar3455[(2'h3):(1'h0)]);
                      reg3556 <= {(~{$signed(forvar3524)})};
                    end
                end
              reg3557 <= reg3516;
              reg3558 <= $unsigned({reg3444[(1'h1):(1'h1)]});
            end
          else
            begin
              for (forvar3547 = (1'h0); (forvar3547 < (2'h3)); forvar3547 = (forvar3547 + (1'h1)))
                begin
                  if ({(($signed(reg3499) && forvar3398) ?
                          $signed((forvar3398 ~^ forvar3508)) : (forvar3474 > (reg3388 != (8'hb2))))})
                    begin
                      reg3548 <= $signed(({{wire3369}} > ((8'hb7) ^ (reg3384 | reg3516))));
                      reg3549 <= forvar3383[(4'h8):(4'h8)];
                    end
                  else
                    begin
                      reg3548 <= (^~$unsigned((~&{forvar3441})));
                      reg3549 <= (|(8'ha0));
                      reg3550 <= forvar3440[(3'h6):(2'h2)];
                    end
                  for (forvar3551 = (1'h0); (forvar3551 < (2'h2)); forvar3551 = (forvar3551 + (1'h1)))
                    begin
                      reg3552 <= reg3404;
                      reg3553 <= reg3499[(3'h4):(3'h4)];
                      reg3554 <= (((~^reg3502[(1'h1):(1'h0)]) ?
                          (8'hb8) : forvar3448) << (8'hb1));
                      reg3555 <= ({$unsigned((^forvar3405))} == $signed((-reg3463[(1'h1):(1'h1)])));
                    end
                end
              reg3556 <= ($signed(forvar3481[(3'h6):(3'h5)]) || reg3516);
              reg3557 <= (((reg3534[(1'h1):(1'h1)] ?
                      (~^reg3457) : reg3491[(3'h6):(3'h4)]) ?
                  $unsigned(reg3502) : $signed($signed(reg3476))) || {reg3476[(3'h6):(3'h6)]});
              if (((reg3535 ?
                  $signed((reg3557 <= reg3404)) : forvar3499[(4'hd):(4'hc)]) >>> ($signed(forvar3498) ?
                  reg3538[(4'ha):(3'h5)] : (reg3555[(3'h4):(1'h1)] ?
                      reg3547[(4'h8):(1'h0)] : forvar3478))))
                begin
                  reg3558 <= forvar3440[(2'h2):(1'h1)];
                  for (forvar3559 = (1'h0); (forvar3559 < (2'h3)); forvar3559 = (forvar3559 + (1'h1)))
                    begin
                      reg3560 <= $signed($signed(reg3543[(1'h1):(1'h1)]));
                      reg3561 <= (reg3460 & $signed($signed({reg3400})));
                      reg3562 <= $signed(reg3385);
                    end
                  for (forvar3563 = (1'h0); (forvar3563 < (2'h3)); forvar3563 = (forvar3563 + (1'h1)))
                    begin
                      reg3564 <= $signed((~|$signed((~|reg3481))));
                      reg3565 <= forvar3498;
                      reg3566 <= {(8'haf)};
                    end
                end
              else
                begin
                  for (forvar3558 = (1'h0); (forvar3558 < (1'h1)); forvar3558 = (forvar3558 + (1'h1)))
                    begin
                      reg3559 <= $unsigned($signed((8'hae)));
                      reg3560 <= reg3495;
                    end
                end
            end
          for (forvar3567 = (1'h0); (forvar3567 < (2'h3)); forvar3567 = (forvar3567 + (1'h1)))
            begin
              if (((^forvar3469) & wire3374))
                begin
                  for (forvar3568 = (1'h0); (forvar3568 < (1'h0)); forvar3568 = (forvar3568 + (1'h1)))
                    begin
                      reg3569 <= $signed(reg3527[(3'h6):(2'h3)]);
                      reg3570 <= $signed($unsigned(forvar3386[(1'h0):(1'h0)]));
                      reg3571 <= $unsigned((((reg3560 - reg3517) < forvar3469[(2'h3):(1'h1)]) <<< $unsigned($unsigned((8'ha5)))));
                      reg3572 <= (((8'ha4) ?
                          $signed((reg3494 | forvar3476)) : (+reg3390[(1'h0):(1'h0)])) >> ((^$unsigned(reg3450)) ?
                          forvar3480[(4'h9):(4'h8)] : (&(reg3491 ?
                              forvar3398 : reg3479))));
                    end
                  reg3573 <= reg3535[(4'h9):(3'h6)];
                  if (($unsigned((reg3516 ^~ (8'ha0))) ~^ (~&(&$signed(forvar3567)))))
                    begin
                      reg3574 <= (+{(forvar3455[(3'h6):(1'h0)] ^ reg3556[(3'h5):(3'h4)])});
                    end
                  else
                    begin
                      reg3574 <= $signed(reg3451);
                      reg3575 <= reg3562;
                    end
                end
              else
                begin
                  if ($unsigned((~&($unsigned(reg3406) ?
                      $unsigned(reg3377) : {(8'haa)}))))
                    begin
                      reg3568 <= (&(~&($unsigned(reg3483) ?
                          (reg3507 ?
                              forvar3464 : reg3548) : $unsigned(reg3401))));
                      reg3569 <= {(8'hb1)};
                      reg3570 <= ((reg3503 ?
                              (reg3385[(1'h1):(1'h0)] ?
                                  reg3458[(2'h2):(2'h2)] : (forvar3511 ^ forvar3563)) : (|(wire3414 ^ reg3553))) ?
                          $signed($signed($signed(reg3447))) : (reg3390[(2'h2):(1'h1)] ?
                              {$unsigned(reg3465)} : ((forvar3495 >>> reg3408) ?
                                  (reg3486 ?
                                      reg3552 : (8'ha1)) : {forvar3481})));
                      reg3571 <= ($unsigned($signed(forvar3480[(1'h0):(1'h0)])) >= $signed($signed((~|reg3385))));
                    end
                  else
                    begin
                      reg3568 <= (^($unsigned((reg3554 ? wire3437 : reg3478)) ?
                          $signed((^~reg3575)) : (~(~|wire3371))));
                      reg3569 <= (8'hb7);
                    end
                  for (forvar3572 = (1'h0); (forvar3572 < (1'h1)); forvar3572 = (forvar3572 + (1'h1)))
                    begin
                      reg3573 <= {$signed((8'hb5))};
                      reg3574 <= ($unsigned(forvar3503[(2'h3):(2'h3)]) + (wire3368[(2'h3):(2'h2)] == {{reg3565}}));
                      reg3575 <= $unsigned($signed($unsigned(reg3471[(1'h0):(1'h0)])));
                    end
                end
            end
          for (forvar3576 = (1'h0); (forvar3576 < (2'h3)); forvar3576 = (forvar3576 + (1'h1)))
            begin
              if ((^~($unsigned($unsigned(reg3377)) ?
                  $signed(forvar3485[(3'h5):(3'h4)]) : ($signed(reg3389) == (reg3466 ?
                      (8'hb1) : reg3450)))))
                begin
                  for (forvar3577 = (1'h0); (forvar3577 < (2'h3)); forvar3577 = (forvar3577 + (1'h1)))
                    begin
                      reg3578 <= $unsigned(wire3437[(1'h1):(1'h0)]);
                      reg3579 <= (({(reg3477 == forvar3522)} != {reg3551[(1'h1):(1'h0)]}) | ((^$signed(reg3502)) <<< ((forvar3506 <<< forvar3443) ?
                          reg3466[(1'h0):(1'h0)] : (reg3531 + reg3384))));
                      reg3580 <= $unsigned(((~forvar3524) ?
                          (&(wire3370 > (8'h9e))) : ((reg3478 >= forvar3465) ?
                              (forvar3495 << reg3496) : (reg3500 >> (8'ha7)))));
                      reg3581 <= forvar3490;
                    end
                end
              else
                begin
                  for (forvar3577 = (1'h0); (forvar3577 < (1'h0)); forvar3577 = (forvar3577 + (1'h1)))
                    begin
                      reg3578 <= $signed((+(^~{forvar3442})));
                      reg3579 <= $signed((^~reg3532));
                      reg3580 <= $signed((&(~^reg3504[(1'h0):(1'h0)])));
                      reg3581 <= {((forvar3469 ^ reg3482) || (reg3572 ?
                              (8'ha5) : $unsigned((8'ha2))))};
                    end
                end
              reg3582 <= $signed($unsigned(($signed(wire3414) >= forvar3456)));
              for (forvar3583 = (1'h0); (forvar3583 < (1'h1)); forvar3583 = (forvar3583 + (1'h1)))
                begin
                  for (forvar3584 = (1'h0); (forvar3584 < (1'h0)); forvar3584 = (forvar3584 + (1'h1)))
                    begin
                      reg3585 <= $signed({reg3571});
                      reg3586 <= ((reg3527[(1'h1):(1'h1)] ?
                              forvar3552 : $unsigned((&forvar3376))) ?
                          {{((8'h9c) ?
                                      (8'hae) : reg3534)}} : $unsigned(reg3468));
                    end
                  for (forvar3587 = (1'h0); (forvar3587 < (2'h2)); forvar3587 = (forvar3587 + (1'h1)))
                    begin
                      reg3588 <= forvar3478[(2'h2):(1'h1)];
                      reg3589 <= reg3535[(4'h9):(1'h0)];
                    end
                  if (reg3534)
                    begin
                      reg3590 <= $signed((reg3381 ?
                          $signed(((8'h9d) ? wire3374 : reg3532)) : ((reg3495 ?
                                  reg3465 : wire3375) ?
                              reg3547[(4'hc):(4'h8)] : (reg3460 ?
                                  reg3566 : reg3384))));
                      reg3591 <= ($unsigned({(!reg3488)}) - ({(forvar3587 ?
                              reg3535 : reg3503)} <= ((~&forvar3577) ?
                          $signed(reg3511) : (reg3536 ?
                              reg3459 : forvar3510))));
                      reg3592 <= forvar3500[(2'h2):(1'h0)];
                      reg3593 <= forvar3587;
                    end
                  else
                    begin
                      reg3590 <= ($unsigned((reg3480[(2'h2):(1'h0)] ?
                              ((8'hb9) ?
                                  forvar3458 : forvar3522) : $unsigned(reg3558))) ?
                          forvar3576[(1'h0):(1'h0)] : reg3388[(4'ha):(1'h1)]);
                      reg3591 <= $unsigned($unsigned(reg3408[(2'h2):(2'h2)]));
                      reg3592 <= ($unsigned($signed(((8'hb0) <<< (8'had)))) ?
                          $unsigned($unsigned($unsigned(reg3580))) : $signed($signed((reg3497 ?
                              (8'hb0) : forvar3455))));
                    end
                end
              reg3594 <= {{(^(reg3590 && forvar3558))}};
            end
          if ((|reg3594[(3'h5):(3'h4)]))
            begin
              for (forvar3595 = (1'h0); (forvar3595 < (2'h3)); forvar3595 = (forvar3595 + (1'h1)))
                begin
                  for (forvar3596 = (1'h0); (forvar3596 < (1'h0)); forvar3596 = (forvar3596 + (1'h1)))
                    begin
                      reg3597 <= $signed(reg3534);
                      reg3598 <= ({forvar3500} ?
                          forvar3595[(3'h5):(1'h0)] : $signed($unsigned({reg3464})));
                      reg3599 <= (&(((forvar3442 ? forvar3448 : forvar3530) ?
                              wire3370[(1'h0):(1'h0)] : $signed(reg3573)) ?
                          (8'ha6) : ((reg3565 == wire3375) & (~|reg3594))));
                      reg3600 <= $unsigned(reg3401[(1'h0):(1'h0)]);
                    end
                  if (($unsigned($unsigned(((8'hab) ^~ reg3528))) & (((|reg3389) | $signed((8'hb1))) * reg3553)))
                    begin
                      reg3601 <= ($signed((-(reg3447 >>> forvar3495))) == ($unsigned(wire3375) <= wire3370));
                    end
                  else
                    begin
                      reg3601 <= (^$signed(($signed(reg3586) ?
                          (~^reg3478) : $signed(reg3494))));
                    end
                end
              reg3602 <= (~^$unsigned((~|reg3589)));
            end
          else
            begin
              if ({((-(forvar3465 ?
                      forvar3495 : (8'h9c))) <= $unsigned(forvar3587[(3'h5):(3'h4)]))})
                begin
                  for (forvar3595 = (1'h0); (forvar3595 < (2'h3)); forvar3595 = (forvar3595 + (1'h1)))
                    begin
                      reg3596 <= ((8'h9e) * (!((forvar3499 != reg3461) ?
                          $unsigned(reg3470) : {reg3589})));
                    end
                  for (forvar3597 = (1'h0); (forvar3597 < (1'h0)); forvar3597 = (forvar3597 + (1'h1)))
                    begin
                      reg3598 <= reg3464;
                    end
                  reg3599 <= wire3372;
                end
              else
                begin
                  for (forvar3595 = (1'h0); (forvar3595 < (1'h0)); forvar3595 = (forvar3595 + (1'h1)))
                    begin
                      reg3596 <= $unsigned(($signed($unsigned(wire3373)) ?
                          (|(forvar3491 + forvar3454)) : $unsigned($signed(reg3493))));
                      reg3597 <= $signed((reg3411 ?
                          reg3500[(2'h2):(1'h0)] : forvar3469));
                      reg3598 <= (&(!reg3570[(2'h2):(1'h1)]));
                      reg3599 <= reg3382;
                    end
                  for (forvar3600 = (1'h0); (forvar3600 < (1'h0)); forvar3600 = (forvar3600 + (1'h1)))
                    begin
                      reg3601 <= (reg3453[(3'h5):(2'h3)] < reg3553[(1'h1):(1'h1)]);
                    end
                  reg3602 <= $unsigned($unsigned((reg3514[(1'h0):(1'h0)] ?
                      ((8'had) & reg3516) : (forvar3522 <= reg3499))));
                end
              for (forvar3603 = (1'h0); (forvar3603 < (2'h3)); forvar3603 = (forvar3603 + (1'h1)))
                begin
                  for (forvar3604 = (1'h0); (forvar3604 < (1'h1)); forvar3604 = (forvar3604 + (1'h1)))
                    begin
                      reg3605 <= $signed(reg3385);
                      reg3606 <= (reg3520[(3'h4):(3'h4)] ?
                          ((~|(!(8'haf))) | forvar3376[(4'hd):(3'h7)]) : $unsigned(((reg3475 && forvar3604) ?
                              $unsigned(reg3377) : wire3371[(3'h4):(1'h0)])));
                      reg3607 <= $signed(forvar3547[(3'h4):(2'h3)]);
                    end
                end
              reg3608 <= ({reg3555[(2'h3):(1'h0)]} ?
                  ((!$signed(reg3488)) ?
                      $unsigned($signed((8'ha6))) : ((forvar3503 == forvar3480) ?
                          forvar3522[(2'h3):(1'h0)] : reg3469[(3'h5):(1'h1)])) : $unsigned((((8'hac) & reg3494) ?
                      $signed(reg3501) : $signed(reg3497))));
            end
        end
      else
        begin
          if ($signed((reg3513[(4'hb):(3'h5)] ? forvar3440 : reg3412)))
            begin
              if ($signed(reg3411))
                begin
                  for (forvar3547 = (1'h0); (forvar3547 < (2'h2)); forvar3547 = (forvar3547 + (1'h1)))
                    begin
                      reg3548 <= $signed($signed((forvar3446 >= reg3488[(1'h1):(1'h1)])));
                      reg3549 <= $signed((-$unsigned($signed(forvar3446))));
                      reg3550 <= (({(forvar3440 && forvar3506)} >= ({reg3389} | reg3596[(4'hb):(3'h6)])) ?
                          {wire3374} : ($unsigned($unsigned(reg3529)) ?
                              $signed((^~forvar3576)) : $signed(reg3542)));
                      reg3551 <= (~reg3495);
                    end
                  for (forvar3552 = (1'h0); (forvar3552 < (1'h0)); forvar3552 = (forvar3552 + (1'h1)))
                    begin
                      reg3553 <= reg3541;
                      reg3554 <= reg3467;
                    end
                end
              else
                begin
                  reg3547 <= (+{(8'hb1)});
                  for (forvar3548 = (1'h0); (forvar3548 < (1'h0)); forvar3548 = (forvar3548 + (1'h1)))
                    begin
                      reg3549 <= $unsigned(forvar3576);
                      reg3550 <= $unsigned($signed($unsigned($signed(reg3594))));
                    end
                  for (forvar3551 = (1'h0); (forvar3551 < (2'h3)); forvar3551 = (forvar3551 + (1'h1)))
                    begin
                      reg3552 <= ($signed((reg3413 ?
                          $unsigned(reg3507) : $unsigned(forvar3441))) >>> (!reg3509));
                      reg3553 <= (wire3372 ?
                          forvar3454 : $unsigned({(reg3464 ?
                                  reg3564 : forvar3485)}));
                      reg3554 <= $signed($signed((8'hab)));
                    end
                end
              for (forvar3555 = (1'h0); (forvar3555 < (2'h2)); forvar3555 = (forvar3555 + (1'h1)))
                begin
                  for (forvar3556 = (1'h0); (forvar3556 < (2'h2)); forvar3556 = (forvar3556 + (1'h1)))
                    begin
                      reg3557 <= $unsigned((8'ha2));
                      reg3558 <= forvar3597;
                      reg3559 <= $unsigned(forvar3563);
                    end
                end
              for (forvar3560 = (1'h0); (forvar3560 < (2'h2)); forvar3560 = (forvar3560 + (1'h1)))
                begin
                  reg3561 <= forvar3563[(1'h0):(1'h0)];
                  for (forvar3562 = (1'h0); (forvar3562 < (1'h0)); forvar3562 = (forvar3562 + (1'h1)))
                    begin
                      reg3563 <= $signed($signed({reg3502[(2'h2):(2'h2)]}));
                      reg3564 <= $unsigned(forvar3522[(1'h1):(1'h0)]);
                      reg3565 <= $signed({(reg3467[(1'h0):(1'h0)] ?
                              (reg3589 == reg3439) : forvar3556[(1'h1):(1'h1)])});
                    end
                end
              if (reg3463[(1'h1):(1'h1)])
                begin
                  for (forvar3566 = (1'h0); (forvar3566 < (2'h2)); forvar3566 = (forvar3566 + (1'h1)))
                    begin
                      reg3567 <= reg3572[(3'h4):(1'h1)];
                      reg3568 <= (reg3535[(3'h4):(3'h4)] <= $signed($unsigned(reg3558)));
                    end
                  for (forvar3569 = (1'h0); (forvar3569 < (2'h2)); forvar3569 = (forvar3569 + (1'h1)))
                    begin
                      reg3570 <= $unsigned($unsigned($signed((wire3373 + reg3452))));
                      reg3571 <= (forvar3521[(1'h1):(1'h1)] ?
                          (^reg3481[(4'hc):(4'hc)]) : $unsigned({(forvar3443 ?
                                  forvar3556 : reg3572)}));
                    end
                  for (forvar3572 = (1'h0); (forvar3572 < (1'h0)); forvar3572 = (forvar3572 + (1'h1)))
                    begin
                      reg3573 <= reg3500;
                      reg3574 <= (&((~|reg3460) ?
                          (reg3386 <= (&reg3456)) : ((~&reg3593) >= reg3413)));
                      reg3575 <= reg3381[(4'ha):(4'ha)];
                    end
                end
              else
                begin
                  for (forvar3566 = (1'h0); (forvar3566 < (1'h0)); forvar3566 = (forvar3566 + (1'h1)))
                    begin
                      reg3567 <= $unsigned({forvar3510});
                      reg3568 <= $unsigned({$unsigned((reg3541 & reg3507))});
                    end
                  for (forvar3569 = (1'h0); (forvar3569 < (1'h0)); forvar3569 = (forvar3569 + (1'h1)))
                    begin
                      reg3570 <= $unsigned((((reg3532 <<< reg3556) ?
                              $unsigned((8'h9c)) : $signed(reg3394)) ?
                          $signed($unsigned((8'hae))) : $unsigned((^~(8'ha5)))));
                      reg3571 <= $signed($signed(($signed(reg3386) || wire3415)));
                      reg3572 <= (((~$signed(forvar3600)) >> $signed(forvar3455)) & (reg3585[(4'h9):(3'h5)] ?
                          $signed((!forvar3600)) : forvar3454));
                      reg3573 <= $signed((({forvar3395} ?
                          ((8'had) ?
                              forvar3562 : reg3568) : $unsigned(reg3477)) ~^ ((reg3485 ?
                              forvar3506 : reg3544) ?
                          $unsigned(wire3437) : (|reg3380))));
                    end
                  for (forvar3574 = (1'h0); (forvar3574 < (2'h2)); forvar3574 = (forvar3574 + (1'h1)))
                    begin
                      reg3575 <= $signed((~((~reg3464) * (reg3439 ?
                          forvar3587 : wire3415))));
                    end
                end
            end
          else
            begin
              if ($unsigned((~&$unsigned({(8'h9c)}))))
                begin
                  reg3547 <= (((~$unsigned(reg3489)) ?
                      $unsigned(forvar3485) : ((forvar3476 ?
                              reg3559 : reg3384) ?
                          {forvar3491} : (reg3594 ?
                              reg3397 : reg3406))) & ((~reg3534[(3'h5):(1'h1)]) ?
                      {$signed(reg3588)} : reg3602));
                end
              else
                begin
                  for (forvar3547 = (1'h0); (forvar3547 < (1'h1)); forvar3547 = (forvar3547 + (1'h1)))
                    begin
                      reg3548 <= reg3407[(1'h0):(1'h0)];
                      reg3549 <= ($unsigned($signed(((8'hba) >> reg3565))) ?
                          (~{(|forvar3490)}) : $signed(reg3607[(1'h0):(1'h0)]));
                    end
                  reg3550 <= $unsigned({(~^$unsigned((8'ha8)))});
                  reg3551 <= {(-$unsigned($signed((8'ha4))))};
                  if (($signed((&{forvar3560})) * {(!$unsigned(reg3498))}))
                    begin
                      reg3552 <= (forvar3515[(1'h1):(1'h0)] ?
                          forvar3448 : $signed($unsigned((+reg3504))));
                      reg3553 <= wire3374[(2'h3):(1'h1)];
                      reg3554 <= ($unsigned((reg3540 ?
                              (forvar3548 ? forvar3604 : reg3525) : (reg3566 ?
                                  forvar3469 : reg3459))) ?
                          forvar3469[(1'h0):(1'h0)] : (reg3529 * (~&{forvar3386})));
                    end
                  else
                    begin
                      reg3552 <= (&(((reg3535 ?
                          reg3413 : reg3408) <= (+(8'ha4))) >>> ((reg3569 ?
                          reg3500 : reg3506) != forvar3508)));
                      reg3553 <= (wire3375 ?
                          {forvar3499[(3'h7):(3'h6)]} : $unsigned((~&(wire3375 ?
                              reg3546 : reg3381))));
                      reg3554 <= reg3555;
                      reg3555 <= (reg3404 | $signed((~^reg3549)));
                    end
                end
              reg3556 <= (~^reg3401[(1'h1):(1'h0)]);
            end
          if (({$unsigned($unsigned(forvar3499))} ?
              ($signed($signed(forvar3508)) ?
                  forvar3491 : $signed($signed(reg3482))) : $unsigned(((&forvar3574) > (reg3558 <= reg3475)))))
            begin
              for (forvar3576 = (1'h0); (forvar3576 < (2'h3)); forvar3576 = (forvar3576 + (1'h1)))
                begin
                  if (((reg3450[(1'h1):(1'h0)] ^~ reg3496) ?
                      forvar3521[(4'h9):(4'h8)] : $signed(reg3557[(3'h4):(2'h3)])))
                    begin
                      reg3577 <= forvar3503[(1'h1):(1'h1)];
                      reg3578 <= ($signed(((reg3548 ?
                              forvar3481 : forvar3441) ^ $unsigned(wire3370))) ?
                          $signed($signed(forvar3387)) : ((~^(~^reg3551)) <= (+reg3413)));
                    end
                  else
                    begin
                      reg3577 <= (^reg3519[(2'h2):(1'h1)]);
                      reg3578 <= (($unsigned({wire3368}) ?
                              $unsigned((~^reg3592)) : $unsigned($signed(wire3373))) ?
                          $signed($unsigned($signed(forvar3574))) : ($unsigned({reg3489}) ?
                              reg3392 : $signed((forvar3559 && reg3450))));
                      reg3579 <= $unsigned(((&forvar3448) > (+$unsigned(reg3386))));
                    end
                  for (forvar3580 = (1'h0); (forvar3580 < (1'h1)); forvar3580 = (forvar3580 + (1'h1)))
                    begin
                      reg3581 <= reg3459[(4'h8):(4'h8)];
                    end
                end
              if (((+reg3558) ?
                  $unsigned(forvar3515) : (reg3397[(2'h3):(1'h1)] < reg3387)))
                begin
                  for (forvar3582 = (1'h0); (forvar3582 < (1'h0)); forvar3582 = (forvar3582 + (1'h1)))
                    begin
                      reg3583 <= reg3572[(1'h1):(1'h0)];
                      reg3584 <= reg3529;
                      reg3585 <= reg3572;
                      reg3586 <= ((~(~^(reg3574 ? forvar3455 : forvar3595))) ?
                          $signed((!$signed(forvar3568))) : (8'haa));
                    end
                  reg3587 <= $signed($unsigned(reg3512));
                  if ($unsigned((|(forvar3595[(3'h6):(3'h5)] * (reg3484 ?
                      forvar3600 : forvar3395)))))
                    begin
                      reg3588 <= (reg3550[(2'h3):(1'h0)] ?
                          (&reg3458[(2'h2):(1'h1)]) : reg3410);
                    end
                  else
                    begin
                      reg3588 <= (reg3495[(4'h8):(2'h2)] ^~ $signed($unsigned($unsigned(forvar3398))));
                      reg3589 <= ($unsigned(forvar3545[(1'h1):(1'h0)]) ~^ $signed($signed((forvar3443 ~^ reg3399))));
                      reg3590 <= ((^~$unsigned($signed(reg3549))) ?
                          (&(|forvar3582)) : reg3534[(2'h2):(1'h0)]);
                      reg3591 <= (!(^(-forvar3522[(1'h0):(1'h0)])));
                    end
                end
              else
                begin
                  reg3582 <= $unsigned({(forvar3500 + forvar3508)});
                  for (forvar3583 = (1'h0); (forvar3583 < (2'h2)); forvar3583 = (forvar3583 + (1'h1)))
                    begin
                      reg3584 <= (~|({(forvar3580 ? reg3497 : reg3445)} ?
                          ($unsigned(reg3400) ?
                              $unsigned(reg3505) : $signed(reg3581)) : ({reg3491} ?
                              reg3467 : (reg3477 ^ forvar3405))));
                    end
                end
              if (reg3399)
                begin
                  reg3592 <= (forvar3530 ?
                      ($unsigned(reg3529) & $signed(reg3395)) : (8'ha3));
                end
              else
                begin
                  for (forvar3592 = (1'h0); (forvar3592 < (2'h3)); forvar3592 = (forvar3592 + (1'h1)))
                    begin
                      reg3593 <= ((8'ha0) ?
                          reg3377[(4'ha):(1'h1)] : forvar3388[(3'h5):(1'h0)]);
                      reg3594 <= (8'ha7);
                      reg3595 <= forvar3398;
                      reg3596 <= $unsigned((-{reg3483[(4'hc):(3'h7)]}));
                    end
                  for (forvar3597 = (1'h0); (forvar3597 < (2'h2)); forvar3597 = (forvar3597 + (1'h1)))
                    begin
                      reg3598 <= ((reg3486 < $signed((^forvar3568))) ?
                          reg3396 : $signed(reg3565[(2'h2):(2'h2)]));
                      reg3599 <= ((~&($signed(reg3482) << $unsigned(forvar3458))) ^ forvar3600);
                      reg3600 <= reg3484;
                    end
                  if ((^~(|$unsigned($unsigned(reg3569)))))
                    begin
                      reg3601 <= $signed($unsigned({(~&wire3371)}));
                      reg3602 <= $signed(forvar3510);
                      reg3603 <= $signed($signed((!forvar3595)));
                    end
                  else
                    begin
                      reg3601 <= ((~^{$signed(reg3485)}) << $signed({(reg3582 ?
                              reg3551 : reg3484)}));
                      reg3602 <= $signed(reg3523);
                      reg3603 <= (8'hb8);
                      reg3604 <= wire3437;
                    end
                end
            end
          else
            begin
              if (reg3473)
                begin
                  reg3576 <= reg3381[(3'h5):(1'h1)];
                  for (forvar3577 = (1'h0); (forvar3577 < (1'h0)); forvar3577 = (forvar3577 + (1'h1)))
                    begin
                      reg3578 <= reg3550;
                      reg3579 <= reg3606;
                    end
                  for (forvar3580 = (1'h0); (forvar3580 < (2'h2)); forvar3580 = (forvar3580 + (1'h1)))
                    begin
                      reg3581 <= $signed(((~^$signed(reg3471)) == reg3606));
                      reg3582 <= $unsigned($unsigned({reg3593[(2'h2):(2'h2)]}));
                      reg3583 <= $unsigned($signed(($signed(reg3570) >> $signed(forvar3545))));
                      reg3584 <= (~&$signed($signed((reg3593 == reg3598))));
                    end
                  for (forvar3585 = (1'h0); (forvar3585 < (1'h1)); forvar3585 = (forvar3585 + (1'h1)))
                    begin
                      reg3586 <= reg3486[(3'h4):(1'h1)];
                      reg3587 <= ({$unsigned((forvar3454 ?
                              reg3514 : forvar3387))} ~^ reg3603[(2'h2):(1'h1)]);
                      reg3588 <= forvar3506[(3'h4):(1'h1)];
                      reg3589 <= ((forvar3511 ?
                          reg3501[(4'h9):(3'h4)] : (|forvar3574[(1'h0):(1'h0)])) | reg3461);
                    end
                end
              else
                begin
                  for (forvar3576 = (1'h0); (forvar3576 < (1'h1)); forvar3576 = (forvar3576 + (1'h1)))
                    begin
                      reg3577 <= (~^$signed(reg3483));
                    end
                  reg3578 <= {((&reg3498) ?
                          $unsigned($signed(reg3599)) : reg3466)};
                  reg3579 <= forvar3480;
                  reg3580 <= forvar3399[(3'h6):(1'h1)];
                end
              for (forvar3590 = (1'h0); (forvar3590 < (1'h0)); forvar3590 = (forvar3590 + (1'h1)))
                begin
                  if ($signed(reg3499[(1'h0):(1'h0)]))
                    begin
                      reg3591 <= ($signed($unsigned($signed(reg3472))) ?
                          reg3593 : forvar3518[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg3591 <= {$unsigned((^reg3540[(4'h9):(3'h5)]))};
                      reg3592 <= $signed((^~(forvar3464[(1'h1):(1'h0)] - ((8'ha0) >> reg3469))));
                    end
                  if ((~^(forvar3524[(3'h4):(3'h4)] ?
                      (~&(forvar3511 ?
                          reg3538 : reg3557)) : forvar3574[(2'h2):(1'h1)])))
                    begin
                      reg3593 <= $unsigned($signed(($signed(reg3599) <<< reg3391[(1'h1):(1'h1)])));
                      reg3594 <= forvar3395[(3'h5):(1'h0)];
                      reg3595 <= $unsigned(($unsigned($signed(reg3585)) ^ forvar3559[(1'h0):(1'h0)]));
                      reg3596 <= (8'ha7);
                    end
                  else
                    begin
                      reg3593 <= reg3562[(2'h3):(2'h2)];
                      reg3594 <= (~&reg3562);
                    end
                end
              for (forvar3597 = (1'h0); (forvar3597 < (1'h0)); forvar3597 = (forvar3597 + (1'h1)))
                begin
                  for (forvar3598 = (1'h0); (forvar3598 < (2'h3)); forvar3598 = (forvar3598 + (1'h1)))
                    begin
                      reg3599 <= reg3461[(1'h1):(1'h1)];
                      reg3600 <= $unsigned($signed($signed(reg3406[(2'h2):(1'h0)])));
                      reg3601 <= ($unsigned((reg3554 || (^reg3572))) ?
                          reg3509 : $unsigned(((reg3581 ?
                              wire3372 : (8'hba)) >> (reg3447 ?
                              reg3526 : reg3544))));
                      reg3602 <= $unsigned($unsigned((~$signed(reg3514))));
                    end
                  reg3603 <= $signed($signed((^~(reg3546 ?
                      (8'ha2) : forvar3515))));
                  for (forvar3604 = (1'h0); (forvar3604 < (2'h2)); forvar3604 = (forvar3604 + (1'h1)))
                    begin
                      reg3605 <= ((~&($unsigned(reg3477) & $unsigned(reg3547))) ^ (forvar3567[(3'h4):(1'h1)] && {(8'hae)}));
                      reg3606 <= $signed((-{((8'h9f) > forvar3545)}));
                    end
                  reg3607 <= ($unsigned(reg3445[(3'h7):(2'h3)]) ?
                      wire3368[(4'ha):(3'h5)] : ($unsigned($unsigned(reg3604)) ?
                          {$signed(forvar3551)} : reg3481));
                end
            end
          for (forvar3608 = (1'h0); (forvar3608 < (1'h1)); forvar3608 = (forvar3608 + (1'h1)))
            begin
              reg3609 <= forvar3577;
            end
          reg3610 <= $unsigned(forvar3555);
        end
      reg3611 <= {reg3548};
      reg3612 <= (reg3517 >>> (($unsigned(reg3472) == $unsigned(reg3468)) ?
          ($unsigned(reg3561) >>> forvar3567) : $unsigned((reg3592 ?
              reg3519 : reg3599))));
    end
  assign wire3613 = $signed(((~|$unsigned(forvar3442)) ?
                        ($unsigned(forvar3577) ?
                            {reg3477} : (forvar3458 <= reg3388)) : (^(reg3484 == forvar3443))));
  assign wire3614 = ((forvar3383 & (8'hb8)) ?
                        $signed($unsigned((~^reg3596))) : forvar3440);
  assign wire3615 = (reg3596 ?
                        $signed($signed((reg3608 ^ reg3585))) : $signed($signed(reg3531)));
  always
    @(posedge clk) begin
      for (forvar3616 = (1'h0); (forvar3616 < (2'h3)); forvar3616 = (forvar3616 + (1'h1)))
        begin
          for (forvar3617 = (1'h0); (forvar3617 < (1'h1)); forvar3617 = (forvar3617 + (1'h1)))
            begin
              for (forvar3618 = (1'h0); (forvar3618 < (1'h0)); forvar3618 = (forvar3618 + (1'h1)))
                begin
                  for (forvar3619 = (1'h0); (forvar3619 < (2'h3)); forvar3619 = (forvar3619 + (1'h1)))
                    begin
                      reg3620 <= (reg3504 ?
                          ($signed(reg3485[(4'hb):(3'h5)]) || forvar3582[(3'h4):(1'h1)]) : (forvar3617[(2'h2):(1'h0)] <= {(reg3393 - forvar3508)}));
                    end
                  if ($unsigned($signed((~|(~reg3583)))))
                    begin
                      reg3621 <= {((~(|forvar3583)) >>> forvar3485)};
                    end
                  else
                    begin
                      reg3621 <= (+forvar3500);
                    end
                  for (forvar3622 = (1'h0); (forvar3622 < (2'h2)); forvar3622 = (forvar3622 + (1'h1)))
                    begin
                      reg3623 <= (^~(8'had));
                    end
                  for (forvar3624 = (1'h0); (forvar3624 < (1'h0)); forvar3624 = (forvar3624 + (1'h1)))
                    begin
                      reg3625 <= reg3452[(4'h8):(3'h6)];
                      reg3626 <= ((^~(|reg3497[(3'h5):(2'h3)])) ?
                          forvar3576[(4'he):(4'hb)] : $signed((reg3410 ?
                              (forvar3377 ~^ reg3557) : reg3382[(1'h1):(1'h1)])));
                      reg3627 <= wire3614[(2'h3):(2'h3)];
                    end
                end
            end
        end
    end
  assign wire3628 = reg3564;
  assign wire3629 = reg3400;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2168  (y, clk, wire2173, wire2172, wire2171, wire2170, wire2169);
  output wire [(32'hbf8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire2173;
  input wire signed [(4'hf):(1'h0)] wire2172;
  input wire [(4'he):(1'h0)] wire2171;
  input wire [(4'hd):(1'h0)] wire2170;
  input wire [(3'h6):(1'h0)] wire2169;
  reg signed [(2'h3):(1'h0)] reg3364 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3363 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3359 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3362 = (1'h0);
  reg [(4'hb):(1'h0)] reg3361 = (1'h0);
  reg [(3'h7):(1'h0)] reg3360 = (1'h0);
  reg [(3'h7):(1'h0)] reg3359 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3358 = (1'h0);
  reg [(3'h4):(1'h0)] reg3357 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3356 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3355 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3354 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3353 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3352 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3351 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3350 = (1'h0);
  reg [(3'h6):(1'h0)] reg3349 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3348 = (1'h0);
  reg [(2'h3):(1'h0)] reg3347 = (1'h0);
  reg [(2'h2):(1'h0)] reg3346 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3345 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3344 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3343 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3342 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3341 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3340 = (1'h0);
  reg [(4'hb):(1'h0)] reg3339 = (1'h0);
  reg [(3'h5):(1'h0)] reg3338 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3337 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3336 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3335 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3333 = (1'h0);
  reg [(2'h3):(1'h0)] reg3332 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3331 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3330 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3329 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3328 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3327 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3326 = (1'h0);
  reg [(4'h8):(1'h0)] reg3325 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3324 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3323 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3322 = (1'h0);
  reg [(4'hf):(1'h0)] reg3321 = (1'h0);
  reg [(2'h2):(1'h0)] reg3320 = (1'h0);
  reg [(3'h4):(1'h0)] reg3319 = (1'h0);
  reg [(4'hb):(1'h0)] reg3318 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3317 = (1'h0);
  reg [(2'h2):(1'h0)] reg3316 = (1'h0);
  reg [(4'h9):(1'h0)] reg3315 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3314 = (1'h0);
  reg [(3'h7):(1'h0)] reg3313 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3312 = (1'h0);
  reg [(5'h10):(1'h0)] reg3311 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3310 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3309 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3308 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3307 = (1'h0);
  reg [(4'h9):(1'h0)] reg3306 = (1'h0);
  reg [(4'hc):(1'h0)] reg3305 = (1'h0);
  reg [(2'h2):(1'h0)] reg3304 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3303 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3302 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3301 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3300 = (1'h0);
  reg [(4'h9):(1'h0)] reg3299 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3298 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3297 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3296 = (1'h0);
  reg [(2'h2):(1'h0)] reg3295 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3294 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3293 = (1'h0);
  reg [(4'hb):(1'h0)] reg3292 = (1'h0);
  reg [(5'h10):(1'h0)] reg3291 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3290 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3289 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3288 = (1'h0);
  reg [(4'hd):(1'h0)] reg3287 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3286 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3285 = (1'h0);
  reg [(4'h8):(1'h0)] reg3284 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3283 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3282 = (1'h0);
  reg [(5'h10):(1'h0)] reg3269 = (1'h0);
  reg [(4'hd):(1'h0)] reg3281 = (1'h0);
  reg [(4'ha):(1'h0)] reg3280 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3279 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3274 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3279 = (1'h0);
  reg [(4'hd):(1'h0)] reg3278 = (1'h0);
  reg [(4'he):(1'h0)] reg3277 = (1'h0);
  reg [(2'h3):(1'h0)] reg3276 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3275 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3274 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3273 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3272 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3271 = (1'h0);
  reg [(4'ha):(1'h0)] reg3270 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3269 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3268 = (1'h0);
  reg [(4'hb):(1'h0)] reg3267 = (1'h0);
  reg [(4'ha):(1'h0)] reg3252 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3248 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3245 = (1'h0);
  reg [(4'hf):(1'h0)] reg3266 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3265 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3263 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3264 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3263 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3262 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3261 = (1'h0);
  reg [(4'hb):(1'h0)] reg3260 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3259 = (1'h0);
  reg [(4'ha):(1'h0)] reg3244 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3258 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3257 = (1'h0);
  reg [(4'hb):(1'h0)] reg3256 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3255 = (1'h0);
  reg [(4'hd):(1'h0)] reg3254 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3253 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3252 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3251 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3250 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3249 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3248 = (1'h0);
  reg [(4'h8):(1'h0)] reg3247 = (1'h0);
  reg [(3'h5):(1'h0)] reg3246 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3245 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3244 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3243 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3242 = (1'h0);
  reg [(4'h9):(1'h0)] reg3241 = (1'h0);
  reg [(3'h5):(1'h0)] reg3240 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3239 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3238 = (1'h0);
  reg [(2'h2):(1'h0)] reg3237 = (1'h0);
  reg [(4'ha):(1'h0)] reg3236 = (1'h0);
  reg [(4'ha):(1'h0)] reg3235 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3234 = (1'h0);
  reg [(4'hd):(1'h0)] reg3233 = (1'h0);
  reg [(3'h4):(1'h0)] reg3232 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3231 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3230 = (1'h0);
  reg [(3'h6):(1'h0)] reg3229 = (1'h0);
  reg [(4'hc):(1'h0)] reg3228 = (1'h0);
  reg [(5'h10):(1'h0)] reg3227 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3226 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3225 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3224 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3199 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3223 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3222 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3221 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3220 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3217 = (1'h0);
  reg [(4'ha):(1'h0)] reg3219 = (1'h0);
  reg [(4'h8):(1'h0)] reg3218 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3217 = (1'h0);
  reg [(4'he):(1'h0)] reg3216 = (1'h0);
  reg [(4'hb):(1'h0)] reg3215 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3214 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3213 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3212 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3211 = (1'h0);
  reg [(3'h6):(1'h0)] reg3210 = (1'h0);
  reg [(2'h2):(1'h0)] reg3209 = (1'h0);
  reg [(4'hc):(1'h0)] reg3208 = (1'h0);
  reg [(4'hd):(1'h0)] reg3207 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3206 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3204 = (1'h0);
  reg [(2'h3):(1'h0)] reg3203 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3201 = (1'h0);
  reg [(4'h9):(1'h0)] reg3205 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3204 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3203 = (1'h0);
  reg [(3'h5):(1'h0)] reg3202 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3201 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3200 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3199 = (1'h0);
  reg [(3'h4):(1'h0)] reg3198 = (1'h0);
  reg [(5'h10):(1'h0)] reg3197 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3196 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3195 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3194 = (1'h0);
  reg [(4'h8):(1'h0)] reg3193 = (1'h0);
  reg [(5'h10):(1'h0)] reg3192 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3191 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3190 = (1'h0);
  reg [(4'hd):(1'h0)] reg3189 = (1'h0);
  reg [(4'ha):(1'h0)] reg3188 = (1'h0);
  reg [(3'h4):(1'h0)] reg3187 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3186 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3185 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3184 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3183 = (1'h0);
  reg [(2'h2):(1'h0)] reg3182 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3181 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3180 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3179 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3178 = (1'h0);
  reg [(2'h3):(1'h0)] reg3177 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3176 = (1'h0);
  reg [(2'h2):(1'h0)] reg3175 = (1'h0);
  reg [(4'he):(1'h0)] forvar3174 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3173 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3172 = (1'h0);
  reg [(3'h6):(1'h0)] reg3171 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3170 = (1'h0);
  reg [(2'h2):(1'h0)] reg3169 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3168 = (1'h0);
  reg [(3'h7):(1'h0)] reg3167 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3166 = (1'h0);
  reg [(3'h7):(1'h0)] reg3165 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3164 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3163 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3162 = (1'h0);
  reg [(4'ha):(1'h0)] reg3161 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3160 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3159 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3152 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3151 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3146 = (1'h0);
  reg [(4'he):(1'h0)] reg3142 = (1'h0);
  reg [(4'hd):(1'h0)] reg3158 = (1'h0);
  reg [(4'hf):(1'h0)] reg3157 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3156 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3155 = (1'h0);
  reg [(2'h3):(1'h0)] reg3154 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3153 = (1'h0);
  reg [(3'h7):(1'h0)] reg3152 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3151 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3150 = (1'h0);
  reg [(4'hc):(1'h0)] reg3149 = (1'h0);
  reg [(4'he):(1'h0)] reg3148 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3147 = (1'h0);
  reg [(3'h5):(1'h0)] reg3146 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3145 = (1'h0);
  reg [(4'hb):(1'h0)] reg3144 = (1'h0);
  reg [(4'ha):(1'h0)] reg3143 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3142 = (1'h0);
  reg [(4'hd):(1'h0)] reg3141 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3140 = (1'h0);
  reg [(3'h5):(1'h0)] reg3140 = (1'h0);
  reg [(4'hb):(1'h0)] reg3139 = (1'h0);
  reg [(3'h7):(1'h0)] reg3138 = (1'h0);
  reg [(4'ha):(1'h0)] reg3137 = (1'h0);
  reg [(4'hb):(1'h0)] reg3136 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3135 = (1'h0);
  reg [(4'hb):(1'h0)] reg3134 = (1'h0);
  reg [(4'hc):(1'h0)] reg3133 = (1'h0);
  reg [(3'h7):(1'h0)] reg3132 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3131 = (1'h0);
  reg [(4'ha):(1'h0)] reg3130 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3129 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3128 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3127 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3126 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3125 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3124 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3123 = (1'h0);
  reg [(2'h2):(1'h0)] reg3122 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3121 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3120 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3119 = (1'h0);
  reg [(4'ha):(1'h0)] reg3118 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3117 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3116 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3115 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3114 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3113 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3112 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire3110;
  wire [(3'h7):(1'h0)] wire2224;
  reg [(3'h5):(1'h0)] reg2223 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2186 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2184 = (1'h0);
  reg [(3'h5):(1'h0)] reg2182 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2181 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2221 = (1'h0);
  reg [(2'h2):(1'h0)] reg2217 = (1'h0);
  reg [(3'h4):(1'h0)] reg2222 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2221 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2220 = (1'h0);
  reg [(4'hd):(1'h0)] reg2219 = (1'h0);
  reg [(4'he):(1'h0)] reg2218 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2217 = (1'h0);
  reg [(3'h5):(1'h0)] reg2216 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2215 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2214 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2213 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2212 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2208 = (1'h0);
  reg [(4'hd):(1'h0)] reg2212 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2211 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2210 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2209 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2208 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2207 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2206 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2205 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2204 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2203 = (1'h0);
  reg [(3'h5):(1'h0)] reg2202 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2201 = (1'h0);
  reg [(4'ha):(1'h0)] reg2200 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2199 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2198 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2197 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2196 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2193 = (1'h0);
  reg [(4'h9):(1'h0)] reg2197 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2196 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2195 = (1'h0);
  reg [(4'ha):(1'h0)] reg2194 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2193 = (1'h0);
  reg [(4'he):(1'h0)] reg2192 = (1'h0);
  reg [(3'h7):(1'h0)] reg2191 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2190 = (1'h0);
  reg [(2'h2):(1'h0)] reg2189 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2188 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2187 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2186 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2185 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2184 = (1'h0);
  reg [(3'h4):(1'h0)] reg2183 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2182 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2181 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2180 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2179 = (1'h0);
  reg [(3'h6):(1'h0)] reg2178 = (1'h0);
  reg [(3'h6):(1'h0)] reg2177 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2176 = (1'h0);
  wire [(4'ha):(1'h0)] wire2175;
  wire signed [(4'h9):(1'h0)] wire2174;
  assign y = {reg3364,
                 forvar3363,
                 forvar3359,
                 reg3362,
                 reg3361,
                 reg3360,
                 reg3359,
                 reg3358,
                 reg3357,
                 reg3356,
                 reg3355,
                 reg3354,
                 forvar3353,
                 forvar3352,
                 reg3351,
                 reg3350,
                 reg3349,
                 forvar3348,
                 reg3347,
                 reg3346,
                 forvar3345,
                 reg3344,
                 reg3343,
                 reg3342,
                 reg3341,
                 forvar3340,
                 reg3339,
                 reg3338,
                 reg3337,
                 forvar3336,
                 forvar3335,
                 reg3334,
                 reg3333,
                 reg3332,
                 forvar3331,
                 reg3330,
                 reg3329,
                 reg3328,
                 forvar3327,
                 forvar3326,
                 reg3325,
                 forvar3324,
                 reg3323,
                 forvar3322,
                 reg3321,
                 reg3320,
                 reg3319,
                 reg3318,
                 reg3317,
                 reg3316,
                 reg3315,
                 reg3314,
                 reg3313,
                 reg3312,
                 reg3311,
                 reg3310,
                 reg3309,
                 forvar3308,
                 forvar3307,
                 reg3306,
                 reg3305,
                 reg3304,
                 reg3303,
                 forvar3302,
                 reg3301,
                 reg3300,
                 reg3299,
                 reg3298,
                 forvar3297,
                 forvar3296,
                 reg3295,
                 forvar3294,
                 reg3293,
                 reg3292,
                 reg3291,
                 reg3290,
                 reg3289,
                 reg3288,
                 reg3287,
                 reg3286,
                 reg3285,
                 reg3284,
                 forvar3283,
                 forvar3282,
                 reg3269,
                 reg3281,
                 reg3280,
                 forvar3279,
                 forvar3274,
                 reg3279,
                 reg3278,
                 reg3277,
                 reg3276,
                 reg3275,
                 reg3274,
                 reg3273,
                 reg3272,
                 reg3271,
                 reg3270,
                 forvar3269,
                 forvar3268,
                 reg3267,
                 reg3252,
                 forvar3248,
                 forvar3245,
                 reg3266,
                 reg3265,
                 forvar3263,
                 reg3264,
                 reg3263,
                 reg3262,
                 reg3261,
                 reg3260,
                 forvar3259,
                 reg3244,
                 reg3258,
                 forvar3257,
                 reg3256,
                 reg3255,
                 reg3254,
                 reg3253,
                 forvar3252,
                 reg3251,
                 reg3250,
                 reg3249,
                 reg3248,
                 reg3247,
                 reg3246,
                 reg3245,
                 forvar3244,
                 reg3243,
                 forvar3242,
                 reg3241,
                 reg3240,
                 reg3239,
                 reg3238,
                 reg3237,
                 reg3236,
                 reg3235,
                 reg3234,
                 reg3233,
                 reg3232,
                 forvar3231,
                 reg3230,
                 reg3229,
                 reg3228,
                 reg3227,
                 forvar3226,
                 forvar3225,
                 forvar3224,
                 reg3199,
                 reg3223,
                 reg3222,
                 forvar3221,
                 forvar3220,
                 reg3217,
                 reg3219,
                 reg3218,
                 forvar3217,
                 reg3216,
                 reg3215,
                 reg3214,
                 reg3213,
                 forvar3212,
                 reg3211,
                 reg3210,
                 reg3209,
                 reg3208,
                 reg3207,
                 reg3206,
                 forvar3204,
                 reg3203,
                 forvar3201,
                 reg3205,
                 reg3204,
                 forvar3203,
                 reg3202,
                 reg3201,
                 reg3200,
                 forvar3199,
                 reg3198,
                 reg3197,
                 reg3196,
                 reg3195,
                 reg3194,
                 reg3193,
                 reg3192,
                 forvar3191,
                 reg3190,
                 reg3189,
                 reg3188,
                 reg3187,
                 reg3186,
                 reg3185,
                 reg3184,
                 reg3183,
                 reg3182,
                 forvar3181,
                 reg3180,
                 reg3179,
                 forvar3178,
                 reg3177,
                 reg3176,
                 reg3175,
                 forvar3174,
                 reg3173,
                 forvar3172,
                 reg3171,
                 reg3170,
                 reg3169,
                 reg3168,
                 reg3167,
                 reg3166,
                 reg3165,
                 reg3164,
                 forvar3163,
                 forvar3162,
                 reg3161,
                 reg3160,
                 forvar3159,
                 forvar3152,
                 reg3151,
                 forvar3146,
                 reg3142,
                 reg3158,
                 reg3157,
                 reg3156,
                 reg3155,
                 reg3154,
                 reg3153,
                 reg3152,
                 forvar3151,
                 reg3150,
                 reg3149,
                 reg3148,
                 reg3147,
                 reg3146,
                 reg3145,
                 reg3144,
                 reg3143,
                 forvar3142,
                 reg3141,
                 forvar3140,
                 reg3140,
                 reg3139,
                 reg3138,
                 reg3137,
                 reg3136,
                 reg3135,
                 reg3134,
                 reg3133,
                 reg3132,
                 reg3131,
                 reg3130,
                 reg3129,
                 forvar3128,
                 forvar3127,
                 reg3126,
                 forvar3125,
                 forvar3124,
                 forvar3123,
                 reg3122,
                 reg3121,
                 reg3120,
                 reg3119,
                 reg3118,
                 reg3117,
                 reg3116,
                 reg3115,
                 reg3114,
                 forvar3113,
                 forvar3112,
                 wire3110,
                 wire2224,
                 reg2223,
                 reg2186,
                 reg2184,
                 reg2182,
                 forvar2181,
                 reg2221,
                 reg2217,
                 reg2222,
                 forvar2221,
                 reg2220,
                 reg2219,
                 reg2218,
                 forvar2217,
                 reg2216,
                 reg2215,
                 reg2214,
                 reg2213,
                 forvar2212,
                 reg2208,
                 reg2212,
                 reg2211,
                 reg2210,
                 reg2209,
                 forvar2208,
                 reg2207,
                 reg2206,
                 reg2205,
                 reg2204,
                 forvar2203,
                 reg2202,
                 forvar2201,
                 reg2200,
                 reg2199,
                 reg2198,
                 forvar2197,
                 reg2196,
                 reg2193,
                 reg2197,
                 forvar2196,
                 reg2195,
                 reg2194,
                 forvar2193,
                 reg2192,
                 reg2191,
                 reg2190,
                 reg2189,
                 reg2188,
                 forvar2187,
                 forvar2186,
                 reg2185,
                 forvar2184,
                 reg2183,
                 forvar2182,
                 reg2181,
                 forvar2180,
                 reg2179,
                 reg2178,
                 reg2177,
                 forvar2176,
                 wire2175,
                 wire2174,
                 (1'h0)};
  assign wire2174 = wire2171;
  assign wire2175 = (8'h9e);
  always
    @(posedge clk) begin
      for (forvar2176 = (1'h0); (forvar2176 < (1'h0)); forvar2176 = (forvar2176 + (1'h1)))
        begin
          reg2177 <= ((~&(~^(wire2170 ^~ wire2169))) ?
              $unsigned($signed((8'hae))) : $unsigned($unsigned((~&(8'hae)))));
          reg2178 <= (wire2173 * {((-wire2169) ?
                  wire2175[(3'h7):(2'h2)] : wire2171[(1'h1):(1'h0)])});
        end
      reg2179 <= $unsigned((-reg2178[(2'h2):(2'h2)]));
      if (wire2171[(3'h5):(2'h3)])
        begin
          for (forvar2180 = (1'h0); (forvar2180 < (1'h0)); forvar2180 = (forvar2180 + (1'h1)))
            begin
              reg2181 <= wire2173[(4'hc):(3'h6)];
            end
          for (forvar2182 = (1'h0); (forvar2182 < (1'h0)); forvar2182 = (forvar2182 + (1'h1)))
            begin
              reg2183 <= $signed($unsigned($signed((forvar2176 ?
                  wire2174 : forvar2182))));
            end
          for (forvar2184 = (1'h0); (forvar2184 < (2'h3)); forvar2184 = (forvar2184 + (1'h1)))
            begin
              reg2185 <= $unsigned(wire2172);
              for (forvar2186 = (1'h0); (forvar2186 < (2'h2)); forvar2186 = (forvar2186 + (1'h1)))
                begin
                  for (forvar2187 = (1'h0); (forvar2187 < (1'h0)); forvar2187 = (forvar2187 + (1'h1)))
                    begin
                      reg2188 <= reg2178[(3'h6):(3'h4)];
                      reg2189 <= reg2181;
                      reg2190 <= (+(forvar2180 ?
                          $unsigned(forvar2184) : ((wire2172 ?
                                  (8'hb1) : forvar2187) ?
                              (~&(8'hb4)) : (&(8'ha4)))));
                    end
                  reg2191 <= (reg2177[(3'h6):(3'h4)] ?
                      $signed($unsigned($signed((8'hb3)))) : ((&(wire2173 ^~ forvar2180)) ?
                          (forvar2182[(2'h3):(2'h3)] ?
                              forvar2182 : reg2181) : $signed($unsigned(reg2188))));
                end
              if ($unsigned((wire2174 || reg2179[(2'h3):(2'h2)])))
                begin
                  reg2192 <= (forvar2180[(2'h2):(1'h0)] ?
                      $signed(((forvar2182 ? reg2177 : reg2181) ?
                          $unsigned(reg2185) : ((8'hb1) * reg2189))) : (forvar2182 && (forvar2180 ?
                          reg2190 : ((8'haa) ? wire2172 : reg2189))));
                  for (forvar2193 = (1'h0); (forvar2193 < (2'h3)); forvar2193 = (forvar2193 + (1'h1)))
                    begin
                      reg2194 <= forvar2182[(3'h5):(1'h0)];
                      reg2195 <= $unsigned(forvar2176);
                    end
                  for (forvar2196 = (1'h0); (forvar2196 < (2'h2)); forvar2196 = (forvar2196 + (1'h1)))
                    begin
                      reg2197 <= reg2189[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  reg2192 <= reg2190;
                  if (forvar2196)
                    begin
                      reg2193 <= (wire2174[(4'h8):(3'h5)] ?
                          (({reg2178} ? (forvar2186 == reg2178) : {reg2191}) ?
                              (!$unsigned(reg2191)) : ((reg2191 | reg2177) ?
                                  $signed(forvar2176) : (reg2197 * reg2181))) : (8'h9d));
                      reg2194 <= ((reg2190[(2'h3):(2'h3)] ^~ $signed(forvar2187[(2'h2):(1'h0)])) ?
                          {($unsigned(forvar2196) ?
                                  wire2175 : wire2173[(4'h9):(2'h2)])} : (~(wire2174 >= (~reg2194))));
                    end
                  else
                    begin
                      reg2193 <= reg2191[(1'h1):(1'h0)];
                      reg2194 <= (((|(reg2191 ?
                          forvar2187 : reg2178)) < ({wire2172} <= wire2175[(4'h9):(3'h6)])) <= ($unsigned($unsigned(reg2183)) ?
                          ({reg2177} ?
                              {wire2171} : reg2191[(2'h2):(2'h2)]) : (~|(~|reg2190))));
                      reg2195 <= $unsigned((($signed(forvar2186) << $unsigned(reg2188)) > ($unsigned((8'ha8)) <<< (forvar2176 ?
                          wire2173 : (8'hb9)))));
                      reg2196 <= $signed($signed((|(wire2169 ?
                          reg2183 : (8'hba)))));
                    end
                  for (forvar2197 = (1'h0); (forvar2197 < (1'h0)); forvar2197 = (forvar2197 + (1'h1)))
                    begin
                      reg2198 <= (|($unsigned((reg2191 ? reg2189 : reg2192)) ?
                          $unsigned($unsigned(reg2196)) : (-(reg2196 || reg2190))));
                      reg2199 <= $unsigned($unsigned($signed($unsigned(forvar2184))));
                      reg2200 <= $unsigned(reg2194);
                    end
                  for (forvar2201 = (1'h0); (forvar2201 < (2'h3)); forvar2201 = (forvar2201 + (1'h1)))
                    begin
                      reg2202 <= reg2194[(1'h0):(1'h0)];
                    end
                end
            end
          for (forvar2203 = (1'h0); (forvar2203 < (1'h0)); forvar2203 = (forvar2203 + (1'h1)))
            begin
              if (wire2174)
                begin
                  if (reg2192[(4'ha):(4'h9)])
                    begin
                      reg2204 <= forvar2187[(1'h0):(1'h0)];
                      reg2205 <= $signed(reg2197[(3'h5):(3'h4)]);
                      reg2206 <= {reg2200};
                    end
                  else
                    begin
                      reg2204 <= $unsigned(forvar2187[(1'h0):(1'h0)]);
                      reg2205 <= $unsigned(forvar2186);
                      reg2206 <= $signed(({$signed(wire2169)} <= (~&(|reg2193))));
                      reg2207 <= (^~$unsigned({wire2175[(4'ha):(3'h6)]}));
                    end
                  for (forvar2208 = (1'h0); (forvar2208 < (1'h1)); forvar2208 = (forvar2208 + (1'h1)))
                    begin
                      reg2209 <= reg2191[(3'h4):(1'h0)];
                      reg2210 <= (~&wire2175[(3'h6):(2'h3)]);
                      reg2211 <= (~|(~^$signed((8'ha0))));
                      reg2212 <= (~^$unsigned((^~reg2196[(2'h2):(2'h2)])));
                    end
                end
              else
                begin
                  if ($unsigned((($unsigned((8'hb0)) ~^ forvar2176[(4'h9):(3'h6)]) ?
                      reg2196 : (^~$signed(forvar2203)))))
                    begin
                      reg2204 <= ((((reg2197 < wire2171) ?
                          reg2185 : (forvar2196 ?
                              reg2199 : wire2175)) > $unsigned({wire2175})) ~^ $unsigned($signed((reg2211 ?
                          reg2192 : reg2189))));
                      reg2205 <= $signed(wire2174);
                      reg2206 <= (~^$unsigned((~|(8'ha2))));
                    end
                  else
                    begin
                      reg2204 <= $signed(reg2205[(1'h1):(1'h0)]);
                      reg2205 <= forvar2208;
                      reg2206 <= $unsigned(reg2205[(2'h3):(2'h3)]);
                      reg2207 <= $signed(reg2209[(4'h9):(4'h9)]);
                    end
                  if (reg2185[(4'hd):(4'hc)])
                    begin
                      reg2208 <= $signed($unsigned($signed(reg2211[(1'h0):(1'h0)])));
                      reg2209 <= (|$unsigned({reg2209[(1'h0):(1'h0)]}));
                      reg2210 <= {reg2178[(3'h4):(1'h0)]};
                    end
                  else
                    begin
                      reg2208 <= reg2188;
                      reg2209 <= reg2197;
                      reg2210 <= (&$signed($signed((+reg2189))));
                    end
                  reg2211 <= ({(reg2200[(3'h6):(1'h1)] > $signed(reg2200))} ?
                      reg2194 : reg2212);
                  for (forvar2212 = (1'h0); (forvar2212 < (1'h1)); forvar2212 = (forvar2212 + (1'h1)))
                    begin
                      reg2213 <= ($unsigned(reg2179) ? reg2194 : (8'ha9));
                      reg2214 <= {$signed($unsigned((~&reg2210)))};
                      reg2215 <= reg2191[(3'h6):(2'h3)];
                      reg2216 <= ($signed($signed((^reg2205))) ^ reg2195[(4'ha):(4'h8)]);
                    end
                end
              if (reg2208[(3'h4):(3'h4)])
                begin
                  for (forvar2217 = (1'h0); (forvar2217 < (1'h0)); forvar2217 = (forvar2217 + (1'h1)))
                    begin
                      reg2218 <= $signed((((8'hb6) ?
                              (reg2179 ? reg2211 : reg2207) : (reg2191 ?
                                  wire2173 : reg2198)) ?
                          (|wire2175) : (~&(reg2215 != forvar2212))));
                      reg2219 <= reg2183[(1'h1):(1'h1)];
                      reg2220 <= (~&{((reg2218 ? (8'ha7) : reg2208) ?
                              reg2192 : {(8'h9d)})});
                    end
                  for (forvar2221 = (1'h0); (forvar2221 < (2'h3)); forvar2221 = (forvar2221 + (1'h1)))
                    begin
                      reg2222 <= (reg2188[(4'h8):(3'h7)] == $unsigned({$unsigned(forvar2176)}));
                    end
                end
              else
                begin
                  reg2217 <= (8'ha1);
                  if ({forvar2197[(3'h7):(3'h7)]})
                    begin
                      reg2218 <= $unsigned(reg2210);
                      reg2219 <= (reg2213[(4'hf):(4'h8)] <<< (forvar2186 & forvar2208[(4'ha):(2'h2)]));
                    end
                  else
                    begin
                      reg2218 <= (8'ha1);
                      reg2219 <= $unsigned($unsigned((~|$unsigned(reg2217))));
                    end
                  reg2220 <= $signed((~($signed(wire2174) ?
                      reg2215 : $unsigned(reg2190))));
                  reg2221 <= $signed(reg2210);
                end
            end
        end
      else
        begin
          for (forvar2180 = (1'h0); (forvar2180 < (2'h2)); forvar2180 = (forvar2180 + (1'h1)))
            begin
              for (forvar2181 = (1'h0); (forvar2181 < (2'h3)); forvar2181 = (forvar2181 + (1'h1)))
                begin
                  if (($signed(reg2217[(2'h2):(1'h0)]) ?
                      reg2195 : $signed({(reg2190 ? reg2189 : reg2208)})))
                    begin
                      reg2182 <= $signed(reg2216[(1'h0):(1'h0)]);
                      reg2183 <= reg2210;
                      reg2184 <= {((8'hb0) * $signed(forvar2184[(2'h3):(2'h3)]))};
                      reg2185 <= (8'hb6);
                    end
                  else
                    begin
                      reg2182 <= {(-(-wire2172[(2'h2):(1'h0)]))};
                    end
                end
            end
          reg2186 <= (((~^((8'ha6) ? reg2207 : forvar2184)) * (reg2204 ?
                  $signed(reg2178) : reg2209[(3'h7):(2'h2)])) ?
              (((reg2198 <<< reg2188) ?
                  ((8'ha4) ?
                      forvar2221 : forvar2217) : $signed(reg2189)) >>> $signed(reg2189)) : ($unsigned($signed(reg2202)) ?
                  (!{reg2215}) : reg2200));
        end
      reg2223 <= reg2191[(2'h3):(2'h2)];
    end
  assign wire2224 = (($unsigned(reg2202[(3'h4):(1'h1)]) ?
                        (^~(!(8'hb2))) : reg2217[(1'h0):(1'h0)]) & {((reg2206 ?
                                reg2214 : (8'h9f)) ?
                            reg2214[(3'h6):(3'h5)] : $unsigned(reg2222))});
  module2225 modinst3111 (wire3110, clk, reg2205, wire2173, forvar2176, reg2195);
  always
    @(posedge clk) begin
      for (forvar3112 = (1'h0); (forvar3112 < (2'h2)); forvar3112 = (forvar3112 + (1'h1)))
        begin
          for (forvar3113 = (1'h0); (forvar3113 < (2'h3)); forvar3113 = (forvar3113 + (1'h1)))
            begin
              if (($unsigned({(^reg2186)}) ?
                  ($signed($signed(forvar2182)) > ($unsigned(reg2193) << $signed(reg2200))) : $unsigned(($unsigned(reg2215) & {forvar2201}))))
                begin
                  reg3114 <= reg2223[(3'h4):(1'h1)];
                  if (((+(reg2209 ?
                      reg2212 : (wire2172 ?
                          reg2193 : reg2189))) >= $signed(((~&reg2184) + $signed(forvar2176)))))
                    begin
                      reg3115 <= (-(+$unsigned(reg2202[(2'h2):(2'h2)])));
                      reg3116 <= forvar3113[(2'h3):(1'h1)];
                      reg3117 <= $signed((~&(^~forvar2221[(1'h0):(1'h0)])));
                      reg3118 <= (~&(wire2170[(4'hc):(1'h1)] >= ((!forvar2197) + (!(8'ha1)))));
                    end
                  else
                    begin
                      reg3115 <= ($unsigned(reg2205[(4'hc):(4'hc)]) <= ($signed(reg2211) == ((reg2221 ?
                              reg2212 : forvar3113) ?
                          $unsigned(reg3115) : $unsigned(reg2204))));
                    end
                  reg3119 <= $unsigned({(reg2223 ?
                          $signed(wire2169) : (!reg3115))});
                end
              else
                begin
                  if ($signed($unsigned(($signed(forvar3112) ?
                      reg2207 : $unsigned(reg2204)))))
                    begin
                      reg3114 <= {$unsigned(($signed(reg2182) ?
                              (forvar2193 ? reg2210 : forvar2212) : reg2220))};
                      reg3115 <= (reg2220 && $signed((+$unsigned(wire2175))));
                    end
                  else
                    begin
                      reg3114 <= (!$signed($signed($unsigned(wire2224))));
                    end
                  if ((((reg2218[(4'ha):(3'h6)] ?
                      reg2191 : forvar3112[(3'h7):(3'h6)]) < $signed($unsigned(reg2199))) || wire2171))
                    begin
                      reg3116 <= $unsigned(reg2213);
                      reg3117 <= forvar2182;
                      reg3118 <= (($signed($signed(reg2178)) + (!((8'haf) ?
                              reg2178 : reg2205))) ?
                          {((reg2185 ?
                                  forvar2184 : reg2223) == (~&reg2197))} : (wire2174[(3'h5):(3'h4)] <= (forvar2181 ?
                              reg2216 : (reg2192 & reg2206))));
                    end
                  else
                    begin
                      reg3116 <= (8'ha8);
                      reg3117 <= reg2178[(1'h0):(1'h0)];
                      reg3118 <= (~(~^((^forvar2212) && (reg2195 ?
                          reg3118 : forvar2208))));
                    end
                  if (wire2170[(4'ha):(2'h3)])
                    begin
                      reg3119 <= ({{$signed(reg2197)}} <<< ((&$signed(forvar2221)) ?
                          ($signed(forvar2221) ?
                              (8'ha7) : reg2222[(2'h2):(1'h1)]) : $signed((forvar2217 ?
                              reg2191 : reg2212))));
                      reg3120 <= (((^~$unsigned(forvar2184)) * wire2174[(1'h0):(1'h0)]) < (~&forvar2212[(3'h4):(1'h0)]));
                      reg3121 <= (reg2196 ?
                          $signed(({wire2224} ?
                              (reg2223 & reg2195) : $unsigned(reg2193))) : $unsigned(reg2207[(2'h3):(2'h3)]));
                      reg3122 <= (reg2181[(1'h1):(1'h1)] >>> ({(^reg2217)} << (^(wire2175 + reg2213))));
                    end
                  else
                    begin
                      reg3119 <= (({((8'ha3) - reg2208)} ?
                              ($signed(reg3121) >= (~^(8'hb3))) : (|forvar2180[(2'h2):(1'h1)])) ?
                          {($unsigned(reg2217) != (|(8'hba)))} : $signed({(wire2174 || reg2184)}));
                      reg3120 <= $signed({{$signed((8'hb8))}});
                      reg3121 <= ($signed(reg2193[(3'h4):(2'h2)]) | (($unsigned(reg3120) ?
                          $signed(forvar2201) : $unsigned((8'ha4))) <= $unsigned((^reg2210))));
                    end
                end
            end
          for (forvar3123 = (1'h0); (forvar3123 < (1'h1)); forvar3123 = (forvar3123 + (1'h1)))
            begin
              for (forvar3124 = (1'h0); (forvar3124 < (2'h2)); forvar3124 = (forvar3124 + (1'h1)))
                begin
                  for (forvar3125 = (1'h0); (forvar3125 < (1'h0)); forvar3125 = (forvar3125 + (1'h1)))
                    begin
                      reg3126 <= $signed((({forvar2208} ?
                          (reg2217 ?
                              forvar2176 : reg2199) : reg3121) << ((reg2219 >> reg2204) > (reg2190 <<< reg2190))));
                    end
                end
              for (forvar3127 = (1'h0); (forvar3127 < (1'h1)); forvar3127 = (forvar3127 + (1'h1)))
                begin
                  for (forvar3128 = (1'h0); (forvar3128 < (1'h1)); forvar3128 = (forvar3128 + (1'h1)))
                    begin
                      reg3129 <= (($signed($unsigned((8'hab))) ?
                              (reg2179[(1'h1):(1'h0)] <<< (forvar3125 ?
                                  (8'haf) : forvar2181)) : wire2170) ?
                          {$unsigned(forvar3112[(3'h7):(1'h1)])} : reg3126[(1'h0):(1'h0)]);
                      reg3130 <= (($unsigned((reg2193 ? reg2215 : wire2175)) ?
                              reg2200[(2'h2):(2'h2)] : ((reg2200 ?
                                      wire2170 : reg2195) ?
                                  (reg2186 & wire2173) : {wire2170})) ?
                          reg2188[(3'h5):(3'h5)] : ((forvar2176 ?
                              $unsigned(wire2224) : (reg3126 >>> (8'h9e))) <<< $signed((+(8'haf)))));
                    end
                  if (reg2223)
                    begin
                      reg3131 <= reg2193;
                      reg3132 <= $unsigned($unsigned(forvar2184[(2'h3):(1'h1)]));
                      reg3133 <= (((~^((8'hae) - (8'hb2))) ?
                              $unsigned(reg2192[(1'h1):(1'h1)]) : (!wire2169[(2'h3):(2'h3)])) ?
                          {{(8'had)}} : $signed($unsigned($signed(reg2222))));
                    end
                  else
                    begin
                      reg3131 <= (~{(reg2220[(3'h6):(3'h5)] && {(8'ha1)})});
                      reg3132 <= $unsigned($unsigned((~|reg2210)));
                      reg3133 <= $signed(reg3121[(4'he):(3'h5)]);
                      reg3134 <= (wire2175 != (((reg3115 ^~ (8'h9f)) ?
                          $signed(reg2221) : $unsigned(reg2216)) - $signed((8'ha8))));
                    end
                  if ({$signed({$signed(forvar2186)})})
                    begin
                      reg3135 <= reg2189;
                      reg3136 <= reg2211;
                    end
                  else
                    begin
                      reg3135 <= $signed($unsigned({wire2224}));
                      reg3136 <= (reg2191[(3'h4):(1'h0)] ?
                          $unsigned(reg2177[(1'h0):(1'h0)]) : (8'h9e));
                      reg3137 <= (~forvar2193[(3'h4):(3'h4)]);
                      reg3138 <= (&reg3118);
                    end
                  reg3139 <= reg2196;
                end
              if ($unsigned((reg3139 ?
                  ($signed(reg2181) ?
                      {forvar2203} : $signed((8'haf))) : ($unsigned(wire2169) * forvar3112))))
                begin
                  reg3140 <= ({$signed(((8'hb3) ^~ (8'had)))} ?
                      (((reg2188 + reg2221) >= (~^forvar3128)) ?
                          forvar2212[(1'h1):(1'h1)] : (^$signed(reg3131))) : (^$unsigned((reg2199 ^ forvar2184))));
                end
              else
                begin
                  for (forvar3140 = (1'h0); (forvar3140 < (1'h1)); forvar3140 = (forvar3140 + (1'h1)))
                    begin
                      reg3141 <= reg2220[(3'h7):(2'h2)];
                    end
                end
              if ($signed($unsigned(($unsigned(reg3126) && ((8'hb9) ?
                  forvar3125 : (8'hac))))))
                begin
                  for (forvar3142 = (1'h0); (forvar3142 < (2'h2)); forvar3142 = (forvar3142 + (1'h1)))
                    begin
                      reg3143 <= reg2178;
                      reg3144 <= ({forvar3142[(3'h5):(1'h1)]} ?
                          $signed(forvar3112[(3'h7):(3'h7)]) : (^~($unsigned(wire2171) ?
                              (reg2219 ?
                                  forvar2197 : reg2207) : ((8'hb3) | (8'h9f)))));
                      reg3145 <= ((((reg3143 <<< reg2199) ?
                              (reg3138 <= (8'hb2)) : reg2189) != (reg2212[(4'hb):(1'h1)] >= reg2210[(1'h0):(1'h0)])) ?
                          {{forvar3113[(1'h0):(1'h0)]}} : reg2184[(1'h1):(1'h1)]);
                      reg3146 <= ((((reg2210 ? reg2195 : forvar3142) ?
                          ((8'hb7) ?
                              reg2222 : forvar3128) : (-forvar2217)) | reg2218[(3'h7):(3'h7)]) + reg3141[(2'h2):(2'h2)]);
                    end
                  if ($unsigned(reg3116[(3'h7):(1'h0)]))
                    begin
                      reg3147 <= reg2197;
                      reg3148 <= (^~$unsigned(reg3144[(3'h4):(1'h0)]));
                    end
                  else
                    begin
                      reg3147 <= (~&reg3115[(1'h0):(1'h0)]);
                      reg3148 <= forvar3127;
                      reg3149 <= (!$signed($unsigned((forvar3124 <<< reg2194))));
                      reg3150 <= (-wire2224);
                    end
                  for (forvar3151 = (1'h0); (forvar3151 < (1'h1)); forvar3151 = (forvar3151 + (1'h1)))
                    begin
                      reg3152 <= {$unsigned($signed(forvar2201))};
                      reg3153 <= $signed($unsigned(reg3140[(3'h5):(2'h3)]));
                      reg3154 <= (((!$signed(reg3115)) >> (8'ha1)) ?
                          $unsigned($signed((&reg3144))) : {reg2184});
                    end
                  if ((~&$unsigned(((reg3138 << reg3119) >= (~&(8'ha5))))))
                    begin
                      reg3155 <= (~reg3116);
                      reg3156 <= $unsigned(($signed({forvar3113}) == ($unsigned(wire2173) ?
                          (8'hba) : (-reg2193))));
                      reg3157 <= forvar2181[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3155 <= (|reg2207);
                      reg3156 <= ($signed($signed((reg2220 ?
                          reg3130 : forvar3140))) - $unsigned($signed((reg3116 & reg2202))));
                      reg3157 <= forvar2176;
                      reg3158 <= {(&reg3114[(3'h4):(1'h0)])};
                    end
                end
              else
                begin
                  if (((|$unsigned($signed(reg3135))) && $unsigned((-(reg2198 ?
                      forvar2208 : reg2219)))))
                    begin
                      reg3142 <= $signed({$unsigned(wire2174)});
                      reg3143 <= (-$signed(reg2216));
                      reg3144 <= (($unsigned((reg2184 ^~ (8'hb0))) - $unsigned({reg3116})) ?
                          reg2219 : (reg2199[(1'h0):(1'h0)] ?
                              $unsigned((reg3118 ?
                                  reg2186 : reg3144)) : (~&$signed(reg2188))));
                      reg3145 <= (^~{$unsigned((reg2189 ^ reg3144))});
                    end
                  else
                    begin
                      reg3142 <= $unsigned(($signed($unsigned(reg2206)) ?
                          ((reg3115 ~^ reg3132) ?
                              reg2200[(1'h1):(1'h1)] : $unsigned((8'ha2))) : $signed({reg2216})));
                      reg3143 <= wire3110;
                      reg3144 <= $unsigned(reg3141[(4'hd):(4'hd)]);
                      reg3145 <= reg3142[(4'ha):(2'h3)];
                    end
                  for (forvar3146 = (1'h0); (forvar3146 < (1'h0)); forvar3146 = (forvar3146 + (1'h1)))
                    begin
                      reg3147 <= (reg2186 ?
                          (&(^~(reg3148 <<< reg3156))) : $signed(reg3139[(3'h7):(3'h6)]));
                      reg3148 <= $signed(reg3145);
                    end
                  if ((reg2222 ^~ reg3145[(4'hb):(4'h8)]))
                    begin
                      reg3149 <= (~&reg3136);
                      reg3150 <= reg2177[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg3149 <= $unsigned(((~reg3119) ?
                          ((~^reg2198) ? reg2216 : (^~reg2190)) : reg2211));
                      reg3150 <= (wire2171 & reg3132);
                      reg3151 <= ($signed(((!reg3156) ?
                          (reg2192 ?
                              reg3130 : reg2192) : $signed((8'ha2)))) <= {$signed(((8'ha1) >= reg2216))});
                    end
                  for (forvar3152 = (1'h0); (forvar3152 < (2'h2)); forvar3152 = (forvar3152 + (1'h1)))
                    begin
                      reg3153 <= ((|{$signed(reg2212)}) != reg2197[(2'h3):(2'h2)]);
                    end
                end
            end
        end
      for (forvar3159 = (1'h0); (forvar3159 < (1'h0)); forvar3159 = (forvar3159 + (1'h1)))
        begin
          reg3160 <= $unsigned(({$signed(reg3114)} <<< forvar2212[(3'h4):(1'h0)]));
        end
      reg3161 <= {($signed((^~wire2175)) > $signed((forvar2187 ?
              reg3156 : reg2179)))};
      for (forvar3162 = (1'h0); (forvar3162 < (2'h2)); forvar3162 = (forvar3162 + (1'h1)))
        begin
          for (forvar3163 = (1'h0); (forvar3163 < (1'h0)); forvar3163 = (forvar3163 + (1'h1)))
            begin
              if (($signed(((8'hb5) ~^ (reg3122 ? reg3139 : reg3153))) ?
                  forvar2221 : (!$unsigned($signed(reg2185)))))
                begin
                  reg3164 <= (forvar3152[(4'h8):(3'h7)] >= $unsigned($signed(reg3153)));
                end
              else
                begin
                  reg3164 <= $unsigned(wire2170);
                  reg3165 <= ({(8'hb3)} ?
                      reg2205[(4'hd):(4'hb)] : $signed($unsigned(((8'hb1) || wire2169))));
                  if (reg2191[(3'h7):(3'h6)])
                    begin
                      reg3166 <= $unsigned((~&(^forvar2201[(3'h7):(1'h0)])));
                      reg3167 <= $unsigned($signed((-reg3150[(1'h0):(1'h0)])));
                      reg3168 <= wire2174[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3166 <= (($signed((wire2171 ^~ forvar3113)) ?
                              (((8'hb0) ? reg3119 : forvar2212) ?
                                  (+reg2221) : (reg2189 ?
                                      reg3131 : reg3158)) : wire2224[(1'h0):(1'h0)]) ?
                          ($unsigned(wire2174[(3'h4):(1'h1)]) != $unsigned({reg2208})) : (+$signed((reg3143 ^ (8'ha6)))));
                      reg3167 <= reg3120;
                    end
                end
              if ($signed($signed(({reg3115} >> (|reg3119)))))
                begin
                  if ($unsigned(((((8'hb6) <= (8'ha0)) ?
                          (reg2202 <<< forvar3162) : (forvar2193 < wire2175)) ?
                      reg2189[(1'h1):(1'h0)] : wire2171[(4'h9):(3'h7)])))
                    begin
                      reg3169 <= wire2171;
                    end
                  else
                    begin
                      reg3169 <= $unsigned($signed(($unsigned(reg3156) <<< $unsigned(forvar2197))));
                      reg3170 <= $unsigned((-(((8'h9e) ? (8'h9c) : forvar2193) ?
                          reg3160[(1'h1):(1'h1)] : (forvar2212 || reg2195))));
                    end
                end
              else
                begin
                  if (({(forvar3127 ^~ $unsigned(reg2218))} ?
                      (reg3129[(1'h1):(1'h1)] ?
                          (reg3129 ?
                              {reg2182} : $signed(forvar2186)) : (&forvar2201)) : $signed(forvar2187)))
                    begin
                      reg3169 <= reg3135;
                    end
                  else
                    begin
                      reg3169 <= ($signed(reg2183) ?
                          $signed(forvar3127) : (^(~|$unsigned(reg3167))));
                      reg3170 <= ((^~{$signed(wire2169)}) | (((reg2214 ^ reg3150) < forvar3151) & (((8'hb9) | wire2169) << $signed(reg3116))));
                      reg3171 <= {(~|(!reg2213))};
                    end
                  for (forvar3172 = (1'h0); (forvar3172 < (2'h3)); forvar3172 = (forvar3172 + (1'h1)))
                    begin
                      reg3173 <= (((reg2184[(1'h0):(1'h0)] * reg2186[(4'ha):(3'h4)]) ?
                              ($unsigned(reg3116) <<< {forvar3152}) : ($signed(reg2192) * reg3139)) ?
                          reg3154[(1'h1):(1'h0)] : wire2175[(4'h8):(3'h6)]);
                    end
                  for (forvar3174 = (1'h0); (forvar3174 < (1'h1)); forvar3174 = (forvar3174 + (1'h1)))
                    begin
                      reg3175 <= (~&($signed((reg3114 ? reg2195 : reg3143)) ?
                          forvar2193[(4'h9):(3'h6)] : $unsigned($signed(forvar3152))));
                      reg3176 <= ((!(~|(|reg2196))) - $signed(reg2223[(2'h2):(2'h2)]));
                      reg3177 <= ($unsigned($unsigned(reg3138[(3'h7):(3'h5)])) - forvar3151[(2'h3):(2'h2)]);
                    end
                  for (forvar3178 = (1'h0); (forvar3178 < (1'h0)); forvar3178 = (forvar3178 + (1'h1)))
                    begin
                      reg3179 <= ({forvar2196[(4'hd):(3'h6)]} ?
                          $signed((8'hab)) : $unsigned(reg3142[(3'h5):(3'h5)]));
                      reg3180 <= reg3154;
                    end
                end
              for (forvar3181 = (1'h0); (forvar3181 < (1'h1)); forvar3181 = (forvar3181 + (1'h1)))
                begin
                  if ((reg3121[(5'h10):(4'he)] * $unsigned((forvar3142[(3'h5):(1'h1)] + ((8'ha4) ?
                      forvar3159 : forvar3163)))))
                    begin
                      reg3182 <= (~((!$unsigned(wire2170)) ?
                          ($unsigned(reg2217) ?
                              (reg2208 ?
                                  forvar2212 : reg3140) : $unsigned(forvar2203)) : (reg3141 ?
                              $signed(reg2218) : reg3153)));
                    end
                  else
                    begin
                      reg3182 <= reg3165[(3'h4):(1'h1)];
                      reg3183 <= reg3157;
                      reg3184 <= $signed((&reg3138));
                    end
                  if ($unsigned(reg2202))
                    begin
                      reg3185 <= $unsigned((forvar3112 != {{reg3132}}));
                      reg3186 <= (^reg3161[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg3185 <= {$unsigned(reg3143[(3'h7):(1'h0)])};
                    end
                  if ({((-$signed(forvar2197)) == (~|(reg2216 ?
                          wire2174 : (8'ha9))))})
                    begin
                      reg3187 <= {reg3122};
                      reg3188 <= (forvar3162 ?
                          reg2221[(2'h3):(1'h1)] : reg2216);
                    end
                  else
                    begin
                      reg3187 <= ((reg3180[(4'h8):(2'h2)] ?
                              (^~reg3168) : (~&reg3169)) ?
                          {($signed(reg3188) - (reg3183 ?
                                  reg3131 : (8'had)))} : (~^$unsigned(reg3116[(4'he):(3'h4)])));
                      reg3188 <= reg3182;
                      reg3189 <= (~^(~(&$unsigned(reg2211))));
                      reg3190 <= (8'hb5);
                    end
                end
              for (forvar3191 = (1'h0); (forvar3191 < (1'h0)); forvar3191 = (forvar3191 + (1'h1)))
                begin
                  if (((reg3145[(2'h3):(2'h3)] == {$signed(reg2183)}) < reg3115[(3'h7):(2'h3)]))
                    begin
                      reg3192 <= reg3166;
                      reg3193 <= reg3118[(4'h8):(4'h8)];
                      reg3194 <= reg2193[(3'h4):(1'h0)];
                      reg3195 <= forvar3163[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg3192 <= {forvar3174[(3'h7):(2'h2)]};
                    end
                  if (reg3151[(3'h7):(1'h1)])
                    begin
                      reg3196 <= reg3126;
                      reg3197 <= reg2207;
                      reg3198 <= $unsigned({(-reg3186[(1'h1):(1'h0)])});
                    end
                  else
                    begin
                      reg3196 <= $unsigned($signed($unsigned($unsigned((8'h9f)))));
                      reg3197 <= reg3131[(3'h4):(1'h1)];
                      reg3198 <= forvar3112[(4'h9):(3'h4)];
                    end
                end
            end
          if (forvar3178)
            begin
              if ((&$signed(((!reg2202) ?
                  (~&(8'ha6)) : forvar3191[(3'h4):(1'h1)]))))
                begin
                  for (forvar3199 = (1'h0); (forvar3199 < (2'h2)); forvar3199 = (forvar3199 + (1'h1)))
                    begin
                      reg3200 <= (((8'h9e) & $unsigned(forvar2212[(3'h4):(2'h2)])) >>> reg3170[(2'h2):(1'h0)]);
                      reg3201 <= reg3147;
                      reg3202 <= (reg3168 ?
                          forvar3152[(3'h4):(1'h1)] : forvar3162[(2'h2):(2'h2)]);
                    end
                  for (forvar3203 = (1'h0); (forvar3203 < (2'h3)); forvar3203 = (forvar3203 + (1'h1)))
                    begin
                      reg3204 <= reg3185;
                      reg3205 <= (~|(forvar2212[(1'h0):(1'h0)] && {$signed(forvar3152)}));
                    end
                end
              else
                begin
                  for (forvar3199 = (1'h0); (forvar3199 < (1'h0)); forvar3199 = (forvar3199 + (1'h1)))
                    begin
                      reg3200 <= $unsigned((~^((~|forvar2217) ?
                          (reg3155 ?
                              reg3144 : forvar3163) : $signed(forvar3191))));
                    end
                  for (forvar3201 = (1'h0); (forvar3201 < (1'h1)); forvar3201 = (forvar3201 + (1'h1)))
                    begin
                      reg3202 <= forvar2187;
                      reg3203 <= reg3179;
                    end
                  for (forvar3204 = (1'h0); (forvar3204 < (1'h0)); forvar3204 = (forvar3204 + (1'h1)))
                    begin
                      reg3205 <= ((reg3168[(1'h1):(1'h0)] - ((|reg3160) ?
                              $unsigned(reg3166) : $unsigned(reg3202))) ?
                          ($signed((^reg3116)) ?
                              (8'hb7) : reg3182[(2'h2):(1'h1)]) : $unsigned(forvar2212[(1'h1):(1'h0)]));
                      reg3206 <= $unsigned(reg3139);
                      reg3207 <= forvar2208[(3'h4):(1'h1)];
                    end
                  if (reg3170[(2'h2):(2'h2)])
                    begin
                      reg3208 <= {$signed({(reg2178 - forvar2182)})};
                      reg3209 <= (&$signed((reg3115 | (8'ha4))));
                    end
                  else
                    begin
                      reg3208 <= {reg3203};
                      reg3209 <= $unsigned(reg2188[(2'h3):(2'h2)]);
                      reg3210 <= {$signed({{reg3193}})};
                      reg3211 <= {(&(~^forvar2217[(4'h8):(3'h5)]))};
                    end
                end
              if ($signed(reg2186))
                begin
                  for (forvar3212 = (1'h0); (forvar3212 < (1'h0)); forvar3212 = (forvar3212 + (1'h1)))
                    begin
                      reg3213 <= (reg3141[(3'h5):(2'h3)] != $signed((reg2219[(3'h7):(1'h0)] >> $unsigned(reg2192))));
                      reg3214 <= (reg3154[(2'h2):(2'h2)] ?
                          (({reg2202} >= $signed(forvar3203)) && ($unsigned(reg2193) != (forvar2201 > reg3149))) : ((+(reg2181 ?
                              reg2222 : reg2217)) ^~ (8'ha3)));
                      reg3215 <= {$unsigned($unsigned((~&forvar3113)))};
                      reg3216 <= ($signed($unsigned($unsigned(reg3188))) ^ forvar3127[(3'h5):(1'h0)]);
                    end
                  for (forvar3217 = (1'h0); (forvar3217 < (2'h2)); forvar3217 = (forvar3217 + (1'h1)))
                    begin
                      reg3218 <= (8'haf);
                      reg3219 <= reg2198[(2'h3):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar3212 = (1'h0); (forvar3212 < (2'h2)); forvar3212 = (forvar3212 + (1'h1)))
                    begin
                      reg3213 <= reg3120;
                    end
                  reg3214 <= $unsigned(($signed(forvar3159) ?
                      ($signed(reg3147) == reg3138) : $signed((~reg2196))));
                  if ((8'hb9))
                    begin
                      reg3215 <= (+(~^reg3132[(1'h0):(1'h0)]));
                      reg3216 <= (~|forvar2197);
                      reg3217 <= {reg2220};
                    end
                  else
                    begin
                      reg3215 <= forvar3123[(1'h1):(1'h1)];
                      reg3216 <= (reg2194 ? reg2216 : forvar3203);
                      reg3217 <= reg3142;
                      reg3218 <= (($unsigned(reg3202[(2'h2):(1'h1)]) ?
                              reg3194[(1'h0):(1'h0)] : (!(~&reg3179))) ?
                          reg3138[(1'h1):(1'h1)] : ((8'hb3) < $signed($unsigned(reg3196))));
                    end
                end
              for (forvar3220 = (1'h0); (forvar3220 < (2'h3)); forvar3220 = (forvar3220 + (1'h1)))
                begin
                  for (forvar3221 = (1'h0); (forvar3221 < (1'h1)); forvar3221 = (forvar3221 + (1'h1)))
                    begin
                      reg3222 <= $signed($signed(reg2220[(1'h1):(1'h0)]));
                      reg3223 <= $unsigned((reg3142[(2'h2):(2'h2)] - $signed($unsigned(reg3152))));
                    end
                end
            end
          else
            begin
              if (($unsigned($unsigned(forvar3212)) ?
                  $unsigned($signed((reg2190 ?
                      reg2178 : forvar3152))) : reg2193))
                begin
                  if (reg3184[(2'h2):(2'h2)])
                    begin
                      reg3199 <= (8'hb1);
                      reg3200 <= $unsigned($signed((+reg2188)));
                      reg3201 <= $unsigned(((reg3205[(3'h4):(2'h2)] | (reg3194 * forvar3191)) > $unsigned((^~(8'ha1)))));
                      reg3202 <= $signed(((8'hb2) ?
                          {$signed(reg3184)} : $signed($unsigned(forvar3174))));
                    end
                  else
                    begin
                      reg3199 <= $unsigned(wire2224);
                      reg3200 <= (~^$signed(reg3195[(1'h1):(1'h0)]));
                      reg3201 <= reg3177[(1'h1):(1'h1)];
                      reg3202 <= ((wire2170 >= ((reg3167 - reg3190) ?
                          $unsigned(reg3203) : (reg3145 ?
                              reg3194 : reg2207))) < (&reg2218));
                    end
                end
              else
                begin
                  for (forvar3199 = (1'h0); (forvar3199 < (2'h3)); forvar3199 = (forvar3199 + (1'h1)))
                    begin
                      reg3200 <= $signed(reg3198[(2'h3):(1'h0)]);
                      reg3201 <= forvar2176[(1'h1):(1'h0)];
                      reg3202 <= ($signed($unsigned(((8'haf) <<< forvar3203))) ?
                          (^((|reg3122) ?
                              (reg2218 <= reg3156) : $signed((8'h9d)))) : forvar2196[(2'h2):(1'h1)]);
                    end
                  if ($unsigned((^{{reg2189}})))
                    begin
                      reg3203 <= $signed($unsigned((&reg3213[(1'h1):(1'h0)])));
                      reg3204 <= $signed({reg3198});
                    end
                  else
                    begin
                      reg3203 <= {{(!$signed(forvar2201))}};
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar3224 = (1'h0); (forvar3224 < (1'h0)); forvar3224 = (forvar3224 + (1'h1)))
        begin
          for (forvar3225 = (1'h0); (forvar3225 < (2'h3)); forvar3225 = (forvar3225 + (1'h1)))
            begin
              for (forvar3226 = (1'h0); (forvar3226 < (1'h0)); forvar3226 = (forvar3226 + (1'h1)))
                begin
                  if ((reg3211[(3'h5):(2'h3)] != reg2214[(1'h1):(1'h0)]))
                    begin
                      reg3227 <= {(((forvar3163 * reg3135) ?
                              forvar3127 : {(8'ha4)}) || $signed(reg3213[(3'h4):(1'h1)]))};
                    end
                  else
                    begin
                      reg3227 <= reg2191;
                      reg3228 <= reg2217;
                      reg3229 <= forvar2221;
                      reg3230 <= ($signed(((reg3114 ? (8'ha9) : reg3152) ?
                          (8'hb7) : ((8'ha1) ^~ forvar3174))) * reg2213);
                    end
                  for (forvar3231 = (1'h0); (forvar3231 < (2'h2)); forvar3231 = (forvar3231 + (1'h1)))
                    begin
                      reg3232 <= reg3148;
                    end
                  if ($signed((($unsigned(reg3131) > ((8'ha9) >> reg3158)) ^ forvar2203)))
                    begin
                      reg3233 <= forvar3162;
                      reg3234 <= ($signed((^~reg3130)) ?
                          reg2218 : reg2221[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg3233 <= reg2193;
                      reg3234 <= wire3110[(2'h3):(2'h3)];
                      reg3235 <= {$signed(reg2189)};
                      reg3236 <= (8'hb7);
                    end
                  if (($signed((8'ha6)) == {(8'hb1)}))
                    begin
                      reg3237 <= forvar3151[(1'h1):(1'h0)];
                      reg3238 <= (reg3130[(3'h7):(3'h5)] == ((~^(forvar3151 ?
                          forvar3174 : reg3229)) << $unsigned($unsigned((8'hb9)))));
                      reg3239 <= (8'hba);
                      reg3240 <= (~((|reg3164[(2'h2):(1'h0)]) == reg3214[(4'hb):(4'ha)]));
                    end
                  else
                    begin
                      reg3237 <= (~|$signed(reg3154[(2'h3):(2'h3)]));
                    end
                end
            end
        end
      reg3241 <= ((8'hac) ?
          (((reg2223 > reg2222) ?
                  $unsigned(forvar2187) : (reg3161 + forvar2180)) ?
              (~|(wire2171 ?
                  reg3222 : reg2215)) : $signed(reg3165[(2'h2):(1'h1)])) : (&(-reg3187[(1'h0):(1'h0)])));
      for (forvar3242 = (1'h0); (forvar3242 < (2'h2)); forvar3242 = (forvar3242 + (1'h1)))
        begin
          reg3243 <= $unsigned($signed(reg3232[(2'h3):(1'h0)]));
          if ({(8'ha6)})
            begin
              if (reg3199)
                begin
                  for (forvar3244 = (1'h0); (forvar3244 < (1'h1)); forvar3244 = (forvar3244 + (1'h1)))
                    begin
                      reg3245 <= $unsigned({((forvar2180 ~^ reg2223) ?
                              $unsigned(forvar2203) : (^reg2194))});
                      reg3246 <= wire2170;
                      reg3247 <= (!$signed(forvar2197));
                    end
                  if (reg3246[(2'h3):(1'h1)])
                    begin
                      reg3248 <= {reg3138[(1'h0):(1'h0)]};
                      reg3249 <= reg3157;
                      reg3250 <= ($unsigned($unsigned((reg3232 <<< forvar2181))) ?
                          $unsigned((~reg3116)) : $unsigned($signed((^~reg2219))));
                      reg3251 <= ($signed(reg3234) <<< ((^(reg3187 ^ reg3133)) ?
                          ($unsigned(reg3248) << $signed(forvar3174)) : ($signed(reg2196) < {reg3122})));
                    end
                  else
                    begin
                      reg3248 <= reg2221[(1'h0):(1'h0)];
                      reg3249 <= $unsigned(((8'hb9) <= $signed((forvar3162 >= reg3116))));
                      reg3250 <= wire2224;
                    end
                  for (forvar3252 = (1'h0); (forvar3252 < (1'h1)); forvar3252 = (forvar3252 + (1'h1)))
                    begin
                      reg3253 <= (~|(^~{{(8'hae)}}));
                      reg3254 <= {$signed(({(8'hb5)} ?
                              {forvar2196} : (reg2221 < reg2204)))};
                      reg3255 <= $signed($unsigned(forvar3112));
                      reg3256 <= (8'ha3);
                    end
                  for (forvar3257 = (1'h0); (forvar3257 < (1'h0)); forvar3257 = (forvar3257 + (1'h1)))
                    begin
                      reg3258 <= (($signed(reg2194[(3'h6):(3'h4)]) ?
                          $unsigned($unsigned(reg3137)) : $unsigned((|reg3196))) < (($unsigned(forvar2193) ?
                              forvar2201[(1'h1):(1'h0)] : {forvar3163}) ?
                          (-forvar3174[(4'hb):(1'h0)]) : (forvar3252 * reg3134)));
                    end
                end
              else
                begin
                  if ({((~^(|reg2213)) ?
                          $signed((~forvar2187)) : forvar2180[(1'h1):(1'h0)])})
                    begin
                      reg3244 <= (!({$unsigned(reg3197)} << forvar3162[(3'h7):(3'h4)]));
                      reg3245 <= (forvar3174 ?
                          (((reg3228 ^~ reg3156) ^~ (forvar3204 >> reg3177)) > {(reg3228 ?
                                  reg3170 : reg3216)}) : $signed((-(reg3146 != reg2215))));
                      reg3246 <= $signed((!reg2188));
                    end
                  else
                    begin
                      reg3244 <= $unsigned((reg3160[(1'h1):(1'h0)] ?
                          {((8'hac) ?
                                  (8'ha7) : reg3183)} : reg3227[(1'h0):(1'h0)]));
                      reg3245 <= (|$signed($unsigned({reg3218})));
                    end
                  if (forvar3123[(3'h7):(3'h6)])
                    begin
                      reg3247 <= (reg3216[(4'ha):(3'h6)] ?
                          forvar3231[(4'h8):(3'h4)] : (^~({(8'hab)} ?
                              $signed(forvar3152) : reg2207[(3'h4):(3'h4)])));
                      reg3248 <= {$signed(reg3240)};
                    end
                  else
                    begin
                      reg3247 <= reg3188;
                      reg3248 <= reg3173;
                      reg3249 <= $unsigned($unsigned(reg3165[(1'h0):(1'h0)]));
                    end
                  reg3250 <= $unsigned(forvar2187);
                end
              for (forvar3259 = (1'h0); (forvar3259 < (2'h2)); forvar3259 = (forvar3259 + (1'h1)))
                begin
                  reg3260 <= ((!$signed(reg3246)) ^~ reg3179[(4'he):(4'h9)]);
                  reg3261 <= (-(|{$unsigned(reg2205)}));
                  if ((((forvar3124[(2'h3):(1'h0)] >> (reg3192 ?
                          reg3160 : forvar2187)) ?
                      forvar3163[(3'h7):(3'h4)] : $signed(forvar2193)) && (reg3214[(4'ha):(4'ha)] ?
                      $unsigned($unsigned(forvar3231)) : {(reg3215 ^~ reg2210)})))
                    begin
                      reg3262 <= ((($unsigned(reg2192) + reg2206[(4'h8):(3'h6)]) >= {((8'haf) ?
                                  (8'hb2) : forvar2193)}) ?
                          reg3136[(3'h5):(2'h3)] : {reg2200[(2'h2):(1'h1)]});
                    end
                  else
                    begin
                      reg3262 <= ($signed(reg2189) ?
                          (+$unsigned($signed(reg3133))) : (~^forvar2184[(1'h0):(1'h0)]));
                    end
                end
              if (reg3173[(4'h8):(4'h8)])
                begin
                  reg3263 <= reg2195;
                  reg3264 <= ($unsigned(forvar2181) <<< (|(8'hb6)));
                end
              else
                begin
                  for (forvar3263 = (1'h0); (forvar3263 < (1'h1)); forvar3263 = (forvar3263 + (1'h1)))
                    begin
                      reg3264 <= (reg3248[(1'h0):(1'h0)] ?
                          $unsigned((reg3118[(4'h9):(3'h4)] ?
                              (reg2212 & reg2219) : (reg3215 + reg3193))) : reg2197);
                      reg3265 <= reg3251[(3'h4):(1'h1)];
                      reg3266 <= $unsigned((reg3193[(3'h5):(1'h0)] == $signed((reg3167 ?
                          (8'hb4) : reg2217))));
                    end
                end
            end
          else
            begin
              for (forvar3244 = (1'h0); (forvar3244 < (1'h1)); forvar3244 = (forvar3244 + (1'h1)))
                begin
                  for (forvar3245 = (1'h0); (forvar3245 < (2'h2)); forvar3245 = (forvar3245 + (1'h1)))
                    begin
                      reg3246 <= ((^~((forvar2208 ? (8'hba) : reg3158) ?
                              $unsigned(reg3192) : reg3176)) ?
                          $signed((((8'ha5) == reg3228) & $signed(reg3188))) : $unsigned($unsigned($signed(reg2205))));
                      reg3247 <= {{reg3208}};
                    end
                  for (forvar3248 = (1'h0); (forvar3248 < (2'h3)); forvar3248 = (forvar3248 + (1'h1)))
                    begin
                      reg3249 <= reg3209[(2'h2):(1'h0)];
                      reg3250 <= reg3210[(3'h5):(2'h3)];
                      reg3251 <= {reg2220};
                    end
                  if (reg3149[(2'h3):(2'h2)])
                    begin
                      reg3252 <= {$unsigned(reg3183)};
                      reg3253 <= {(^~$unsigned(reg2177[(2'h3):(1'h1)]))};
                      reg3254 <= $unsigned((forvar2182[(3'h5):(1'h1)] && $unsigned(reg3149)));
                    end
                  else
                    begin
                      reg3252 <= ((($unsigned(reg2210) ?
                                  $unsigned(reg3114) : $unsigned(reg3233)) ?
                              reg2222[(1'h1):(1'h1)] : $signed(reg3150)) ?
                          $signed(forvar3191) : forvar2193);
                      reg3253 <= $unsigned($unsigned(reg3222));
                      reg3254 <= ((^~{(^reg3118)}) ?
                          (&$unsigned(((8'h9e) ?
                              forvar3127 : (8'hb3)))) : $unsigned(((|reg2207) ?
                              {reg3251} : (reg2218 ? reg3247 : reg2219))));
                    end
                end
            end
          reg3267 <= reg2197;
        end
      for (forvar3268 = (1'h0); (forvar3268 < (1'h1)); forvar3268 = (forvar3268 + (1'h1)))
        begin
          if ($unsigned(forvar3128[(1'h1):(1'h0)]))
            begin
              for (forvar3269 = (1'h0); (forvar3269 < (1'h1)); forvar3269 = (forvar3269 + (1'h1)))
                begin
                  if ($unsigned($unsigned(((forvar2193 >>> (8'hba)) ^ (8'hb3)))))
                    begin
                      reg3270 <= $unsigned(reg2191[(3'h6):(3'h6)]);
                    end
                  else
                    begin
                      reg3270 <= $unsigned((~|wire2224));
                      reg3271 <= reg2199[(2'h2):(1'h0)];
                    end
                  if ($unsigned(((forvar2193 ? $unsigned(reg2218) : wire2170) ?
                      ((8'hb2) ?
                          $unsigned(reg3240) : $unsigned(wire2172)) : $signed($signed(reg3202)))))
                    begin
                      reg3272 <= reg2204[(3'h6):(3'h6)];
                    end
                  else
                    begin
                      reg3272 <= $unsigned(reg3217);
                      reg3273 <= ((+$signed($signed(reg3215))) != $unsigned((((8'h9d) <= reg3214) ?
                          {reg3247} : (reg3194 ? reg2185 : reg3236))));
                      reg3274 <= reg2208;
                      reg3275 <= (({(reg2211 ? (8'hab) : reg3248)} ?
                              ({reg2197} != (reg3190 ?
                                  reg3238 : reg3222)) : (^~forvar3159)) ?
                          reg2184[(2'h3):(1'h1)] : $unsigned({(reg3234 && reg3216)}));
                    end
                  if (({{(reg3215 >> forvar2212)}} ?
                      reg3121[(4'ha):(4'h9)] : (reg2200 * forvar3127[(1'h0):(1'h0)])))
                    begin
                      reg3276 <= (forvar3125[(2'h3):(1'h1)] * $unsigned($signed(reg3201)));
                      reg3277 <= forvar3152;
                      reg3278 <= $signed($signed($signed((^reg3152))));
                      reg3279 <= ($signed($unsigned($signed(reg2210))) ?
                          reg3230 : $signed(reg3256[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg3276 <= (reg3277[(4'h9):(1'h1)] ?
                          reg3238[(4'ha):(1'h1)] : $unsigned(reg3121));
                      reg3277 <= (~reg2179[(1'h1):(1'h1)]);
                      reg3278 <= (((^~(reg3270 ? reg3188 : forvar3142)) ?
                          $unsigned(reg3238) : $unsigned((reg2202 ?
                              (8'hb9) : reg2198))) <<< (~forvar2186));
                    end
                end
            end
          else
            begin
              if (($unsigned((+(^forvar3226))) || $signed(reg3211)))
                begin
                  for (forvar3269 = (1'h0); (forvar3269 < (2'h3)); forvar3269 = (forvar3269 + (1'h1)))
                    begin
                      reg3270 <= reg3144;
                      reg3271 <= ((^(&wire2174)) - forvar3151[(4'h8):(2'h2)]);
                      reg3272 <= (|(!{$unsigned(reg3198)}));
                      reg3273 <= forvar3178[(1'h1):(1'h0)];
                    end
                  for (forvar3274 = (1'h0); (forvar3274 < (1'h1)); forvar3274 = (forvar3274 + (1'h1)))
                    begin
                      reg3275 <= reg2181[(3'h7):(1'h0)];
                      reg3276 <= reg3274[(3'h5):(3'h4)];
                      reg3277 <= (($unsigned(reg3254) ?
                          (~$signed(reg2192)) : $signed((reg2178 + reg2205))) | $unsigned(forvar3199));
                      reg3278 <= reg3180[(2'h3):(1'h0)];
                    end
                  for (forvar3279 = (1'h0); (forvar3279 < (1'h0)); forvar3279 = (forvar3279 + (1'h1)))
                    begin
                      reg3280 <= (8'hae);
                      reg3281 <= reg3222;
                    end
                end
              else
                begin
                  if ($signed($signed($unsigned(forvar2196[(4'hd):(1'h0)]))))
                    begin
                      reg3269 <= $signed($signed(($signed(reg3161) ?
                          $unsigned((8'hb3)) : (&reg3241))));
                      reg3270 <= (reg3269[(1'h1):(1'h1)] - (!$unsigned((wire2175 ^~ reg3167))));
                      reg3271 <= ((((+forvar3125) >> (forvar3140 > forvar3217)) != ($signed((8'h9e)) ?
                          (reg2220 ?
                              reg2204 : (8'h9e)) : reg3196[(3'h7):(2'h3)])) <= (!$signed((~&reg2222))));
                      reg3272 <= $signed($unsigned(reg3177[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg3269 <= $unsigned(($unsigned($signed(reg2183)) | (reg3184 ?
                          forvar3212 : $signed(reg3171))));
                      reg3270 <= $unsigned(((8'hb7) ?
                          $signed((8'hb4)) : forvar3113));
                      reg3271 <= reg3117;
                    end
                end
              for (forvar3282 = (1'h0); (forvar3282 < (2'h2)); forvar3282 = (forvar3282 + (1'h1)))
                begin
                  for (forvar3283 = (1'h0); (forvar3283 < (2'h3)); forvar3283 = (forvar3283 + (1'h1)))
                    begin
                      reg3284 <= $signed(reg3219[(1'h0):(1'h0)]);
                      reg3285 <= wire2175;
                    end
                  if (forvar2187[(2'h2):(2'h2)])
                    begin
                      reg3286 <= ((^$unsigned(reg2189)) ?
                          {$signed(reg3246[(3'h5):(2'h2)])} : reg3153[(1'h0):(1'h0)]);
                      reg3287 <= ($signed($signed($signed(reg3264))) ?
                          (+$signed(reg2194)) : ((-(reg2183 ?
                                  reg3253 : forvar3259)) ?
                              reg3141 : (reg2222 ~^ (forvar3199 & reg3203))));
                    end
                  else
                    begin
                      reg3286 <= ($unsigned($unsigned((reg2207 <<< forvar3242))) ?
                          {{((8'hb3) >= reg3177)}} : (8'ha5));
                      reg3287 <= reg3202[(3'h4):(1'h1)];
                      reg3288 <= (8'h9c);
                    end
                  reg3289 <= (reg3288[(3'h6):(2'h2)] ?
                      ({(reg3197 ? (8'ha6) : reg3210)} ?
                          reg2195[(1'h0):(1'h0)] : ((reg2205 << reg3237) ?
                              reg3120[(4'h8):(1'h0)] : reg3192[(4'hf):(4'hc)])) : (-(reg3117[(1'h1):(1'h0)] >= $unsigned(forvar2176))));
                end
              if (reg3155)
                begin
                  if ((reg3250 | reg3267[(4'h8):(1'h1)]))
                    begin
                      reg3290 <= (~^$signed((forvar3127 == $signed(reg3243))));
                      reg3291 <= (!$signed((^~$unsigned(forvar2217))));
                      reg3292 <= reg2179;
                      reg3293 <= ($unsigned($unsigned($unsigned((8'h9f)))) & (reg3139[(4'h9):(2'h2)] ?
                          {$unsigned(forvar3212)} : ({reg2218} > (^forvar3181))));
                    end
                  else
                    begin
                      reg3290 <= (!(forvar3151[(4'h8):(3'h7)] ~^ ((reg3213 & reg3233) ?
                          (~^reg2188) : forvar2212)));
                      reg3291 <= wire2170;
                      reg3292 <= forvar3201;
                    end
                  for (forvar3294 = (1'h0); (forvar3294 < (1'h1)); forvar3294 = (forvar3294 + (1'h1)))
                    begin
                      reg3295 <= {(~^$signed(reg2189[(2'h2):(1'h0)]))};
                    end
                end
              else
                begin
                  reg3290 <= reg3199[(2'h3):(2'h2)];
                  if ((^~reg3248))
                    begin
                      reg3291 <= $signed(forvar3142[(3'h4):(1'h0)]);
                      reg3292 <= reg3263[(1'h0):(1'h0)];
                      reg3293 <= $signed($unsigned(forvar3191));
                    end
                  else
                    begin
                      reg3291 <= ((reg3230 ?
                              $signed((reg3261 ?
                                  wire3110 : reg2179)) : ({reg3260} ?
                                  (reg3255 > reg2192) : $signed(forvar3220))) ?
                          ($unsigned(reg2182[(3'h5):(3'h4)]) | reg3120[(4'hb):(3'h4)]) : (|((reg3223 || reg3245) ?
                              $unsigned(forvar3203) : reg2200[(4'ha):(4'h8)])));
                      reg3292 <= ($unsigned($unsigned($signed(forvar3225))) ?
                          $signed({(reg3241 ?
                                  reg2205 : forvar3159)}) : {$signed((~&forvar2212))});
                      reg3293 <= (reg3168[(1'h1):(1'h0)] ?
                          $unsigned((~{(8'ha6)})) : forvar2208);
                    end
                end
              for (forvar3296 = (1'h0); (forvar3296 < (2'h3)); forvar3296 = (forvar3296 + (1'h1)))
                begin
                  for (forvar3297 = (1'h0); (forvar3297 < (2'h2)); forvar3297 = (forvar3297 + (1'h1)))
                    begin
                      reg3298 <= reg3156;
                      reg3299 <= (~reg3272);
                      reg3300 <= $signed(reg3284);
                      reg3301 <= (!(~&$unsigned(wire2171[(2'h2):(2'h2)])));
                    end
                  for (forvar3302 = (1'h0); (forvar3302 < (2'h3)); forvar3302 = (forvar3302 + (1'h1)))
                    begin
                      reg3303 <= (^~($signed((reg3160 ?
                          (8'hb3) : wire2224)) == {$unsigned(reg2222)}));
                      reg3304 <= ($unsigned($unsigned((reg2217 > forvar3244))) != ($signed(((8'ha0) ?
                          forvar2187 : reg2199)) == $unsigned($signed(reg3260))));
                      reg3305 <= $signed((!reg3194));
                      reg3306 <= (reg3261 ? (8'h9f) : {$unsigned(forvar2212)});
                    end
                end
            end
          for (forvar3307 = (1'h0); (forvar3307 < (1'h0)); forvar3307 = (forvar3307 + (1'h1)))
            begin
              for (forvar3308 = (1'h0); (forvar3308 < (2'h3)); forvar3308 = (forvar3308 + (1'h1)))
                begin
                  if ((~&(&forvar3225[(1'h0):(1'h0)])))
                    begin
                      reg3309 <= reg2188;
                      reg3310 <= (~^(|(~^reg2197[(3'h6):(3'h4)])));
                    end
                  else
                    begin
                      reg3309 <= forvar3308[(1'h0):(1'h0)];
                      reg3310 <= (reg3293 ?
                          (reg2210[(4'ha):(3'h5)] - (~|$unsigned(forvar3302))) : {{(forvar3242 ?
                                      (8'hb3) : forvar2196)}});
                      reg3311 <= ($signed(($unsigned(reg2190) < $signed(forvar3191))) >> forvar3178[(4'hb):(4'hb)]);
                      reg3312 <= reg3214;
                    end
                  reg3313 <= (^~$signed($unsigned((~^(8'h9e)))));
                  if ((reg3309[(3'h6):(1'h0)] ?
                      {$unsigned($unsigned(reg3208))} : forvar3259))
                    begin
                      reg3314 <= (~|(+$signed($unsigned((8'hb1)))));
                      reg3315 <= {reg3143};
                      reg3316 <= ({$unsigned(reg2179)} >= ($unsigned($signed(reg2197)) & forvar3162[(3'h4):(1'h1)]));
                    end
                  else
                    begin
                      reg3314 <= $unsigned(reg3274[(4'h9):(3'h6)]);
                      reg3315 <= $signed(($unsigned((8'ha4)) ?
                          reg3288[(1'h0):(1'h0)] : $unsigned((reg2202 ?
                              reg3189 : reg2216))));
                      reg3316 <= ({(~&{forvar3127})} <<< {(forvar3140[(3'h7):(1'h0)] ?
                              $unsigned(reg3304) : (~(8'ha6)))});
                      reg3317 <= forvar3128;
                    end
                  if ({forvar3245[(1'h1):(1'h0)]})
                    begin
                      reg3318 <= $signed(reg2217);
                    end
                  else
                    begin
                      reg3318 <= reg3233[(4'h8):(2'h2)];
                      reg3319 <= reg3201[(4'ha):(2'h3)];
                      reg3320 <= $signed((reg3137[(3'h6):(3'h6)] && $unsigned((reg3264 ?
                          forvar3163 : reg3202))));
                      reg3321 <= $unsigned(reg3232[(2'h3):(1'h0)]);
                    end
                end
              for (forvar3322 = (1'h0); (forvar3322 < (2'h3)); forvar3322 = (forvar3322 + (1'h1)))
                begin
                  reg3323 <= (($signed($signed(reg3169)) * $signed(reg2198[(3'h7):(2'h3)])) ?
                      ((((8'hab) >>> forvar3282) & $unsigned(reg3148)) >= ((&reg3184) ?
                          reg3136 : $unsigned((8'ha2)))) : (8'hb3));
                  for (forvar3324 = (1'h0); (forvar3324 < (2'h3)); forvar3324 = (forvar3324 + (1'h1)))
                    begin
                      reg3325 <= $unsigned(reg3264[(1'h1):(1'h1)]);
                    end
                end
              for (forvar3326 = (1'h0); (forvar3326 < (2'h3)); forvar3326 = (forvar3326 + (1'h1)))
                begin
                  for (forvar3327 = (1'h0); (forvar3327 < (2'h3)); forvar3327 = (forvar3327 + (1'h1)))
                    begin
                      reg3328 <= (|{(~|(8'ha9))});
                      reg3329 <= (-forvar3140);
                      reg3330 <= ($unsigned((-$unsigned(reg2197))) | (|(reg2177 ?
                          $unsigned((8'hb8)) : forvar3252)));
                    end
                  for (forvar3331 = (1'h0); (forvar3331 < (2'h3)); forvar3331 = (forvar3331 + (1'h1)))
                    begin
                      reg3332 <= reg3320[(1'h0):(1'h0)];
                      reg3333 <= $signed($signed($unsigned((reg3237 << forvar3203))));
                    end
                  reg3334 <= ($signed((~(8'hb1))) && reg3167);
                end
            end
          if ({{$unsigned((+reg3201))}})
            begin
              for (forvar3335 = (1'h0); (forvar3335 < (2'h2)); forvar3335 = (forvar3335 + (1'h1)))
                begin
                  for (forvar3336 = (1'h0); (forvar3336 < (2'h3)); forvar3336 = (forvar3336 + (1'h1)))
                    begin
                      reg3337 <= ((((reg3152 == reg3173) ?
                              (reg3219 * reg3293) : ((8'hb1) < reg3193)) ?
                          ($unsigned(reg3147) ^~ {reg3131}) : $unsigned($unsigned((8'hb7)))) || ($unsigned($signed(reg2184)) | {{forvar3199}}));
                      reg3338 <= $unsigned(forvar3181[(1'h1):(1'h0)]);
                      reg3339 <= ((~^$signed((reg3139 ?
                          (8'ha6) : forvar2208))) ~^ ($unsigned((&forvar2180)) ?
                          reg2209 : $unsigned($unsigned(reg3250))));
                    end
                  for (forvar3340 = (1'h0); (forvar3340 < (1'h0)); forvar3340 = (forvar3340 + (1'h1)))
                    begin
                      reg3341 <= (reg3237[(1'h0):(1'h0)] <= (^$signed($signed(reg3233))));
                      reg3342 <= ((reg2217 | (forvar2203[(4'h8):(4'h8)] ?
                          (reg3233 ?
                              reg2179 : reg2186) : forvar2182)) - $unsigned($signed({forvar3331})));
                      reg3343 <= $signed(forvar3225[(2'h2):(2'h2)]);
                      reg3344 <= {((reg3120 < reg2192) | ((reg3333 ?
                              reg3200 : reg2186) << (wire2171 ?
                              reg2188 : reg3229)))};
                    end
                  for (forvar3345 = (1'h0); (forvar3345 < (1'h0)); forvar3345 = (forvar3345 + (1'h1)))
                    begin
                      reg3346 <= reg2184[(1'h0):(1'h0)];
                      reg3347 <= (&{forvar3257});
                    end
                  for (forvar3348 = (1'h0); (forvar3348 < (2'h2)); forvar3348 = (forvar3348 + (1'h1)))
                    begin
                      reg3349 <= reg3271[(2'h2):(1'h0)];
                      reg3350 <= forvar3268;
                    end
                end
              reg3351 <= (reg3169[(1'h1):(1'h1)] != reg3287);
              for (forvar3352 = (1'h0); (forvar3352 < (2'h2)); forvar3352 = (forvar3352 + (1'h1)))
                begin
                  for (forvar3353 = (1'h0); (forvar3353 < (1'h1)); forvar3353 = (forvar3353 + (1'h1)))
                    begin
                      reg3354 <= $signed($unsigned(forvar3353[(1'h1):(1'h0)]));
                      reg3355 <= forvar3231[(3'h5):(2'h3)];
                      reg3356 <= (-($signed(reg3338) ?
                          reg3343[(3'h7):(3'h7)] : $unsigned({reg3156})));
                      reg3357 <= ((|reg3234) ? (8'had) : $signed((~(8'ha9))));
                    end
                  reg3358 <= reg3205[(3'h5):(3'h4)];
                end
              if (((^(|forvar3353[(2'h2):(2'h2)])) * {reg3215[(2'h2):(1'h1)]}))
                begin
                  if (reg3138[(2'h2):(1'h1)])
                    begin
                      reg3359 <= $signed(reg3311[(4'ha):(3'h4)]);
                      reg3360 <= ((8'ha1) - (wire2173[(4'hd):(4'ha)] ?
                          reg3122 : (-(forvar3159 ~^ reg3171))));
                      reg3361 <= (~$unsigned(reg3175));
                    end
                  else
                    begin
                      reg3359 <= (8'hb1);
                    end
                  reg3362 <= ($signed($signed(reg3115)) >= reg3160[(2'h2):(2'h2)]);
                end
              else
                begin
                  for (forvar3359 = (1'h0); (forvar3359 < (2'h2)); forvar3359 = (forvar3359 + (1'h1)))
                    begin
                      reg3360 <= (~reg2217[(1'h0):(1'h0)]);
                      reg3361 <= (~$unsigned(reg3185[(4'hb):(4'ha)]));
                      reg3362 <= (^(|(reg2178[(3'h5):(1'h1)] ?
                          $signed(reg3122) : (8'hb2))));
                    end
                  for (forvar3363 = (1'h0); (forvar3363 < (2'h3)); forvar3363 = (forvar3363 + (1'h1)))
                    begin
                      reg3364 <= {(|(8'h9c))};
                    end
                end
            end
          else
            begin
              for (forvar3335 = (1'h0); (forvar3335 < (2'h2)); forvar3335 = (forvar3335 + (1'h1)))
                begin
                  for (forvar3336 = (1'h0); (forvar3336 < (1'h0)); forvar3336 = (forvar3336 + (1'h1)))
                    begin
                      reg3337 <= $unsigned(((!((8'ha1) ?
                              forvar3191 : forvar3336)) ?
                          $unsigned({forvar3225}) : reg3233));
                      reg3338 <= ((8'h9c) & (~&($unsigned(reg3316) ?
                          (^reg2221) : forvar3242)));
                      reg3339 <= ($unsigned(((reg2209 ?
                          reg3204 : forvar3348) << reg3245[(2'h3):(1'h1)])) > reg3160);
                    end
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1160  (y, clk, wire1161, wire1162, wire1163, wire1164);
  output wire [(32'h3bd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire1161;
  input wire signed [(3'h4):(1'h0)] wire1162;
  input wire signed [(4'hb):(1'h0)] wire1163;
  input wire signed [(4'hb):(1'h0)] wire1164;
  wire signed [(3'h6):(1'h0)] wire2161;
  wire [(3'h7):(1'h0)] wire1165;
  wire signed [(4'h8):(1'h0)] wire1166;
  wire signed [(3'h6):(1'h0)] wire1697;
  reg [(4'hc):(1'h0)] reg1699 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1700 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1701 = (1'h0);
  reg [(3'h4):(1'h0)] reg1702 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1703 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1704 = (1'h0);
  reg [(5'h10):(1'h0)] reg1705 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1706 = (1'h0);
  reg [(4'h8):(1'h0)] reg1707 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1708 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1709 = (1'h0);
  reg [(4'h8):(1'h0)] reg1710 = (1'h0);
  reg [(4'hc):(1'h0)] reg1711 = (1'h0);
  reg [(3'h6):(1'h0)] reg1712 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1713 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1714 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1715 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1716 = (1'h0);
  reg [(4'ha):(1'h0)] reg1717 = (1'h0);
  reg [(2'h3):(1'h0)] reg1718 = (1'h0);
  reg [(4'he):(1'h0)] reg1719 = (1'h0);
  reg [(4'he):(1'h0)] reg1720 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1721 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1722 = (1'h0);
  reg [(4'ha):(1'h0)] reg1723 = (1'h0);
  reg [(4'ha):(1'h0)] reg1724 = (1'h0);
  reg [(4'hd):(1'h0)] reg1725 = (1'h0);
  reg [(3'h6):(1'h0)] reg1716 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1726 = (1'h0);
  reg [(4'he):(1'h0)] reg1727 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1728 = (1'h0);
  reg [(4'h8):(1'h0)] reg1729 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1730 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1731 = (1'h0);
  reg [(2'h2):(1'h0)] reg1732 = (1'h0);
  reg [(4'hf):(1'h0)] reg1733 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1734 = (1'h0);
  reg [(3'h5):(1'h0)] reg1735 = (1'h0);
  reg [(4'h8):(1'h0)] reg1736 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1737 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1738 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1739 = (1'h0);
  reg [(3'h5):(1'h0)] reg1740 = (1'h0);
  reg [(3'h6):(1'h0)] reg1741 = (1'h0);
  reg [(3'h7):(1'h0)] reg1742 = (1'h0);
  reg [(4'hd):(1'h0)] reg1743 = (1'h0);
  reg [(4'hc):(1'h0)] reg1744 = (1'h0);
  reg [(4'h8):(1'h0)] reg1745 = (1'h0);
  reg [(4'hd):(1'h0)] reg1746 = (1'h0);
  reg [(4'hb):(1'h0)] reg1747 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1748 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1749 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1750 = (1'h0);
  reg [(3'h4):(1'h0)] reg1751 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1752 = (1'h0);
  reg [(5'h10):(1'h0)] reg1753 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1754 = (1'h0);
  reg [(5'h10):(1'h0)] reg1755 = (1'h0);
  reg [(4'hf):(1'h0)] reg1756 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1757 = (1'h0);
  reg [(2'h3):(1'h0)] reg1758 = (1'h0);
  reg [(4'hf):(1'h0)] reg1759 = (1'h0);
  reg [(2'h3):(1'h0)] reg1760 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1761 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1762 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1763 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1764 = (1'h0);
  reg [(2'h2):(1'h0)] reg1765 = (1'h0);
  reg [(5'h10):(1'h0)] reg1766 = (1'h0);
  reg [(2'h2):(1'h0)] reg1767 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1768 = (1'h0);
  reg [(2'h2):(1'h0)] reg1769 = (1'h0);
  reg [(2'h2):(1'h0)] reg1770 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1771 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1772 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1773 = (1'h0);
  reg [(4'h8):(1'h0)] reg1774 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1775 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1776 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1777 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1778 = (1'h0);
  reg [(3'h6):(1'h0)] reg1779 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1780 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1777 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1779 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1781 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1782 = (1'h0);
  reg [(5'h10):(1'h0)] reg1783 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1784 = (1'h0);
  reg [(3'h6):(1'h0)] reg1776 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1778 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1780 = (1'h0);
  reg [(3'h5):(1'h0)] reg1785 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1786 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1787 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1788 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1789 = (1'h0);
  reg [(2'h2):(1'h0)] reg1790 = (1'h0);
  reg [(3'h6):(1'h0)] reg1791 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire1792;
  wire signed [(3'h6):(1'h0)] wire1793;
  wire signed [(3'h5):(1'h0)] wire2159;
  assign y = {wire2161,
                 wire1165,
                 wire1166,
                 wire1697,
                 reg1699,
                 forvar1700,
                 forvar1701,
                 reg1702,
                 forvar1703,
                 forvar1704,
                 reg1705,
                 reg1706,
                 reg1707,
                 reg1708,
                 reg1709,
                 reg1710,
                 reg1711,
                 reg1712,
                 reg1713,
                 reg1714,
                 reg1715,
                 forvar1716,
                 reg1717,
                 reg1718,
                 reg1719,
                 reg1720,
                 reg1721,
                 reg1722,
                 reg1723,
                 reg1724,
                 reg1725,
                 reg1716,
                 forvar1726,
                 reg1727,
                 forvar1728,
                 reg1729,
                 reg1730,
                 reg1731,
                 reg1732,
                 reg1733,
                 forvar1734,
                 reg1735,
                 reg1736,
                 forvar1737,
                 forvar1738,
                 forvar1739,
                 reg1740,
                 reg1741,
                 reg1742,
                 reg1743,
                 reg1744,
                 reg1745,
                 reg1746,
                 reg1747,
                 reg1748,
                 reg1749,
                 reg1750,
                 reg1751,
                 reg1752,
                 reg1753,
                 forvar1754,
                 reg1755,
                 reg1756,
                 forvar1757,
                 reg1758,
                 reg1759,
                 reg1760,
                 reg1761,
                 forvar1762,
                 forvar1763,
                 reg1764,
                 reg1765,
                 reg1766,
                 reg1767,
                 forvar1768,
                 reg1769,
                 reg1770,
                 reg1771,
                 forvar1772,
                 forvar1773,
                 reg1774,
                 reg1775,
                 forvar1776,
                 forvar1777,
                 reg1778,
                 reg1779,
                 reg1780,
                 reg1777,
                 forvar1779,
                 reg1781,
                 reg1782,
                 reg1783,
                 reg1784,
                 reg1776,
                 forvar1778,
                 forvar1780,
                 reg1785,
                 reg1786,
                 forvar1787,
                 forvar1788,
                 reg1789,
                 reg1790,
                 reg1791,
                 wire1792,
                 wire1793,
                 wire2159,
                 (1'h0)};
  assign wire1165 = $signed(((wire1162[(1'h1):(1'h0)] && wire1162[(1'h1):(1'h0)]) ^~ $signed($unsigned((8'hb5)))));
  assign wire1166 = $signed(wire1162);
  module1167 modinst1698 (.clk(clk), .wire1171(wire1165), .y(wire1697), .wire1169(wire1164), .wire1168(wire1163), .wire1170(wire1161));
  always
    @(posedge clk) begin
      reg1699 <= (!wire1161);
      for (forvar1700 = (1'h0); (forvar1700 < (2'h3)); forvar1700 = (forvar1700 + (1'h1)))
        begin
          for (forvar1701 = (1'h0); (forvar1701 < (2'h3)); forvar1701 = (forvar1701 + (1'h1)))
            begin
              reg1702 <= (8'ha6);
              for (forvar1703 = (1'h0); (forvar1703 < (2'h3)); forvar1703 = (forvar1703 + (1'h1)))
                begin
                  for (forvar1704 = (1'h0); (forvar1704 < (1'h0)); forvar1704 = (forvar1704 + (1'h1)))
                    begin
                      reg1705 <= wire1161;
                      reg1706 <= $signed(((^wire1165) || $unsigned($unsigned(wire1164))));
                      reg1707 <= (($signed(reg1702[(2'h2):(1'h0)]) <<< wire1165[(3'h6):(3'h4)]) ?
                          ($unsigned((8'hb2)) << $unsigned(wire1162)) : ($signed(reg1706[(3'h4):(2'h3)]) & ((forvar1701 ?
                              forvar1703 : reg1699) || {wire1166})));
                      reg1708 <= {wire1697};
                    end
                  if ((reg1702 != forvar1701[(4'hc):(3'h5)]))
                    begin
                      reg1709 <= (reg1699 ?
                          (!(8'h9c)) : ((wire1165[(1'h1):(1'h1)] <<< wire1697[(3'h4):(2'h3)]) ?
                              wire1162[(2'h2):(2'h2)] : {forvar1703[(1'h0):(1'h0)]}));
                      reg1710 <= forvar1701[(4'hf):(3'h5)];
                      reg1711 <= (forvar1700 ?
                          $unsigned($unsigned(reg1705)) : (~^$signed((wire1166 ?
                              wire1161 : wire1164))));
                      reg1712 <= reg1707;
                    end
                  else
                    begin
                      reg1709 <= reg1705;
                      reg1710 <= $unsigned($unsigned(wire1166));
                    end
                  if ((((forvar1700 ?
                          wire1165 : $unsigned(wire1164)) || $unsigned(reg1712)) ?
                      (^~{$signed((8'h9d))}) : ((~reg1709[(4'h8):(2'h3)]) ?
                          $signed((reg1707 ? wire1161 : wire1163)) : reg1707)))
                    begin
                      reg1713 <= ($signed($signed((forvar1703 ?
                              reg1711 : reg1710))) ?
                          (~&$unsigned((8'ha2))) : ($unsigned($signed(wire1165)) ?
                              $unsigned((~(8'hb0))) : $signed({forvar1701})));
                      reg1714 <= $unsigned($signed($signed($signed(reg1713))));
                    end
                  else
                    begin
                      reg1713 <= {$signed({((8'hab) ^~ wire1166)})};
                      reg1714 <= ({wire1164} << (!{(&wire1161)}));
                      reg1715 <= (~^reg1711);
                    end
                end
              if (reg1712[(2'h2):(1'h1)])
                begin
                  for (forvar1716 = (1'h0); (forvar1716 < (1'h0)); forvar1716 = (forvar1716 + (1'h1)))
                    begin
                      reg1717 <= $signed(($unsigned($unsigned((8'hb0))) <= reg1714));
                      reg1718 <= (reg1706 != $unsigned(({reg1706} || $signed(reg1717))));
                      reg1719 <= {((&$signed(wire1163)) >> $signed(reg1708))};
                    end
                  if (wire1162[(1'h0):(1'h0)])
                    begin
                      reg1720 <= reg1702[(1'h1):(1'h1)];
                      reg1721 <= forvar1716[(5'h10):(5'h10)];
                    end
                  else
                    begin
                      reg1720 <= forvar1701;
                    end
                  reg1722 <= (wire1163 ?
                      (((~^reg1717) != (^wire1697)) <= ((reg1718 <= wire1163) && {wire1164})) : reg1707[(3'h6):(1'h0)]);
                  if ((~|(reg1712 ? {reg1706} : forvar1716[(1'h0):(1'h0)])))
                    begin
                      reg1723 <= {(wire1163 ?
                              ((8'ha6) >= ((8'haf) ?
                                  reg1713 : wire1166)) : (~^(reg1709 ?
                                  wire1166 : forvar1703)))};
                    end
                  else
                    begin
                      reg1723 <= (&$unsigned($unsigned($unsigned(reg1717))));
                      reg1724 <= $unsigned($signed(reg1719[(2'h3):(1'h0)]));
                      reg1725 <= wire1697[(3'h5):(2'h2)];
                    end
                end
              else
                begin
                  reg1716 <= reg1702[(2'h3):(2'h3)];
                  if (($signed(($unsigned(reg1709) - $unsigned(wire1165))) ?
                      $unsigned(($signed(reg1699) ^~ $unsigned(reg1715))) : ($unsigned((~^forvar1703)) <= $signed((reg1715 && forvar1703)))))
                    begin
                      reg1717 <= reg1718[(2'h2):(1'h0)];
                      reg1718 <= (reg1721 ?
                          ((reg1707 ?
                                  reg1707[(3'h7):(1'h0)] : forvar1701[(3'h4):(3'h4)]) ?
                              {(reg1710 ?
                                      (8'ha4) : reg1715)} : (wire1163[(4'hb):(3'h6)] + (forvar1701 ?
                                  reg1702 : forvar1700))) : (+$signed((reg1715 ?
                              reg1699 : wire1164))));
                    end
                  else
                    begin
                      reg1717 <= (~(-(|$signed(wire1161))));
                      reg1718 <= (wire1163[(3'h7):(2'h3)] ?
                          (+(~&$unsigned(reg1716))) : $signed(((reg1705 >> reg1711) ?
                              (wire1165 >> forvar1701) : (reg1702 ?
                                  (8'hae) : (8'hb5)))));
                      reg1719 <= ((((+wire1697) ?
                                  (8'hb7) : (reg1702 > wire1165)) ?
                              (~&wire1165[(1'h0):(1'h0)]) : ((!reg1722) ?
                                  forvar1703 : $unsigned(reg1723))) ?
                          (($signed((8'h9c)) != reg1707) >>> (|(wire1163 >>> reg1719))) : reg1721[(3'h4):(2'h2)]);
                      reg1720 <= reg1708[(1'h1):(1'h1)];
                    end
                  if (($unsigned($signed(reg1714[(4'h9):(3'h7)])) ?
                      wire1165 : wire1165))
                    begin
                      reg1721 <= $signed((~|reg1724));
                      reg1722 <= ($unsigned(((wire1165 | reg1715) - reg1724[(3'h4):(2'h3)])) > (8'hb4));
                      reg1723 <= (wire1163[(1'h0):(1'h0)] ?
                          $signed(forvar1701) : ({$unsigned(reg1718)} ?
                              (&$signed(reg1716)) : ((+wire1164) ?
                                  $signed(wire1166) : (forvar1703 ?
                                      reg1717 : forvar1716))));
                      reg1724 <= (({reg1710[(3'h4):(2'h3)]} >= (|(!wire1697))) ?
                          ((&wire1166) ?
                              {$signed(reg1707)} : reg1709[(1'h0):(1'h0)]) : $unsigned((^~{wire1697})));
                    end
                  else
                    begin
                      reg1721 <= ($unsigned(({reg1712} ?
                              reg1708[(3'h7):(3'h4)] : wire1164[(3'h5):(3'h5)])) ?
                          {(reg1711[(1'h0):(1'h0)] ?
                                  {(8'hb6)} : (reg1719 ?
                                      reg1709 : reg1699))} : (-(8'ha4)));
                      reg1722 <= (forvar1703[(1'h1):(1'h0)] ~^ $unsigned(((!reg1719) ?
                          $unsigned(reg1705) : $unsigned(reg1717))));
                    end
                end
              for (forvar1726 = (1'h0); (forvar1726 < (1'h1)); forvar1726 = (forvar1726 + (1'h1)))
                begin
                  reg1727 <= wire1166;
                  for (forvar1728 = (1'h0); (forvar1728 < (2'h2)); forvar1728 = (forvar1728 + (1'h1)))
                    begin
                      reg1729 <= $signed(reg1722[(4'hf):(4'h8)]);
                      reg1730 <= $signed((forvar1700[(2'h3):(1'h0)] ?
                          ($signed(forvar1728) ?
                              reg1710 : (reg1714 ?
                                  forvar1703 : reg1709)) : reg1711[(4'h8):(2'h2)]));
                      reg1731 <= $unsigned(($unsigned((reg1714 > forvar1701)) > $unsigned((reg1702 + forvar1703))));
                      reg1732 <= wire1163;
                    end
                  reg1733 <= $unsigned(reg1725);
                  for (forvar1734 = (1'h0); (forvar1734 < (2'h2)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= ($unsigned(reg1725) ?
                          $signed($unsigned((reg1721 ?
                              (8'hb8) : reg1708))) : (!(forvar1703[(1'h0):(1'h0)] ?
                              $signed(reg1699) : (~|reg1712))));
                      reg1736 <= {({$unsigned((8'haa))} ?
                              (!reg1735[(2'h2):(1'h1)]) : $unsigned($unsigned(reg1721)))};
                    end
                end
            end
          for (forvar1737 = (1'h0); (forvar1737 < (2'h2)); forvar1737 = (forvar1737 + (1'h1)))
            begin
              for (forvar1738 = (1'h0); (forvar1738 < (2'h2)); forvar1738 = (forvar1738 + (1'h1)))
                begin
                  for (forvar1739 = (1'h0); (forvar1739 < (2'h3)); forvar1739 = (forvar1739 + (1'h1)))
                    begin
                      reg1740 <= ($unsigned(reg1707) ?
                          forvar1716[(2'h3):(1'h1)] : (^~($signed(wire1161) == (reg1713 ?
                              forvar1700 : forvar1703))));
                    end
                  if ((($signed($signed(reg1707)) ?
                      ((~|forvar1703) ?
                          reg1720 : {reg1740}) : ({forvar1738} ^~ $signed(reg1719))) > (((-forvar1704) + reg1699) ?
                      $signed($unsigned((8'hb9))) : $signed((reg1712 ?
                          reg1727 : forvar1739)))))
                    begin
                      reg1741 <= reg1714;
                      reg1742 <= (reg1714 & $unsigned((|forvar1738[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg1741 <= (~&((~|(reg1722 <<< reg1712)) ?
                          (8'hb2) : reg1725));
                      reg1742 <= (+($unsigned((reg1742 < reg1706)) | ($unsigned(forvar1700) ?
                          reg1718 : reg1727)));
                    end
                  if ($signed(((reg1713[(3'h5):(2'h2)] ?
                      reg1707[(2'h2):(2'h2)] : $unsigned(reg1740)) ~^ (8'ha0))))
                    begin
                      reg1743 <= reg1741;
                      reg1744 <= forvar1716;
                      reg1745 <= forvar1700[(3'h4):(1'h0)];
                      reg1746 <= (~&reg1699);
                    end
                  else
                    begin
                      reg1743 <= (wire1164 ?
                          (((reg1740 ?
                              (8'ha7) : reg1732) | reg1735[(1'h1):(1'h1)]) + $signed(reg1711[(4'hc):(4'ha)])) : {forvar1716[(3'h5):(1'h1)]});
                      reg1744 <= $unsigned(reg1712[(1'h0):(1'h0)]);
                    end
                  if ((~^reg1719[(4'hd):(4'hc)]))
                    begin
                      reg1747 <= (^~reg1712);
                      reg1748 <= ((reg1705[(3'h4):(1'h1)] ?
                              ((reg1745 ? reg1736 : forvar1716) <<< ((8'ha7) ?
                                  reg1707 : reg1743)) : reg1699) ?
                          ({$signed(reg1724)} ~^ {(wire1697 & forvar1737)}) : (&{reg1708}));
                      reg1749 <= ($signed(($unsigned(forvar1701) ?
                          reg1715 : (reg1713 ?
                              forvar1700 : forvar1700))) || reg1720[(4'ha):(4'h8)]);
                      reg1750 <= (^~$unsigned(((reg1749 <<< (8'ha7)) ?
                          $signed((8'hae)) : ((8'hb4) ? wire1165 : (8'ha0)))));
                    end
                  else
                    begin
                      reg1747 <= {((^$signed(reg1714)) ?
                              {(~&forvar1734)} : $signed($unsigned((8'ha1))))};
                      reg1748 <= {(~|(|{reg1743}))};
                    end
                end
              if ($signed((|$signed((reg1713 && reg1743)))))
                begin
                  if ({$unsigned({(forvar1737 != forvar1734)})})
                    begin
                      reg1751 <= $unsigned((((&reg1745) ?
                          (reg1716 ?
                              forvar1701 : wire1162) : $signed(wire1165)) + ($signed(wire1162) <= reg1710)));
                      reg1752 <= ($unsigned((forvar1701[(1'h0):(1'h0)] ^ (reg1740 ?
                          (8'ha9) : reg1748))) * $unsigned(reg1715));
                      reg1753 <= wire1163;
                    end
                  else
                    begin
                      reg1751 <= (($unsigned($unsigned(reg1727)) | $unsigned((reg1702 ?
                              reg1736 : (8'ha6)))) ?
                          ($signed({reg1712}) == forvar1738) : reg1741);
                    end
                  for (forvar1754 = (1'h0); (forvar1754 < (1'h0)); forvar1754 = (forvar1754 + (1'h1)))
                    begin
                      reg1755 <= ($unsigned({(8'hb9)}) ?
                          reg1705[(5'h10):(5'h10)] : $unsigned(wire1165[(1'h1):(1'h1)]));
                      reg1756 <= (((~&$unsigned(reg1714)) ?
                              reg1744[(4'h9):(1'h0)] : reg1716) ?
                          (reg1705[(2'h2):(1'h1)] <<< $unsigned($unsigned(reg1711))) : $signed($unsigned((reg1730 ?
                              wire1162 : (8'h9c)))));
                    end
                  for (forvar1757 = (1'h0); (forvar1757 < (1'h0)); forvar1757 = (forvar1757 + (1'h1)))
                    begin
                      reg1758 <= $unsigned((($signed(reg1709) >>> {reg1720}) ?
                          (~^{reg1732}) : ((-reg1729) ^~ (~|reg1707))));
                      reg1759 <= $unsigned((reg1725 ?
                          (forvar1726[(2'h3):(2'h3)] ?
                              (^reg1706) : (reg1745 << reg1752)) : $unsigned(wire1162)));
                      reg1760 <= ((reg1724 << (^((8'ha6) ?
                          (8'ha5) : reg1743))) << (reg1755 - (reg1707 ?
                          forvar1739 : $unsigned(reg1742))));
                    end
                  reg1761 <= ((~^((reg1756 ?
                      reg1725 : forvar1737) == reg1748[(3'h5):(1'h1)])) > $signed((forvar1734[(3'h6):(1'h0)] ?
                      (reg1731 < (8'hb3)) : (reg1731 ? reg1718 : (8'had)))));
                end
              else
                begin
                  if ($signed({$signed({reg1722})}))
                    begin
                      reg1751 <= ($signed(reg1745[(1'h1):(1'h0)]) ~^ ((-(reg1707 ?
                          reg1743 : reg1743)) <<< $unsigned((&reg1740))));
                      reg1752 <= {forvar1701};
                      reg1753 <= reg1711[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1751 <= {(8'h9e)};
                      reg1752 <= ($unsigned(reg1716) * $signed($signed((reg1712 ?
                          (8'h9f) : wire1161))));
                    end
                end
              for (forvar1762 = (1'h0); (forvar1762 < (1'h0)); forvar1762 = (forvar1762 + (1'h1)))
                begin
                  for (forvar1763 = (1'h0); (forvar1763 < (1'h1)); forvar1763 = (forvar1763 + (1'h1)))
                    begin
                      reg1764 <= forvar1738[(3'h7):(3'h5)];
                      reg1765 <= $unsigned($unsigned(((forvar1716 ?
                          reg1724 : reg1735) & reg1756[(4'hb):(3'h7)])));
                      reg1766 <= reg1761;
                    end
                  reg1767 <= $unsigned($signed((!(~^reg1699))));
                  for (forvar1768 = (1'h0); (forvar1768 < (2'h2)); forvar1768 = (forvar1768 + (1'h1)))
                    begin
                      reg1769 <= $unsigned(reg1752[(1'h1):(1'h1)]);
                      reg1770 <= (((~^reg1705[(1'h0):(1'h0)]) != reg1745[(4'h8):(3'h6)]) ?
                          forvar1704[(4'h8):(4'h8)] : reg1730[(1'h0):(1'h0)]);
                      reg1771 <= {forvar1728[(1'h1):(1'h1)]};
                    end
                end
              for (forvar1772 = (1'h0); (forvar1772 < (1'h0)); forvar1772 = (forvar1772 + (1'h1)))
                begin
                  for (forvar1773 = (1'h0); (forvar1773 < (2'h3)); forvar1773 = (forvar1773 + (1'h1)))
                    begin
                      reg1774 <= ((((8'hb8) ?
                              $unsigned(reg1720) : (!(8'hac))) == reg1730[(4'h8):(3'h5)]) ?
                          (^~reg1751[(1'h0):(1'h0)]) : $signed($unsigned((~&reg1718))));
                      reg1775 <= reg1767[(1'h0):(1'h0)];
                    end
                end
            end
          if ($signed($signed(((reg1731 ? (8'ha6) : forvar1716) ?
              (reg1743 >>> reg1711) : (reg1735 >>> reg1713)))))
            begin
              for (forvar1776 = (1'h0); (forvar1776 < (1'h0)); forvar1776 = (forvar1776 + (1'h1)))
                begin
                  for (forvar1777 = (1'h0); (forvar1777 < (1'h1)); forvar1777 = (forvar1777 + (1'h1)))
                    begin
                      reg1778 <= forvar1768;
                      reg1779 <= (8'ha1);
                    end
                end
              reg1780 <= reg1731;
            end
          else
            begin
              if (reg1735[(1'h0):(1'h0)])
                begin
                  for (forvar1776 = (1'h0); (forvar1776 < (1'h1)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 <= reg1729;
                      reg1778 <= (^(~|({reg1761} ?
                          $signed(reg1742) : ((8'ha8) ?
                              (8'hb0) : forvar1776))));
                    end
                  for (forvar1779 = (1'h0); (forvar1779 < (2'h3)); forvar1779 = (forvar1779 + (1'h1)))
                    begin
                      reg1780 <= $unsigned(forvar1763[(2'h3):(2'h3)]);
                      reg1781 <= (^forvar1773[(1'h1):(1'h1)]);
                      reg1782 <= $unsigned(({$unsigned(reg1708)} ?
                          ($signed(forvar1773) ^~ reg1727[(1'h0):(1'h0)]) : $unsigned({wire1161})));
                    end
                  if ($signed((reg1723[(3'h4):(1'h1)] ?
                      $unsigned(((8'ha4) + forvar1728)) : $unsigned(forvar1701))))
                    begin
                      reg1783 <= reg1712;
                      reg1784 <= (|$unsigned(reg1724));
                    end
                  else
                    begin
                      reg1783 <= reg1756;
                      reg1784 <= $unsigned(reg1710);
                    end
                end
              else
                begin
                  if ((8'h9e))
                    begin
                      reg1776 <= reg1765[(1'h0):(1'h0)];
                      reg1777 <= $unsigned((^~(8'hb3)));
                    end
                  else
                    begin
                      reg1776 <= {(($signed(reg1776) | $unsigned(reg1764)) == $signed((~&reg1749)))};
                      reg1777 <= $signed((((-reg1764) ?
                              (|reg1730) : (reg1745 <<< (8'hae))) ?
                          reg1719 : $unsigned($signed(reg1749))));
                    end
                  for (forvar1778 = (1'h0); (forvar1778 < (1'h1)); forvar1778 = (forvar1778 + (1'h1)))
                    begin
                      reg1779 <= wire1163;
                    end
                  for (forvar1780 = (1'h0); (forvar1780 < (1'h1)); forvar1780 = (forvar1780 + (1'h1)))
                    begin
                      reg1781 <= {(^(8'ha6))};
                      reg1782 <= $signed({reg1725[(4'hd):(2'h2)]});
                      reg1783 <= (&$unsigned((reg1778[(3'h4):(1'h0)] ?
                          $unsigned(wire1165) : (~&(8'hb5)))));
                    end
                  if (reg1731[(4'h8):(1'h1)])
                    begin
                      reg1784 <= (~&((!reg1699[(4'h9):(1'h1)]) ?
                          ((~&reg1705) <= $unsigned(reg1732)) : (reg1713 | (reg1750 ?
                              reg1702 : (8'h9d)))));
                      reg1785 <= reg1777;
                    end
                  else
                    begin
                      reg1784 <= (((~reg1746[(4'hc):(2'h2)]) >> {reg1777[(1'h1):(1'h1)]}) >= (|(!(reg1720 ?
                          forvar1773 : reg1779))));
                      reg1785 <= reg1743[(3'h4):(3'h4)];
                      reg1786 <= (-(8'ha6));
                    end
                end
            end
          for (forvar1787 = (1'h0); (forvar1787 < (2'h2)); forvar1787 = (forvar1787 + (1'h1)))
            begin
              for (forvar1788 = (1'h0); (forvar1788 < (1'h1)); forvar1788 = (forvar1788 + (1'h1)))
                begin
                  if (((reg1744 ?
                          (&reg1744[(4'hc):(3'h6)]) : reg1785[(2'h2):(1'h1)]) ?
                      reg1767 : $signed(((forvar1780 ? reg1776 : reg1786) ?
                          $unsigned(forvar1734) : (forvar1777 ^ reg1748)))))
                    begin
                      reg1789 <= {reg1717};
                    end
                  else
                    begin
                      reg1789 <= (!(8'ha8));
                      reg1790 <= $signed((~&($signed(reg1716) ?
                          reg1759[(1'h1):(1'h1)] : reg1729)));
                    end
                end
              reg1791 <= reg1771;
            end
        end
    end
  assign wire1792 = ($unsigned(($signed(reg1714) == (8'had))) ?
                        ($signed(forvar1780[(1'h1):(1'h0)]) <= (~|(forvar1773 ?
                            forvar1763 : forvar1701))) : reg1730);
  assign wire1793 = (^$unsigned(((reg1789 ^ reg1759) > $unsigned(forvar1734))));
  module1794 modinst2160 (wire2159, clk, reg1721, wire1166, reg1761, reg1764, reg1752);
  assign wire2161 = ((~^reg1752[(3'h5):(1'h0)]) << $unsigned($signed(reg1720[(4'hb):(3'h6)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1794
#( parameter param2158 = ((+(((8'hb2) ? (8'h9d) : (8'ha8)) ? ((8'hac) ? (8'ha2) : (8'ha2)) : ((8'hb0) | (8'hab)))) ^~ (~^((^(8'hac)) * (+(8'hba))))) )
(y, clk, wire1795, wire1796, wire1797, wire1798, wire1799);
  output wire [(32'h33):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h5):(1'h0)] wire1795;
  input wire [(3'h7):(1'h0)] wire1796;
  input wire [(4'hd):(1'h0)] wire1797;
  input wire [(4'hc):(1'h0)] wire1798;
  input wire signed [(4'he):(1'h0)] wire1799;
  wire [(4'h8):(1'h0)] wire2157;
  wire signed [(5'h10):(1'h0)] wire1800;
  wire [(4'ha):(1'h0)] wire1801;
  wire [(4'h8):(1'h0)] wire1802;
  wire signed [(4'h8):(1'h0)] wire2155;
  assign y = {wire2157, wire1800, wire1801, wire1802, wire2155, (1'h0)};
  assign wire1800 = (-wire1796[(2'h2):(1'h0)]);
  assign wire1801 = (8'haf);
  assign wire1802 = (((8'h9c) ? wire1801 : {$signed(wire1795)}) ?
                        {$unsigned($signed(wire1801))} : ((8'hab) ^ wire1800));
  module1803 modinst2156 (.wire1808(wire1799), .wire1806(wire1797), .wire1804(wire1796), .y(wire2155), .wire1805(wire1802), .clk(clk), .wire1807(wire1800));
  assign wire2157 = $unsigned((wire2155 & (^(~wire1798))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1167  (y, clk, wire1168, wire1169, wire1170, wire1171);
  output wire [(32'hdf5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire1168;
  input wire [(4'hb):(1'h0)] wire1169;
  input wire [(3'h5):(1'h0)] wire1170;
  input wire [(3'h7):(1'h0)] wire1171;
  wire signed [(2'h2):(1'h0)] wire1696;
  wire [(4'hf):(1'h0)] wire1695;
  wire [(4'h9):(1'h0)] wire1694;
  reg [(3'h5):(1'h0)] forvar1675 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1673 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1669 = (1'h0);
  reg [(2'h2):(1'h0)] reg1668 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1663 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1659 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1648 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1647 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1636 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1625 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1623 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1643 = (1'h0);
  reg [(2'h3):(1'h0)] reg1642 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1639 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1631 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1630 = (1'h0);
  reg [(2'h2):(1'h0)] reg1629 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1627 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1693 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1692 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1691 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1690 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1689 = (1'h0);
  reg [(4'he):(1'h0)] reg1688 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1687 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1687 = (1'h0);
  reg [(4'hf):(1'h0)] reg1686 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1685 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1684 = (1'h0);
  reg [(3'h4):(1'h0)] reg1683 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1682 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1678 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1682 = (1'h0);
  reg [(4'hb):(1'h0)] reg1681 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1680 = (1'h0);
  reg [(3'h5):(1'h0)] reg1679 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1677 = (1'h0);
  reg [(3'h7):(1'h0)] reg1676 = (1'h0);
  reg [(4'hb):(1'h0)] reg1675 = (1'h0);
  reg [(2'h3):(1'h0)] reg1674 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1671 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1670 = (1'h0);
  reg [(2'h2):(1'h0)] reg1673 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1672 = (1'h0);
  reg [(4'hf):(1'h0)] reg1671 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1670 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1669 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1668 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1667 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1666 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1665 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1664 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1663 = (1'h0);
  reg [(3'h4):(1'h0)] reg1662 = (1'h0);
  reg [(3'h7):(1'h0)] reg1661 = (1'h0);
  reg [(4'h9):(1'h0)] reg1660 = (1'h0);
  reg [(4'h8):(1'h0)] reg1659 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1658 = (1'h0);
  reg [(4'hd):(1'h0)] reg1657 = (1'h0);
  reg [(5'h10):(1'h0)] reg1656 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1655 = (1'h0);
  reg [(2'h2):(1'h0)] reg1654 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1653 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1652 = (1'h0);
  reg [(4'hf):(1'h0)] reg1651 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1650 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1649 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1648 = (1'h0);
  reg [(2'h3):(1'h0)] reg1647 = (1'h0);
  reg [(2'h3):(1'h0)] reg1646 = (1'h0);
  reg [(4'hd):(1'h0)] reg1645 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1644 = (1'h0);
  reg [(4'ha):(1'h0)] reg1643 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1642 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1641 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1640 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1639 = (1'h0);
  reg [(4'ha):(1'h0)] reg1638 = (1'h0);
  reg [(4'hc):(1'h0)] reg1637 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1636 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1635 = (1'h0);
  reg [(2'h2):(1'h0)] reg1634 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1633 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1632 = (1'h0);
  reg [(3'h5):(1'h0)] reg1631 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1630 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1629 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1628 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1624 = (1'h0);
  reg [(4'hc):(1'h0)] reg1627 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1626 = (1'h0);
  reg [(3'h4):(1'h0)] reg1625 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1624 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1623 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire1622;
  reg signed [(4'h8):(1'h0)] forvar1605 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1607 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1598 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1621 = (1'h0);
  reg [(4'hb):(1'h0)] reg1620 = (1'h0);
  reg [(4'ha):(1'h0)] reg1619 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1618 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1617 = (1'h0);
  reg [(3'h7):(1'h0)] reg1613 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1609 = (1'h0);
  reg [(3'h6):(1'h0)] reg1608 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1604 = (1'h0);
  reg [(2'h3):(1'h0)] reg1616 = (1'h0);
  reg [(3'h6):(1'h0)] reg1615 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1614 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1613 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1612 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1611 = (1'h0);
  reg [(3'h7):(1'h0)] reg1610 = (1'h0);
  reg [(4'hb):(1'h0)] reg1609 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1608 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1607 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1606 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1605 = (1'h0);
  reg [(3'h7):(1'h0)] reg1604 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1601 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1603 = (1'h0);
  reg [(2'h3):(1'h0)] reg1602 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1601 = (1'h0);
  reg [(4'he):(1'h0)] reg1600 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1599 = (1'h0);
  reg [(3'h5):(1'h0)] reg1598 = (1'h0);
  reg [(4'he):(1'h0)] forvar1597 = (1'h0);
  reg [(4'ha):(1'h0)] reg1596 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1595 = (1'h0);
  reg [(4'hd):(1'h0)] reg1594 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1593 = (1'h0);
  reg [(4'hd):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1591 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1590 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1590 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1589 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1588 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1576 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1568 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1567 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1565 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1564 = (1'h0);
  reg [(4'hb):(1'h0)] reg1587 = (1'h0);
  reg [(3'h6):(1'h0)] reg1586 = (1'h0);
  reg [(4'he):(1'h0)] forvar1585 = (1'h0);
  reg [(2'h2):(1'h0)] reg1584 = (1'h0);
  reg [(4'hf):(1'h0)] reg1583 = (1'h0);
  reg [(2'h2):(1'h0)] reg1582 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1581 = (1'h0);
  reg [(3'h7):(1'h0)] reg1580 = (1'h0);
  reg [(2'h3):(1'h0)] reg1579 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1578 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1577 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1576 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1575 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1574 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1573 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1572 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1571 = (1'h0);
  reg [(4'h8):(1'h0)] reg1570 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1569 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1568 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1567 = (1'h0);
  reg [(4'h9):(1'h0)] reg1566 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1565 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1564 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1563 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1562 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1561 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1560 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1559 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1558 = (1'h0);
  reg [(4'hd):(1'h0)] reg1557 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1556 = (1'h0);
  reg [(3'h4):(1'h0)] reg1555 = (1'h0);
  reg [(4'he):(1'h0)] reg1553 = (1'h0);
  reg [(4'he):(1'h0)] forvar1552 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1547 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1544 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1549 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1548 = (1'h0);
  reg [(4'h9):(1'h0)] reg1554 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1553 = (1'h0);
  reg [(4'hf):(1'h0)] reg1552 = (1'h0);
  reg [(2'h2):(1'h0)] reg1551 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1550 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1549 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1548 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1547 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1546 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1545 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1544 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1543 = (1'h0);
  reg [(3'h5):(1'h0)] reg1542 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1541 = (1'h0);
  reg [(4'hc):(1'h0)] reg1540 = (1'h0);
  reg [(4'hb):(1'h0)] reg1539 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1538 = (1'h0);
  reg [(3'h4):(1'h0)] reg1537 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1536 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1535 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1534 = (1'h0);
  reg [(3'h4):(1'h0)] reg1533 = (1'h0);
  reg [(3'h6):(1'h0)] reg1532 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1531 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1530 = (1'h0);
  reg [(2'h2):(1'h0)] reg1525 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1529 = (1'h0);
  reg [(5'h10):(1'h0)] reg1528 = (1'h0);
  reg [(3'h6):(1'h0)] reg1527 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1526 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1525 = (1'h0);
  reg [(4'hb):(1'h0)] reg1524 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1523 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1522 = (1'h0);
  reg [(3'h5):(1'h0)] reg1521 = (1'h0);
  reg [(4'hc):(1'h0)] reg1520 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1519 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1518 = (1'h0);
  reg [(4'hb):(1'h0)] reg1517 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1516 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1515 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1514 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1513 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1512 = (1'h0);
  reg [(4'ha):(1'h0)] reg1511 = (1'h0);
  reg [(4'hb):(1'h0)] reg1510 = (1'h0);
  reg [(4'he):(1'h0)] forvar1509 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1508 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1507 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1506 = (1'h0);
  reg [(4'ha):(1'h0)] reg1505 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1504 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1502 = (1'h0);
  reg [(4'hb):(1'h0)] reg1497 = (1'h0);
  reg [(2'h3):(1'h0)] reg1496 = (1'h0);
  reg [(4'he):(1'h0)] forvar1494 = (1'h0);
  reg [(4'hf):(1'h0)] reg1485 = (1'h0);
  reg [(3'h5):(1'h0)] reg1484 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1482 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1481 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1503 = (1'h0);
  reg [(4'hf):(1'h0)] reg1502 = (1'h0);
  reg [(3'h5):(1'h0)] reg1501 = (1'h0);
  reg [(3'h6):(1'h0)] reg1500 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1499 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1498 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1497 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1496 = (1'h0);
  reg [(4'h9):(1'h0)] reg1495 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1494 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1492 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1490 = (1'h0);
  reg [(3'h5):(1'h0)] reg1489 = (1'h0);
  reg [(5'h10):(1'h0)] reg1493 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1492 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1491 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1490 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1489 = (1'h0);
  reg [(3'h4):(1'h0)] reg1488 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1487 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1486 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1485 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1484 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1479 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1473 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1483 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1482 = (1'h0);
  reg [(2'h2):(1'h0)] reg1481 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1480 = (1'h0);
  reg [(4'hb):(1'h0)] reg1479 = (1'h0);
  reg [(4'he):(1'h0)] reg1478 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1477 = (1'h0);
  reg [(3'h4):(1'h0)] reg1476 = (1'h0);
  reg [(4'h8):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1474 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1473 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1472 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1471 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1470 = (1'h0);
  reg [(3'h7):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1468 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1467 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1461 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1457 = (1'h0);
  reg [(4'h8):(1'h0)] reg1456 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1466 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1465 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1464 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1463 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1462 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1461 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1460 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1459 = (1'h0);
  reg [(4'h9):(1'h0)] reg1458 = (1'h0);
  reg [(3'h7):(1'h0)] reg1457 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1456 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1455 = (1'h0);
  reg [(4'ha):(1'h0)] reg1454 = (1'h0);
  reg [(2'h2):(1'h0)] reg1453 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1452 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1451 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1450 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1449 = (1'h0);
  reg [(4'hd):(1'h0)] reg1448 = (1'h0);
  reg [(5'h10):(1'h0)] reg1447 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1446 = (1'h0);
  reg [(4'hb):(1'h0)] reg1442 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1438 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1445 = (1'h0);
  reg [(4'hf):(1'h0)] reg1444 = (1'h0);
  reg [(4'hb):(1'h0)] reg1443 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1442 = (1'h0);
  reg [(5'h10):(1'h0)] reg1441 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1440 = (1'h0);
  reg [(4'he):(1'h0)] reg1439 = (1'h0);
  reg [(4'ha):(1'h0)] reg1438 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1437 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1436 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1396 = (1'h0);
  reg [(3'h4):(1'h0)] reg1395 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1390 = (1'h0);
  reg [(4'hd):(1'h0)] reg1387 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1385 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1381 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1435 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1434 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1433 = (1'h0);
  reg [(3'h4):(1'h0)] reg1432 = (1'h0);
  reg [(4'h8):(1'h0)] reg1431 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1430 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1429 = (1'h0);
  reg [(4'hb):(1'h0)] reg1428 = (1'h0);
  reg [(4'hf):(1'h0)] reg1427 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1426 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1425 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1424 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1423 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1422 = (1'h0);
  reg [(5'h10):(1'h0)] reg1421 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1420 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1419 = (1'h0);
  reg [(2'h3):(1'h0)] reg1418 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1417 = (1'h0);
  reg [(4'ha):(1'h0)] reg1416 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1415 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1414 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1413 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1412 = (1'h0);
  reg [(4'ha):(1'h0)] reg1411 = (1'h0);
  reg [(4'h8):(1'h0)] reg1410 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1409 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1408 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1407 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1406 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1405 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1404 = (1'h0);
  reg [(4'hc):(1'h0)] reg1403 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1402 = (1'h0);
  reg [(4'hb):(1'h0)] reg1401 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1400 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1399 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1398 = (1'h0);
  reg [(5'h10):(1'h0)] reg1397 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1396 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1395 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1394 = (1'h0);
  reg [(4'ha):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1392 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1391 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1390 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1379 = (1'h0);
  reg [(4'he):(1'h0)] reg1389 = (1'h0);
  reg [(4'hf):(1'h0)] reg1388 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1387 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1386 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1385 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1384 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1383 = (1'h0);
  reg [(3'h7):(1'h0)] reg1382 = (1'h0);
  reg [(4'h9):(1'h0)] reg1381 = (1'h0);
  reg [(4'he):(1'h0)] forvar1380 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1380 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1379 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire1172;
  wire [(3'h4):(1'h0)] wire1377;
  assign y = {wire1696,
                 wire1695,
                 wire1694,
                 forvar1675,
                 forvar1673,
                 forvar1669,
                 reg1668,
                 forvar1663,
                 forvar1659,
                 forvar1648,
                 forvar1647,
                 reg1636,
                 forvar1625,
                 reg1623,
                 forvar1643,
                 reg1642,
                 reg1639,
                 forvar1631,
                 forvar1630,
                 reg1629,
                 forvar1627,
                 reg1693,
                 reg1692,
                 reg1691,
                 reg1690,
                 forvar1689,
                 reg1688,
                 forvar1687,
                 reg1687,
                 reg1686,
                 reg1685,
                 reg1684,
                 reg1683,
                 forvar1682,
                 forvar1678,
                 reg1682,
                 reg1681,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1674,
                 forvar1671,
                 reg1670,
                 reg1673,
                 reg1672,
                 reg1671,
                 forvar1670,
                 reg1669,
                 forvar1668,
                 reg1667,
                 reg1666,
                 reg1665,
                 reg1664,
                 reg1663,
                 reg1662,
                 reg1661,
                 reg1660,
                 reg1659,
                 reg1658,
                 reg1657,
                 reg1656,
                 forvar1655,
                 reg1654,
                 forvar1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 forvar1642,
                 forvar1641,
                 reg1640,
                 forvar1639,
                 reg1638,
                 reg1637,
                 forvar1636,
                 reg1635,
                 reg1634,
                 forvar1633,
                 reg1632,
                 reg1631,
                 reg1630,
                 forvar1629,
                 reg1628,
                 forvar1624,
                 reg1627,
                 reg1626,
                 reg1625,
                 reg1624,
                 forvar1623,
                 wire1622,
                 forvar1605,
                 forvar1607,
                 forvar1598,
                 reg1621,
                 reg1620,
                 reg1619,
                 reg1618,
                 forvar1617,
                 reg1613,
                 forvar1609,
                 reg1608,
                 forvar1604,
                 reg1616,
                 reg1615,
                 reg1614,
                 forvar1613,
                 reg1612,
                 reg1611,
                 reg1610,
                 reg1609,
                 forvar1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1601,
                 reg1603,
                 reg1602,
                 forvar1601,
                 reg1600,
                 reg1599,
                 reg1598,
                 forvar1597,
                 reg1596,
                 reg1595,
                 reg1594,
                 reg1593,
                 reg1592,
                 forvar1591,
                 forvar1590,
                 reg1590,
                 reg1589,
                 forvar1588,
                 forvar1576,
                 reg1568,
                 forvar1567,
                 reg1565,
                 reg1564,
                 reg1587,
                 reg1586,
                 forvar1585,
                 reg1584,
                 reg1583,
                 reg1582,
                 forvar1581,
                 reg1580,
                 reg1579,
                 reg1578,
                 reg1577,
                 reg1576,
                 reg1575,
                 reg1574,
                 reg1573,
                 forvar1572,
                 forvar1571,
                 reg1570,
                 reg1569,
                 forvar1568,
                 reg1567,
                 reg1566,
                 forvar1565,
                 forvar1564,
                 reg1563,
                 forvar1562,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1558,
                 reg1557,
                 forvar1556,
                 reg1555,
                 reg1553,
                 forvar1552,
                 forvar1547,
                 forvar1544,
                 reg1549,
                 forvar1548,
                 reg1554,
                 forvar1553,
                 reg1552,
                 reg1551,
                 reg1550,
                 forvar1549,
                 reg1548,
                 reg1547,
                 reg1546,
                 reg1545,
                 reg1544,
                 reg1543,
                 reg1542,
                 reg1541,
                 reg1540,
                 reg1539,
                 forvar1538,
                 reg1537,
                 reg1536,
                 forvar1535,
                 forvar1534,
                 reg1533,
                 reg1532,
                 forvar1531,
                 reg1530,
                 reg1525,
                 reg1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 forvar1525,
                 reg1524,
                 forvar1523,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 reg1518,
                 reg1517,
                 reg1516,
                 forvar1515,
                 forvar1514,
                 forvar1513,
                 reg1512,
                 reg1511,
                 reg1510,
                 forvar1509,
                 reg1508,
                 reg1507,
                 reg1506,
                 reg1505,
                 reg1504,
                 forvar1502,
                 reg1497,
                 reg1496,
                 forvar1494,
                 reg1485,
                 reg1484,
                 reg1482,
                 forvar1481,
                 reg1503,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1499,
                 reg1498,
                 forvar1497,
                 forvar1496,
                 reg1495,
                 reg1494,
                 forvar1492,
                 forvar1490,
                 reg1489,
                 reg1493,
                 reg1492,
                 reg1491,
                 reg1490,
                 forvar1489,
                 reg1488,
                 reg1487,
                 reg1486,
                 forvar1485,
                 forvar1484,
                 forvar1479,
                 reg1473,
                 reg1483,
                 forvar1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1475,
                 reg1474,
                 forvar1473,
                 forvar1472,
                 reg1471,
                 reg1470,
                 reg1469,
                 forvar1468,
                 reg1467,
                 reg1461,
                 forvar1457,
                 reg1456,
                 reg1466,
                 reg1465,
                 reg1464,
                 reg1463,
                 reg1462,
                 forvar1461,
                 reg1460,
                 reg1459,
                 reg1458,
                 reg1457,
                 forvar1456,
                 reg1455,
                 reg1454,
                 reg1453,
                 reg1452,
                 reg1451,
                 reg1450,
                 forvar1449,
                 reg1448,
                 reg1447,
                 reg1446,
                 reg1442,
                 forvar1438,
                 reg1445,
                 reg1444,
                 reg1443,
                 forvar1442,
                 reg1441,
                 reg1440,
                 reg1439,
                 reg1438,
                 forvar1437,
                 forvar1436,
                 forvar1396,
                 reg1395,
                 reg1390,
                 reg1387,
                 forvar1385,
                 forvar1381,
                 reg1435,
                 reg1434,
                 forvar1433,
                 reg1432,
                 reg1431,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 forvar1425,
                 forvar1424,
                 forvar1423,
                 reg1422,
                 reg1421,
                 reg1420,
                 reg1419,
                 reg1418,
                 forvar1417,
                 reg1416,
                 reg1415,
                 forvar1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 reg1410,
                 reg1409,
                 reg1408,
                 forvar1407,
                 forvar1406,
                 reg1405,
                 reg1404,
                 reg1403,
                 reg1402,
                 reg1401,
                 reg1400,
                 reg1399,
                 reg1398,
                 reg1397,
                 reg1396,
                 forvar1395,
                 reg1394,
                 reg1393,
                 reg1392,
                 reg1391,
                 forvar1390,
                 forvar1379,
                 reg1389,
                 reg1388,
                 forvar1387,
                 reg1386,
                 reg1385,
                 reg1384,
                 forvar1383,
                 reg1382,
                 reg1381,
                 forvar1380,
                 reg1380,
                 reg1379,
                 wire1172,
                 wire1377,
                 (1'h0)};
  assign wire1172 = $unsigned($unsigned(wire1168));
  module1173 modinst1378 (wire1377, clk, wire1168, wire1169, wire1171, wire1172, wire1170);
  always
    @(posedge clk) begin
      if ((($unsigned($unsigned(wire1377)) == $unsigned((wire1168 ?
          wire1172 : wire1168))) <= (~(~|$unsigned(wire1377)))))
        begin
          if (wire1169[(3'h4):(1'h1)])
            begin
              reg1379 <= $signed($unsigned($signed($unsigned(wire1171))));
              if ($signed(($signed({(8'hab)}) >>> (^{wire1168}))))
                begin
                  reg1380 <= ($unsigned(((~wire1169) ?
                      wire1377 : {reg1379})) == ((-$signed(wire1170)) ?
                      wire1377 : ((reg1379 ? wire1172 : wire1172) ?
                          (wire1172 ? wire1172 : wire1169) : (~|(8'h9d)))));
                end
              else
                begin
                  for (forvar1380 = (1'h0); (forvar1380 < (2'h3)); forvar1380 = (forvar1380 + (1'h1)))
                    begin
                      reg1381 <= wire1170;
                      reg1382 <= ($signed((8'hb4)) ?
                          ((reg1380 ?
                                  (wire1172 ?
                                      reg1380 : wire1168) : $signed(forvar1380)) ?
                              wire1377[(1'h1):(1'h0)] : {wire1168}) : reg1380);
                    end
                  for (forvar1383 = (1'h0); (forvar1383 < (1'h0)); forvar1383 = (forvar1383 + (1'h1)))
                    begin
                      reg1384 <= wire1168;
                      reg1385 <= (reg1379[(2'h2):(1'h0)] | $unsigned({((8'hab) && wire1169)}));
                    end
                  if ($unsigned((~{{reg1384}})))
                    begin
                      reg1386 <= ((((~&reg1380) ?
                                  $unsigned(wire1171) : (&reg1379)) ?
                              (~&(reg1385 ?
                                  forvar1380 : wire1168)) : $signed($signed(wire1172))) ?
                          $signed((wire1377[(1'h1):(1'h0)] | wire1377)) : wire1169);
                    end
                  else
                    begin
                      reg1386 <= (~(wire1172 >>> $signed((^wire1172))));
                    end
                end
              for (forvar1387 = (1'h0); (forvar1387 < (1'h0)); forvar1387 = (forvar1387 + (1'h1)))
                begin
                  reg1388 <= ((($unsigned(wire1172) ?
                      reg1384[(1'h1):(1'h1)] : (forvar1387 + reg1382)) >> $signed((8'ha8))) <= $unsigned((~wire1171[(3'h4):(2'h2)])));
                end
              reg1389 <= {wire1172[(4'ha):(4'h9)]};
            end
          else
            begin
              if (reg1385)
                begin
                  reg1379 <= (wire1170[(3'h5):(3'h5)] || $signed(($signed(forvar1380) >> (8'h9d))));
                  reg1380 <= ($unsigned(reg1382[(1'h1):(1'h1)]) ~^ (~&reg1386));
                end
              else
                begin
                  for (forvar1379 = (1'h0); (forvar1379 < (1'h1)); forvar1379 = (forvar1379 + (1'h1)))
                    begin
                      reg1380 <= (((~|(forvar1379 << forvar1387)) & ((8'ha5) || $unsigned(wire1171))) ?
                          ((^{forvar1380}) <= wire1169) : (!$unsigned($signed(reg1382))));
                    end
                end
            end
          if ($signed({$signed($unsigned(reg1389))}))
            begin
              for (forvar1390 = (1'h0); (forvar1390 < (2'h2)); forvar1390 = (forvar1390 + (1'h1)))
                begin
                  if (({$signed((wire1170 ? (8'hb4) : (8'ha8)))} ?
                      reg1389 : (8'h9f)))
                    begin
                      reg1391 <= $unsigned((reg1386[(2'h2):(2'h2)] ?
                          forvar1379 : reg1381[(4'h8):(1'h1)]));
                      reg1392 <= $unsigned((reg1384[(4'hb):(3'h7)] ?
                          (~&$signed(wire1170)) : $signed((wire1170 >>> reg1379))));
                    end
                  else
                    begin
                      reg1391 <= $unsigned((reg1381[(4'h9):(4'h8)] ^ (reg1385 ?
                          (~^reg1388) : (wire1172 ? reg1389 : reg1386))));
                      reg1392 <= forvar1379[(3'h4):(2'h2)];
                      reg1393 <= ((reg1392 ?
                          (reg1385[(4'hc):(3'h5)] ?
                              (reg1381 ? (8'haf) : forvar1380) : (reg1380 ?
                                  forvar1390 : reg1388)) : $signed(wire1168[(3'h6):(3'h4)])) + (&(reg1385 ?
                          ((8'h9c) <= forvar1379) : reg1385[(1'h1):(1'h0)])));
                      reg1394 <= $unsigned(wire1170[(1'h1):(1'h0)]);
                    end
                end
            end
          else
            begin
              for (forvar1390 = (1'h0); (forvar1390 < (1'h1)); forvar1390 = (forvar1390 + (1'h1)))
                begin
                  if (wire1377)
                    begin
                      reg1391 <= {reg1384};
                    end
                  else
                    begin
                      reg1391 <= $signed((reg1380 ?
                          reg1384 : ((reg1379 == reg1381) ?
                              $signed(wire1172) : (+reg1388))));
                      reg1392 <= $unsigned((reg1391 ?
                          (|reg1382) : wire1171[(1'h1):(1'h0)]));
                      reg1393 <= reg1385;
                    end
                  reg1394 <= {wire1171};
                end
              for (forvar1395 = (1'h0); (forvar1395 < (2'h2)); forvar1395 = (forvar1395 + (1'h1)))
                begin
                  if ((reg1379[(1'h1):(1'h0)] ?
                      wire1172 : {$unsigned(reg1381)}))
                    begin
                      reg1396 <= (^~reg1380[(3'h5):(3'h4)]);
                      reg1397 <= wire1168;
                      reg1398 <= (forvar1395 ?
                          (reg1381 ?
                              ($signed(forvar1390) <= $signed((8'hb4))) : {$signed(reg1391)}) : (wire1169 < $unsigned({(8'hba)})));
                    end
                  else
                    begin
                      reg1396 <= ((wire1169 ~^ forvar1390[(3'h4):(2'h3)]) ^ ({$signed(wire1170)} ?
                          (~|$unsigned(reg1388)) : $signed(wire1168[(4'h9):(1'h1)])));
                    end
                  if ($signed(($signed(reg1380) && $signed($signed(reg1385)))))
                    begin
                      reg1399 <= $signed(({$unsigned((8'ha7))} ?
                          reg1384 : (reg1381[(2'h3):(1'h0)] & $signed(reg1388))));
                      reg1400 <= $unsigned($unsigned((^~{reg1382})));
                      reg1401 <= $signed(((~&(&reg1386)) ^~ $signed(reg1399)));
                    end
                  else
                    begin
                      reg1399 <= reg1398[(3'h4):(2'h3)];
                    end
                  if ({(^reg1380[(3'h4):(2'h2)])})
                    begin
                      reg1402 <= (~&$signed($unsigned($signed(reg1384))));
                      reg1403 <= ({((wire1170 ?
                              forvar1379 : wire1171) >= $unsigned(forvar1379))} - $unsigned({(reg1400 ?
                              reg1396 : forvar1390)}));
                      reg1404 <= ($signed(reg1402[(1'h1):(1'h1)]) ?
                          $signed($signed((~^reg1379))) : {($unsigned(forvar1379) && reg1380[(4'h8):(4'h8)])});
                    end
                  else
                    begin
                      reg1402 <= (wire1170[(2'h2):(1'h0)] && $unsigned(forvar1383[(2'h3):(2'h3)]));
                      reg1403 <= ((reg1393[(4'h9):(4'h9)] < (wire1172[(3'h5):(2'h3)] | {reg1394})) ?
                          reg1400 : $signed((~^wire1377[(1'h0):(1'h0)])));
                    end
                  reg1405 <= $signed(wire1171);
                end
              for (forvar1406 = (1'h0); (forvar1406 < (1'h0)); forvar1406 = (forvar1406 + (1'h1)))
                begin
                  for (forvar1407 = (1'h0); (forvar1407 < (1'h0)); forvar1407 = (forvar1407 + (1'h1)))
                    begin
                      reg1408 <= ((8'hb8) & (-($unsigned(forvar1380) || (reg1391 <<< reg1405))));
                      reg1409 <= reg1405;
                      reg1410 <= reg1402[(4'ha):(2'h3)];
                    end
                  if ($unsigned((reg1393 <<< forvar1395)))
                    begin
                      reg1411 <= forvar1379[(4'h9):(1'h1)];
                      reg1412 <= (~|($unsigned(forvar1395) ?
                          reg1392 : {(!reg1386)}));
                    end
                  else
                    begin
                      reg1411 <= {$unsigned(((reg1386 == (8'h9e)) ?
                              (reg1397 ?
                                  reg1398 : reg1380) : $unsigned((8'hb6))))};
                      reg1412 <= {({reg1396[(1'h0):(1'h0)]} ?
                              ({forvar1387} ?
                                  $signed(wire1377) : $unsigned(wire1170)) : $unsigned(reg1402[(3'h7):(3'h7)]))};
                      reg1413 <= {(wire1169[(3'h7):(2'h2)] ?
                              (reg1410 ?
                                  $signed((8'haf)) : $unsigned(forvar1380)) : $signed((wire1171 ?
                                  reg1389 : reg1399)))};
                    end
                  for (forvar1414 = (1'h0); (forvar1414 < (1'h1)); forvar1414 = (forvar1414 + (1'h1)))
                    begin
                      reg1415 <= (($signed(forvar1383) || wire1170[(3'h5):(3'h5)]) > ({$unsigned(reg1411)} ^ $unsigned(forvar1395)));
                      reg1416 <= (^wire1377[(2'h3):(1'h0)]);
                    end
                  for (forvar1417 = (1'h0); (forvar1417 < (2'h2)); forvar1417 = (forvar1417 + (1'h1)))
                    begin
                      reg1418 <= reg1415[(2'h3):(2'h2)];
                      reg1419 <= reg1405;
                      reg1420 <= reg1381;
                      reg1421 <= $signed((8'ha4));
                    end
                end
              reg1422 <= ((8'h9e) <= reg1394[(4'he):(4'ha)]);
            end
          for (forvar1423 = (1'h0); (forvar1423 < (1'h1)); forvar1423 = (forvar1423 + (1'h1)))
            begin
              for (forvar1424 = (1'h0); (forvar1424 < (1'h1)); forvar1424 = (forvar1424 + (1'h1)))
                begin
                  for (forvar1425 = (1'h0); (forvar1425 < (2'h2)); forvar1425 = (forvar1425 + (1'h1)))
                    begin
                      reg1426 <= reg1400;
                      reg1427 <= (reg1405 <<< $signed(reg1394[(3'h4):(1'h1)]));
                      reg1428 <= (reg1421[(3'h6):(3'h6)] ?
                          $signed(reg1389) : (wire1377 ?
                              reg1391 : reg1391[(4'h8):(3'h7)]));
                      reg1429 <= ((+wire1377) ?
                          (|reg1427[(4'ha):(2'h3)]) : $unsigned((8'hb4)));
                    end
                  if ((^reg1402))
                    begin
                      reg1430 <= ((~^{((8'ha8) + (8'ha7))}) >> $unsigned(({reg1412} ?
                          reg1418[(1'h0):(1'h0)] : ((8'hae) ?
                              reg1429 : (8'ha9)))));
                      reg1431 <= reg1391;
                      reg1432 <= {$unsigned(reg1380[(4'h8):(4'h8)])};
                    end
                  else
                    begin
                      reg1430 <= reg1386[(2'h3):(1'h1)];
                      reg1431 <= $unsigned($unsigned(forvar1424[(1'h1):(1'h0)]));
                    end
                  for (forvar1433 = (1'h0); (forvar1433 < (1'h1)); forvar1433 = (forvar1433 + (1'h1)))
                    begin
                      reg1434 <= (&({{reg1402}} ?
                          forvar1395 : (~&$signed(wire1377))));
                      reg1435 <= reg1396;
                    end
                end
            end
        end
      else
        begin
          for (forvar1379 = (1'h0); (forvar1379 < (2'h3)); forvar1379 = (forvar1379 + (1'h1)))
            begin
              for (forvar1380 = (1'h0); (forvar1380 < (1'h0)); forvar1380 = (forvar1380 + (1'h1)))
                begin
                  for (forvar1381 = (1'h0); (forvar1381 < (1'h1)); forvar1381 = (forvar1381 + (1'h1)))
                    begin
                      reg1382 <= ((^$signed({(8'hac)})) * (forvar1387[(1'h0):(1'h0)] ^ reg1427[(4'hd):(1'h0)]));
                    end
                  for (forvar1383 = (1'h0); (forvar1383 < (1'h0)); forvar1383 = (forvar1383 + (1'h1)))
                    begin
                      reg1384 <= $unsigned($signed({$signed(wire1170)}));
                    end
                end
              if (reg1410[(3'h6):(3'h6)])
                begin
                  for (forvar1385 = (1'h0); (forvar1385 < (1'h0)); forvar1385 = (forvar1385 + (1'h1)))
                    begin
                      reg1386 <= $unsigned((reg1431 ?
                          (reg1410 ^ (~reg1389)) : (~wire1170[(3'h4):(1'h0)])));
                      reg1387 <= (($unsigned(reg1420[(1'h1):(1'h1)]) ?
                          {{forvar1387}} : (^wire1377)) * {(~^(^reg1389))});
                      reg1388 <= $signed({{(reg1394 ? reg1386 : reg1397)}});
                    end
                  reg1389 <= (((~^$unsigned(forvar1381)) ?
                      {(+wire1172)} : $signed((|reg1413))) + $unsigned($unsigned(reg1432)));
                end
              else
                begin
                  for (forvar1385 = (1'h0); (forvar1385 < (2'h2)); forvar1385 = (forvar1385 + (1'h1)))
                    begin
                      reg1386 <= reg1394;
                      reg1387 <= $signed($unsigned($signed($unsigned((8'had)))));
                    end
                  if ($unsigned(reg1387))
                    begin
                      reg1388 <= $unsigned((+$unsigned((reg1391 > reg1388))));
                    end
                  else
                    begin
                      reg1388 <= ((~{$signed(reg1393)}) ?
                          reg1388 : (|$signed($signed(reg1404))));
                      reg1389 <= reg1435;
                      reg1390 <= (($unsigned(reg1380) < ((reg1418 >= (8'hb8)) >= $unsigned(forvar1433))) ?
                          reg1411[(3'h7):(3'h6)] : (8'haa));
                    end
                  reg1391 <= $unsigned((forvar1433 ?
                      (reg1422 && $signed(forvar1406)) : $unsigned((reg1386 ?
                          reg1390 : forvar1423))));
                  if (((&((wire1170 ?
                      reg1418 : reg1380) || reg1413)) <<< (^~$signed((reg1409 & reg1411)))))
                    begin
                      reg1392 <= {({$signed(reg1387)} ?
                              $signed($unsigned((8'hb8))) : reg1387[(3'h7):(2'h3)])};
                    end
                  else
                    begin
                      reg1392 <= reg1428;
                      reg1393 <= {$unsigned((reg1429[(3'h5):(1'h1)] ~^ (reg1408 << (8'ha9))))};
                    end
                end
              reg1394 <= reg1384[(3'h6):(3'h6)];
            end
          if (wire1172)
            begin
              reg1395 <= ($signed($signed((~&forvar1407))) ?
                  $signed(reg1418[(1'h0):(1'h0)]) : reg1431);
              for (forvar1396 = (1'h0); (forvar1396 < (1'h1)); forvar1396 = (forvar1396 + (1'h1)))
                begin
                  reg1397 <= ($unsigned(reg1420) ?
                      (($signed(reg1422) | (reg1415 >>> wire1168)) || $unsigned(forvar1407)) : $unsigned(reg1415[(1'h0):(1'h0)]));
                  if ((!$unsigned((forvar1423 ^~ (forvar1387 ?
                      (8'hb4) : reg1435)))))
                    begin
                      reg1398 <= ($unsigned((~&(~|reg1432))) ?
                          $signed(((reg1395 < reg1427) + reg1434[(3'h7):(2'h3)])) : reg1405[(4'hb):(1'h0)]);
                    end
                  else
                    begin
                      reg1398 <= reg1413;
                      reg1399 <= wire1168;
                      reg1400 <= (($unsigned(((8'ha2) & (8'hb8))) << (reg1382 ?
                              $signed(reg1408) : (reg1419 | forvar1407))) ?
                          (^~$signed((+(8'ha6)))) : $signed($signed((~^reg1400))));
                      reg1401 <= (wire1172[(4'h9):(2'h3)] ?
                          reg1412[(1'h1):(1'h0)] : (~reg1393[(2'h3):(1'h1)]));
                    end
                end
            end
          else
            begin
              reg1395 <= (!(forvar1423[(4'h8):(3'h5)] >= (forvar1390 ?
                  (forvar1433 ^~ forvar1433) : (~^reg1389))));
            end
        end
      for (forvar1436 = (1'h0); (forvar1436 < (1'h1)); forvar1436 = (forvar1436 + (1'h1)))
        begin
          for (forvar1437 = (1'h0); (forvar1437 < (1'h0)); forvar1437 = (forvar1437 + (1'h1)))
            begin
              if (reg1394[(2'h2):(1'h1)])
                begin
                  if (forvar1387[(1'h0):(1'h0)])
                    begin
                      reg1438 <= forvar1407[(3'h7):(1'h0)];
                      reg1439 <= (reg1394[(3'h6):(1'h1)] > reg1382[(2'h3):(2'h2)]);
                      reg1440 <= reg1429;
                      reg1441 <= $signed((wire1168 ?
                          ((-forvar1423) << $unsigned(reg1393)) : (reg1408 ?
                              reg1409[(4'h8):(2'h3)] : reg1408[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg1438 <= {forvar1390};
                      reg1439 <= $signed(forvar1424[(2'h2):(1'h1)]);
                      reg1440 <= ($unsigned(reg1411[(3'h4):(3'h4)]) - (+reg1385[(4'hc):(3'h6)]));
                      reg1441 <= (((~^(reg1408 - (8'hb7))) ?
                          reg1401[(2'h2):(2'h2)] : reg1389) ^~ $signed((8'ha9)));
                    end
                  for (forvar1442 = (1'h0); (forvar1442 < (1'h0)); forvar1442 = (forvar1442 + (1'h1)))
                    begin
                      reg1443 <= forvar1436;
                      reg1444 <= reg1411[(3'h5):(3'h5)];
                      reg1445 <= ((((reg1394 * reg1410) ?
                          (reg1380 ?
                              reg1402 : forvar1396) : $unsigned(forvar1406)) + $signed($signed(reg1389))) || reg1430[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar1438 = (1'h0); (forvar1438 < (2'h3)); forvar1438 = (forvar1438 + (1'h1)))
                    begin
                      reg1439 <= (reg1441[(2'h3):(1'h0)] ?
                          reg1401 : forvar1390);
                      reg1440 <= {reg1405};
                      reg1441 <= (reg1380 && $unsigned(reg1379));
                      reg1442 <= reg1404[(1'h0):(1'h0)];
                    end
                  if (reg1427[(2'h2):(1'h1)])
                    begin
                      reg1443 <= reg1405;
                      reg1444 <= {$signed($unsigned($signed((8'ha6))))};
                      reg1445 <= reg1390[(4'h9):(4'h9)];
                      reg1446 <= $unsigned((8'ha0));
                    end
                  else
                    begin
                      reg1443 <= $signed(forvar1406);
                      reg1444 <= wire1170;
                      reg1445 <= (reg1444 ?
                          (($unsigned(reg1397) + reg1410) >>> ((reg1418 ?
                              (8'ha7) : (8'hb3)) + reg1427[(4'hd):(4'hb)])) : (reg1384[(4'hb):(3'h4)] ?
                              ((reg1443 ?
                                  reg1389 : (8'ha9)) >>> $unsigned(wire1168)) : ($unsigned(reg1420) ^~ (reg1416 != forvar1424))));
                      reg1446 <= $signed((({reg1416} >= $unsigned((8'ha7))) && ((8'haf) ?
                          $signed(reg1384) : (-reg1446))));
                    end
                  reg1447 <= $unsigned(reg1384);
                  reg1448 <= forvar1433[(3'h6):(1'h0)];
                end
              for (forvar1449 = (1'h0); (forvar1449 < (2'h3)); forvar1449 = (forvar1449 + (1'h1)))
                begin
                  reg1450 <= ($signed($unsigned(forvar1406)) & $unsigned((reg1430[(3'h5):(2'h2)] ^ {(8'hac)})));
                  if ((8'ha7))
                    begin
                      reg1451 <= (((~|(reg1440 & reg1409)) ?
                              wire1169[(2'h3):(1'h1)] : {(reg1396 * reg1402)}) ?
                          $unsigned({$signed(reg1400)}) : (~^wire1171));
                      reg1452 <= $unsigned({((reg1403 ?
                              reg1432 : reg1430) != (reg1402 || reg1412))});
                    end
                  else
                    begin
                      reg1451 <= (forvar1379[(3'h4):(3'h4)] ?
                          reg1432[(3'h4):(1'h0)] : ({forvar1417[(4'h9):(2'h2)]} ?
                              {(reg1427 ? reg1440 : reg1429)} : (~(reg1422 ?
                                  reg1438 : reg1403))));
                      reg1452 <= (-{reg1386[(2'h3):(2'h3)]});
                      reg1453 <= $signed({$signed(forvar1438[(1'h0):(1'h0)])});
                      reg1454 <= $signed(reg1403);
                    end
                  reg1455 <= (|((((8'haa) | reg1413) ^ $signed(reg1392)) ?
                      $signed(forvar1436[(3'h7):(3'h5)]) : reg1409));
                end
              if ((~&({$signed(reg1439)} ?
                  ((reg1396 - reg1398) ?
                      forvar1396[(3'h6):(3'h6)] : $unsigned(reg1440)) : $signed((reg1445 ?
                      reg1403 : reg1422)))))
                begin
                  for (forvar1456 = (1'h0); (forvar1456 < (1'h1)); forvar1456 = (forvar1456 + (1'h1)))
                    begin
                      reg1457 <= (~&reg1410[(2'h3):(1'h1)]);
                    end
                  if (($signed((|(reg1392 * wire1172))) & ((reg1443 <<< wire1172) ?
                      ($signed(forvar1437) ^ $unsigned(reg1420)) : ((reg1379 << (8'hb4)) ?
                          reg1429 : {forvar1387}))))
                    begin
                      reg1458 <= $unsigned($signed(reg1390[(3'h4):(2'h2)]));
                      reg1459 <= (&$unsigned(((forvar1424 < reg1448) ?
                          (~forvar1417) : (^reg1430))));
                      reg1460 <= reg1421[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg1458 <= forvar1379;
                    end
                  for (forvar1461 = (1'h0); (forvar1461 < (2'h2)); forvar1461 = (forvar1461 + (1'h1)))
                    begin
                      reg1462 <= {reg1447[(3'h5):(1'h1)]};
                    end
                  if (((|(~&$unsigned(reg1393))) <<< {(|reg1418[(1'h1):(1'h0)])}))
                    begin
                      reg1463 <= $signed(((reg1382 << reg1430[(4'h8):(3'h5)]) * ((wire1170 ?
                              reg1398 : reg1379) ?
                          $unsigned(reg1418) : $signed(forvar1424))));
                      reg1464 <= $signed(reg1434);
                      reg1465 <= forvar1417;
                    end
                  else
                    begin
                      reg1463 <= $signed((^~reg1381[(2'h2):(2'h2)]));
                      reg1464 <= ((($signed(reg1418) ?
                          $unsigned(reg1397) : $unsigned(forvar1395)) ~^ $signed((reg1384 || reg1384))) * forvar1456[(2'h3):(2'h3)]);
                      reg1465 <= $unsigned(($signed((reg1440 ?
                              forvar1385 : (8'hb4))) ?
                          reg1447[(1'h0):(1'h0)] : (^~forvar1442)));
                      reg1466 <= ($unsigned(($signed(reg1460) ?
                          reg1386 : $unsigned(reg1426))) >= $unsigned($unsigned(reg1442[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  if (forvar1390)
                    begin
                      reg1456 <= $unsigned((8'ha7));
                    end
                  else
                    begin
                      reg1456 <= (forvar1456[(2'h3):(1'h1)] ?
                          reg1402 : (|(reg1404[(2'h3):(2'h3)] ?
                              (reg1429 ?
                                  reg1408 : (8'hae)) : $unsigned(reg1415))));
                    end
                  for (forvar1457 = (1'h0); (forvar1457 < (1'h1)); forvar1457 = (forvar1457 + (1'h1)))
                    begin
                      reg1458 <= ((^~reg1455[(4'hc):(3'h4)]) ?
                          (~((&reg1394) | (reg1393 ?
                              reg1418 : forvar1395))) : $signed(reg1400[(2'h2):(1'h0)]));
                    end
                  if ($signed(($unsigned($unsigned(wire1170)) >= $unsigned($signed(forvar1424)))))
                    begin
                      reg1459 <= $signed((reg1446[(3'h4):(1'h1)] <<< ({reg1456} < (~^(8'ha7)))));
                      reg1460 <= (forvar1383[(3'h5):(1'h1)] | $unsigned((((8'hb4) ?
                          forvar1442 : forvar1424) >>> (-reg1387))));
                      reg1461 <= (reg1386 ~^ $unsigned(reg1439));
                      reg1462 <= (^(((wire1171 ? reg1461 : reg1462) ?
                          (reg1466 ?
                              forvar1380 : reg1409) : reg1434[(3'h5):(2'h2)]) && reg1441[(4'ha):(3'h5)]));
                    end
                  else
                    begin
                      reg1459 <= ((reg1459 | {(forvar1379 ?
                                  forvar1407 : reg1450)}) ?
                          wire1170[(2'h3):(1'h0)] : (reg1461 ?
                              $signed(reg1451[(3'h4):(1'h1)]) : {forvar1425[(3'h4):(1'h0)]}));
                      reg1460 <= {$signed({reg1463[(4'h9):(1'h1)]})};
                      reg1461 <= ($unsigned(reg1457[(2'h2):(1'h0)]) >>> (~|{(~^reg1438)}));
                    end
                end
              reg1467 <= $unsigned($signed(((forvar1380 ? reg1381 : reg1432) ?
                  (~|wire1169) : $signed(reg1401))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1468 = (1'h0); (forvar1468 < (2'h2)); forvar1468 = (forvar1468 + (1'h1)))
        begin
          reg1469 <= reg1458;
          reg1470 <= $signed(reg1393);
        end
    end
  always
    @(posedge clk) begin
      reg1471 <= reg1415[(2'h2):(2'h2)];
      if ((forvar1381 * $signed(forvar1438)))
        begin
          for (forvar1472 = (1'h0); (forvar1472 < (1'h0)); forvar1472 = (forvar1472 + (1'h1)))
            begin
              if (((8'ha3) ?
                  $signed(reg1404[(2'h3):(2'h2)]) : ((|$unsigned(reg1463)) ^~ ((~reg1400) < {reg1462}))))
                begin
                  for (forvar1473 = (1'h0); (forvar1473 < (2'h3)); forvar1473 = (forvar1473 + (1'h1)))
                    begin
                      reg1474 <= $unsigned(reg1397[(5'h10):(3'h7)]);
                      reg1475 <= (8'hb2);
                      reg1476 <= reg1443[(2'h3):(1'h1)];
                      reg1477 <= reg1462[(2'h2):(2'h2)];
                    end
                  if ($signed(reg1428))
                    begin
                      reg1478 <= forvar1449[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg1478 <= ($signed($unsigned((reg1429 ~^ forvar1457))) ?
                          $unsigned((-{reg1416})) : $signed((!(reg1388 ?
                              reg1401 : (8'h9d)))));
                      reg1479 <= (forvar1438[(1'h1):(1'h1)] == $unsigned(((^~forvar1417) ?
                          reg1450[(2'h2):(2'h2)] : (~(8'ha8)))));
                      reg1480 <= (forvar1417[(4'hd):(3'h5)] ?
                          (~&reg1405[(3'h7):(1'h1)]) : forvar1449[(1'h1):(1'h1)]);
                      reg1481 <= (forvar1457[(4'h8):(1'h1)] ?
                          {(^~(&reg1429))} : forvar1385);
                    end
                  for (forvar1482 = (1'h0); (forvar1482 < (1'h0)); forvar1482 = (forvar1482 + (1'h1)))
                    begin
                      reg1483 <= (8'hb6);
                    end
                end
              else
                begin
                  if ((forvar1482 && ($signed(reg1431) + ((~&reg1458) ?
                      forvar1456 : (^reg1409)))))
                    begin
                      reg1473 <= (reg1398[(4'ha):(1'h0)] ?
                          forvar1457 : reg1455);
                      reg1474 <= (((((8'hb5) || reg1413) ?
                              (reg1397 ^ reg1411) : (8'haa)) ?
                          reg1401 : reg1393) << $unsigned($unsigned(((8'ha1) ?
                          reg1435 : reg1459))));
                      reg1475 <= {$signed(($signed(reg1415) | reg1451[(4'ha):(3'h5)]))};
                    end
                  else
                    begin
                      reg1473 <= (reg1464 ~^ (wire1171[(2'h3):(2'h2)] ?
                          (((8'ha4) ? (8'h9f) : reg1465) ?
                              {(8'haa)} : $unsigned((8'h9e))) : $unsigned((~^reg1392))));
                      reg1474 <= {$unsigned(reg1386[(2'h2):(1'h0)])};
                    end
                  if ((($signed(forvar1383[(3'h4):(2'h3)]) >>> (&$unsigned(reg1427))) >= reg1386[(1'h1):(1'h0)]))
                    begin
                      reg1476 <= {{(!wire1170)}};
                      reg1477 <= (~|((^(8'hac)) ^ (|wire1169)));
                    end
                  else
                    begin
                      reg1476 <= reg1405[(4'h8):(1'h1)];
                      reg1477 <= reg1447[(4'hb):(3'h7)];
                      reg1478 <= $signed((((|reg1481) ?
                              reg1429[(2'h3):(2'h2)] : reg1428[(3'h4):(1'h1)]) ?
                          (~^(reg1454 <<< forvar1417)) : $signed(reg1415)));
                    end
                  for (forvar1479 = (1'h0); (forvar1479 < (1'h0)); forvar1479 = (forvar1479 + (1'h1)))
                    begin
                      reg1480 <= (|(~&forvar1390));
                    end
                end
              for (forvar1484 = (1'h0); (forvar1484 < (1'h1)); forvar1484 = (forvar1484 + (1'h1)))
                begin
                  for (forvar1485 = (1'h0); (forvar1485 < (2'h3)); forvar1485 = (forvar1485 + (1'h1)))
                    begin
                      reg1486 <= ($signed(reg1444[(3'h5):(2'h3)]) ?
                          ($signed($signed((8'ha4))) <= ($unsigned(reg1480) ~^ (reg1415 || reg1386))) : ({forvar1433} & forvar1457));
                      reg1487 <= $signed(reg1479);
                    end
                end
              if (reg1447[(4'h8):(3'h7)])
                begin
                  reg1488 <= (({(^~reg1416)} ?
                      ($signed(reg1475) ?
                          $signed((8'h9e)) : (reg1453 ?
                              forvar1484 : reg1439)) : $unsigned(reg1487[(3'h5):(1'h1)])) ^~ (^~(forvar1482 - $unsigned(reg1444))));
                  for (forvar1489 = (1'h0); (forvar1489 < (1'h0)); forvar1489 = (forvar1489 + (1'h1)))
                    begin
                      reg1490 <= ($unsigned($unsigned(((8'hb7) | forvar1438))) ?
                          wire1170 : forvar1395);
                      reg1491 <= reg1391[(3'h5):(3'h5)];
                      reg1492 <= ((8'h9c) && reg1457);
                      reg1493 <= (reg1420 ?
                          ((reg1477[(1'h1):(1'h1)] ^~ (reg1481 ?
                                  reg1479 : (8'hb9))) ?
                              ($signed(reg1413) << reg1381[(3'h5):(2'h3)]) : forvar1383) : (($unsigned((8'ha2)) | (reg1467 <= reg1453)) ?
                              (forvar1468 + $unsigned(forvar1438)) : $signed((reg1396 >= reg1442))));
                    end
                end
              else
                begin
                  if ((^~$signed($unsigned(forvar1472))))
                    begin
                      reg1488 <= ((~|(&(reg1387 ?
                          forvar1485 : (8'hae)))) || $unsigned($signed((^~(8'hb8)))));
                      reg1489 <= $unsigned({$unsigned((^forvar1406))});
                    end
                  else
                    begin
                      reg1488 <= (8'hac);
                      reg1489 <= reg1446[(4'h9):(1'h1)];
                    end
                  for (forvar1490 = (1'h0); (forvar1490 < (1'h1)); forvar1490 = (forvar1490 + (1'h1)))
                    begin
                      reg1491 <= $signed(forvar1436);
                    end
                  for (forvar1492 = (1'h0); (forvar1492 < (2'h3)); forvar1492 = (forvar1492 + (1'h1)))
                    begin
                      reg1493 <= (-(reg1415 && $unsigned((forvar1482 <<< reg1469))));
                      reg1494 <= forvar1482[(4'h8):(3'h4)];
                      reg1495 <= (~^{($unsigned(reg1459) >= forvar1396)});
                    end
                end
              for (forvar1496 = (1'h0); (forvar1496 < (2'h3)); forvar1496 = (forvar1496 + (1'h1)))
                begin
                  for (forvar1497 = (1'h0); (forvar1497 < (2'h2)); forvar1497 = (forvar1497 + (1'h1)))
                    begin
                      reg1498 <= {$signed($signed(((8'ha4) <<< forvar1425)))};
                    end
                  if ($signed($unsigned(((reg1443 ? (8'hb3) : forvar1437) ?
                      $signed(reg1395) : $signed(reg1395)))))
                    begin
                      reg1499 <= (^$signed($signed(reg1390)));
                      reg1500 <= ($signed((^~(forvar1425 & reg1481))) >> $signed((reg1459[(4'hd):(3'h7)] ?
                          reg1458 : {reg1403})));
                    end
                  else
                    begin
                      reg1499 <= {{((~reg1430) + (forvar1485 >> reg1469))}};
                      reg1500 <= reg1478;
                    end
                  reg1501 <= forvar1437;
                  if (($unsigned($signed((reg1421 ?
                      reg1461 : reg1400))) - ($unsigned($unsigned(reg1483)) >= ((|forvar1387) <<< ((8'h9d) << reg1434)))))
                    begin
                      reg1502 <= $unsigned($unsigned((^(reg1409 ?
                          reg1389 : reg1395))));
                      reg1503 <= (&(!(&(forvar1417 <<< reg1405))));
                    end
                  else
                    begin
                      reg1502 <= $unsigned((|((reg1393 ?
                          reg1447 : forvar1485) ^~ reg1386)));
                    end
                end
            end
        end
      else
        begin
          for (forvar1472 = (1'h0); (forvar1472 < (2'h3)); forvar1472 = (forvar1472 + (1'h1)))
            begin
              if ($unsigned(forvar1383))
                begin
                  for (forvar1473 = (1'h0); (forvar1473 < (1'h0)); forvar1473 = (forvar1473 + (1'h1)))
                    begin
                      reg1474 <= ($unsigned($unsigned($unsigned(reg1403))) >>> (reg1470[(4'hb):(4'ha)] ?
                          reg1402 : $signed((forvar1457 || reg1447))));
                      reg1475 <= $signed(reg1457[(1'h1):(1'h0)]);
                      reg1476 <= ({$unsigned(reg1410[(3'h6):(3'h4)])} <= reg1446[(4'hc):(3'h7)]);
                      reg1477 <= $signed(reg1503[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar1473 = (1'h0); (forvar1473 < (1'h0)); forvar1473 = (forvar1473 + (1'h1)))
                    begin
                      reg1474 <= (~^$signed((reg1501 ?
                          (forvar1485 ?
                              reg1387 : reg1498) : (wire1168 >>> forvar1433))));
                    end
                  if ((reg1381 ?
                      $signed({$unsigned((8'hb3))}) : $signed($signed((~&forvar1437)))))
                    begin
                      reg1475 <= reg1381[(2'h2):(1'h1)];
                      reg1476 <= {reg1390[(4'ha):(1'h0)]};
                      reg1477 <= forvar1442;
                      reg1478 <= (-{$unsigned((~forvar1380))});
                    end
                  else
                    begin
                      reg1475 <= reg1492[(4'hd):(4'hd)];
                    end
                end
              if ((^~(~(+$signed(forvar1437)))))
                begin
                  if (forvar1482)
                    begin
                      reg1479 <= reg1476;
                      reg1480 <= $unsigned($signed(reg1458[(1'h1):(1'h0)]));
                      reg1481 <= {$signed((~&(8'hb4)))};
                    end
                  else
                    begin
                      reg1479 <= $signed(($signed({reg1381}) ?
                          $unsigned(reg1408[(1'h0):(1'h0)]) : $unsigned($signed(reg1421))));
                      reg1480 <= $signed((wire1171 & ((forvar1424 >> (8'hb8)) ?
                          (~^reg1489) : forvar1461[(2'h3):(2'h2)])));
                    end
                end
              else
                begin
                  for (forvar1479 = (1'h0); (forvar1479 < (1'h0)); forvar1479 = (forvar1479 + (1'h1)))
                    begin
                      reg1480 <= $unsigned(((-(reg1379 ? reg1380 : reg1462)) ?
                          (-$unsigned(reg1388)) : $signed((~|forvar1456))));
                    end
                  for (forvar1481 = (1'h0); (forvar1481 < (2'h2)); forvar1481 = (forvar1481 + (1'h1)))
                    begin
                      reg1482 <= $unsigned($signed(reg1409));
                      reg1483 <= reg1397;
                      reg1484 <= (~&({forvar1387} ?
                          (forvar1436 ?
                              (~|(8'hae)) : (reg1390 ?
                                  (8'h9d) : forvar1490)) : $signed(reg1399[(3'h6):(3'h5)])));
                      reg1485 <= $signed(reg1501[(2'h2):(1'h1)]);
                    end
                  if ($signed((8'ha1)))
                    begin
                      reg1486 <= (reg1478 <<< (-(^~$signed(forvar1383))));
                      reg1487 <= (reg1458[(4'h9):(2'h2)] ?
                          (+reg1415) : $unsigned((reg1494[(3'h4):(3'h4)] ?
                              $signed(reg1415) : reg1403)));
                      reg1488 <= forvar1414[(3'h5):(2'h3)];
                      reg1489 <= (forvar1456[(1'h0):(1'h0)] | reg1442[(4'h8):(2'h3)]);
                    end
                  else
                    begin
                      reg1486 <= $unsigned((reg1434 - $unsigned(reg1485[(2'h3):(2'h3)])));
                      reg1487 <= (((~reg1491[(2'h2):(1'h1)]) ?
                              (reg1478[(3'h4):(2'h2)] ?
                                  (forvar1457 | reg1467) : (reg1478 ?
                                      reg1384 : forvar1438)) : $unsigned((~|reg1480))) ?
                          {(reg1411 ?
                                  reg1403 : {reg1478})} : reg1434[(2'h2):(1'h1)]);
                      reg1488 <= (reg1384[(4'hd):(4'hd)] ?
                          $unsigned($unsigned((^~reg1501))) : {reg1410[(3'h5):(2'h3)]});
                    end
                  if ($signed((^$signed((!reg1400)))))
                    begin
                      reg1490 <= $signed(reg1411[(1'h0):(1'h0)]);
                      reg1491 <= $unsigned($signed((~&reg1431[(3'h5):(2'h3)])));
                    end
                  else
                    begin
                      reg1490 <= reg1393[(4'h9):(1'h1)];
                      reg1491 <= ($unsigned({(~forvar1390)}) ?
                          ((~^reg1459[(4'h8):(3'h4)]) < (8'hb4)) : reg1393);
                      reg1492 <= ((((reg1385 | forvar1461) ?
                              {(8'hb8)} : $signed(forvar1449)) | (~|$signed(reg1452))) ?
                          (~^(8'ha9)) : reg1404);
                      reg1493 <= ((~&reg1405) ?
                          ({((8'ha8) ? reg1450 : reg1445)} ?
                              $signed($signed(forvar1414)) : reg1381[(3'h5):(3'h5)]) : (&(~(~reg1486))));
                    end
                end
              for (forvar1494 = (1'h0); (forvar1494 < (1'h0)); forvar1494 = (forvar1494 + (1'h1)))
                begin
                  if ((($unsigned((reg1380 ? forvar1490 : (8'hba))) ?
                      ($signed(reg1487) > reg1481[(1'h0):(1'h0)]) : forvar1383) >> ($signed($unsigned((8'ha0))) >>> $signed(reg1418))))
                    begin
                      reg1495 <= {reg1490};
                      reg1496 <= (^$signed({$unsigned(forvar1456)}));
                      reg1497 <= (~&reg1467);
                      reg1498 <= (~|($signed(forvar1473[(2'h3):(1'h1)]) ?
                          (+(^~reg1405)) : ((~&reg1488) ?
                              reg1494[(2'h2):(2'h2)] : $signed(reg1394))));
                    end
                  else
                    begin
                      reg1495 <= $signed($unsigned($unsigned((~reg1466))));
                      reg1496 <= (+$signed($unsigned((forvar1380 ^ forvar1381))));
                      reg1497 <= ((wire1172[(1'h0):(1'h0)] << (|$unsigned(forvar1472))) ^ {(!(reg1499 << forvar1407))});
                      reg1498 <= reg1413;
                    end
                  if (reg1463)
                    begin
                      reg1499 <= $signed(forvar1482[(4'hc):(4'h9)]);
                      reg1500 <= reg1452[(1'h0):(1'h0)];
                      reg1501 <= {reg1440};
                    end
                  else
                    begin
                      reg1499 <= $signed((&(~&(8'hb7))));
                      reg1500 <= (reg1439 >> $unsigned({(&reg1483)}));
                      reg1501 <= $signed((~^$unsigned($unsigned((8'h9f)))));
                    end
                end
              if (((reg1487 ?
                  (~^(reg1439 | reg1385)) : ((forvar1396 ~^ (8'hb8)) ?
                      reg1447 : (8'ha3))) && $signed($unsigned((forvar1383 ?
                  reg1441 : wire1377)))))
                begin
                  for (forvar1502 = (1'h0); (forvar1502 < (1'h1)); forvar1502 = (forvar1502 + (1'h1)))
                    begin
                      reg1503 <= reg1441[(3'h4):(1'h1)];
                      reg1504 <= (!{(8'ha7)});
                      reg1505 <= (~&$signed({$unsigned(forvar1490)}));
                      reg1506 <= $signed(reg1460);
                    end
                end
              else
                begin
                  for (forvar1502 = (1'h0); (forvar1502 < (1'h1)); forvar1502 = (forvar1502 + (1'h1)))
                    begin
                      reg1503 <= (($signed((+(8'ha8))) <<< $signed((reg1405 ?
                              reg1487 : reg1455))) ?
                          ($signed((reg1385 ?
                              (8'ha4) : forvar1485)) & (+$signed(reg1402))) : ({reg1456} ?
                              reg1493 : (~^(&forvar1496))));
                    end
                  if (reg1464[(2'h2):(1'h1)])
                    begin
                      reg1504 <= $unsigned(forvar1407);
                      reg1505 <= (($signed((forvar1379 ? reg1401 : reg1462)) ?
                              reg1492[(4'hc):(2'h3)] : {(|reg1392)}) ?
                          reg1432 : $unsigned($unsigned((reg1431 ?
                              reg1483 : reg1477))));
                    end
                  else
                    begin
                      reg1504 <= forvar1484[(3'h5):(3'h5)];
                      reg1505 <= forvar1380;
                      reg1506 <= reg1442[(2'h2):(2'h2)];
                      reg1507 <= reg1471[(2'h3):(1'h0)];
                    end
                  reg1508 <= $unsigned({(reg1381[(4'h8):(4'h8)] | wire1172[(4'hb):(2'h2)])});
                  for (forvar1509 = (1'h0); (forvar1509 < (2'h2)); forvar1509 = (forvar1509 + (1'h1)))
                    begin
                      reg1510 <= $unsigned(reg1466);
                      reg1511 <= (+reg1426[(2'h3):(2'h3)]);
                      reg1512 <= reg1422[(4'h8):(2'h3)];
                    end
                end
            end
        end
      for (forvar1513 = (1'h0); (forvar1513 < (2'h2)); forvar1513 = (forvar1513 + (1'h1)))
        begin
          for (forvar1514 = (1'h0); (forvar1514 < (2'h2)); forvar1514 = (forvar1514 + (1'h1)))
            begin
              for (forvar1515 = (1'h0); (forvar1515 < (2'h3)); forvar1515 = (forvar1515 + (1'h1)))
                begin
                  if (reg1395[(1'h1):(1'h0)])
                    begin
                      reg1516 <= $signed(reg1467);
                      reg1517 <= (~reg1398[(1'h1):(1'h0)]);
                      reg1518 <= $unsigned((reg1397 ?
                          reg1502[(4'hc):(4'ha)] : (~^(reg1403 ?
                              reg1506 : reg1418))));
                      reg1519 <= reg1421;
                    end
                  else
                    begin
                      reg1516 <= $signed(forvar1515[(2'h3):(1'h1)]);
                      reg1517 <= reg1519;
                      reg1518 <= $unsigned($unsigned((8'hb1)));
                      reg1519 <= {(~&$unsigned({forvar1497}))};
                    end
                  if ({reg1455[(3'h4):(1'h1)]})
                    begin
                      reg1520 <= (forvar1379[(1'h0):(1'h0)] ?
                          ($unsigned(((8'hb1) && wire1171)) ~^ {(wire1168 ?
                                  reg1381 : forvar1481)}) : ({(~|(8'hb0))} ?
                              ((~&reg1475) >>> $signed(reg1518)) : reg1494));
                    end
                  else
                    begin
                      reg1520 <= (reg1439[(2'h2):(2'h2)] ?
                          {reg1390[(4'hc):(4'hc)]} : $unsigned(($unsigned(reg1396) <= $unsigned((8'h9f)))));
                      reg1521 <= ($signed(forvar1407[(5'h10):(4'hb)]) ?
                          reg1396[(2'h2):(2'h2)] : ($signed((reg1507 + reg1455)) ?
                              $unsigned(forvar1407[(4'h8):(2'h2)]) : ($signed(reg1395) ?
                                  reg1507 : (reg1416 ? (8'hb0) : reg1431))));
                      reg1522 <= (~reg1489[(2'h2):(1'h0)]);
                    end
                  for (forvar1523 = (1'h0); (forvar1523 < (1'h1)); forvar1523 = (forvar1523 + (1'h1)))
                    begin
                      reg1524 <= {(8'ha0)};
                    end
                end
              if (($unsigned((+(forvar1479 >> reg1498))) - $unsigned(reg1411[(3'h6):(3'h6)])))
                begin
                  for (forvar1525 = (1'h0); (forvar1525 < (1'h1)); forvar1525 = (forvar1525 + (1'h1)))
                    begin
                      reg1526 <= forvar1456;
                      reg1527 <= (|({(forvar1515 <= forvar1406)} != $signed($unsigned((8'h9e)))));
                      reg1528 <= $signed((8'hba));
                      reg1529 <= (-((8'h9f) && $signed($signed(forvar1497))));
                    end
                end
              else
                begin
                  if ($signed($signed(forvar1490)))
                    begin
                      reg1525 <= (~&{reg1391[(5'h10):(4'he)]});
                      reg1526 <= $signed(((^~(forvar1515 + wire1169)) <<< $unsigned({reg1455})));
                    end
                  else
                    begin
                      reg1525 <= (+(|($unsigned(reg1402) ?
                          (!(8'ha0)) : reg1440[(1'h1):(1'h0)])));
                      reg1526 <= reg1385[(3'h6):(3'h6)];
                      reg1527 <= reg1447[(4'he):(4'ha)];
                      reg1528 <= (~|($signed(reg1476) ?
                          reg1474[(3'h4):(2'h3)] : ($signed(reg1398) >> (8'had))));
                    end
                  reg1529 <= $signed((8'hb7));
                  reg1530 <= ((reg1508 != ($signed(reg1386) ?
                      (reg1463 ? reg1443 : reg1474) : (reg1465 ?
                          forvar1424 : reg1405))) > reg1386[(1'h0):(1'h0)]);
                  for (forvar1531 = (1'h0); (forvar1531 < (2'h2)); forvar1531 = (forvar1531 + (1'h1)))
                    begin
                      reg1532 <= $signed((|($signed(reg1525) > $unsigned(reg1391))));
                      reg1533 <= (^~reg1440[(3'h5):(3'h5)]);
                    end
                end
              for (forvar1534 = (1'h0); (forvar1534 < (1'h1)); forvar1534 = (forvar1534 + (1'h1)))
                begin
                  for (forvar1535 = (1'h0); (forvar1535 < (1'h0)); forvar1535 = (forvar1535 + (1'h1)))
                    begin
                      reg1536 <= $signed((^~reg1411));
                    end
                  reg1537 <= forvar1390;
                end
            end
          if ($signed(({(&reg1518)} ? ((!reg1486) >>> {reg1421}) : forvar1406)))
            begin
              for (forvar1538 = (1'h0); (forvar1538 < (2'h2)); forvar1538 = (forvar1538 + (1'h1)))
                begin
                  if ((reg1518 * (+reg1525)))
                    begin
                      reg1539 <= reg1393[(1'h1):(1'h0)];
                      reg1540 <= ($signed(({reg1441} || reg1470[(2'h2):(2'h2)])) ?
                          reg1524 : forvar1385[(4'h8):(4'h8)]);
                    end
                  else
                    begin
                      reg1539 <= ((((forvar1479 <<< reg1429) ?
                          forvar1485 : $unsigned(reg1390)) <= $unsigned($signed(forvar1407))) || $signed(reg1527));
                      reg1540 <= {$unsigned($unsigned((reg1443 >= reg1459)))};
                      reg1541 <= reg1461;
                    end
                  reg1542 <= {$unsigned((-$signed(forvar1484)))};
                  if (($signed({(reg1432 != reg1405)}) ?
                      forvar1489 : {$signed(reg1536)}))
                    begin
                      reg1543 <= (((reg1516 | $signed((8'hb0))) || reg1396) ?
                          (!((reg1440 ? reg1474 : reg1490) ?
                              reg1411 : $signed(forvar1494))) : reg1479);
                      reg1544 <= $unsigned(($unsigned((reg1426 >> reg1537)) >> {(forvar1473 ^~ reg1517)}));
                      reg1545 <= reg1498;
                      reg1546 <= ((~&($unsigned(reg1475) >>> reg1495)) || reg1544[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1543 <= ((((+forvar1479) == $unsigned(reg1396)) ?
                              ($unsigned(reg1435) ?
                                  {(8'hb7)} : reg1473[(3'h5):(2'h2)]) : ((^~reg1440) < (|reg1388))) ?
                          $signed(($unsigned(reg1527) ^ (forvar1442 ?
                              reg1427 : forvar1468))) : $unsigned(((~|forvar1482) <<< $signed(forvar1417))));
                    end
                end
              reg1547 <= ((^~$signed((|reg1507))) * ($unsigned(forvar1379[(4'hf):(2'h2)]) & $unsigned((8'ha3))));
              if ($unsigned(forvar1497))
                begin
                  reg1548 <= $signed(($signed((^forvar1525)) | ((forvar1514 ?
                          reg1410 : (8'hb7)) ?
                      $signed((8'haa)) : $unsigned(reg1540))));
                  for (forvar1549 = (1'h0); (forvar1549 < (2'h3)); forvar1549 = (forvar1549 + (1'h1)))
                    begin
                      reg1550 <= $unsigned($unsigned(((reg1476 ?
                              reg1539 : reg1503) ?
                          (reg1381 == reg1491) : (8'ha2))));
                      reg1551 <= reg1539;
                      reg1552 <= reg1429[(3'h4):(2'h3)];
                    end
                  for (forvar1553 = (1'h0); (forvar1553 < (1'h0)); forvar1553 = (forvar1553 + (1'h1)))
                    begin
                      reg1554 <= reg1440[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar1548 = (1'h0); (forvar1548 < (1'h0)); forvar1548 = (forvar1548 + (1'h1)))
                    begin
                      reg1549 <= (reg1491 * (reg1498 <<< reg1479));
                      reg1550 <= reg1451[(2'h3):(1'h0)];
                      reg1551 <= (forvar1494[(4'hd):(4'ha)] ?
                          ($unsigned(reg1390[(4'hb):(3'h5)]) ?
                              (reg1408[(1'h0):(1'h0)] * (8'hb6)) : {reg1552}) : $signed(($signed(reg1452) ?
                              reg1549[(1'h0):(1'h0)] : $unsigned(wire1170))));
                      reg1552 <= (-$unsigned($signed((reg1429 ^ (8'had)))));
                    end
                end
            end
          else
            begin
              for (forvar1538 = (1'h0); (forvar1538 < (1'h0)); forvar1538 = (forvar1538 + (1'h1)))
                begin
                  if ({$unsigned((((8'hb9) && reg1512) * (~&wire1169)))})
                    begin
                      reg1539 <= (($signed($signed((8'hb9))) ?
                          $signed({forvar1449}) : (+forvar1523[(1'h1):(1'h1)])) || reg1539[(4'ha):(4'h8)]);
                      reg1540 <= ($unsigned($unsigned(reg1478[(2'h2):(1'h1)])) ?
                          forvar1423[(4'h9):(3'h7)] : {$signed((reg1548 ?
                                  reg1443 : reg1487))});
                      reg1541 <= $unsigned((~|reg1520));
                      reg1542 <= (-$unsigned({(!(8'hb0))}));
                    end
                  else
                    begin
                      reg1539 <= ((~&$unsigned((reg1537 + forvar1473))) ~^ (&$signed($signed(reg1489))));
                    end
                  reg1543 <= (((forvar1534 * (8'hb3)) ?
                      (reg1404[(2'h3):(2'h3)] ?
                          (8'haf) : reg1382[(3'h4):(2'h3)]) : forvar1456) + ($signed(forvar1387[(1'h0):(1'h0)]) ?
                      $signed(reg1405[(2'h2):(1'h1)]) : {(reg1539 > forvar1456)}));
                  for (forvar1544 = (1'h0); (forvar1544 < (1'h0)); forvar1544 = (forvar1544 + (1'h1)))
                    begin
                      reg1545 <= $signed(($signed((reg1456 ?
                          reg1435 : reg1521)) && reg1482[(4'hc):(2'h2)]));
                      reg1546 <= {(((8'h9c) ?
                              reg1413[(2'h2):(2'h2)] : (wire1171 && reg1464)) != forvar1390[(1'h0):(1'h0)])};
                    end
                end
              for (forvar1547 = (1'h0); (forvar1547 < (2'h2)); forvar1547 = (forvar1547 + (1'h1)))
                begin
                  if ((({reg1506[(3'h5):(1'h0)]} != reg1476[(3'h4):(2'h3)]) ?
                      $signed(((reg1389 ^~ reg1490) ?
                          {reg1438} : reg1427[(4'hf):(4'hf)])) : forvar1472[(1'h1):(1'h1)]))
                    begin
                      reg1548 <= (reg1447 == $signed(((reg1459 ?
                              wire1169 : reg1544) ?
                          $signed(reg1466) : {forvar1496})));
                      reg1549 <= (~&($unsigned({reg1413}) ?
                          forvar1535[(4'hb):(1'h0)] : reg1494[(2'h3):(1'h0)]));
                      reg1550 <= {(8'ha7)};
                    end
                  else
                    begin
                      reg1548 <= ((!reg1456[(3'h6):(3'h5)]) ?
                          $signed({reg1461[(1'h1):(1'h1)]}) : reg1487);
                      reg1549 <= ((reg1460 ?
                              $signed($signed(reg1452)) : $unsigned(wire1169)) ?
                          (($unsigned(reg1533) != (~^reg1485)) ?
                              reg1546 : {$signed(reg1493)}) : forvar1489);
                      reg1550 <= ($signed((reg1463 ^~ $signed(reg1499))) <<< ((^(^~reg1485)) < (~|reg1421)));
                      reg1551 <= $signed(reg1464);
                    end
                  for (forvar1552 = (1'h0); (forvar1552 < (2'h2)); forvar1552 = (forvar1552 + (1'h1)))
                    begin
                      reg1553 <= ($unsigned($unsigned(reg1398)) ?
                          ($signed((~|reg1494)) ?
                              forvar1442 : (~$unsigned(forvar1534))) : (~&(((8'hac) ~^ reg1470) ?
                              $unsigned(reg1439) : {(8'ha0)})));
                      reg1554 <= (((+$unsigned(reg1445)) <= (~$unsigned(forvar1407))) ?
                          $unsigned($unsigned($unsigned(reg1518))) : ((^{forvar1489}) ?
                              $unsigned((reg1455 ?
                                  forvar1494 : reg1458)) : ($unsigned(reg1455) > reg1529[(2'h2):(1'h1)])));
                    end
                  reg1555 <= (reg1411[(3'h5):(2'h3)] << (^~$signed(reg1459)));
                  for (forvar1556 = (1'h0); (forvar1556 < (1'h1)); forvar1556 = (forvar1556 + (1'h1)))
                    begin
                      reg1557 <= ((reg1504 > ($signed(reg1466) * $signed((8'hac)))) ?
                          reg1477 : {(&(&reg1517))});
                      reg1558 <= (&reg1516[(1'h0):(1'h0)]);
                      reg1559 <= $signed((((reg1442 ? reg1553 : forvar1425) ?
                              {reg1522} : $unsigned(reg1461)) ?
                          reg1553 : ((^reg1464) ? (~^forvar1461) : {reg1489})));
                      reg1560 <= forvar1502;
                    end
                end
              reg1561 <= {{$unsigned(forvar1383[(3'h6):(1'h0)])}};
            end
        end
      for (forvar1562 = (1'h0); (forvar1562 < (1'h0)); forvar1562 = (forvar1562 + (1'h1)))
        begin
          if (reg1390)
            begin
              reg1563 <= {$unsigned($unsigned(reg1471[(2'h3):(2'h2)]))};
              for (forvar1564 = (1'h0); (forvar1564 < (1'h1)); forvar1564 = (forvar1564 + (1'h1)))
                begin
                  for (forvar1565 = (1'h0); (forvar1565 < (1'h1)); forvar1565 = (forvar1565 + (1'h1)))
                    begin
                      reg1566 <= reg1502;
                    end
                  reg1567 <= ($signed(reg1505) ?
                      $signed((reg1398[(2'h2):(1'h1)] ?
                          $signed(reg1421) : $signed((8'h9f)))) : $unsigned(forvar1482[(3'h4):(1'h0)]));
                  for (forvar1568 = (1'h0); (forvar1568 < (1'h1)); forvar1568 = (forvar1568 + (1'h1)))
                    begin
                      reg1569 <= reg1435[(4'h8):(2'h3)];
                      reg1570 <= (&$unsigned(reg1408[(1'h0):(1'h0)]));
                    end
                end
              for (forvar1571 = (1'h0); (forvar1571 < (2'h2)); forvar1571 = (forvar1571 + (1'h1)))
                begin
                  for (forvar1572 = (1'h0); (forvar1572 < (2'h2)); forvar1572 = (forvar1572 + (1'h1)))
                    begin
                      reg1573 <= $unsigned((~^$unsigned((reg1438 ?
                          reg1460 : forvar1472))));
                    end
                  if (($unsigned(reg1485[(4'h9):(4'h9)]) * (+((reg1541 ?
                          (8'ha1) : forvar1385) ?
                      (reg1569 ?
                          forvar1485 : forvar1548) : reg1504[(1'h0):(1'h0)]))))
                    begin
                      reg1574 <= ((((&reg1387) ?
                              (|reg1386) : $signed(reg1516)) ?
                          $unsigned(reg1480) : (^{reg1501})) && {(~^reg1527)});
                    end
                  else
                    begin
                      reg1574 <= forvar1381;
                      reg1575 <= $signed((reg1475[(1'h1):(1'h1)] < $unsigned(forvar1457[(3'h5):(2'h3)])));
                      reg1576 <= reg1442;
                    end
                end
              if (($signed($signed((~^reg1524))) * forvar1496))
                begin
                  if ($signed({((forvar1442 << reg1508) <= $signed(reg1503))}))
                    begin
                      reg1577 <= forvar1383[(1'h1):(1'h0)];
                      reg1578 <= $unsigned(reg1486);
                      reg1579 <= $signed($unsigned((&$signed((8'ha4)))));
                    end
                  else
                    begin
                      reg1577 <= ((|$signed((~(8'hb2)))) && ((reg1462 > reg1458) ?
                          ((reg1469 << reg1508) ?
                              (reg1494 ?
                                  forvar1436 : reg1511) : reg1455[(1'h0):(1'h0)]) : forvar1538));
                      reg1578 <= forvar1385;
                    end
                end
              else
                begin
                  reg1577 <= wire1377;
                  if (forvar1481[(3'h5):(1'h1)])
                    begin
                      reg1578 <= reg1442[(3'h6):(3'h4)];
                      reg1579 <= (~|$signed(((reg1566 << (8'had)) ?
                          $signed(reg1399) : (~^forvar1497))));
                      reg1580 <= forvar1381[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1578 <= (reg1399 ?
                          $unsigned(((+reg1491) ?
                              $unsigned(forvar1383) : (~^reg1454))) : forvar1414[(4'hc):(1'h1)]);
                      reg1579 <= ($unsigned($unsigned(reg1559)) ?
                          reg1413 : wire1168);
                    end
                  for (forvar1581 = (1'h0); (forvar1581 < (1'h0)); forvar1581 = (forvar1581 + (1'h1)))
                    begin
                      reg1582 <= (^~($signed(reg1440) ?
                          ((8'hac) < $signed(reg1574)) : reg1489));
                      reg1583 <= (|reg1552);
                      reg1584 <= (({$unsigned(reg1557)} ?
                          {$unsigned(reg1427)} : (~{(8'hba)})) ^~ forvar1549[(4'hb):(4'ha)]);
                    end
                  for (forvar1585 = (1'h0); (forvar1585 < (2'h3)); forvar1585 = (forvar1585 + (1'h1)))
                    begin
                      reg1586 <= ($signed((!reg1446[(2'h2):(1'h0)])) <<< forvar1433);
                      reg1587 <= $signed(reg1577);
                    end
                end
            end
          else
            begin
              if (reg1493[(4'ha):(2'h2)])
                begin
                  if ((reg1517[(1'h1):(1'h0)] << (8'hb4)))
                    begin
                      reg1563 <= {{reg1403}};
                      reg1564 <= ({(~&reg1510[(4'h8):(2'h2)])} ?
                          $signed((8'hb3)) : $signed($signed((reg1525 & reg1389))));
                      reg1565 <= ((~^$signed((|(8'hb6)))) || (((reg1545 ?
                                  reg1458 : reg1537) ?
                              (forvar1481 ? reg1466 : reg1530) : (reg1573 ?
                                  reg1467 : wire1170)) ?
                          (~|(~(8'ha9))) : reg1578[(3'h6):(3'h4)]));
                      reg1566 <= $unsigned(((&(~|reg1397)) ?
                          $unsigned(reg1476) : $unsigned((forvar1552 ~^ (8'had)))));
                    end
                  else
                    begin
                      reg1563 <= (^~$signed(($signed(reg1524) ?
                          forvar1562[(2'h2):(2'h2)] : reg1578)));
                    end
                  for (forvar1567 = (1'h0); (forvar1567 < (1'h0)); forvar1567 = (forvar1567 + (1'h1)))
                    begin
                      reg1568 <= {((^reg1389[(4'he):(4'h8)]) <<< $signed((8'hb7)))};
                      reg1569 <= $signed((($unsigned(reg1396) ~^ $signed(reg1564)) ?
                          $signed({reg1452}) : (^(reg1505 ?
                              reg1477 : reg1427))));
                      reg1570 <= ($unsigned(reg1415) > (forvar1425 ?
                          $signed((reg1441 ? (8'hba) : reg1536)) : (8'hb2)));
                    end
                end
              else
                begin
                  if (forvar1449)
                    begin
                      reg1563 <= $signed((((reg1519 ?
                          (8'ha8) : reg1454) ^~ $unsigned((8'hac))) ~^ (~&$unsigned(reg1408))));
                    end
                  else
                    begin
                      reg1563 <= $unsigned(reg1536[(1'h1):(1'h0)]);
                    end
                end
              for (forvar1571 = (1'h0); (forvar1571 < (2'h2)); forvar1571 = (forvar1571 + (1'h1)))
                begin
                  for (forvar1572 = (1'h0); (forvar1572 < (2'h2)); forvar1572 = (forvar1572 + (1'h1)))
                    begin
                      reg1573 <= (^reg1385[(1'h1):(1'h0)]);
                      reg1574 <= $unsigned({$unsigned((forvar1548 ?
                              reg1427 : reg1389))});
                      reg1575 <= (($unsigned(forvar1482) ?
                          $signed(reg1463) : {(reg1533 < (8'hba))}) & ((8'ha2) != (^(~|reg1573))));
                    end
                  for (forvar1576 = (1'h0); (forvar1576 < (2'h3)); forvar1576 = (forvar1576 + (1'h1)))
                    begin
                      reg1577 <= $signed(forvar1562);
                    end
                end
            end
          for (forvar1588 = (1'h0); (forvar1588 < (1'h0)); forvar1588 = (forvar1588 + (1'h1)))
            begin
              reg1589 <= ($unsigned($unsigned($signed(reg1456))) ^~ reg1452);
            end
          if (forvar1468)
            begin
              reg1590 <= $signed(reg1528[(4'hc):(1'h0)]);
            end
          else
            begin
              for (forvar1590 = (1'h0); (forvar1590 < (2'h2)); forvar1590 = (forvar1590 + (1'h1)))
                begin
                  for (forvar1591 = (1'h0); (forvar1591 < (2'h3)); forvar1591 = (forvar1591 + (1'h1)))
                    begin
                      reg1592 <= (8'h9c);
                      reg1593 <= ((8'hae) <<< reg1583);
                      reg1594 <= reg1557[(1'h0):(1'h0)];
                      reg1595 <= $signed({reg1401[(1'h1):(1'h1)]});
                    end
                end
            end
          if ((8'h9e))
            begin
              if ($unsigned((-$unsigned((~^wire1377)))))
                begin
                  reg1596 <= $signed($signed(forvar1513));
                  for (forvar1597 = (1'h0); (forvar1597 < (2'h3)); forvar1597 = (forvar1597 + (1'h1)))
                    begin
                      reg1598 <= $signed(forvar1379);
                      reg1599 <= {(($signed(reg1569) ?
                                  forvar1406[(1'h0):(1'h0)] : forvar1424) ?
                              $unsigned($signed(reg1590)) : (reg1488[(1'h1):(1'h1)] ?
                                  (forvar1383 ?
                                      reg1451 : reg1446) : {reg1502}))};
                      reg1600 <= (($signed($signed((8'ha6))) ?
                              $signed({reg1519}) : ((reg1526 ?
                                  reg1547 : reg1477) ^~ reg1418[(2'h3):(2'h2)])) ?
                          (-(reg1543[(3'h5):(2'h2)] ^~ forvar1515[(3'h7):(2'h3)])) : ($signed(forvar1385) ?
                              $unsigned($unsigned(reg1530)) : {reg1496}));
                    end
                  for (forvar1601 = (1'h0); (forvar1601 < (1'h1)); forvar1601 = (forvar1601 + (1'h1)))
                    begin
                      reg1602 <= (~|reg1496[(2'h2):(1'h0)]);
                      reg1603 <= $signed($signed($unsigned((forvar1571 * forvar1484))));
                    end
                end
              else
                begin
                  reg1596 <= forvar1535[(4'hc):(2'h2)];
                  for (forvar1597 = (1'h0); (forvar1597 < (1'h0)); forvar1597 = (forvar1597 + (1'h1)))
                    begin
                      reg1598 <= forvar1564;
                      reg1599 <= wire1171;
                      reg1600 <= ((-reg1530) ?
                          ((^~reg1553) | {$unsigned(reg1501)}) : (((reg1400 ?
                                      wire1377 : (8'hab)) ?
                                  (reg1578 ^ reg1439) : (&(8'h9f))) ?
                              reg1459 : $signed((reg1400 > reg1548))));
                    end
                  if (forvar1597)
                    begin
                      reg1601 <= (8'ha6);
                    end
                  else
                    begin
                      reg1601 <= (+$signed((8'h9d)));
                      reg1602 <= ((|$unsigned((8'h9f))) ?
                          {($unsigned(forvar1485) | {reg1578})} : {{((8'hb1) > reg1460)}});
                      reg1603 <= $unsigned($signed((reg1600[(4'hc):(1'h0)] - reg1429[(1'h0):(1'h0)])));
                    end
                end
              if ($signed($signed($signed($signed(forvar1514)))))
                begin
                  if (($signed($unsigned(reg1568[(3'h7):(3'h7)])) ?
                      (!(^~(reg1558 <<< reg1580))) : (((reg1506 ?
                              (8'h9e) : reg1490) | reg1598) ?
                          (8'hac) : (reg1447 > reg1594))))
                    begin
                      reg1604 <= $unsigned($signed($unsigned($signed((8'hac)))));
                      reg1605 <= reg1550;
                      reg1606 <= reg1549[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1604 <= ($signed(($signed(reg1443) != reg1456)) <= forvar1597);
                      reg1605 <= $signed((8'hb3));
                      reg1606 <= forvar1396[(1'h0):(1'h0)];
                      reg1607 <= (($unsigned(reg1432) || $unsigned($unsigned((8'ha2)))) != reg1392);
                    end
                  for (forvar1608 = (1'h0); (forvar1608 < (1'h0)); forvar1608 = (forvar1608 + (1'h1)))
                    begin
                      reg1609 <= {({reg1444[(3'h7):(3'h4)]} ?
                              (!(forvar1406 ?
                                  (8'ha3) : reg1439)) : (^~reg1528[(3'h7):(3'h5)]))};
                      reg1610 <= reg1412;
                      reg1611 <= ($signed((^$unsigned(reg1466))) + forvar1425[(3'h4):(2'h2)]);
                      reg1612 <= reg1594;
                    end
                  for (forvar1613 = (1'h0); (forvar1613 < (1'h0)); forvar1613 = (forvar1613 + (1'h1)))
                    begin
                      reg1614 <= (8'ha5);
                      reg1615 <= reg1570;
                      reg1616 <= ((-$signed((8'hb1))) ?
                          {((^~reg1504) && $unsigned(wire1172))} : forvar1531);
                    end
                end
              else
                begin
                  for (forvar1604 = (1'h0); (forvar1604 < (1'h1)); forvar1604 = (forvar1604 + (1'h1)))
                    begin
                      reg1605 <= {reg1600};
                      reg1606 <= {(forvar1597 >> ((8'hb2) ?
                              reg1445[(3'h6):(3'h6)] : ((8'h9f) != forvar1461)))};
                      reg1607 <= $unsigned((&((!forvar1395) ?
                          reg1380[(3'h7):(1'h0)] : {reg1491})));
                      reg1608 <= ((+(forvar1588[(4'hb):(4'hb)] ?
                              (reg1548 >= reg1440) : reg1451[(2'h2):(2'h2)])) ?
                          {$unsigned((reg1497 >>> (8'hb5)))} : (8'hb1));
                    end
                  for (forvar1609 = (1'h0); (forvar1609 < (1'h0)); forvar1609 = (forvar1609 + (1'h1)))
                    begin
                      reg1610 <= $unsigned({reg1593});
                      reg1611 <= forvar1601[(2'h3):(2'h2)];
                      reg1612 <= $unsigned((forvar1390[(2'h2):(1'h1)] | (!(~&forvar1562))));
                    end
                  if (reg1614[(2'h2):(1'h1)])
                    begin
                      reg1613 <= forvar1407[(4'hd):(3'h7)];
                    end
                  else
                    begin
                      reg1613 <= reg1458;
                      reg1614 <= (-reg1394);
                    end
                  reg1615 <= reg1584;
                end
              for (forvar1617 = (1'h0); (forvar1617 < (2'h2)); forvar1617 = (forvar1617 + (1'h1)))
                begin
                  reg1618 <= (($signed((reg1474 <= reg1499)) ?
                      $signed(((8'ha8) ?
                          reg1593 : reg1429)) : {{reg1386}}) == ({(reg1410 ?
                          reg1576 : (8'hba))} < reg1586[(3'h4):(2'h2)]));
                  if (reg1567[(2'h3):(2'h2)])
                    begin
                      reg1619 <= reg1612[(2'h2):(1'h1)];
                      reg1620 <= reg1512;
                    end
                  else
                    begin
                      reg1619 <= ({reg1558} + {$unsigned((-(8'h9d)))});
                      reg1620 <= $unsigned(($unsigned($unsigned(reg1380)) ?
                          ((reg1506 ?
                              (8'hb3) : reg1418) <<< $signed((8'h9c))) : reg1410[(3'h5):(3'h4)]));
                      reg1621 <= (reg1527[(3'h6):(1'h1)] || $unsigned(((!reg1567) ?
                          (^~reg1580) : $unsigned(forvar1567))));
                    end
                end
            end
          else
            begin
              reg1596 <= (^(~&$unsigned($signed(reg1420))));
              for (forvar1597 = (1'h0); (forvar1597 < (2'h2)); forvar1597 = (forvar1597 + (1'h1)))
                begin
                  for (forvar1598 = (1'h0); (forvar1598 < (1'h0)); forvar1598 = (forvar1598 + (1'h1)))
                    begin
                      reg1599 <= ((~&($signed((8'h9d)) ?
                          forvar1437 : ((8'h9e) ?
                              (8'ha2) : reg1455))) * (((8'hae) ?
                          (forvar1423 ?
                              reg1587 : forvar1608) : $signed(reg1458)) ~^ ($signed(forvar1479) ?
                          reg1443 : $unsigned(reg1577))));
                      reg1600 <= $signed($signed($signed(((8'ha5) ?
                          forvar1576 : reg1422))));
                    end
                  for (forvar1601 = (1'h0); (forvar1601 < (2'h2)); forvar1601 = (forvar1601 + (1'h1)))
                    begin
                      reg1602 <= reg1565[(2'h3):(1'h0)];
                    end
                  reg1603 <= reg1493;
                end
              if ($signed((reg1445[(4'hb):(4'hb)] >> forvar1591[(1'h0):(1'h0)])))
                begin
                  for (forvar1604 = (1'h0); (forvar1604 < (1'h1)); forvar1604 = (forvar1604 + (1'h1)))
                    begin
                      reg1605 <= reg1452;
                      reg1606 <= {$unsigned((wire1170[(1'h1):(1'h0)] ?
                              $unsigned(reg1552) : {forvar1538}))};
                    end
                  for (forvar1607 = (1'h0); (forvar1607 < (2'h2)); forvar1607 = (forvar1607 + (1'h1)))
                    begin
                      reg1608 <= reg1391;
                      reg1609 <= $signed($signed(($unsigned(reg1429) ?
                          $signed((8'hb3)) : (!wire1170))));
                      reg1610 <= $signed({reg1589[(3'h6):(3'h6)]});
                    end
                end
              else
                begin
                  reg1604 <= reg1454;
                  for (forvar1605 = (1'h0); (forvar1605 < (1'h0)); forvar1605 = (forvar1605 + (1'h1)))
                    begin
                      reg1606 <= $unsigned($signed($unsigned((-(8'haa)))));
                      reg1607 <= ($signed(forvar1576[(4'h9):(3'h7)]) * (~&(~^reg1405)));
                    end
                  for (forvar1608 = (1'h0); (forvar1608 < (1'h1)); forvar1608 = (forvar1608 + (1'h1)))
                    begin
                      reg1609 <= {reg1614};
                      reg1610 <= forvar1549[(4'h8):(2'h3)];
                      reg1611 <= $unsigned(forvar1515);
                      reg1612 <= $signed($unsigned(((wire1171 & wire1377) && reg1557[(4'hd):(4'hb)])));
                    end
                  for (forvar1613 = (1'h0); (forvar1613 < (1'h0)); forvar1613 = (forvar1613 + (1'h1)))
                    begin
                      reg1614 <= reg1610[(3'h7):(1'h0)];
                      reg1615 <= $unsigned($signed((reg1524[(1'h0):(1'h0)] >>> {reg1599})));
                    end
                end
            end
        end
    end
  assign wire1622 = (-forvar1438[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      if ({{reg1616}})
        begin
          for (forvar1623 = (1'h0); (forvar1623 < (1'h1)); forvar1623 = (forvar1623 + (1'h1)))
            begin
              if ($signed(reg1428[(3'h6):(2'h3)]))
                begin
                  reg1624 <= {$signed(reg1461)};
                  if (reg1486)
                    begin
                      reg1625 <= (&((reg1586[(1'h1):(1'h0)] + (reg1610 | (8'hb3))) ?
                          (^reg1456) : reg1476[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg1625 <= (reg1447 || $unsigned((^~(+reg1395))));
                      reg1626 <= $unsigned(($signed(forvar1576) ^ $signed({reg1578})));
                    end
                  reg1627 <= (~^((8'ha9) << (|(8'hb8))));
                end
              else
                begin
                  for (forvar1624 = (1'h0); (forvar1624 < (2'h3)); forvar1624 = (forvar1624 + (1'h1)))
                    begin
                      reg1625 <= (^~reg1558);
                      reg1626 <= (({reg1381} ?
                              $unsigned(reg1626[(4'hb):(3'h7)]) : reg1566[(3'h7):(2'h3)]) ?
                          (($unsigned(reg1427) ? {reg1390} : {forvar1457}) ?
                              ((reg1476 ?
                                  reg1532 : forvar1514) < {(8'ha7)}) : ($signed(reg1400) ?
                                  reg1438 : (-(8'ha8)))) : $signed((~forvar1433)));
                      reg1627 <= reg1402[(4'he):(3'h5)];
                    end
                end
              reg1628 <= forvar1604;
            end
          for (forvar1629 = (1'h0); (forvar1629 < (1'h1)); forvar1629 = (forvar1629 + (1'h1)))
            begin
              if (((-$signed({reg1396})) ? reg1530[(4'h8):(3'h4)] : forvar1549))
                begin
                  if (reg1402)
                    begin
                      reg1630 <= reg1418[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg1630 <= $signed((reg1569 ?
                          ({reg1520} && reg1422[(3'h6):(3'h6)]) : $signed($signed(forvar1617))));
                      reg1631 <= reg1384[(3'h4):(3'h4)];
                      reg1632 <= forvar1406;
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h2)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= reg1616[(1'h1):(1'h0)];
                      reg1635 <= ((&(forvar1417 ^~ $signed((8'hb9)))) ~^ reg1440);
                    end
                  for (forvar1636 = (1'h0); (forvar1636 < (1'h1)); forvar1636 = (forvar1636 + (1'h1)))
                    begin
                      reg1637 <= $signed($signed($signed(reg1539[(3'h4):(1'h0)])));
                      reg1638 <= reg1445;
                    end
                  for (forvar1639 = (1'h0); (forvar1639 < (2'h3)); forvar1639 = (forvar1639 + (1'h1)))
                    begin
                      reg1640 <= ($unsigned((~|(reg1497 ? (8'hb4) : reg1616))) ?
                          (reg1530[(4'ha):(3'h6)] ?
                              reg1488[(3'h4):(1'h0)] : $signed($signed((8'h9d)))) : ($unsigned((~|forvar1379)) && ($signed((8'hae)) ?
                              reg1611 : $signed(reg1520))));
                    end
                end
              else
                begin
                  if ({$unsigned(reg1499)})
                    begin
                      reg1630 <= (((~$unsigned(reg1580)) ?
                          $unsigned($signed(reg1564)) : (|{(8'hba)})) ^~ $unsigned((!(forvar1502 == reg1548))));
                      reg1631 <= ($unsigned((!(reg1638 ? reg1567 : reg1640))) ?
                          ((-forvar1639) || ((|forvar1502) ?
                              ((8'ha6) ^~ forvar1438) : forvar1629[(3'h5):(3'h5)])) : $unsigned(reg1634));
                      reg1632 <= ($unsigned((8'hba)) ?
                          ($unsigned({reg1427}) | reg1482) : ((((8'h9e) ?
                              (8'ha7) : reg1484) >>> reg1429) > wire1622));
                    end
                  else
                    begin
                      reg1630 <= $unsigned(reg1391);
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (1'h1)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= {{(~^{reg1457})}};
                    end
                end
              for (forvar1641 = (1'h0); (forvar1641 < (2'h3)); forvar1641 = (forvar1641 + (1'h1)))
                begin
                  for (forvar1642 = (1'h0); (forvar1642 < (2'h3)); forvar1642 = (forvar1642 + (1'h1)))
                    begin
                      reg1643 <= $signed((reg1561[(3'h4):(1'h1)] ?
                          (^$unsigned(forvar1623)) : forvar1562));
                      reg1644 <= $unsigned(reg1415[(1'h0):(1'h0)]);
                      reg1645 <= (~&$unsigned({(|(8'hab))}));
                      reg1646 <= $signed($signed(reg1602[(1'h0):(1'h0)]));
                    end
                  if (reg1615[(3'h4):(3'h4)])
                    begin
                      reg1647 <= $unsigned($signed(reg1539[(4'h9):(4'h9)]));
                      reg1648 <= (forvar1581[(1'h0):(1'h0)] ?
                          $unsigned({(^~reg1467)}) : (^{$unsigned((8'ha4))}));
                    end
                  else
                    begin
                      reg1647 <= reg1428;
                      reg1648 <= $signed($unsigned({$unsigned((8'ha3))}));
                    end
                  if ($signed($unsigned($unsigned((forvar1534 ?
                      reg1448 : reg1475)))))
                    begin
                      reg1649 <= $signed((forvar1552 ?
                          {(~^forvar1414)} : reg1565));
                      reg1650 <= $unsigned($signed(forvar1639[(1'h0):(1'h0)]));
                      reg1651 <= $signed((($signed(reg1640) >= (forvar1437 ?
                          forvar1383 : reg1396)) & $unsigned($signed(reg1422))));
                    end
                  else
                    begin
                      reg1649 <= reg1574[(2'h2):(2'h2)];
                      reg1650 <= ($signed($signed((reg1495 ?
                          reg1554 : reg1634))) - $signed(reg1577));
                      reg1651 <= {(wire1622[(1'h1):(1'h1)] | forvar1571[(4'h8):(2'h2)])};
                      reg1652 <= $unsigned((|(-((8'hba) ? reg1458 : reg1401))));
                    end
                  for (forvar1653 = (1'h0); (forvar1653 < (1'h1)); forvar1653 = (forvar1653 + (1'h1)))
                    begin
                      reg1654 <= ($signed(((reg1551 >= (8'h9d)) ^ $unsigned(reg1557))) <<< (8'ha0));
                    end
                end
              for (forvar1655 = (1'h0); (forvar1655 < (2'h3)); forvar1655 = (forvar1655 + (1'h1)))
                begin
                  if ($signed($unsigned(forvar1562)))
                    begin
                      reg1656 <= {(~|$unsigned((reg1630 * reg1491)))};
                      reg1657 <= (~&$unsigned(reg1397[(4'h8):(4'h8)]));
                      reg1658 <= reg1596;
                      reg1659 <= reg1520;
                    end
                  else
                    begin
                      reg1656 <= (~&(^~(-reg1387[(3'h6):(2'h2)])));
                      reg1657 <= reg1380;
                    end
                  if (($unsigned(reg1441) * (8'h9c)))
                    begin
                      reg1660 <= ($unsigned($unsigned({reg1640})) ?
                          ($unsigned((+reg1557)) ?
                              ($signed((8'ha2)) ?
                                  wire1171 : (-forvar1442)) : $signed($signed(reg1568))) : (~&forvar1485[(3'h6):(1'h1)]));
                    end
                  else
                    begin
                      reg1660 <= {({(forvar1502 ? reg1560 : (8'ha1))} ?
                              reg1620[(4'h8):(3'h5)] : $unsigned((reg1660 | reg1466)))};
                      reg1661 <= (^~$unsigned(reg1506[(4'h9):(3'h7)]));
                      reg1662 <= reg1431[(1'h0):(1'h0)];
                      reg1663 <= (($signed(reg1521) - $signed($unsigned(reg1605))) ?
                          $signed($signed((forvar1572 ?
                              forvar1608 : forvar1549))) : (reg1390[(3'h6):(3'h5)] ?
                              reg1611[(2'h3):(2'h2)] : $signed(reg1557)));
                    end
                  if ((forvar1591 ?
                      ((-forvar1461) << (^~forvar1624)) : reg1528))
                    begin
                      reg1664 <= reg1532;
                      reg1665 <= ($unsigned($unsigned(reg1506[(4'hf):(4'ha)])) ?
                          $unsigned($unsigned(reg1516[(2'h2):(1'h0)])) : (($signed(forvar1568) ?
                                  (reg1548 >= forvar1502) : $signed(forvar1556)) ?
                              ((forvar1379 ?
                                  reg1554 : forvar1417) != reg1402) : reg1603[(4'h9):(2'h2)]));
                    end
                  else
                    begin
                      reg1664 <= reg1643[(3'h7):(1'h1)];
                      reg1665 <= (~{($signed(reg1646) + reg1416[(4'h9):(3'h6)])});
                      reg1666 <= (-($unsigned(forvar1490) | $unsigned((reg1502 ?
                          reg1471 : forvar1567))));
                      reg1667 <= reg1421;
                    end
                end
            end
          for (forvar1668 = (1'h0); (forvar1668 < (1'h0)); forvar1668 = (forvar1668 + (1'h1)))
            begin
              reg1669 <= $signed(reg1470[(3'h5):(3'h5)]);
              if ((~^(^($unsigned(reg1412) ?
                  reg1457[(3'h4):(1'h0)] : reg1397))))
                begin
                  for (forvar1670 = (1'h0); (forvar1670 < (1'h1)); forvar1670 = (forvar1670 + (1'h1)))
                    begin
                      reg1671 <= (~{reg1552});
                      reg1672 <= (forvar1655[(2'h2):(1'h0)] + reg1627[(3'h7):(3'h5)]);
                      reg1673 <= reg1511[(3'h7):(3'h7)];
                    end
                end
              else
                begin
                  reg1670 <= (^reg1428);
                  for (forvar1671 = (1'h0); (forvar1671 < (1'h1)); forvar1671 = (forvar1671 + (1'h1)))
                    begin
                      reg1672 <= $signed((8'h9c));
                      reg1673 <= ($signed(((~|reg1440) >> (~&reg1478))) ~^ (forvar1379 ?
                          reg1561 : $signed(reg1463[(1'h0):(1'h0)])));
                    end
                  if ($signed({$unsigned({reg1552})}))
                    begin
                      reg1674 <= $unsigned(({$unsigned(reg1661)} <<< $signed(forvar1538[(3'h4):(1'h1)])));
                      reg1675 <= forvar1601;
                    end
                  else
                    begin
                      reg1674 <= ((reg1403 * (|(&reg1644))) >= (forvar1564[(4'h8):(3'h6)] & (^reg1428)));
                      reg1675 <= reg1532;
                      reg1676 <= forvar1449;
                    end
                  reg1677 <= ($signed($unsigned((reg1599 ?
                      forvar1636 : reg1573))) && reg1620[(3'h4):(1'h0)]);
                end
              if (reg1555)
                begin
                  reg1678 <= (reg1662[(3'h4):(2'h2)] ^~ reg1479[(3'h7):(2'h3)]);
                  if ({$signed({(~&forvar1485)})})
                    begin
                      reg1679 <= $unsigned(reg1626);
                    end
                  else
                    begin
                      reg1679 <= (+{$signed($signed((8'haa)))});
                      reg1680 <= (-forvar1552);
                      reg1681 <= reg1507;
                      reg1682 <= $unsigned((|reg1527[(3'h6):(3'h5)]));
                    end
                end
              else
                begin
                  for (forvar1678 = (1'h0); (forvar1678 < (2'h2)); forvar1678 = (forvar1678 + (1'h1)))
                    begin
                      reg1679 <= reg1537[(2'h3):(1'h1)];
                      reg1680 <= reg1451;
                      reg1681 <= ((&$signed($signed(reg1434))) - forvar1514[(3'h6):(3'h5)]);
                    end
                  for (forvar1682 = (1'h0); (forvar1682 < (2'h3)); forvar1682 = (forvar1682 + (1'h1)))
                    begin
                      reg1683 <= $unsigned(reg1567);
                      reg1684 <= (8'ha5);
                      reg1685 <= ($signed(reg1440[(2'h3):(2'h2)]) ?
                          reg1521 : $unsigned($unsigned({(8'h9e)})));
                      reg1686 <= {(((~reg1463) ?
                                  (forvar1548 ^ reg1674) : (^~reg1493)) ?
                              $unsigned({reg1576}) : wire1377)};
                    end
                end
              if ($unsigned({$signed($unsigned(reg1540))}))
                begin
                  reg1687 <= (^~(^$unsigned((reg1678 || forvar1514))));
                end
              else
                begin
                  for (forvar1687 = (1'h0); (forvar1687 < (2'h2)); forvar1687 = (forvar1687 + (1'h1)))
                    begin
                      reg1688 <= ((&forvar1687[(2'h2):(2'h2)]) ?
                          $unsigned($unsigned((8'hb3))) : {{$unsigned(forvar1479)}});
                    end
                  for (forvar1689 = (1'h0); (forvar1689 < (1'h0)); forvar1689 = (forvar1689 + (1'h1)))
                    begin
                      reg1690 <= reg1510;
                      reg1691 <= $signed((forvar1613 ^ $unsigned($signed(reg1647))));
                      reg1692 <= forvar1534[(3'h4):(1'h1)];
                      reg1693 <= ((8'hb9) & (($signed(reg1614) ?
                          (forvar1438 ?
                              reg1637 : reg1688) : $unsigned(reg1676)) <= $signed($unsigned(reg1487))));
                    end
                end
            end
        end
      else
        begin
          if ($unsigned(reg1654))
            begin
              if ({({(forvar1668 <= reg1537)} && (+(reg1469 ?
                      reg1603 : (8'ha1))))})
                begin
                  for (forvar1623 = (1'h0); (forvar1623 < (1'h0)); forvar1623 = (forvar1623 + (1'h1)))
                    begin
                      reg1624 <= reg1519;
                      reg1625 <= $unsigned(reg1532);
                      reg1626 <= (((reg1654[(1'h1):(1'h1)] ?
                              reg1646[(1'h0):(1'h0)] : reg1672[(1'h1):(1'h1)]) < $signed({reg1679})) ?
                          (reg1555 ?
                              $unsigned({reg1580}) : (~&reg1498)) : (+forvar1472));
                    end
                end
              else
                begin
                  for (forvar1623 = (1'h0); (forvar1623 < (2'h3)); forvar1623 = (forvar1623 + (1'h1)))
                    begin
                      reg1624 <= $unsigned($signed($unsigned((reg1602 ?
                          reg1584 : reg1518))));
                      reg1625 <= (reg1416 ?
                          ($signed($unsigned(reg1645)) & (8'ha3)) : reg1384[(3'h6):(3'h6)]);
                      reg1626 <= $signed($signed((~|{forvar1379})));
                    end
                  for (forvar1627 = (1'h0); (forvar1627 < (1'h0)); forvar1627 = (forvar1627 + (1'h1)))
                    begin
                      reg1628 <= reg1441[(3'h4):(1'h0)];
                      reg1629 <= ((($signed(reg1630) && (reg1410 ?
                              reg1441 : reg1502)) ?
                          $unsigned($signed(forvar1605)) : forvar1671[(1'h0):(1'h0)]) >>> (($unsigned(reg1489) - (reg1539 ?
                          wire1172 : reg1690)) >= $unsigned((reg1630 * forvar1442))));
                    end
                end
              for (forvar1630 = (1'h0); (forvar1630 < (1'h1)); forvar1630 = (forvar1630 + (1'h1)))
                begin
                  for (forvar1631 = (1'h0); (forvar1631 < (1'h0)); forvar1631 = (forvar1631 + (1'h1)))
                    begin
                      reg1632 <= reg1648[(3'h4):(1'h0)];
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (1'h1)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= ($signed(reg1582[(1'h1):(1'h1)]) <<< $signed(forvar1425));
                      reg1635 <= (~$signed((~&(forvar1424 ?
                          reg1465 : forvar1572))));
                    end
                end
              for (forvar1636 = (1'h0); (forvar1636 < (1'h1)); forvar1636 = (forvar1636 + (1'h1)))
                begin
                  if ((reg1397[(4'hc):(3'h6)] ?
                      {reg1392} : (($unsigned((8'ha0)) ?
                          reg1474[(4'ha):(4'h9)] : $unsigned(forvar1531)) << reg1574)))
                    begin
                      reg1637 <= reg1690;
                    end
                  else
                    begin
                      reg1637 <= reg1578[(4'h8):(3'h6)];
                      reg1638 <= forvar1571;
                      reg1639 <= (!reg1600[(4'h9):(2'h3)]);
                      reg1640 <= $unsigned((-$signed(reg1418[(2'h3):(1'h0)])));
                    end
                end
              for (forvar1641 = (1'h0); (forvar1641 < (2'h2)); forvar1641 = (forvar1641 + (1'h1)))
                begin
                  reg1642 <= {reg1444[(3'h7):(1'h1)]};
                  for (forvar1643 = (1'h0); (forvar1643 < (2'h3)); forvar1643 = (forvar1643 + (1'h1)))
                    begin
                      reg1644 <= reg1510[(3'h7):(1'h1)];
                      reg1645 <= reg1479[(4'ha):(3'h7)];
                      reg1646 <= {(forvar1556[(2'h2):(1'h1)] ?
                              {(reg1473 ? reg1549 : (8'hb3))} : reg1497)};
                    end
                end
            end
          else
            begin
              if ((^reg1530))
                begin
                  if (reg1395[(1'h0):(1'h0)])
                    begin
                      reg1623 <= reg1438[(4'h8):(3'h7)];
                      reg1624 <= {{(~|reg1426)}};
                      reg1625 <= forvar1381;
                      reg1626 <= reg1601[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1623 <= (&$signed(($signed(reg1570) ?
                          ((8'ha4) * reg1496) : ((8'hae) ?
                              forvar1552 : reg1640))));
                      reg1624 <= (reg1384[(4'hd):(2'h3)] - reg1587[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar1623 = (1'h0); (forvar1623 < (2'h2)); forvar1623 = (forvar1623 + (1'h1)))
                    begin
                      reg1624 <= (~reg1666[(2'h3):(1'h0)]);
                    end
                  for (forvar1625 = (1'h0); (forvar1625 < (2'h2)); forvar1625 = (forvar1625 + (1'h1)))
                    begin
                      reg1626 <= (|(&reg1589));
                      reg1627 <= $unsigned({(~(reg1594 ?
                              forvar1387 : reg1542))});
                      reg1628 <= {((reg1410[(3'h7):(1'h1)] ?
                                  (reg1667 && reg1688) : (-(8'ha7))) ?
                              reg1409[(1'h0):(1'h0)] : $unsigned(forvar1609))};
                    end
                  if ($unsigned({($unsigned(forvar1576) ?
                          $unsigned(forvar1437) : (8'hb1))}))
                    begin
                      reg1629 <= (~|reg1478[(4'h8):(3'h6)]);
                      reg1630 <= (-(reg1613 ?
                          $signed(forvar1456) : (reg1619 ^~ (reg1601 >>> reg1452))));
                      reg1631 <= reg1502;
                      reg1632 <= reg1595[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg1629 <= reg1618[(2'h2):(1'h0)];
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h2)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= (!(8'ha0));
                      reg1635 <= (reg1488[(2'h3):(2'h2)] ~^ (~^reg1393[(4'h8):(3'h7)]));
                    end
                end
              reg1636 <= $unsigned($unsigned((reg1590[(3'h4):(1'h1)] * $unsigned(reg1589))));
            end
          for (forvar1647 = (1'h0); (forvar1647 < (2'h3)); forvar1647 = (forvar1647 + (1'h1)))
            begin
              if (((reg1508 ?
                  reg1469[(3'h4):(1'h0)] : $unsigned((&(8'ha2)))) <= (~|($signed(reg1421) ?
                  (wire1622 ? forvar1438 : (8'hb5)) : (~|forvar1531)))))
                begin
                  reg1648 <= $unsigned((8'hac));
                end
              else
                begin
                  for (forvar1648 = (1'h0); (forvar1648 < (2'h3)); forvar1648 = (forvar1648 + (1'h1)))
                    begin
                      reg1649 <= forvar1461[(2'h3):(1'h1)];
                      reg1650 <= (-(^(|(reg1564 ? forvar1629 : forvar1383))));
                      reg1651 <= $signed({(!forvar1564[(1'h1):(1'h1)])});
                      reg1652 <= $unsigned(forvar1642);
                    end
                end
              for (forvar1653 = (1'h0); (forvar1653 < (1'h0)); forvar1653 = (forvar1653 + (1'h1)))
                begin
                  if (forvar1556)
                    begin
                      reg1654 <= $unsigned($signed($signed((8'had))));
                    end
                  else
                    begin
                      reg1654 <= reg1431;
                    end
                  for (forvar1655 = (1'h0); (forvar1655 < (1'h0)); forvar1655 = (forvar1655 + (1'h1)))
                    begin
                      reg1656 <= {{(~^(forvar1601 ? wire1171 : reg1453))}};
                      reg1657 <= $signed(reg1640);
                      reg1658 <= ({forvar1442} || $unsigned((8'ha4)));
                    end
                  for (forvar1659 = (1'h0); (forvar1659 < (2'h3)); forvar1659 = (forvar1659 + (1'h1)))
                    begin
                      reg1660 <= ($signed((reg1670 * forvar1601)) ?
                          $signed(reg1686[(3'h5):(2'h2)]) : $signed(((~reg1544) ?
                              {reg1454} : reg1678)));
                      reg1661 <= $signed($signed(reg1390[(3'h4):(2'h2)]));
                      reg1662 <= {($signed({forvar1496}) ?
                              reg1643[(3'h6):(2'h2)] : (reg1488 || $signed(reg1593)))};
                    end
                end
              if (((reg1627[(2'h3):(2'h3)] ?
                      (~&(8'hb0)) : ($unsigned(reg1393) ?
                          ((8'hae) ?
                              forvar1624 : reg1567) : reg1382[(2'h2):(1'h0)])) ?
                  {{(reg1435 >= reg1566)}} : reg1654))
                begin
                  if (($unsigned({{wire1377}}) <<< ((reg1524 ?
                          forvar1523[(2'h3):(1'h1)] : reg1686) ?
                      (8'hb5) : $unsigned((reg1573 != forvar1538)))))
                    begin
                      reg1663 <= forvar1588[(4'h8):(1'h0)];
                      reg1664 <= $signed((+reg1483));
                      reg1665 <= (-$unsigned({reg1493}));
                    end
                  else
                    begin
                      reg1663 <= $signed((+$signed(reg1661)));
                      reg1664 <= reg1392;
                    end
                end
              else
                begin
                  for (forvar1663 = (1'h0); (forvar1663 < (1'h0)); forvar1663 = (forvar1663 + (1'h1)))
                    begin
                      reg1664 <= ({{reg1453[(1'h0):(1'h0)]}} + (((reg1579 ?
                                  reg1386 : (8'ha9)) ?
                              $unsigned(reg1462) : ((8'hb4) ?
                                  reg1557 : forvar1547)) ?
                          {(reg1529 ?
                                  forvar1572 : reg1541)} : (~|$signed((8'hb6)))));
                      reg1665 <= (+(^($signed((8'ha8)) ?
                          $unsigned(forvar1576) : (reg1608 ?
                              forvar1489 : reg1421))));
                    end
                  if ((((&$unsigned(reg1626)) ?
                      $unsigned((-forvar1379)) : reg1459) != ({forvar1423} >>> (forvar1531 ?
                      (~^reg1592) : reg1550[(3'h4):(1'h1)]))))
                    begin
                      reg1666 <= $signed({$unsigned(forvar1468)});
                      reg1667 <= (((reg1527 - (&reg1530)) ?
                              (forvar1509 ?
                                  (reg1623 ?
                                      (8'ha4) : (8'ha5)) : $unsigned(reg1498)) : (~|{(8'ha7)})) ?
                          $unsigned((8'ha3)) : ($unsigned($unsigned(reg1543)) & (-(reg1460 ?
                              forvar1485 : reg1500))));
                    end
                  else
                    begin
                      reg1666 <= $signed(reg1665[(3'h6):(2'h2)]);
                      reg1667 <= (~^{reg1408[(1'h1):(1'h1)]});
                      reg1668 <= (~^$unsigned(reg1601[(1'h1):(1'h1)]));
                    end
                end
              if ((($unsigned((reg1624 > forvar1624)) << (&(reg1593 ?
                      reg1474 : forvar1605))) ?
                  reg1400[(2'h3):(1'h0)] : (&{$unsigned((8'ha9))})))
                begin
                  for (forvar1669 = (1'h0); (forvar1669 < (2'h3)); forvar1669 = (forvar1669 + (1'h1)))
                    begin
                      reg1670 <= (((-forvar1414) & $signed($signed(forvar1473))) ?
                          $signed($unsigned({reg1657})) : (-forvar1655));
                      reg1671 <= $signed({{reg1512}});
                      reg1672 <= (((^~$unsigned(forvar1572)) ?
                              reg1583 : (~{forvar1682})) ?
                          (^~{(forvar1395 ?
                                  reg1447 : reg1662)}) : $signed(({reg1642} ~^ $signed((8'hb9)))));
                    end
                end
              else
                begin
                  reg1669 <= (($unsigned((~^reg1458)) <<< $unsigned(forvar1682[(1'h0):(1'h0)])) ?
                      ((8'had) ?
                          ((|reg1502) <<< forvar1585) : $signed(reg1678)) : forvar1642);
                end
            end
          for (forvar1673 = (1'h0); (forvar1673 < (1'h0)); forvar1673 = (forvar1673 + (1'h1)))
            begin
              if (reg1520[(4'ha):(3'h7)])
                begin
                  reg1674 <= reg1494[(1'h1):(1'h0)];
                end
              else
                begin
                  reg1674 <= ((8'hb3) & ((~|reg1528) ^~ $signed(reg1444[(1'h0):(1'h0)])));
                  for (forvar1675 = (1'h0); (forvar1675 < (2'h2)); forvar1675 = (forvar1675 + (1'h1)))
                    begin
                      reg1676 <= $signed((~&((8'had) ?
                          $signed(forvar1380) : $unsigned((8'ha2)))));
                    end
                end
              reg1677 <= $signed($unsigned({$unsigned(reg1680)}));
              for (forvar1678 = (1'h0); (forvar1678 < (2'h2)); forvar1678 = (forvar1678 + (1'h1)))
                begin
                  if ((|forvar1617[(1'h1):(1'h0)]))
                    begin
                      reg1679 <= (({$unsigned(forvar1564)} ?
                              $signed(((8'hb7) ~^ (8'ha4))) : (|$signed(forvar1639))) ?
                          forvar1497 : {(forvar1468 >= forvar1552[(3'h4):(3'h4)])});
                    end
                  else
                    begin
                      reg1679 <= {(|({reg1551} <= $signed(reg1379)))};
                      reg1680 <= $signed(forvar1490[(1'h0):(1'h0)]);
                      reg1681 <= reg1495[(3'h5):(3'h4)];
                    end
                  reg1682 <= ($signed($unsigned($signed(reg1500))) << ((^$unsigned(reg1427)) ?
                      ($signed(forvar1668) ?
                          $unsigned(reg1478) : reg1402[(4'hb):(1'h0)]) : $unsigned((&forvar1468))));
                end
            end
        end
    end
  assign wire1694 = $unsigned(reg1657);
  assign wire1695 = forvar1502;
  assign wire1696 = (^~reg1594);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1173
#( parameter param1376 = (((8'ha8) ? (((8'hb2) ? (8'hb2) : (8'hac)) ? ((8'hac) <= (8'hb5)) : {(8'h9f)}) : ((~(8'had)) ? (^~(8'hb5)) : ((8'ha6) & (8'hb7)))) || {(!(-(8'hb2)))}) )
(y, clk, wire1178, wire1177, wire1176, wire1175, wire1174);
  output wire [(32'h8d5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire1178;
  input wire signed [(4'hb):(1'h0)] wire1177;
  input wire [(3'h4):(1'h0)] wire1176;
  input wire [(4'hb):(1'h0)] wire1175;
  input wire [(3'h5):(1'h0)] wire1174;
  reg signed [(4'he):(1'h0)] reg1375 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1374 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1359 = (1'h0);
  reg [(2'h2):(1'h0)] reg1373 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1372 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1366 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1364 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1371 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1370 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1369 = (1'h0);
  reg [(4'h9):(1'h0)] reg1368 = (1'h0);
  reg [(4'h8):(1'h0)] reg1367 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1366 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1365 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1364 = (1'h0);
  reg [(4'h8):(1'h0)] reg1363 = (1'h0);
  reg [(3'h6):(1'h0)] reg1362 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1361 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1360 = (1'h0);
  reg [(2'h2):(1'h0)] reg1359 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1358 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1356 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1354 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1348 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1338 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1343 = (1'h0);
  reg [(2'h3):(1'h0)] reg1341 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1337 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1320 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1334 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1329 = (1'h0);
  reg [(2'h2):(1'h0)] reg1328 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1326 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1322 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1319 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1345 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1344 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1358 = (1'h0);
  reg [(3'h7):(1'h0)] reg1357 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1356 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1352 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1350 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1347 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1355 = (1'h0);
  reg [(4'hb):(1'h0)] reg1354 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1353 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1352 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1351 = (1'h0);
  reg [(3'h5):(1'h0)] reg1350 = (1'h0);
  reg [(4'h8):(1'h0)] reg1349 = (1'h0);
  reg [(3'h5):(1'h0)] reg1348 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1347 = (1'h0);
  reg [(4'h8):(1'h0)] reg1346 = (1'h0);
  reg [(5'h10):(1'h0)] reg1345 = (1'h0);
  reg [(4'he):(1'h0)] forvar1344 = (1'h0);
  reg [(3'h4):(1'h0)] reg1343 = (1'h0);
  reg [(2'h2):(1'h0)] reg1342 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1341 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1340 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1339 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1338 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1337 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1336 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1335 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1334 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1333 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1332 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1331 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1330 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1329 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1328 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1327 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1326 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1323 = (1'h0);
  reg [(4'hb):(1'h0)] reg1325 = (1'h0);
  reg [(4'h9):(1'h0)] reg1324 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1323 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1322 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1321 = (1'h0);
  reg [(4'ha):(1'h0)] reg1320 = (1'h0);
  reg [(4'he):(1'h0)] forvar1319 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire1318;
  wire [(3'h7):(1'h0)] wire1317;
  wire signed [(4'he):(1'h0)] wire1316;
  reg signed [(3'h6):(1'h0)] reg1315 = (1'h0);
  reg [(4'hd):(1'h0)] reg1314 = (1'h0);
  reg [(4'h9):(1'h0)] reg1313 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1312 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1311 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1310 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1309 = (1'h0);
  reg [(5'h10):(1'h0)] reg1308 = (1'h0);
  reg [(4'h8):(1'h0)] reg1307 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1306 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1305 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1304 = (1'h0);
  reg [(3'h5):(1'h0)] reg1303 = (1'h0);
  reg [(4'h9):(1'h0)] reg1302 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1301 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1300 = (1'h0);
  reg [(3'h6):(1'h0)] reg1299 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1298 = (1'h0);
  reg [(4'he):(1'h0)] reg1297 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1296 = (1'h0);
  reg [(4'hc):(1'h0)] reg1295 = (1'h0);
  reg [(4'h9):(1'h0)] reg1294 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1293 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1292 = (1'h0);
  reg [(4'he):(1'h0)] reg1291 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1290 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1289 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1274 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1273 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1288 = (1'h0);
  reg [(4'h9):(1'h0)] reg1287 = (1'h0);
  reg [(4'h8):(1'h0)] reg1286 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1285 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1284 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1283 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1282 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1281 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1280 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1279 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1278 = (1'h0);
  reg [(4'he):(1'h0)] reg1277 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1276 = (1'h0);
  reg [(4'hb):(1'h0)] reg1275 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1274 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1273 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1272 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1269 = (1'h0);
  reg [(4'hd):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1266 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1265 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1255 = (1'h0);
  reg [(2'h3):(1'h0)] reg1254 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1271 = (1'h0);
  reg [(5'h10):(1'h0)] reg1270 = (1'h0);
  reg [(3'h7):(1'h0)] reg1269 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1268 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1267 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1266 = (1'h0);
  reg [(4'hd):(1'h0)] reg1265 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1264 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1263 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1262 = (1'h0);
  reg [(4'h9):(1'h0)] reg1261 = (1'h0);
  reg [(4'h8):(1'h0)] reg1260 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1259 = (1'h0);
  reg [(4'hb):(1'h0)] reg1258 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1257 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1256 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1255 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1254 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1253 = (1'h0);
  reg [(4'h9):(1'h0)] reg1252 = (1'h0);
  reg [(4'he):(1'h0)] reg1251 = (1'h0);
  reg [(2'h2):(1'h0)] reg1250 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1249 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1248 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1246 = (1'h0);
  reg [(5'h10):(1'h0)] reg1245 = (1'h0);
  reg [(3'h6):(1'h0)] reg1241 = (1'h0);
  reg [(5'h10):(1'h0)] reg1247 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1246 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1245 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1244 = (1'h0);
  reg [(3'h7):(1'h0)] reg1243 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1242 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1241 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1240 = (1'h0);
  reg [(4'h9):(1'h0)] reg1239 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1238 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1237 = (1'h0);
  reg [(2'h3):(1'h0)] reg1236 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1235 = (1'h0);
  reg [(4'he):(1'h0)] forvar1234 = (1'h0);
  reg [(5'h10):(1'h0)] reg1233 = (1'h0);
  reg [(2'h3):(1'h0)] reg1232 = (1'h0);
  reg [(3'h6):(1'h0)] reg1231 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1230 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1229 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1225 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1220 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1224 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1223 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1215 = (1'h0);
  reg [(4'hc):(1'h0)] reg1214 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1230 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1229 = (1'h0);
  reg [(5'h10):(1'h0)] reg1228 = (1'h0);
  reg [(3'h7):(1'h0)] reg1227 = (1'h0);
  reg [(4'he):(1'h0)] reg1226 = (1'h0);
  reg [(4'hb):(1'h0)] reg1225 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1224 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1223 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1222 = (1'h0);
  reg [(4'hc):(1'h0)] reg1221 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1220 = (1'h0);
  reg [(4'ha):(1'h0)] reg1219 = (1'h0);
  reg [(4'hb):(1'h0)] reg1218 = (1'h0);
  reg [(4'hb):(1'h0)] reg1217 = (1'h0);
  reg [(3'h7):(1'h0)] reg1216 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1215 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1214 = (1'h0);
  reg [(5'h10):(1'h0)] reg1213 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1212 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1211 = (1'h0);
  wire [(4'hc):(1'h0)] wire1210;
  wire signed [(5'h10):(1'h0)] wire1209;
  wire signed [(5'h10):(1'h0)] wire1208;
  wire [(3'h7):(1'h0)] wire1207;
  reg signed [(4'ha):(1'h0)] forvar1203 = (1'h0);
  reg [(4'ha):(1'h0)] reg1202 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1198 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1196 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1183 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1188 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1182 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1206 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1205 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1203 = (1'h0);
  reg [(4'he):(1'h0)] forvar1202 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1201 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1200 = (1'h0);
  reg [(3'h6):(1'h0)] reg1197 = (1'h0);
  reg [(4'hd):(1'h0)] reg1195 = (1'h0);
  reg [(3'h6):(1'h0)] reg1194 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1193 = (1'h0);
  reg [(4'hc):(1'h0)] reg1190 = (1'h0);
  reg [(4'h8):(1'h0)] reg1189 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1200 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1199 = (1'h0);
  reg [(2'h2):(1'h0)] reg1198 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1197 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1196 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1195 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1194 = (1'h0);
  reg [(2'h3):(1'h0)] reg1193 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1192 = (1'h0);
  reg [(3'h6):(1'h0)] reg1191 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1190 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1189 = (1'h0);
  reg [(2'h3):(1'h0)] reg1185 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1181 = (1'h0);
  reg [(3'h4):(1'h0)] reg1188 = (1'h0);
  reg [(3'h6):(1'h0)] reg1187 = (1'h0);
  reg [(4'hf):(1'h0)] reg1186 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1185 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1184 = (1'h0);
  reg [(2'h3):(1'h0)] reg1183 = (1'h0);
  reg [(4'h9):(1'h0)] reg1182 = (1'h0);
  reg [(4'hc):(1'h0)] reg1181 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1180 = (1'h0);
  wire [(4'hc):(1'h0)] wire1179;
  assign y = {reg1375,
                 reg1374,
                 forvar1359,
                 reg1373,
                 forvar1372,
                 forvar1366,
                 reg1364,
                 reg1371,
                 forvar1370,
                 reg1369,
                 reg1368,
                 reg1367,
                 reg1366,
                 reg1365,
                 forvar1364,
                 reg1363,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 forvar1358,
                 reg1356,
                 forvar1354,
                 forvar1348,
                 forvar1338,
                 forvar1343,
                 reg1341,
                 forvar1337,
                 forvar1320,
                 reg1334,
                 forvar1329,
                 reg1328,
                 forvar1326,
                 forvar1322,
                 reg1319,
                 forvar1345,
                 reg1344,
                 reg1358,
                 reg1357,
                 forvar1356,
                 forvar1352,
                 forvar1350,
                 reg1347,
                 reg1355,
                 reg1354,
                 reg1353,
                 reg1352,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 forvar1347,
                 reg1346,
                 reg1345,
                 forvar1344,
                 reg1343,
                 reg1342,
                 forvar1341,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1337,
                 reg1336,
                 reg1335,
                 forvar1334,
                 reg1333,
                 reg1332,
                 reg1331,
                 reg1330,
                 reg1329,
                 forvar1328,
                 reg1327,
                 reg1326,
                 forvar1323,
                 reg1325,
                 reg1324,
                 reg1323,
                 reg1322,
                 reg1321,
                 reg1320,
                 forvar1319,
                 wire1318,
                 wire1317,
                 wire1316,
                 reg1315,
                 reg1314,
                 reg1313,
                 reg1312,
                 reg1311,
                 reg1310,
                 forvar1309,
                 reg1308,
                 reg1307,
                 reg1306,
                 reg1305,
                 forvar1304,
                 reg1303,
                 reg1302,
                 forvar1301,
                 reg1300,
                 reg1299,
                 forvar1298,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 reg1293,
                 reg1292,
                 reg1291,
                 reg1290,
                 forvar1289,
                 forvar1274,
                 reg1273,
                 reg1288,
                 reg1287,
                 reg1286,
                 forvar1285,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1280,
                 reg1279,
                 reg1278,
                 reg1277,
                 forvar1276,
                 reg1275,
                 reg1274,
                 forvar1273,
                 forvar1272,
                 forvar1269,
                 reg1267,
                 reg1266,
                 forvar1265,
                 forvar1255,
                 reg1254,
                 reg1271,
                 reg1270,
                 reg1269,
                 reg1268,
                 forvar1267,
                 forvar1266,
                 reg1265,
                 reg1264,
                 reg1263,
                 forvar1262,
                 reg1261,
                 reg1260,
                 forvar1258,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 reg1255,
                 forvar1254,
                 forvar1253,
                 reg1252,
                 reg1251,
                 reg1250,
                 forvar1249,
                 reg1248,
                 forvar1246,
                 reg1245,
                 reg1241,
                 reg1247,
                 reg1246,
                 forvar1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 forvar1241,
                 forvar1240,
                 reg1239,
                 reg1238,
                 reg1237,
                 reg1236,
                 reg1235,
                 forvar1234,
                 reg1233,
                 reg1232,
                 reg1231,
                 forvar1230,
                 forvar1229,
                 forvar1225,
                 reg1220,
                 reg1224,
                 forvar1223,
                 forvar1215,
                 reg1214,
                 reg1230,
                 reg1229,
                 reg1228,
                 reg1227,
                 reg1226,
                 reg1225,
                 forvar1224,
                 reg1223,
                 reg1222,
                 reg1221,
                 forvar1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1216,
                 reg1215,
                 forvar1214,
                 reg1213,
                 forvar1212,
                 reg1211,
                 wire1210,
                 wire1209,
                 wire1208,
                 wire1207,
                 forvar1203,
                 reg1202,
                 forvar1198,
                 forvar1196,
                 forvar1183,
                 forvar1188,
                 forvar1182,
                 reg1206,
                 reg1205,
                 reg1204,
                 reg1203,
                 forvar1202,
                 reg1201,
                 forvar1200,
                 reg1197,
                 reg1195,
                 reg1194,
                 forvar1193,
                 reg1190,
                 reg1189,
                 reg1200,
                 reg1199,
                 reg1198,
                 forvar1197,
                 reg1196,
                 forvar1195,
                 forvar1194,
                 reg1193,
                 reg1192,
                 reg1191,
                 forvar1190,
                 forvar1189,
                 reg1185,
                 forvar1181,
                 reg1188,
                 reg1187,
                 reg1186,
                 forvar1185,
                 reg1184,
                 reg1183,
                 reg1182,
                 reg1181,
                 forvar1180,
                 wire1179,
                 (1'h0)};
  assign wire1179 = ($unsigned($signed((wire1175 ? wire1177 : wire1176))) ?
                        wire1175 : wire1178);
  always
    @(posedge clk) begin
      if ((wire1175[(2'h3):(1'h1)] == ($signed(wire1177[(1'h1):(1'h0)]) ?
          wire1174[(2'h2):(1'h1)] : (^wire1178))))
        begin
          for (forvar1180 = (1'h0); (forvar1180 < (2'h3)); forvar1180 = (forvar1180 + (1'h1)))
            begin
              if ($unsigned($unsigned(wire1176[(2'h2):(1'h0)])))
                begin
                  if ({$signed(((wire1175 ? (8'ha5) : wire1176) ?
                          $unsigned(wire1175) : ((8'ha2) >>> wire1175)))})
                    begin
                      reg1181 <= wire1177;
                      reg1182 <= (8'haa);
                      reg1183 <= wire1175;
                      reg1184 <= ($signed((~(wire1176 << reg1181))) ?
                          $unsigned(($unsigned(wire1177) ?
                              (forvar1180 << reg1182) : wire1174)) : {wire1174});
                    end
                  else
                    begin
                      reg1181 <= ($signed({wire1176[(2'h3):(1'h1)]}) * (8'hb1));
                    end
                  for (forvar1185 = (1'h0); (forvar1185 < (1'h1)); forvar1185 = (forvar1185 + (1'h1)))
                    begin
                      reg1186 <= wire1176;
                      reg1187 <= $signed(($unsigned({reg1181}) <= $signed($signed(reg1181))));
                      reg1188 <= (~|$unsigned((reg1187[(1'h1):(1'h0)] ?
                          $signed(reg1182) : (wire1179 - reg1184))));
                    end
                end
              else
                begin
                  for (forvar1181 = (1'h0); (forvar1181 < (2'h3)); forvar1181 = (forvar1181 + (1'h1)))
                    begin
                      reg1182 <= (&$unsigned($unsigned(reg1188)));
                      reg1183 <= {reg1182};
                      reg1184 <= reg1186;
                    end
                  if ({((8'ha8) ?
                          (wire1175 ?
                              (reg1188 >= reg1187) : $signed(reg1186)) : $signed((~wire1178)))})
                    begin
                      reg1185 <= forvar1181;
                      reg1186 <= $signed((^~$unsigned(reg1185[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg1185 <= (^~reg1181[(1'h1):(1'h1)]);
                      reg1186 <= $signed((wire1174[(1'h0):(1'h0)] ?
                          (+wire1179) : (~&(wire1179 && forvar1180))));
                    end
                end
              for (forvar1189 = (1'h0); (forvar1189 < (1'h1)); forvar1189 = (forvar1189 + (1'h1)))
                begin
                  for (forvar1190 = (1'h0); (forvar1190 < (2'h3)); forvar1190 = (forvar1190 + (1'h1)))
                    begin
                      reg1191 <= (~&reg1183);
                      reg1192 <= $unsigned(wire1176);
                      reg1193 <= {(reg1184[(3'h5):(3'h5)] ?
                              (reg1185[(1'h1):(1'h0)] ^ (8'hb2)) : (&forvar1189[(1'h0):(1'h0)]))};
                    end
                end
              for (forvar1194 = (1'h0); (forvar1194 < (2'h2)); forvar1194 = (forvar1194 + (1'h1)))
                begin
                  for (forvar1195 = (1'h0); (forvar1195 < (1'h1)); forvar1195 = (forvar1195 + (1'h1)))
                    begin
                      reg1196 <= reg1181[(4'hb):(3'h6)];
                    end
                  for (forvar1197 = (1'h0); (forvar1197 < (2'h2)); forvar1197 = (forvar1197 + (1'h1)))
                    begin
                      reg1198 <= {(({reg1181} ?
                                  (reg1182 - forvar1185) : $unsigned(forvar1194)) ?
                              (forvar1181 ?
                                  reg1184 : {wire1178}) : (&(+(8'ha0))))};
                      reg1199 <= (&forvar1194);
                      reg1200 <= {reg1188[(2'h3):(1'h1)]};
                    end
                end
            end
        end
      else
        begin
          if (((wire1178 ? reg1185 : $unsigned(reg1183)) ^ (+(+(~^reg1188)))))
            begin
              for (forvar1180 = (1'h0); (forvar1180 < (1'h0)); forvar1180 = (forvar1180 + (1'h1)))
                begin
                  for (forvar1181 = (1'h0); (forvar1181 < (2'h2)); forvar1181 = (forvar1181 + (1'h1)))
                    begin
                      reg1182 <= reg1193;
                      reg1183 <= forvar1195;
                      reg1184 <= wire1177;
                    end
                  if ($unsigned({$signed($signed(forvar1181))}))
                    begin
                      reg1185 <= $unsigned($unsigned((^$signed((8'hb6)))));
                      reg1186 <= $signed($unsigned(wire1178[(3'h5):(1'h1)]));
                      reg1187 <= $unsigned(reg1188);
                    end
                  else
                    begin
                      reg1185 <= {(+reg1198[(2'h2):(2'h2)])};
                      reg1186 <= $unsigned(({(|reg1199)} > (^(reg1196 <<< forvar1180))));
                      reg1187 <= $signed($unsigned(reg1184[(2'h2):(2'h2)]));
                      reg1188 <= wire1178;
                    end
                  if (forvar1194[(1'h0):(1'h0)])
                    begin
                      reg1189 <= $unsigned($signed($signed((reg1184 == reg1181))));
                    end
                  else
                    begin
                      reg1189 <= forvar1194[(1'h0):(1'h0)];
                      reg1190 <= $unsigned($unsigned(wire1176[(1'h1):(1'h1)]));
                      reg1191 <= (forvar1190 <= ((-(~^wire1179)) ?
                          ((!wire1174) ?
                              (8'ha1) : (&reg1191)) : (~(wire1177 & reg1183))));
                      reg1192 <= ($unsigned(reg1189[(3'h4):(1'h1)]) ?
                          $signed(((~forvar1195) ?
                              (8'hae) : reg1191[(2'h2):(1'h1)])) : (~&$unsigned((reg1185 ?
                              reg1190 : reg1200))));
                    end
                  for (forvar1193 = (1'h0); (forvar1193 < (1'h0)); forvar1193 = (forvar1193 + (1'h1)))
                    begin
                      reg1194 <= $unsigned(($unsigned((wire1179 ?
                              (8'ha4) : reg1193)) ?
                          ((reg1182 ?
                              reg1189 : wire1175) <= reg1192) : $signed($unsigned(reg1187))));
                    end
                end
              if (forvar1181[(1'h0):(1'h0)])
                begin
                  if (forvar1194)
                    begin
                      reg1195 <= $signed({forvar1197});
                      reg1196 <= (reg1193 ?
                          ($unsigned((^wire1175)) < reg1199) : ($unsigned($unsigned(wire1175)) * ($signed(reg1190) ?
                              $signed((8'hb9)) : (reg1188 && wire1177))));
                    end
                  else
                    begin
                      reg1195 <= $signed($unsigned($unsigned($unsigned(reg1185))));
                      reg1196 <= (~|$unsigned($signed($signed(reg1190))));
                    end
                  reg1197 <= (~^{reg1183});
                end
              else
                begin
                  for (forvar1195 = (1'h0); (forvar1195 < (1'h1)); forvar1195 = (forvar1195 + (1'h1)))
                    begin
                      reg1196 <= reg1194[(3'h6):(1'h1)];
                      reg1197 <= $signed(((wire1178[(1'h1):(1'h1)] <<< (reg1189 ?
                              (8'ha9) : wire1177)) ?
                          reg1196 : ((reg1183 ? reg1188 : reg1196) ?
                              forvar1185[(2'h2):(1'h1)] : reg1187[(2'h3):(1'h1)])));
                      reg1198 <= $unsigned(reg1197);
                      reg1199 <= reg1188[(3'h4):(2'h2)];
                    end
                end
              for (forvar1200 = (1'h0); (forvar1200 < (1'h1)); forvar1200 = (forvar1200 + (1'h1)))
                begin
                  if (reg1181[(3'h5):(1'h1)])
                    begin
                      reg1201 <= (8'h9d);
                    end
                  else
                    begin
                      reg1201 <= wire1176;
                    end
                  for (forvar1202 = (1'h0); (forvar1202 < (2'h3)); forvar1202 = (forvar1202 + (1'h1)))
                    begin
                      reg1203 <= $unsigned($signed($unsigned($signed(forvar1200))));
                      reg1204 <= ((|(~^forvar1200)) < ($unsigned(reg1190[(2'h3):(2'h3)]) << (reg1198[(1'h0):(1'h0)] >= reg1187[(2'h2):(1'h1)])));
                      reg1205 <= reg1188;
                    end
                end
              reg1206 <= {wire1179[(3'h4):(2'h3)]};
            end
          else
            begin
              if ((8'hab))
                begin
                  for (forvar1180 = (1'h0); (forvar1180 < (1'h0)); forvar1180 = (forvar1180 + (1'h1)))
                    begin
                      reg1181 <= ((reg1181[(3'h7):(3'h6)] ?
                          wire1176 : ((~wire1179) ?
                              {reg1184} : (forvar1193 ?
                                  wire1177 : reg1188))) >>> ((~&(reg1191 > forvar1200)) == (~&((8'h9d) <= reg1204))));
                    end
                  for (forvar1182 = (1'h0); (forvar1182 < (2'h2)); forvar1182 = (forvar1182 + (1'h1)))
                    begin
                      reg1183 <= $signed($signed(((+reg1192) ?
                          (reg1203 && forvar1193) : (~&reg1187))));
                    end
                  if (($unsigned(((-forvar1195) ? (!reg1186) : reg1198)) ?
                      reg1199 : forvar1185[(1'h1):(1'h0)]))
                    begin
                      reg1184 <= forvar1181;
                      reg1185 <= (!$signed(($unsigned(reg1205) ?
                          reg1187 : {reg1189})));
                      reg1186 <= (reg1206 ?
                          ($signed({forvar1182}) ?
                              (~&(~|wire1174)) : $unsigned($signed((8'h9d)))) : $signed((-forvar1193[(1'h1):(1'h0)])));
                      reg1187 <= ((~&(8'hb7)) * $unsigned(({forvar1193} > forvar1182[(3'h5):(1'h0)])));
                    end
                  else
                    begin
                      reg1184 <= $signed((reg1199[(1'h1):(1'h0)] ^~ reg1198[(1'h1):(1'h0)]));
                      reg1185 <= {(8'ha1)};
                      reg1186 <= forvar1197[(2'h2):(1'h0)];
                      reg1187 <= ($unsigned((+$signed((8'hae)))) ?
                          reg1191 : reg1198);
                    end
                  for (forvar1188 = (1'h0); (forvar1188 < (2'h2)); forvar1188 = (forvar1188 + (1'h1)))
                    begin
                      reg1189 <= (8'hab);
                    end
                end
              else
                begin
                  for (forvar1180 = (1'h0); (forvar1180 < (1'h0)); forvar1180 = (forvar1180 + (1'h1)))
                    begin
                      reg1181 <= $unsigned($signed($signed({wire1178})));
                      reg1182 <= $unsigned(((&(forvar1182 ?
                          reg1188 : wire1176)) && wire1177));
                    end
                  for (forvar1183 = (1'h0); (forvar1183 < (2'h2)); forvar1183 = (forvar1183 + (1'h1)))
                    begin
                      reg1184 <= (forvar1190[(1'h0):(1'h0)] ?
                          ((^((8'ha9) ? reg1188 : reg1204)) >> (+(forvar1189 ?
                              forvar1190 : forvar1188))) : reg1200);
                      reg1185 <= forvar1202[(1'h1):(1'h0)];
                      reg1186 <= (reg1190[(3'h7):(3'h4)] ?
                          $unsigned($unsigned((reg1198 ^~ reg1201))) : ($signed({forvar1194}) ?
                              reg1187 : {$unsigned(forvar1189)}));
                      reg1187 <= forvar1189;
                    end
                  if ($signed(reg1192[(3'h6):(2'h2)]))
                    begin
                      reg1188 <= reg1201;
                      reg1189 <= forvar1194[(2'h2):(2'h2)];
                      reg1190 <= {(-(~|reg1197[(3'h5):(2'h3)]))};
                      reg1191 <= reg1206;
                    end
                  else
                    begin
                      reg1188 <= forvar1189;
                    end
                end
              reg1192 <= reg1194;
              for (forvar1193 = (1'h0); (forvar1193 < (1'h0)); forvar1193 = (forvar1193 + (1'h1)))
                begin
                  for (forvar1194 = (1'h0); (forvar1194 < (2'h3)); forvar1194 = (forvar1194 + (1'h1)))
                    begin
                      reg1195 <= reg1193;
                    end
                end
              if ((!$unsigned($unsigned(reg1198))))
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (1'h0)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= reg1185[(1'h1):(1'h1)];
                    end
                  for (forvar1198 = (1'h0); (forvar1198 < (1'h0)); forvar1198 = (forvar1198 + (1'h1)))
                    begin
                      reg1199 <= $signed(($signed($signed(forvar1198)) >>> ((^reg1190) ?
                          $unsigned(forvar1198) : $unsigned((8'hb5)))));
                      reg1200 <= (|{forvar1196[(3'h4):(2'h2)]});
                      reg1201 <= {{$unsigned($unsigned((8'ha1)))}};
                      reg1202 <= (^~reg1190[(3'h5):(1'h1)]);
                    end
                  for (forvar1203 = (1'h0); (forvar1203 < (2'h3)); forvar1203 = (forvar1203 + (1'h1)))
                    begin
                      reg1204 <= reg1196[(4'h9):(4'h8)];
                      reg1205 <= reg1206[(3'h6):(2'h2)];
                      reg1206 <= reg1184[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (2'h3)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= $signed({(forvar1190 ?
                              $unsigned(reg1191) : reg1192)});
                      reg1198 <= ((~&wire1178) < (forvar1200[(4'hd):(3'h4)] ^ (forvar1197[(2'h2):(2'h2)] ?
                          (^reg1200) : (reg1202 ? reg1181 : (8'had)))));
                      reg1199 <= (^wire1174);
                    end
                  for (forvar1200 = (1'h0); (forvar1200 < (1'h0)); forvar1200 = (forvar1200 + (1'h1)))
                    begin
                      reg1201 <= wire1174[(3'h4):(1'h0)];
                    end
                  for (forvar1202 = (1'h0); (forvar1202 < (1'h0)); forvar1202 = (forvar1202 + (1'h1)))
                    begin
                      reg1203 <= (&$unsigned((forvar1202 ^~ (^~forvar1202))));
                      reg1204 <= reg1201;
                      reg1205 <= (reg1197 ?
                          reg1204[(2'h2):(1'h0)] : (($unsigned(forvar1180) ?
                                  (8'hab) : (+reg1201)) ?
                              ($unsigned(reg1189) << (+(8'hb5))) : reg1182[(1'h1):(1'h0)]));
                    end
                end
            end
        end
    end
  assign wire1207 = forvar1200[(4'ha):(1'h1)];
  assign wire1208 = (~^(forvar1180 >> {forvar1189[(3'h4):(2'h3)]}));
  assign wire1209 = forvar1203;
  assign wire1210 = (((!(reg1193 | forvar1195)) ?
                        $signed($signed(reg1187)) : ($unsigned(reg1199) != ((8'hae) ^ reg1193))) | ((forvar1203 ?
                            reg1206[(4'hc):(3'h7)] : (reg1196 | wire1177)) ?
                        wire1175[(2'h3):(2'h3)] : $signed((~|forvar1198))));
  always
    @(posedge clk) begin
      reg1211 <= (forvar1198 < $signed(forvar1181[(1'h1):(1'h1)]));
    end
  always
    @(posedge clk) begin
      for (forvar1212 = (1'h0); (forvar1212 < (2'h2)); forvar1212 = (forvar1212 + (1'h1)))
        begin
          if (($signed($unsigned($unsigned(forvar1197))) ?
              (forvar1188[(3'h4):(1'h0)] == {wire1174[(3'h5):(1'h0)]}) : reg1201))
            begin
              reg1213 <= reg1200[(3'h4):(1'h1)];
              for (forvar1214 = (1'h0); (forvar1214 < (2'h2)); forvar1214 = (forvar1214 + (1'h1)))
                begin
                  reg1215 <= $unsigned((((wire1210 ? (8'hb4) : reg1189) ?
                          $unsigned(reg1183) : $unsigned(reg1185)) ?
                      {$signed(forvar1195)} : ($unsigned((8'hb3)) >> (reg1211 ^ wire1177))));
                end
              if ($signed($unsigned(wire1179[(4'h9):(4'h9)])))
                begin
                  if (reg1190)
                    begin
                      reg1216 <= {{(-{forvar1202})}};
                      reg1217 <= forvar1203[(4'h9):(1'h1)];
                      reg1218 <= reg1195[(3'h4):(1'h1)];
                      reg1219 <= $signed($unsigned({(forvar1182 ^~ reg1196)}));
                    end
                  else
                    begin
                      reg1216 <= (((!$unsigned((8'hb5))) ^ ($unsigned((8'hb8)) ^~ (&reg1219))) ?
                          forvar1180[(1'h1):(1'h0)] : (forvar1185 ?
                              $signed((reg1194 ?
                                  reg1202 : reg1196)) : ((wire1207 && reg1206) ?
                                  {forvar1181} : forvar1196)));
                      reg1217 <= $signed((~^({reg1203} ?
                          $unsigned((8'hb8)) : $signed(reg1200))));
                      reg1218 <= {$signed((~reg1219[(3'h7):(1'h0)]))};
                      reg1219 <= (8'hb7);
                    end
                  for (forvar1220 = (1'h0); (forvar1220 < (1'h0)); forvar1220 = (forvar1220 + (1'h1)))
                    begin
                      reg1221 <= ((forvar1185[(1'h1):(1'h1)] ?
                          ((~&wire1177) ?
                              (forvar1189 ?
                                  forvar1183 : forvar1188) : reg1185[(2'h3):(1'h0)]) : (forvar1188[(3'h5):(3'h5)] ?
                              reg1213 : (^reg1218))) ^~ wire1174[(1'h0):(1'h0)]);
                      reg1222 <= forvar1185[(1'h0):(1'h0)];
                      reg1223 <= (~^$signed($unsigned($unsigned(wire1177))));
                    end
                end
              else
                begin
                  if ($unsigned(($signed(reg1181[(1'h1):(1'h1)]) << (((8'haa) ?
                          forvar1190 : forvar1200) ?
                      $signed(forvar1180) : $unsigned(forvar1220)))))
                    begin
                      reg1216 <= reg1194;
                      reg1217 <= (forvar1195[(2'h2):(2'h2)] ?
                          (((wire1175 * forvar1198) ?
                                  (8'hae) : (forvar1198 << reg1217)) ?
                              $unsigned({forvar1181}) : $signed(reg1213[(4'h8):(3'h7)])) : ($signed((reg1217 & wire1208)) >> $signed((-reg1213))));
                      reg1218 <= (|$unsigned((&$signed(reg1202))));
                    end
                  else
                    begin
                      reg1216 <= reg1189;
                      reg1217 <= $signed($unsigned(forvar1200));
                    end
                end
              if (reg1198[(1'h0):(1'h0)])
                begin
                  for (forvar1224 = (1'h0); (forvar1224 < (1'h0)); forvar1224 = (forvar1224 + (1'h1)))
                    begin
                      reg1225 <= $unsigned(forvar1195);
                      reg1226 <= $signed($signed(((~&reg1183) ?
                          $signed(forvar1212) : (reg1192 <<< forvar1196))));
                    end
                  if (forvar1194[(2'h2):(2'h2)])
                    begin
                      reg1227 <= (((reg1215[(4'hd):(3'h6)] ^~ forvar1196[(3'h5):(3'h4)]) ?
                              (8'hae) : $signed((wire1208 ^ wire1176))) ?
                          forvar1190[(2'h2):(1'h1)] : (reg1193[(2'h2):(2'h2)] ?
                              ((-reg1219) ?
                                  reg1205[(1'h0):(1'h0)] : wire1207[(3'h5):(2'h2)]) : $unsigned((&forvar1196))));
                      reg1228 <= forvar1185;
                      reg1229 <= reg1202[(3'h6):(1'h0)];
                      reg1230 <= $unsigned($unsigned($signed((reg1199 && reg1229))));
                    end
                  else
                    begin
                      reg1227 <= (reg1185 ?
                          (((8'hae) * (-reg1184)) ~^ forvar1190) : $signed((8'hab)));
                    end
                end
              else
                begin
                  for (forvar1224 = (1'h0); (forvar1224 < (1'h0)); forvar1224 = (forvar1224 + (1'h1)))
                    begin
                      reg1225 <= reg1206[(4'hd):(4'ha)];
                    end
                  if ($signed(reg1186))
                    begin
                      reg1226 <= {(+reg1217[(1'h1):(1'h0)])};
                      reg1227 <= ($signed({forvar1180}) ?
                          (8'ha6) : ($signed((reg1192 >>> forvar1188)) || reg1184[(4'h9):(3'h5)]));
                      reg1228 <= (reg1222[(2'h3):(1'h1)] ?
                          (~$signed(wire1209[(4'hc):(2'h3)])) : reg1216[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1226 <= (((forvar1198 >= (~|wire1175)) ^ {$signed(wire1209)}) ?
                          $signed($unsigned($unsigned(forvar1220))) : $unsigned(($unsigned((8'ha5)) ?
                              {reg1195} : $signed(reg1182))));
                      reg1227 <= (^(|({forvar1202} < reg1218[(1'h1):(1'h0)])));
                    end
                  reg1229 <= ({((reg1227 ?
                          forvar1182 : wire1174) <<< (+wire1178))} <= $unsigned(($unsigned(forvar1214) ?
                      (reg1190 || reg1204) : (wire1208 ? (8'hb0) : reg1216))));
                end
            end
          else
            begin
              if ($signed((~|((reg1219 ? forvar1188 : forvar1203) ?
                  reg1204 : $unsigned(reg1230)))))
                begin
                  reg1213 <= ($signed($unsigned((forvar1224 ?
                          reg1189 : reg1189))) ?
                      $unsigned($signed({reg1197})) : $unsigned(reg1223[(1'h1):(1'h1)]));
                  for (forvar1214 = (1'h0); (forvar1214 < (2'h3)); forvar1214 = (forvar1214 + (1'h1)))
                    begin
                      reg1215 <= $unsigned({((8'hb5) > $signed((8'hb3)))});
                      reg1216 <= reg1198[(2'h2):(1'h0)];
                      reg1217 <= reg1223[(1'h1):(1'h0)];
                      reg1218 <= reg1190;
                    end
                end
              else
                begin
                  if ((reg1185[(1'h0):(1'h0)] ?
                      $signed(((reg1215 << reg1202) ?
                          $signed(wire1177) : (~&(8'hab)))) : (+reg1211)))
                    begin
                      reg1213 <= wire1210;
                      reg1214 <= $signed((reg1219[(3'h7):(3'h4)] << {(wire1179 != wire1208)}));
                    end
                  else
                    begin
                      reg1213 <= $unsigned($unsigned(((!forvar1189) <<< forvar1190)));
                    end
                  for (forvar1215 = (1'h0); (forvar1215 < (2'h2)); forvar1215 = (forvar1215 + (1'h1)))
                    begin
                      reg1216 <= reg1229;
                      reg1217 <= ($unsigned($signed({wire1179})) ?
                          reg1197[(2'h3):(1'h1)] : $signed($unsigned((forvar1197 <<< forvar1196))));
                      reg1218 <= forvar1188[(1'h1):(1'h0)];
                    end
                end
              if (({reg1215[(1'h0):(1'h0)]} ?
                  wire1175 : reg1222[(4'hb):(1'h0)]))
                begin
                  if (((reg1216[(2'h2):(2'h2)] ?
                          {reg1195} : {reg1189[(1'h0):(1'h0)]}) ?
                      ({$signed(forvar1195)} ?
                          $signed((reg1192 & wire1174)) : forvar1188[(3'h4):(1'h0)]) : $signed((~&(reg1202 + reg1192)))))
                    begin
                      reg1219 <= $unsigned($unsigned(($signed(reg1197) ?
                          $signed(forvar1212) : $unsigned(forvar1200))));
                    end
                  else
                    begin
                      reg1219 <= ($signed(((forvar1185 ? forvar1185 : reg1200) ?
                              $signed(reg1215) : $unsigned(wire1176))) ?
                          (reg1184 || $unsigned((8'hb0))) : reg1197[(2'h3):(2'h3)]);
                    end
                  for (forvar1220 = (1'h0); (forvar1220 < (1'h1)); forvar1220 = (forvar1220 + (1'h1)))
                    begin
                      reg1221 <= ((~&$unsigned(reg1228[(4'ha):(4'h9)])) ?
                          $signed(reg1191) : (reg1199 ^ reg1196));
                      reg1222 <= wire1209[(5'h10):(1'h1)];
                    end
                  for (forvar1223 = (1'h0); (forvar1223 < (2'h3)); forvar1223 = (forvar1223 + (1'h1)))
                    begin
                      reg1224 <= wire1178;
                      reg1225 <= reg1202[(4'ha):(2'h3)];
                      reg1226 <= reg1225[(3'h6):(3'h4)];
                      reg1227 <= ($signed({(wire1176 ?
                              (8'h9f) : forvar1181)}) <<< $signed((forvar1188[(2'h2):(1'h0)] != $signed(reg1190))));
                    end
                  if (($signed(reg1191[(2'h3):(1'h0)]) ?
                      (~$unsigned($unsigned((8'ha7)))) : reg1182[(1'h0):(1'h0)]))
                    begin
                      reg1228 <= ($unsigned((^$signed(reg1194))) <= reg1198);
                    end
                  else
                    begin
                      reg1228 <= (forvar1198[(1'h1):(1'h1)] ?
                          reg1219[(3'h7):(3'h7)] : wire1175);
                    end
                end
              else
                begin
                  if (((((reg1185 != reg1186) ?
                      reg1204[(1'h0):(1'h0)] : $unsigned(forvar1198)) >= $signed((wire1208 ~^ (8'hb1)))) <<< ((^wire1175[(1'h0):(1'h0)]) - reg1203)))
                    begin
                      reg1219 <= (($unsigned((reg1184 ^~ (8'ha2))) == $signed(reg1206)) ^ wire1210);
                    end
                  else
                    begin
                      reg1219 <= forvar1220;
                      reg1220 <= {reg1200};
                      reg1221 <= $unsigned({(~&(reg1228 || reg1218))});
                      reg1222 <= $unsigned((+$unsigned($signed((8'ha9)))));
                    end
                  for (forvar1223 = (1'h0); (forvar1223 < (1'h0)); forvar1223 = (forvar1223 + (1'h1)))
                    begin
                      reg1224 <= (($unsigned((reg1186 ~^ (8'hac))) <<< ({reg1198} ?
                          $signed(forvar1195) : forvar1183[(1'h0):(1'h0)])) << forvar1181[(2'h3):(2'h3)]);
                    end
                  for (forvar1225 = (1'h0); (forvar1225 < (2'h2)); forvar1225 = (forvar1225 + (1'h1)))
                    begin
                      reg1226 <= ((~|($signed(reg1206) >> forvar1188)) ?
                          (forvar1189 >= wire1209[(3'h6):(3'h5)]) : ((|(!reg1191)) ?
                              ((reg1191 ?
                                  forvar1215 : reg1194) && (forvar1225 ^ forvar1203)) : (8'ha6)));
                      reg1227 <= (reg1213 ?
                          reg1202[(3'h6):(1'h0)] : reg1190[(3'h6):(1'h0)]);
                      reg1228 <= $unsigned($unsigned((~&{reg1195})));
                    end
                end
              for (forvar1229 = (1'h0); (forvar1229 < (1'h1)); forvar1229 = (forvar1229 + (1'h1)))
                begin
                  for (forvar1230 = (1'h0); (forvar1230 < (2'h2)); forvar1230 = (forvar1230 + (1'h1)))
                    begin
                      reg1231 <= $unsigned((!$unsigned((forvar1229 ?
                          forvar1203 : reg1217))));
                      reg1232 <= $unsigned(reg1220);
                      reg1233 <= (reg1230 ? reg1182[(4'h8):(1'h0)] : reg1232);
                    end
                  for (forvar1234 = (1'h0); (forvar1234 < (2'h2)); forvar1234 = (forvar1234 + (1'h1)))
                    begin
                      reg1235 <= $unsigned(forvar1182);
                      reg1236 <= $unsigned((((reg1188 ? reg1230 : wire1208) ?
                          $signed(forvar1195) : reg1221) >= (~reg1195)));
                      reg1237 <= (~&((wire1179 >> (reg1185 ?
                              reg1214 : wire1209)) ?
                          $unsigned((reg1194 ?
                              reg1231 : reg1191)) : forvar1193));
                    end
                end
            end
          reg1238 <= ((((8'haf) ?
                  (reg1230 || reg1183) : $unsigned(reg1227)) ~^ $signed(reg1232)) ?
              $signed($signed(reg1197)) : reg1197[(1'h0):(1'h0)]);
          if ((($unsigned(reg1217) && (|$signed(forvar1198))) ?
              {($signed(reg1235) >>> ((8'hb5) ?
                      reg1202 : forvar1197))} : (reg1225[(3'h7):(1'h0)] ?
                  {reg1183} : $unsigned({reg1223}))))
            begin
              reg1239 <= (&$unsigned((forvar1182[(1'h0):(1'h0)] && reg1188[(2'h2):(2'h2)])));
              for (forvar1240 = (1'h0); (forvar1240 < (2'h2)); forvar1240 = (forvar1240 + (1'h1)))
                begin
                  for (forvar1241 = (1'h0); (forvar1241 < (1'h0)); forvar1241 = (forvar1241 + (1'h1)))
                    begin
                      reg1242 <= (($signed((!(8'h9e))) & (~|forvar1180[(2'h2):(1'h1)])) >> $signed(reg1221[(4'hc):(4'h8)]));
                      reg1243 <= ((reg1220[(1'h0):(1'h0)] ?
                          $unsigned($unsigned(reg1237)) : (!(forvar1214 ?
                              reg1218 : forvar1195))) != wire1175);
                      reg1244 <= reg1188;
                    end
                  for (forvar1245 = (1'h0); (forvar1245 < (2'h2)); forvar1245 = (forvar1245 + (1'h1)))
                    begin
                      reg1246 <= forvar1197;
                      reg1247 <= forvar1196;
                    end
                end
            end
          else
            begin
              reg1239 <= (8'hba);
              for (forvar1240 = (1'h0); (forvar1240 < (1'h0)); forvar1240 = (forvar1240 + (1'h1)))
                begin
                  if ($unsigned(reg1195[(1'h1):(1'h0)]))
                    begin
                      reg1241 <= ((({(8'hb4)} * reg1244[(3'h4):(2'h3)]) ?
                              ((reg1196 * wire1174) >= reg1247) : ((|(8'ha0)) ?
                                  forvar1196 : reg1191[(3'h4):(2'h2)])) ?
                          $signed(({reg1231} >>> (reg1214 ?
                              reg1202 : reg1226))) : (-(8'hae)));
                    end
                  else
                    begin
                      reg1241 <= $unsigned($signed(($unsigned(reg1244) ?
                          (^~reg1205) : (reg1229 >> wire1177))));
                    end
                  if ($unsigned(forvar1185[(1'h0):(1'h0)]))
                    begin
                      reg1242 <= $unsigned((($unsigned((8'hab)) ?
                          (reg1221 >> reg1181) : $unsigned(reg1185)) | ($signed(reg1222) << $signed(reg1232))));
                      reg1243 <= ($unsigned(reg1200[(3'h4):(2'h3)]) << $signed((forvar1225 ^~ $signed(reg1233))));
                      reg1244 <= $unsigned(reg1218);
                      reg1245 <= reg1185;
                    end
                  else
                    begin
                      reg1242 <= reg1224[(3'h6):(1'h1)];
                      reg1243 <= $signed(reg1182[(1'h0):(1'h0)]);
                    end
                  for (forvar1246 = (1'h0); (forvar1246 < (1'h1)); forvar1246 = (forvar1246 + (1'h1)))
                    begin
                      reg1247 <= {({$signed(reg1231)} ?
                              ($unsigned((8'haf)) ?
                                  reg1238 : (forvar1229 == forvar1189)) : (-(reg1226 && (8'haa))))};
                      reg1248 <= (~|(!reg1203));
                    end
                  for (forvar1249 = (1'h0); (forvar1249 < (1'h0)); forvar1249 = (forvar1249 + (1'h1)))
                    begin
                      reg1250 <= $signed((^~$unsigned((-(8'ha6)))));
                      reg1251 <= (~^reg1197);
                    end
                end
              reg1252 <= $signed((reg1246[(4'hb):(1'h1)] ?
                  reg1202[(1'h1):(1'h0)] : (&((8'ha8) ? reg1232 : reg1218))));
            end
        end
      for (forvar1253 = (1'h0); (forvar1253 < (2'h2)); forvar1253 = (forvar1253 + (1'h1)))
        begin
          if ($unsigned(forvar1234[(4'he):(1'h1)]))
            begin
              if (((reg1204 ?
                      $signed(forvar1190) : $signed($unsigned(reg1191))) ?
                  (+$signed($unsigned(reg1230))) : ((~^(!(8'ha4))) - {(reg1194 ?
                          forvar1203 : reg1247)})))
                begin
                  for (forvar1254 = (1'h0); (forvar1254 < (2'h3)); forvar1254 = (forvar1254 + (1'h1)))
                    begin
                      reg1255 <= {reg1197[(3'h5):(1'h1)]};
                      reg1256 <= ($signed((^~$unsigned(forvar1215))) && $signed(wire1207[(2'h2):(2'h2)]));
                      reg1257 <= {{reg1186[(4'h9):(3'h7)]}};
                      reg1258 <= {(reg1216 ?
                              $unsigned($signed((8'hb6))) : ((reg1257 ?
                                      reg1221 : (8'h9c)) ?
                                  reg1248[(4'hb):(4'ha)] : (reg1187 ?
                                      reg1192 : (8'haa))))};
                    end
                  reg1259 <= forvar1229[(3'h4):(1'h0)];
                end
              else
                begin
                  for (forvar1254 = (1'h0); (forvar1254 < (1'h0)); forvar1254 = (forvar1254 + (1'h1)))
                    begin
                      reg1255 <= reg1244[(2'h3):(1'h1)];
                    end
                  if (($unsigned((-(~^forvar1230))) ?
                      ($signed(forvar1220[(3'h7):(1'h0)]) >>> (forvar1197 ?
                          (8'hba) : {forvar1193})) : reg1256))
                    begin
                      reg1256 <= (|(^~reg1206));
                      reg1257 <= (forvar1202[(4'hc):(3'h7)] ?
                          (((reg1215 != reg1236) ? (-reg1222) : reg1203) ?
                              ($signed(forvar1185) ?
                                  forvar1182 : (reg1226 ?
                                      reg1198 : forvar1214)) : {wire1210[(4'ha):(2'h3)]}) : $unsigned((|$signed(reg1250))));
                    end
                  else
                    begin
                      reg1256 <= (^$signed((reg1186[(2'h3):(2'h3)] ?
                          wire1208 : (^~reg1189))));
                    end
                  for (forvar1258 = (1'h0); (forvar1258 < (1'h0)); forvar1258 = (forvar1258 + (1'h1)))
                    begin
                      reg1259 <= (~|(forvar1258[(2'h3):(1'h0)] ?
                          reg1216 : $unsigned($unsigned(reg1205))));
                      reg1260 <= ((($unsigned(reg1232) || $signed(forvar1215)) << reg1239) ?
                          reg1225[(4'h8):(3'h5)] : reg1230[(2'h2):(1'h0)]);
                      reg1261 <= reg1229[(3'h4):(1'h1)];
                    end
                  for (forvar1262 = (1'h0); (forvar1262 < (1'h1)); forvar1262 = (forvar1262 + (1'h1)))
                    begin
                      reg1263 <= ($unsigned(forvar1185) ?
                          {((reg1242 ?
                                  forvar1203 : forvar1182) ^~ reg1211)} : $unsigned($signed((wire1174 >= reg1236))));
                      reg1264 <= (~^wire1175[(2'h3):(2'h3)]);
                      reg1265 <= $signed((|((~&forvar1249) ?
                          {wire1174} : wire1207)));
                    end
                end
              for (forvar1266 = (1'h0); (forvar1266 < (2'h3)); forvar1266 = (forvar1266 + (1'h1)))
                begin
                  for (forvar1267 = (1'h0); (forvar1267 < (2'h2)); forvar1267 = (forvar1267 + (1'h1)))
                    begin
                      reg1268 <= reg1243[(3'h4):(1'h0)];
                      reg1269 <= reg1259;
                      reg1270 <= ($unsigned({$signed((8'hb5))}) ?
                          wire1178[(3'h4):(1'h1)] : (($unsigned(reg1242) ^ (8'ha1)) >> ((+forvar1183) | (8'hb3))));
                      reg1271 <= (|{$unsigned((~reg1251))});
                    end
                end
            end
          else
            begin
              if ($signed(forvar1189[(4'hd):(2'h3)]))
                begin
                  if ($unsigned({(~^((8'haf) & (8'h9c)))}))
                    begin
                      reg1254 <= (^~forvar1182);
                    end
                  else
                    begin
                      reg1254 <= reg1255;
                    end
                  for (forvar1255 = (1'h0); (forvar1255 < (1'h0)); forvar1255 = (forvar1255 + (1'h1)))
                    begin
                      reg1256 <= (^~reg1239);
                      reg1257 <= {({forvar1195} * ((reg1219 ~^ forvar1220) <= (reg1225 ?
                              reg1217 : (8'h9d))))};
                    end
                  if ({(-((reg1264 ? reg1192 : forvar1249) <= reg1242))})
                    begin
                      reg1258 <= (reg1203 ? reg1197[(3'h5):(3'h4)] : (8'hb6));
                      reg1259 <= $signed(reg1186);
                      reg1260 <= $signed(forvar1180);
                      reg1261 <= (forvar1220[(3'h5):(1'h0)] ?
                          $signed(($unsigned(reg1220) ?
                              $unsigned(forvar1182) : (reg1228 ?
                                  reg1259 : reg1196))) : reg1201);
                    end
                  else
                    begin
                      reg1258 <= $signed(reg1228);
                    end
                  for (forvar1262 = (1'h0); (forvar1262 < (2'h2)); forvar1262 = (forvar1262 + (1'h1)))
                    begin
                      reg1263 <= reg1225[(3'h4):(2'h3)];
                      reg1264 <= forvar1249;
                    end
                end
              else
                begin
                  if (((^$signed({(8'hb8)})) && $unsigned(($signed(wire1178) * forvar1194[(1'h1):(1'h0)]))))
                    begin
                      reg1254 <= forvar1200;
                      reg1255 <= $signed($signed(($signed(wire1178) ?
                          (&wire1176) : (forvar1224 ? forvar1180 : reg1199))));
                      reg1256 <= reg1182[(4'h9):(2'h2)];
                      reg1257 <= (forvar1253 ?
                          $unsigned((!(&(8'hba)))) : (((^~reg1198) ?
                              $unsigned(reg1197) : (reg1193 ?
                                  (8'hb5) : reg1260)) | ((~&forvar1253) ?
                              $unsigned(reg1265) : (reg1219 ?
                                  forvar1185 : reg1261))));
                    end
                  else
                    begin
                      reg1254 <= reg1215[(4'h8):(1'h0)];
                      reg1255 <= ($signed((forvar1224[(3'h4):(3'h4)] + {forvar1188})) <<< $signed({(reg1223 ?
                              (8'haf) : forvar1183)}));
                    end
                end
              for (forvar1265 = (1'h0); (forvar1265 < (2'h3)); forvar1265 = (forvar1265 + (1'h1)))
                begin
                  if ((((((8'hba) ? (8'hba) : reg1187) ^~ reg1263) ?
                      reg1218[(2'h2):(1'h0)] : (reg1206 ?
                          reg1205[(1'h0):(1'h0)] : (reg1191 > reg1233))) && reg1191))
                    begin
                      reg1266 <= (8'hb3);
                      reg1267 <= (reg1269[(3'h4):(2'h3)] ?
                          reg1259[(3'h6):(2'h2)] : ($unsigned($signed(wire1179)) ?
                              $unsigned((8'hb2)) : (&reg1231)));
                      reg1268 <= {(8'haa)};
                    end
                  else
                    begin
                      reg1266 <= (forvar1241 <<< ((8'haa) ?
                          (|(forvar1255 ? reg1271 : (8'haf))) : reg1204));
                      reg1267 <= (~wire1207);
                      reg1268 <= {((^~reg1189) ?
                              (+forvar1224[(3'h4):(1'h0)]) : reg1258[(4'ha):(2'h3)])};
                    end
                  for (forvar1269 = (1'h0); (forvar1269 < (1'h0)); forvar1269 = (forvar1269 + (1'h1)))
                    begin
                      reg1270 <= ($signed((-(reg1201 ? reg1241 : wire1178))) ?
                          {($unsigned(reg1225) ?
                                  forvar1197[(2'h2):(1'h0)] : $unsigned((8'ha3)))} : ({forvar1180} + ($unsigned(reg1237) ?
                              (forvar1185 | reg1246) : (forvar1197 ~^ wire1210))));
                    end
                end
              reg1271 <= ((((^~forvar1195) ?
                      reg1188 : (~^reg1252)) >> {forvar1202}) ?
                  forvar1241 : (reg1261[(2'h2):(1'h0)] ?
                      reg1270[(3'h6):(2'h2)] : (&wire1174)));
            end
          for (forvar1272 = (1'h0); (forvar1272 < (1'h0)); forvar1272 = (forvar1272 + (1'h1)))
            begin
              if (wire1178[(2'h3):(1'h1)])
                begin
                  for (forvar1273 = (1'h0); (forvar1273 < (2'h2)); forvar1273 = (forvar1273 + (1'h1)))
                    begin
                      reg1274 <= (&reg1216);
                      reg1275 <= $signed(forvar1246[(3'h5):(1'h1)]);
                    end
                  for (forvar1276 = (1'h0); (forvar1276 < (2'h2)); forvar1276 = (forvar1276 + (1'h1)))
                    begin
                      reg1277 <= reg1235[(1'h0):(1'h0)];
                      reg1278 <= $signed($unsigned((&forvar1220[(2'h2):(1'h0)])));
                      reg1279 <= $unsigned($unsigned(wire1208[(4'hc):(3'h5)]));
                      reg1280 <= $signed(forvar1258[(2'h3):(2'h2)]);
                    end
                  if (reg1197[(3'h4):(1'h0)])
                    begin
                      reg1281 <= (reg1252 ?
                          $signed((~(-reg1189))) : (reg1193[(1'h0):(1'h0)] ?
                              reg1215[(1'h1):(1'h1)] : $signed(reg1192)));
                      reg1282 <= {{((8'h9d) <= $signed(reg1241))}};
                      reg1283 <= {(~|{{wire1208}})};
                      reg1284 <= {$unsigned((forvar1180 ?
                              (reg1228 ? forvar1267 : (8'haf)) : ((8'ha0) ?
                                  forvar1254 : forvar1181)))};
                    end
                  else
                    begin
                      reg1281 <= forvar1195[(1'h1):(1'h0)];
                    end
                  for (forvar1285 = (1'h0); (forvar1285 < (2'h3)); forvar1285 = (forvar1285 + (1'h1)))
                    begin
                      reg1286 <= $signed(forvar1220[(4'h8):(3'h4)]);
                      reg1287 <= $unsigned((-$signed($signed((8'hba)))));
                      reg1288 <= $signed(forvar1225[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  reg1273 <= $signed($signed($signed((~|reg1256))));
                  for (forvar1274 = (1'h0); (forvar1274 < (2'h2)); forvar1274 = (forvar1274 + (1'h1)))
                    begin
                      reg1275 <= (!{$unsigned($signed(reg1181))});
                    end
                end
              for (forvar1289 = (1'h0); (forvar1289 < (2'h2)); forvar1289 = (forvar1289 + (1'h1)))
                begin
                  reg1290 <= $signed((8'hb5));
                  if ((($signed($unsigned(wire1179)) ?
                      reg1263 : $signed(((8'ha7) | reg1248))) - $signed({$signed(reg1192)})))
                    begin
                      reg1291 <= forvar1185[(1'h0):(1'h0)];
                      reg1292 <= $signed({(-{reg1247})});
                      reg1293 <= $unsigned($signed($signed(reg1193[(1'h1):(1'h1)])));
                      reg1294 <= reg1264[(4'h9):(3'h6)];
                    end
                  else
                    begin
                      reg1291 <= $unsigned($signed($signed((8'haf))));
                    end
                  if ($signed(forvar1185))
                    begin
                      reg1295 <= {(-($unsigned(reg1232) ?
                              forvar1230[(3'h6):(3'h6)] : (!reg1226)))};
                      reg1296 <= (8'ha4);
                      reg1297 <= (reg1266[(3'h6):(2'h2)] ?
                          {(~((8'hb7) ^~ (8'hb3)))} : reg1198);
                    end
                  else
                    begin
                      reg1295 <= $unsigned({((reg1267 - reg1292) * (8'hb5))});
                      reg1296 <= forvar1214[(1'h0):(1'h0)];
                      reg1297 <= (($signed(forvar1193) ^~ $signed((wire1178 ?
                              reg1296 : forvar1289))) ?
                          (reg1254[(1'h0):(1'h0)] ?
                              $unsigned((forvar1182 < forvar1181)) : (~reg1275)) : (^~(~|(forvar1262 ?
                              reg1295 : reg1280))));
                    end
                end
              for (forvar1298 = (1'h0); (forvar1298 < (2'h3)); forvar1298 = (forvar1298 + (1'h1)))
                begin
                  if (reg1269[(2'h3):(2'h2)])
                    begin
                      reg1299 <= ($unsigned((~|(8'ha9))) ?
                          forvar1266[(2'h2):(1'h0)] : forvar1272);
                      reg1300 <= (-(!wire1177[(4'h8):(3'h4)]));
                    end
                  else
                    begin
                      reg1299 <= $unsigned((8'ha2));
                    end
                  for (forvar1301 = (1'h0); (forvar1301 < (1'h0)); forvar1301 = (forvar1301 + (1'h1)))
                    begin
                      reg1302 <= ($signed(wire1174) ^ ((forvar1272 ?
                              reg1224[(1'h1):(1'h0)] : (&(8'h9d))) ?
                          (8'hac) : reg1233[(3'h6):(3'h5)]));
                      reg1303 <= ($unsigned($unsigned($unsigned(reg1288))) && $signed(($signed(reg1183) + $unsigned(reg1241))));
                    end
                  for (forvar1304 = (1'h0); (forvar1304 < (2'h3)); forvar1304 = (forvar1304 + (1'h1)))
                    begin
                      reg1305 <= (((reg1277[(1'h1):(1'h0)] ?
                          $signed(reg1302) : (~(8'hb9))) >= forvar1230) | (($unsigned(reg1226) >>> $signed(forvar1220)) >= reg1238[(2'h3):(1'h1)]));
                      reg1306 <= reg1206;
                      reg1307 <= $signed($signed($signed({reg1277})));
                      reg1308 <= (+$signed(reg1238));
                    end
                end
              for (forvar1309 = (1'h0); (forvar1309 < (2'h3)); forvar1309 = (forvar1309 + (1'h1)))
                begin
                  if ({($signed($signed(reg1243)) ?
                          reg1228 : $signed(forvar1195[(1'h0):(1'h0)]))})
                    begin
                      reg1310 <= (8'ha5);
                      reg1311 <= (~|$unsigned($unsigned(wire1179[(3'h4):(1'h0)])));
                      reg1312 <= $unsigned(forvar1225);
                    end
                  else
                    begin
                      reg1310 <= reg1261[(3'h5):(1'h1)];
                      reg1311 <= forvar1193[(1'h0):(1'h0)];
                      reg1312 <= ($unsigned(($unsigned(reg1310) >> (reg1305 ^~ reg1256))) & ({$signed((8'hb2))} >= (&(^forvar1262))));
                    end
                end
            end
          reg1313 <= (((|$unsigned(reg1273)) ?
                  $signed(reg1254[(1'h1):(1'h0)]) : $unsigned($signed(reg1214))) ?
              (wire1210[(1'h0):(1'h0)] > $signed(((8'ha5) ^~ wire1179))) : (^~($signed(forvar1234) >> ((8'ha5) ^~ reg1227))));
        end
      reg1314 <= forvar1224[(2'h2):(1'h0)];
      reg1315 <= (+((~|(reg1243 >> forvar1190)) ?
          forvar1185 : $signed($signed(reg1243))));
    end
  assign wire1316 = {(((~&reg1213) <= reg1181) | $signed(forvar1269))};
  assign wire1317 = {(reg1252 ? $signed(forvar1274) : reg1191[(3'h4):(2'h3)])};
  assign wire1318 = forvar1215;
  always
    @(posedge clk) begin
      if ($signed(($signed((reg1299 ? forvar1194 : reg1188)) ?
          reg1193[(1'h0):(1'h0)] : $signed($signed(wire1175)))))
        begin
          for (forvar1319 = (1'h0); (forvar1319 < (2'h2)); forvar1319 = (forvar1319 + (1'h1)))
            begin
              if ((reg1281[(1'h0):(1'h0)] != {$signed(forvar1223[(1'h0):(1'h0)])}))
                begin
                  if (($unsigned(($unsigned(wire1208) << $unsigned(reg1216))) <<< reg1296))
                    begin
                      reg1320 <= (wire1178[(1'h0):(1'h0)] ?
                          (({reg1268} > (~|reg1236)) >> $unsigned((~&forvar1309))) : reg1278[(3'h4):(1'h0)]);
                      reg1321 <= {forvar1195[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg1320 <= $signed((-forvar1267[(1'h0):(1'h0)]));
                      reg1321 <= ($unsigned($unsigned(reg1275)) + (-reg1310[(3'h5):(1'h0)]));
                      reg1322 <= (reg1308[(4'hb):(1'h0)] ?
                          (reg1216[(1'h0):(1'h0)] ?
                              (-(forvar1190 ^ wire1210)) : ($unsigned(forvar1220) >>> (+wire1210))) : reg1186[(4'hc):(2'h2)]);
                      reg1323 <= (8'h9e);
                    end
                  reg1324 <= $unsigned((forvar1254 ?
                      (forvar1309 ?
                          $signed(reg1193) : $unsigned(reg1287)) : (reg1185[(1'h1):(1'h1)] && {(8'ha9)})));
                  reg1325 <= {(reg1251[(2'h2):(1'h1)] <= $unsigned(reg1181[(1'h0):(1'h0)]))};
                end
              else
                begin
                  if ($signed((&$signed($unsigned((8'h9e))))))
                    begin
                      reg1320 <= (~(reg1250[(1'h1):(1'h0)] != reg1244[(1'h0):(1'h0)]));
                      reg1321 <= (-{(-(forvar1309 ? reg1255 : (8'had)))});
                    end
                  else
                    begin
                      reg1320 <= reg1256;
                    end
                  reg1322 <= forvar1241;
                  for (forvar1323 = (1'h0); (forvar1323 < (2'h2)); forvar1323 = (forvar1323 + (1'h1)))
                    begin
                      reg1324 <= $signed((($unsigned((8'hba)) ?
                              (8'h9e) : wire1176[(3'h4):(3'h4)]) ?
                          (~(reg1275 ?
                              forvar1274 : reg1255)) : $unsigned((forvar1230 ?
                              (8'ha4) : forvar1189))));
                      reg1325 <= (&reg1187);
                      reg1326 <= (reg1190[(2'h3):(2'h2)] > ((~(wire1318 ?
                              forvar1266 : reg1313)) ?
                          reg1228 : reg1293[(4'h9):(3'h6)]));
                      reg1327 <= $signed($unsigned({(~|reg1247)}));
                    end
                end
              for (forvar1328 = (1'h0); (forvar1328 < (2'h2)); forvar1328 = (forvar1328 + (1'h1)))
                begin
                  if ((wire1177 ?
                      (~&$signed((|reg1203))) : reg1196[(2'h3):(2'h3)]))
                    begin
                      reg1329 <= forvar1253[(2'h3):(1'h1)];
                      reg1330 <= reg1329[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1329 <= wire1317;
                    end
                  if ((+$signed($unsigned((wire1317 ^ forvar1194)))))
                    begin
                      reg1331 <= {$unsigned((wire1176[(1'h1):(1'h1)] << $unsigned(reg1256)))};
                      reg1332 <= ((^~reg1300) ?
                          ($signed((reg1252 ? reg1295 : reg1232)) ?
                              forvar1183 : {(forvar1197 ?
                                      forvar1215 : (8'ha6))}) : (reg1269[(2'h2):(1'h1)] ?
                              (wire1209 * (~^reg1215)) : forvar1183[(3'h5):(1'h1)]));
                      reg1333 <= ((~((~^reg1274) ?
                          (~|reg1226) : forvar1180[(2'h2):(1'h0)])) > (reg1192 ?
                          {(reg1246 | reg1310)} : (reg1294 ?
                              $unsigned((8'hae)) : (&forvar1249))));
                    end
                  else
                    begin
                      reg1331 <= (((forvar1258[(1'h1):(1'h0)] ?
                                  reg1275 : {(8'hb5)}) ?
                              $unsigned((!reg1323)) : {(~&reg1299)}) ?
                          (forvar1214[(3'h5):(3'h4)] != {$unsigned(reg1222)}) : ((reg1266 >>> $signed(reg1238)) << ((&reg1224) ?
                              forvar1197 : $signed(reg1215))));
                    end
                  for (forvar1334 = (1'h0); (forvar1334 < (2'h3)); forvar1334 = (forvar1334 + (1'h1)))
                    begin
                      reg1335 <= $signed(($signed((reg1225 | forvar1190)) ?
                          $signed(reg1264[(4'h9):(1'h0)]) : (+$unsigned(reg1225))));
                      reg1336 <= forvar1274[(3'h5):(1'h0)];
                      reg1337 <= $signed(reg1294);
                      reg1338 <= (($unsigned($unsigned(forvar1220)) ?
                              (^forvar1200[(1'h0):(1'h0)]) : {$unsigned(reg1248)}) ?
                          $signed($unsigned(reg1192)) : ($unsigned((wire1316 & forvar1198)) ?
                              (~&(8'h9e)) : {(forvar1197 ?
                                      reg1324 : reg1197)}));
                    end
                  if (reg1259[(1'h0):(1'h0)])
                    begin
                      reg1339 <= $signed((~|$signed((reg1241 ?
                          reg1267 : (8'h9f)))));
                    end
                  else
                    begin
                      reg1339 <= (wire1317[(2'h2):(1'h0)] ?
                          {({forvar1262} ?
                                  (forvar1273 ?
                                      (8'hb7) : reg1311) : (-forvar1230))} : (!({reg1238} ?
                              reg1247[(3'h5):(2'h2)] : reg1227)));
                      reg1340 <= $unsigned(($unsigned((reg1222 ?
                          reg1181 : reg1252)) | (~^{reg1237})));
                    end
                end
            end
          if ((+$unsigned(wire1316[(4'hd):(3'h5)])))
            begin
              for (forvar1341 = (1'h0); (forvar1341 < (1'h0)); forvar1341 = (forvar1341 + (1'h1)))
                begin
                  if ($unsigned((((reg1326 ?
                          (8'ha0) : reg1236) << reg1196[(4'h8):(3'h7)]) ?
                      ($signed(reg1271) - reg1332) : reg1199[(4'h8):(3'h6)])))
                    begin
                      reg1342 <= (forvar1276[(3'h5):(1'h1)] ^~ reg1239);
                      reg1343 <= (~($signed($unsigned(reg1198)) + (|(&(8'ha3)))));
                    end
                  else
                    begin
                      reg1342 <= reg1258[(1'h1):(1'h1)];
                      reg1343 <= $unsigned(((8'hab) < (wire1178 >= $unsigned(reg1271))));
                    end
                  for (forvar1344 = (1'h0); (forvar1344 < (2'h3)); forvar1344 = (forvar1344 + (1'h1)))
                    begin
                      reg1345 <= $unsigned(wire1316[(3'h6):(3'h5)]);
                      reg1346 <= ($signed(($unsigned(reg1332) ?
                          (+wire1179) : forvar1344[(3'h7):(3'h6)])) && ($signed(reg1315) & (8'haa)));
                    end
                end
              if (reg1286[(2'h2):(1'h0)])
                begin
                  for (forvar1347 = (1'h0); (forvar1347 < (1'h0)); forvar1347 = (forvar1347 + (1'h1)))
                    begin
                      reg1348 <= {(reg1198 >> $unsigned(reg1192))};
                      reg1349 <= (reg1182[(2'h2):(1'h1)] ?
                          ({$signed(forvar1298)} ?
                              reg1197 : $unsigned(forvar1323[(3'h5):(2'h3)])) : forvar1189);
                      reg1350 <= ({(((8'hae) >= (8'h9d)) || {reg1252})} ?
                          ($signed($signed(reg1307)) & reg1256) : $unsigned($unsigned(forvar1246[(4'hc):(4'hb)])));
                    end
                  reg1351 <= (~|$unsigned(reg1197[(3'h5):(3'h5)]));
                  reg1352 <= $unsigned((|($signed(reg1311) ^ {reg1300})));
                  if (reg1287)
                    begin
                      reg1353 <= (^~((wire1175 <= (-reg1238)) ?
                          (~&(forvar1240 + wire1176)) : $unsigned((reg1191 - reg1291))));
                      reg1354 <= (|reg1337);
                      reg1355 <= forvar1194[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg1353 <= reg1215[(3'h6):(1'h1)];
                    end
                end
              else
                begin
                  if (reg1346)
                    begin
                      reg1347 <= reg1198[(1'h0):(1'h0)];
                      reg1348 <= $signed((forvar1262 ?
                          ((~^reg1268) ~^ reg1308) : (^~(reg1259 ?
                              reg1247 : reg1258))));
                    end
                  else
                    begin
                      reg1347 <= wire1207;
                      reg1348 <= (8'ha6);
                      reg1349 <= reg1192[(2'h2):(1'h1)];
                    end
                  for (forvar1350 = (1'h0); (forvar1350 < (2'h2)); forvar1350 = (forvar1350 + (1'h1)))
                    begin
                      reg1351 <= $signed(($signed($unsigned(forvar1272)) && $signed((reg1259 & reg1348))));
                    end
                  for (forvar1352 = (1'h0); (forvar1352 < (1'h1)); forvar1352 = (forvar1352 + (1'h1)))
                    begin
                      reg1353 <= $unsigned((((reg1299 ?
                              reg1231 : reg1215) >= (reg1325 ?
                              reg1290 : reg1192)) ?
                          (!reg1235[(2'h3):(2'h2)]) : $unsigned((-(8'hba)))));
                      reg1354 <= ($signed(($unsigned((8'ha3)) ?
                              {reg1332} : $unsigned(reg1244))) ?
                          $signed({$signed((8'haa))}) : wire1209);
                      reg1355 <= $unsigned((~reg1275[(4'h8):(1'h0)]));
                    end
                  for (forvar1356 = (1'h0); (forvar1356 < (1'h1)); forvar1356 = (forvar1356 + (1'h1)))
                    begin
                      reg1357 <= reg1291[(4'ha):(1'h0)];
                      reg1358 <= reg1292[(4'ha):(4'h8)];
                    end
                end
            end
          else
            begin
              for (forvar1341 = (1'h0); (forvar1341 < (1'h1)); forvar1341 = (forvar1341 + (1'h1)))
                begin
                  if (reg1254)
                    begin
                      reg1342 <= (forvar1195 ^ (((+(8'hb6)) <<< $unsigned(reg1273)) * {reg1305}));
                      reg1343 <= $unsigned((reg1261[(4'h9):(1'h1)] && ($unsigned((8'h9c)) * $signed(forvar1265))));
                      reg1344 <= (8'hb5);
                    end
                  else
                    begin
                      reg1342 <= $signed((~&$signed({reg1196})));
                    end
                  for (forvar1345 = (1'h0); (forvar1345 < (1'h0)); forvar1345 = (forvar1345 + (1'h1)))
                    begin
                      reg1346 <= (+$unsigned(((reg1279 ?
                          reg1235 : forvar1200) + (reg1221 ^~ reg1191))));
                    end
                end
              reg1347 <= (&(|forvar1347[(1'h0):(1'h0)]));
            end
        end
      else
        begin
          if (($signed(((^~reg1290) ?
                  (reg1274 ? reg1218 : reg1190) : {reg1241})) ?
              reg1185 : ((|{reg1216}) >>> (forvar1220[(3'h4):(3'h4)] ?
                  forvar1229 : (forvar1301 ? forvar1197 : reg1195)))))
            begin
              if ($unsigned(reg1248))
                begin
                  if (reg1296)
                    begin
                      reg1319 <= (reg1243 >> ({$unsigned(reg1321)} > reg1308));
                      reg1320 <= (8'h9d);
                      reg1321 <= {reg1205[(1'h1):(1'h0)]};
                    end
                  else
                    begin
                      reg1319 <= ($signed(forvar1269) ?
                          reg1263[(1'h0):(1'h0)] : ($unsigned(((8'ha3) & reg1357)) ?
                              (forvar1350 != (~&reg1319)) : (^~forvar1258[(3'h5):(3'h4)])));
                      reg1320 <= {reg1345[(4'h8):(2'h2)]};
                      reg1321 <= forvar1352[(2'h3):(2'h2)];
                    end
                  for (forvar1322 = (1'h0); (forvar1322 < (2'h2)); forvar1322 = (forvar1322 + (1'h1)))
                    begin
                      reg1323 <= $unsigned((~^((reg1235 - (8'h9c)) - (reg1338 ?
                          (8'hba) : reg1307))));
                      reg1324 <= (reg1293 != $signed(($signed(reg1197) ?
                          reg1308[(4'he):(3'h4)] : (|reg1192))));
                    end
                  reg1325 <= $unsigned(reg1282[(1'h1):(1'h1)]);
                  for (forvar1326 = (1'h0); (forvar1326 < (1'h1)); forvar1326 = (forvar1326 + (1'h1)))
                    begin
                      reg1327 <= ((reg1181[(4'hc):(1'h0)] ?
                          forvar1266 : $signed((~(8'ha5)))) & {{$unsigned(reg1354)}});
                      reg1328 <= $signed($unsigned(reg1183[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  reg1319 <= (forvar1269[(4'ha):(1'h0)] ?
                      $unsigned($signed(reg1345[(3'h6):(2'h3)])) : reg1274);
                  if (($signed(((reg1297 | forvar1322) ?
                      (reg1230 != (8'had)) : $signed(reg1206))) && $signed((forvar1196[(1'h1):(1'h1)] ?
                      $signed(forvar1344) : $unsigned(forvar1253)))))
                    begin
                      reg1320 <= {reg1182};
                    end
                  else
                    begin
                      reg1320 <= $signed($unsigned(reg1269[(3'h7):(1'h0)]));
                    end
                  if ((reg1342 ^ ($unsigned({forvar1328}) ?
                      $unsigned({reg1339}) : ($signed(forvar1190) ?
                          (reg1268 <= reg1214) : $unsigned(reg1319)))))
                    begin
                      reg1321 <= ((8'had) ?
                          $unsigned($unsigned((^reg1196))) : {reg1241});
                    end
                  else
                    begin
                      reg1321 <= (((~$signed(reg1315)) >> reg1192) ?
                          wire1317[(3'h4):(2'h3)] : reg1335);
                      reg1322 <= (~|($unsigned(forvar1225[(4'h8):(1'h0)]) - (~&{forvar1301})));
                      reg1323 <= {$signed(({reg1205} ?
                              $unsigned((8'haa)) : $signed(reg1296)))};
                      reg1324 <= (~^($signed((^~forvar1240)) ^~ (!(reg1295 - reg1211))));
                    end
                  if (reg1191)
                    begin
                      reg1325 <= $signed(({forvar1212[(1'h1):(1'h1)]} >= ((wire1174 ?
                          (8'hb7) : reg1274) * reg1275)));
                      reg1326 <= (8'ha2);
                      reg1327 <= (|reg1205);
                      reg1328 <= $unsigned((|($signed(forvar1212) ?
                          (^~reg1254) : reg1283)));
                    end
                  else
                    begin
                      reg1325 <= {(8'hb6)};
                    end
                end
              if ($signed($unsigned((reg1290 <= (wire1318 >> reg1358)))))
                begin
                  for (forvar1329 = (1'h0); (forvar1329 < (2'h2)); forvar1329 = (forvar1329 + (1'h1)))
                    begin
                      reg1330 <= $signed(({(reg1263 ? reg1225 : (8'h9d))} ?
                          {reg1185} : (+(reg1221 ^ forvar1185))));
                      reg1331 <= {reg1269};
                    end
                end
              else
                begin
                  for (forvar1329 = (1'h0); (forvar1329 < (2'h3)); forvar1329 = (forvar1329 + (1'h1)))
                    begin
                      reg1330 <= $signed($unsigned((reg1270[(3'h4):(1'h0)] ?
                          ((8'ha6) ? reg1204 : reg1342) : $unsigned(reg1231))));
                      reg1331 <= {($signed($unsigned(forvar1350)) ?
                              $unsigned($signed(reg1232)) : reg1284)};
                      reg1332 <= {wire1179};
                    end
                  if ({(-($unsigned(reg1228) != $signed(reg1275)))})
                    begin
                      reg1333 <= $signed($signed((&((8'h9e) ?
                          reg1268 : reg1280))));
                      reg1334 <= reg1217[(1'h0):(1'h0)];
                      reg1335 <= reg1238[(3'h6):(2'h3)];
                      reg1336 <= forvar1240;
                    end
                  else
                    begin
                      reg1333 <= $signed((+(-reg1254[(2'h2):(2'h2)])));
                      reg1334 <= forvar1225;
                      reg1335 <= {reg1195[(4'hd):(1'h0)]};
                    end
                end
            end
          else
            begin
              for (forvar1319 = (1'h0); (forvar1319 < (1'h1)); forvar1319 = (forvar1319 + (1'h1)))
                begin
                  for (forvar1320 = (1'h0); (forvar1320 < (2'h2)); forvar1320 = (forvar1320 + (1'h1)))
                    begin
                      reg1321 <= ((~|forvar1202[(1'h1):(1'h0)]) ?
                          $signed(reg1288) : (((forvar1266 ?
                              reg1251 : (8'ha5)) ^~ (~&reg1196)) > (reg1203[(4'h9):(1'h1)] == (reg1351 ?
                              reg1299 : reg1287))));
                      reg1322 <= $unsigned(((^~(8'hb7)) ?
                          ((reg1221 ?
                              forvar1212 : reg1189) != ((8'hb1) >= (8'ha2))) : {reg1237}));
                      reg1323 <= forvar1193[(1'h1):(1'h0)];
                    end
                end
            end
          for (forvar1337 = (1'h0); (forvar1337 < (2'h3)); forvar1337 = (forvar1337 + (1'h1)))
            begin
              if (((&(&{reg1188})) ? {$unsigned((8'ha6))} : (8'hb0)))
                begin
                  if (reg1273)
                    begin
                      reg1338 <= $unsigned($unsigned(reg1232[(2'h2):(1'h0)]));
                      reg1339 <= (($signed((-reg1247)) ?
                              $unsigned(((8'ha2) ?
                                  (8'hb2) : (8'h9c))) : $signed((forvar1326 ?
                                  forvar1272 : reg1247))) ?
                          forvar1269[(4'hb):(4'hb)] : ({reg1252[(3'h4):(2'h3)]} ?
                              $unsigned({forvar1197}) : $signed((forvar1328 >>> forvar1214))));
                      reg1340 <= forvar1344;
                    end
                  else
                    begin
                      reg1338 <= reg1330[(2'h3):(1'h0)];
                      reg1339 <= (+$unsigned(reg1236[(2'h3):(1'h1)]));
                    end
                  reg1341 <= (&reg1330);
                  reg1342 <= wire1318[(2'h2):(1'h0)];
                  for (forvar1343 = (1'h0); (forvar1343 < (2'h3)); forvar1343 = (forvar1343 + (1'h1)))
                    begin
                      reg1344 <= (!(forvar1272[(2'h3):(1'h0)] ?
                          reg1218[(3'h7):(1'h1)] : $signed(reg1192)));
                    end
                end
              else
                begin
                  for (forvar1338 = (1'h0); (forvar1338 < (1'h0)); forvar1338 = (forvar1338 + (1'h1)))
                    begin
                      reg1339 <= ((((forvar1323 == forvar1224) ?
                          forvar1323 : reg1242) ^ ((+wire1209) >= reg1310)) - (~^reg1252));
                      reg1340 <= reg1293;
                      reg1341 <= $signed(forvar1345);
                      reg1342 <= (+$signed((((8'hb0) << forvar1276) < (forvar1254 ?
                          reg1303 : reg1183))));
                    end
                  if (forvar1190[(3'h7):(2'h3)])
                    begin
                      reg1343 <= $unsigned((forvar1285[(1'h1):(1'h1)] ^ $signed((reg1196 + forvar1240))));
                      reg1344 <= ($signed(((~^reg1248) >= (reg1348 ^ reg1229))) ?
                          reg1218[(3'h7):(2'h2)] : forvar1272[(4'ha):(3'h6)]);
                      reg1345 <= forvar1269[(3'h5):(2'h2)];
                      reg1346 <= {(reg1265 + $unsigned($signed(wire1317)))};
                    end
                  else
                    begin
                      reg1343 <= reg1205[(1'h0):(1'h0)];
                      reg1344 <= reg1246[(3'h4):(1'h1)];
                      reg1345 <= forvar1273;
                    end
                  reg1347 <= {reg1182};
                  for (forvar1348 = (1'h0); (forvar1348 < (2'h3)); forvar1348 = (forvar1348 + (1'h1)))
                    begin
                      reg1349 <= reg1259[(3'h6):(3'h6)];
                      reg1350 <= (^~$signed((~^{reg1200})));
                      reg1351 <= ($signed((~|(&reg1183))) + (+(~|(reg1245 ?
                          forvar1334 : forvar1188))));
                      reg1352 <= (~&forvar1344[(3'h5):(3'h5)]);
                    end
                end
              reg1353 <= (8'h9c);
            end
          if (reg1336[(1'h0):(1'h0)])
            begin
              for (forvar1354 = (1'h0); (forvar1354 < (1'h1)); forvar1354 = (forvar1354 + (1'h1)))
                begin
                  if ((!(~^(~(-reg1313)))))
                    begin
                      reg1355 <= reg1348[(3'h4):(1'h0)];
                      reg1356 <= $unsigned($unsigned(reg1299[(3'h4):(2'h2)]));
                      reg1357 <= ($signed((8'hac)) ?
                          (+$signed(forvar1189)) : (+$signed((^~reg1320))));
                    end
                  else
                    begin
                      reg1355 <= ((&reg1268[(2'h2):(1'h1)]) ?
                          (~&(reg1280[(3'h4):(3'h4)] ?
                              (reg1186 ^ reg1200) : forvar1304[(1'h1):(1'h1)])) : ($signed((8'ha0)) ?
                              $unsigned(reg1200) : reg1231[(2'h2):(2'h2)]));
                    end
                  for (forvar1358 = (1'h0); (forvar1358 < (2'h3)); forvar1358 = (forvar1358 + (1'h1)))
                    begin
                      reg1359 <= ($unsigned((^(&reg1218))) >>> reg1187);
                    end
                  if ($signed((|$unsigned((~&forvar1203)))))
                    begin
                      reg1360 <= $signed((|(~&$unsigned(forvar1350))));
                      reg1361 <= $signed((forvar1195[(2'h2):(2'h2)] >>> reg1244[(2'h3):(1'h1)]));
                      reg1362 <= ((8'hae) < {forvar1193});
                      reg1363 <= ($signed(forvar1229[(3'h7):(2'h3)]) * ({$unsigned(forvar1215)} ?
                          ($signed(reg1196) <<< $unsigned(reg1193)) : $unsigned(forvar1230)));
                    end
                  else
                    begin
                      reg1360 <= (~|$unsigned(reg1347));
                      reg1361 <= reg1251[(4'h9):(2'h2)];
                    end
                end
              if ($unsigned(reg1233))
                begin
                  for (forvar1364 = (1'h0); (forvar1364 < (2'h2)); forvar1364 = (forvar1364 + (1'h1)))
                    begin
                      reg1365 <= ((&reg1267[(3'h6):(3'h6)]) ?
                          (reg1255 ?
                              $signed((|reg1359)) : reg1293[(2'h3):(2'h2)]) : ((!(~forvar1185)) && reg1357));
                      reg1366 <= $signed(((-$signed(reg1235)) ^ $signed(reg1225[(1'h1):(1'h0)])));
                    end
                  if ({$signed($signed(reg1344))})
                    begin
                      reg1367 <= reg1295;
                      reg1368 <= $unsigned($unsigned($unsigned((forvar1347 <<< forvar1265))));
                      reg1369 <= reg1259[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1367 <= forvar1364[(5'h10):(4'h9)];
                    end
                  for (forvar1370 = (1'h0); (forvar1370 < (1'h0)); forvar1370 = (forvar1370 + (1'h1)))
                    begin
                      reg1371 <= reg1187;
                    end
                end
              else
                begin
                  reg1364 <= (^(reg1303 >= reg1266[(4'ha):(2'h2)]));
                  reg1365 <= ($unsigned(reg1197[(2'h2):(2'h2)]) ?
                      $signed($signed($signed(forvar1301))) : reg1323[(2'h3):(2'h3)]);
                  for (forvar1366 = (1'h0); (forvar1366 < (2'h3)); forvar1366 = (forvar1366 + (1'h1)))
                    begin
                      reg1367 <= ((|($signed(forvar1366) ?
                          $signed(forvar1266) : reg1238[(2'h2):(2'h2)])) <<< {$unsigned({reg1242})});
                      reg1368 <= $unsigned(($unsigned({reg1229}) ?
                          ((~^reg1311) ?
                              $unsigned(reg1314) : $signed((8'ha1))) : wire1174));
                      reg1369 <= $unsigned(forvar1343[(4'he):(3'h7)]);
                    end
                end
              for (forvar1372 = (1'h0); (forvar1372 < (2'h3)); forvar1372 = (forvar1372 + (1'h1)))
                begin
                  reg1373 <= ((|{reg1270[(4'ha):(4'h8)]}) <<< reg1270);
                end
            end
          else
            begin
              for (forvar1354 = (1'h0); (forvar1354 < (1'h1)); forvar1354 = (forvar1354 + (1'h1)))
                begin
                  if ((|(~|($signed((8'ha6)) && (reg1187 - reg1181)))))
                    begin
                      reg1355 <= reg1362;
                      reg1356 <= {$unsigned($signed(((8'hb1) - (8'hb3))))};
                      reg1357 <= reg1264[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg1355 <= (reg1323[(3'h4):(3'h4)] ^ $unsigned((((8'ha5) ?
                              (8'hb2) : (8'ha9)) ?
                          (forvar1322 ~^ (8'hba)) : (forvar1200 | reg1250))));
                      reg1356 <= $unsigned((~((reg1325 ? forvar1337 : (8'hb2)) ?
                          reg1271 : forvar1344)));
                      reg1357 <= reg1315[(2'h3):(1'h1)];
                      reg1358 <= (forvar1182 || ({forvar1274[(4'hb):(1'h1)]} ?
                          ((reg1291 ? forvar1323 : reg1283) | (reg1237 ?
                              reg1369 : forvar1245)) : $unsigned(forvar1341)));
                    end
                  for (forvar1359 = (1'h0); (forvar1359 < (2'h2)); forvar1359 = (forvar1359 + (1'h1)))
                    begin
                      reg1360 <= {reg1199[(3'h6):(1'h0)]};
                      reg1361 <= $unsigned(forvar1364);
                      reg1362 <= forvar1348;
                    end
                  reg1363 <= ((8'ha1) ?
                      $unsigned($signed(reg1220[(4'h9):(1'h0)])) : reg1190[(2'h2):(1'h0)]);
                  for (forvar1364 = (1'h0); (forvar1364 < (1'h0)); forvar1364 = (forvar1364 + (1'h1)))
                    begin
                      reg1365 <= ($unsigned($signed($signed((8'hb0)))) ?
                          $unsigned($signed($unsigned(reg1254))) : (reg1211 - (^$signed(wire1210))));
                      reg1366 <= ((8'hba) <<< (~^((~^reg1243) * $signed(forvar1245))));
                      reg1367 <= (((reg1223[(1'h0):(1'h0)] == ((8'ha3) ^ (8'hac))) >= {(&reg1211)}) * ($signed((~^reg1293)) ?
                          $unsigned(forvar1354[(2'h2):(1'h0)]) : (reg1283 ?
                              (reg1288 * forvar1319) : ((8'hb7) ?
                                  reg1247 : (8'h9f)))));
                    end
                end
            end
          reg1374 <= $signed(reg1184[(1'h1):(1'h1)]);
        end
      reg1375 <= reg1345;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1803
#( parameter param2154 = ((({(8'h9e)} + ((8'ha0) >= (8'ha5))) * (&(~^(8'h9e)))) ? ({{(8'hac)}} ? (((8'hb4) ^~ (8'had)) && ((8'hae) + (8'haa))) : ((!(8'haa)) | (+(8'h9f)))) : ({((8'ha0) <<< (8'ha0))} >> (((8'hb8) ? (8'ha7) : (8'hb2)) || ((8'ha8) ~^ (8'h9e))))) )
(y, clk, wire1808, wire1807, wire1806, wire1805, wire1804);
  output wire [(32'he06):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire1808;
  input wire signed [(5'h10):(1'h0)] wire1807;
  input wire [(3'h6):(1'h0)] wire1806;
  input wire signed [(4'h8):(1'h0)] wire1805;
  input wire signed [(3'h7):(1'h0)] wire1804;
  reg signed [(4'h8):(1'h0)] reg2153 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2134 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2133 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2132 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2129 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2128 = (1'h0);
  reg [(4'hc):(1'h0)] reg2127 = (1'h0);
  reg [(4'h8):(1'h0)] reg2124 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2118 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2116 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2111 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2114 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2113 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2109 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2108 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2106 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2152 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2151 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2150 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2149 = (1'h0);
  reg [(5'h10):(1'h0)] reg2148 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2147 = (1'h0);
  reg [(2'h3):(1'h0)] reg2146 = (1'h0);
  reg [(4'h9):(1'h0)] reg2145 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2144 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2143 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2142 = (1'h0);
  reg [(4'ha):(1'h0)] reg2141 = (1'h0);
  reg [(4'h8):(1'h0)] reg2139 = (1'h0);
  reg [(2'h2):(1'h0)] reg2140 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2139 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2138 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2137 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2136 = (1'h0);
  reg [(4'he):(1'h0)] reg2135 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2134 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2133 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2132 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2131 = (1'h0);
  reg [(2'h3):(1'h0)] reg2130 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2129 = (1'h0);
  reg [(4'he):(1'h0)] reg2128 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2127 = (1'h0);
  reg [(3'h4):(1'h0)] reg2126 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2125 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2124 = (1'h0);
  reg [(5'h10):(1'h0)] reg2123 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2122 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2121 = (1'h0);
  reg [(3'h5):(1'h0)] reg2120 = (1'h0);
  reg [(3'h7):(1'h0)] reg2119 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2118 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2117 = (1'h0);
  reg [(2'h2):(1'h0)] reg2116 = (1'h0);
  reg [(3'h4):(1'h0)] reg2115 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2114 = (1'h0);
  reg [(4'he):(1'h0)] reg2113 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2112 = (1'h0);
  reg [(3'h4):(1'h0)] reg2111 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2110 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2109 = (1'h0);
  reg [(4'h8):(1'h0)] reg2108 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2107 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2106 = (1'h0);
  reg [(4'he):(1'h0)] reg2093 = (1'h0);
  reg [(3'h6):(1'h0)] reg2105 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2104 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2103 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2102 = (1'h0);
  reg [(4'hb):(1'h0)] reg2101 = (1'h0);
  reg [(3'h6):(1'h0)] reg2100 = (1'h0);
  reg [(4'ha):(1'h0)] reg2099 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2098 = (1'h0);
  reg [(4'hd):(1'h0)] reg2097 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2096 = (1'h0);
  reg [(4'hd):(1'h0)] reg2095 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2094 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2093 = (1'h0);
  reg [(2'h3):(1'h0)] reg2092 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2091 = (1'h0);
  reg [(4'hc):(1'h0)] reg2090 = (1'h0);
  reg [(2'h3):(1'h0)] reg2089 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2088 = (1'h0);
  reg [(3'h7):(1'h0)] reg2087 = (1'h0);
  reg [(4'ha):(1'h0)] reg2086 = (1'h0);
  reg [(4'h8):(1'h0)] reg2085 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2084 = (1'h0);
  reg [(3'h7):(1'h0)] reg2083 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2082 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2081 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2080 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2079 = (1'h0);
  reg [(4'h8):(1'h0)] reg2078 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2077 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2076 = (1'h0);
  reg [(4'h8):(1'h0)] reg2075 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2074 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2073 = (1'h0);
  reg [(4'he):(1'h0)] forvar2070 = (1'h0);
  reg [(4'h8):(1'h0)] reg2069 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2073 = (1'h0);
  reg [(3'h7):(1'h0)] reg2072 = (1'h0);
  reg [(4'hd):(1'h0)] reg2071 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2070 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2069 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2068 = (1'h0);
  reg [(3'h5):(1'h0)] reg2067 = (1'h0);
  reg [(4'hf):(1'h0)] reg2063 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2056 = (1'h0);
  reg [(3'h5):(1'h0)] reg2066 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2065 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2064 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2063 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2062 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2061 = (1'h0);
  reg [(2'h3):(1'h0)] reg2060 = (1'h0);
  reg [(4'h8):(1'h0)] reg2059 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2058 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2057 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2056 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2055 = (1'h0);
  reg [(2'h3):(1'h0)] reg2054 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2053 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2052 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2051 = (1'h0);
  reg [(4'ha):(1'h0)] reg2050 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2049 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2048 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2047 = (1'h0);
  reg [(4'h8):(1'h0)] reg2046 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2045 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2044 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2043 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2042 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2041 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2040 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire2039;
  wire [(5'h10):(1'h0)] wire2038;
  wire signed [(4'h9):(1'h0)] wire2037;
  wire [(2'h2):(1'h0)] wire2036;
  reg [(3'h5):(1'h0)] reg2035 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2034 = (1'h0);
  reg [(4'hf):(1'h0)] reg2033 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2032 = (1'h0);
  reg [(2'h3):(1'h0)] reg2031 = (1'h0);
  reg [(2'h2):(1'h0)] reg2030 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2029 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2028 = (1'h0);
  reg [(5'h10):(1'h0)] reg2027 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2026 = (1'h0);
  reg [(4'hd):(1'h0)] reg2025 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2024 = (1'h0);
  reg [(4'ha):(1'h0)] reg2023 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2022 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2021 = (1'h0);
  reg [(4'hb):(1'h0)] reg2020 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2019 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2018 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2017 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2016 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2015 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2014 = (1'h0);
  reg [(3'h7):(1'h0)] reg2013 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2012 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2011 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2010 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2009 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2008 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2007 = (1'h0);
  reg [(4'h9):(1'h0)] reg2006 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2005 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2004 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2003 = (1'h0);
  reg [(4'ha):(1'h0)] reg2002 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2001 = (1'h0);
  reg [(3'h7):(1'h0)] reg2000 = (1'h0);
  reg [(3'h7):(1'h0)] reg1999 = (1'h0);
  reg [(2'h3):(1'h0)] reg1998 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1997 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1996 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1995 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1982 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1978 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1976 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1975 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1972 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1970 = (1'h0);
  reg [(4'he):(1'h0)] reg1968 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1967 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1987 = (1'h0);
  reg [(5'h10):(1'h0)] reg1994 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1993 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1992 = (1'h0);
  reg [(2'h2):(1'h0)] reg1991 = (1'h0);
  reg [(3'h5):(1'h0)] reg1990 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1989 = (1'h0);
  reg [(2'h3):(1'h0)] reg1988 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1987 = (1'h0);
  reg [(4'h8):(1'h0)] reg1986 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1985 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1984 = (1'h0);
  reg [(4'he):(1'h0)] reg1983 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1982 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1981 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1980 = (1'h0);
  reg [(4'hd):(1'h0)] reg1979 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1978 = (1'h0);
  reg [(4'h8):(1'h0)] reg1977 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1976 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1975 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1974 = (1'h0);
  reg [(4'hd):(1'h0)] reg1973 = (1'h0);
  reg [(2'h3):(1'h0)] reg1972 = (1'h0);
  reg [(4'hf):(1'h0)] reg1971 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1970 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1969 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1968 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1967 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1966 = (1'h0);
  wire signed [(4'he):(1'h0)] wire1965;
  wire [(3'h6):(1'h0)] wire1964;
  wire signed [(4'hf):(1'h0)] wire1963;
  wire signed [(4'h9):(1'h0)] wire1962;
  wire signed [(4'hd):(1'h0)] wire1961;
  wire signed [(2'h2):(1'h0)] wire1960;
  reg [(3'h7):(1'h0)] reg1886 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1878 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1877 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1931 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1930 = (1'h0);
  reg [(4'hb):(1'h0)] reg1959 = (1'h0);
  reg [(2'h3):(1'h0)] reg1958 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1957 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1956 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1944 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1955 = (1'h0);
  reg [(3'h7):(1'h0)] reg1954 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1953 = (1'h0);
  reg [(2'h3):(1'h0)] reg1952 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1951 = (1'h0);
  reg [(3'h5):(1'h0)] reg1950 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1949 = (1'h0);
  reg [(4'h9):(1'h0)] reg1948 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1947 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1946 = (1'h0);
  reg [(5'h10):(1'h0)] reg1945 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1944 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1943 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1942 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1941 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1940 = (1'h0);
  reg [(4'hc):(1'h0)] reg1939 = (1'h0);
  reg [(4'he):(1'h0)] reg1938 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1937 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1936 = (1'h0);
  reg [(4'hf):(1'h0)] reg1935 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1934 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1933 = (1'h0);
  reg [(5'h10):(1'h0)] reg1932 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1931 = (1'h0);
  reg [(3'h5):(1'h0)] reg1930 = (1'h0);
  reg [(4'he):(1'h0)] reg1929 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1928 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1913 = (1'h0);
  reg [(4'hb):(1'h0)] reg1909 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1906 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1898 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1927 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1926 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1925 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1924 = (1'h0);
  reg [(4'hd):(1'h0)] reg1919 = (1'h0);
  reg [(3'h6):(1'h0)] reg1923 = (1'h0);
  reg [(3'h7):(1'h0)] reg1922 = (1'h0);
  reg [(3'h4):(1'h0)] reg1921 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1920 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1919 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1918 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1917 = (1'h0);
  reg [(4'h9):(1'h0)] reg1916 = (1'h0);
  reg [(3'h7):(1'h0)] reg1915 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1914 = (1'h0);
  reg [(5'h10):(1'h0)] reg1913 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1912 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1911 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1910 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1909 = (1'h0);
  reg [(3'h4):(1'h0)] reg1908 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1902 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1907 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1906 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1905 = (1'h0);
  reg [(3'h5):(1'h0)] reg1904 = (1'h0);
  reg [(3'h6):(1'h0)] reg1903 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1902 = (1'h0);
  reg [(4'hd):(1'h0)] reg1901 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1900 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1899 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1898 = (1'h0);
  reg [(3'h7):(1'h0)] reg1897 = (1'h0);
  reg [(4'h8):(1'h0)] reg1896 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1895 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1894 = (1'h0);
  reg [(4'ha):(1'h0)] reg1893 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1892 = (1'h0);
  reg [(4'ha):(1'h0)] reg1891 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1890 = (1'h0);
  reg [(2'h2):(1'h0)] reg1889 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1888 = (1'h0);
  reg [(3'h4):(1'h0)] reg1887 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1886 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1881 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1879 = (1'h0);
  reg [(4'he):(1'h0)] forvar1876 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1875 = (1'h0);
  reg [(2'h2):(1'h0)] reg1874 = (1'h0);
  reg [(2'h3):(1'h0)] reg1885 = (1'h0);
  reg [(4'hc):(1'h0)] reg1884 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1883 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1882 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1881 = (1'h0);
  reg [(2'h2):(1'h0)] reg1880 = (1'h0);
  reg [(4'ha):(1'h0)] reg1879 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1878 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1877 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1876 = (1'h0);
  reg [(3'h7):(1'h0)] reg1875 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1874 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1873 = (1'h0);
  reg [(4'hb):(1'h0)] reg1872 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1871 = (1'h0);
  reg [(3'h6):(1'h0)] reg1870 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1869 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1868 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1867 = (1'h0);
  reg [(4'h9):(1'h0)] reg1867 = (1'h0);
  reg [(4'hb):(1'h0)] reg1866 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1865 = (1'h0);
  reg [(2'h2):(1'h0)] reg1864 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1863 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1859 = (1'h0);
  reg [(3'h4):(1'h0)] reg1857 = (1'h0);
  reg [(4'he):(1'h0)] reg1862 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1861 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1860 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1859 = (1'h0);
  reg [(3'h5):(1'h0)] reg1858 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1857 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1856 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1855 = (1'h0);
  reg [(2'h3):(1'h0)] reg1854 = (1'h0);
  reg [(4'ha):(1'h0)] reg1853 = (1'h0);
  reg [(4'h8):(1'h0)] reg1852 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1851 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1850 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1849 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1848 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1844 = (1'h0);
  reg [(4'ha):(1'h0)] reg1847 = (1'h0);
  reg [(2'h2):(1'h0)] reg1846 = (1'h0);
  reg [(4'hb):(1'h0)] reg1845 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1844 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1843 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1842 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1841 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1836 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1832 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1823 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1816 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1817 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1838 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1840 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1839 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1838 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1837 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1836 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1835 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1830 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1825 = (1'h0);
  reg [(4'hd):(1'h0)] reg1824 = (1'h0);
  reg [(3'h6):(1'h0)] reg1822 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1821 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1818 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1814 = (1'h0);
  reg [(4'hc):(1'h0)] reg1834 = (1'h0);
  reg [(4'h8):(1'h0)] reg1833 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1831 = (1'h0);
  reg [(4'hc):(1'h0)] reg1828 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1826 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1831 = (1'h0);
  reg [(3'h6):(1'h0)] reg1830 = (1'h0);
  reg [(4'ha):(1'h0)] reg1829 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1828 = (1'h0);
  reg [(2'h3):(1'h0)] reg1827 = (1'h0);
  reg [(3'h6):(1'h0)] reg1826 = (1'h0);
  reg [(4'he):(1'h0)] reg1825 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1824 = (1'h0);
  reg [(5'h10):(1'h0)] reg1823 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1822 = (1'h0);
  reg [(4'hd):(1'h0)] reg1821 = (1'h0);
  reg [(4'hc):(1'h0)] reg1820 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1819 = (1'h0);
  reg [(4'h8):(1'h0)] reg1818 = (1'h0);
  reg [(3'h5):(1'h0)] reg1817 = (1'h0);
  reg [(3'h4):(1'h0)] reg1816 = (1'h0);
  reg [(3'h4):(1'h0)] reg1815 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1814 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire1813;
  wire [(5'h10):(1'h0)] wire1812;
  wire signed [(4'hd):(1'h0)] wire1811;
  wire [(4'he):(1'h0)] wire1810;
  wire [(4'hc):(1'h0)] wire1809;
  assign y = {reg2153,
                 forvar2134,
                 reg2133,
                 reg2132,
                 forvar2129,
                 forvar2128,
                 reg2127,
                 reg2124,
                 reg2118,
                 forvar2116,
                 forvar2111,
                 reg2114,
                 forvar2113,
                 reg2109,
                 forvar2108,
                 reg2106,
                 reg2152,
                 reg2151,
                 reg2150,
                 reg2149,
                 reg2148,
                 reg2147,
                 reg2146,
                 reg2145,
                 forvar2144,
                 reg2143,
                 forvar2142,
                 reg2141,
                 reg2139,
                 reg2140,
                 forvar2139,
                 forvar2138,
                 reg2137,
                 reg2136,
                 reg2135,
                 reg2134,
                 forvar2133,
                 forvar2132,
                 reg2131,
                 reg2130,
                 reg2129,
                 reg2128,
                 forvar2127,
                 reg2126,
                 reg2125,
                 forvar2124,
                 reg2123,
                 reg2122,
                 forvar2121,
                 reg2120,
                 reg2119,
                 forvar2118,
                 reg2117,
                 reg2116,
                 reg2115,
                 forvar2114,
                 reg2113,
                 reg2112,
                 reg2111,
                 reg2110,
                 forvar2109,
                 reg2108,
                 forvar2107,
                 forvar2106,
                 reg2093,
                 reg2105,
                 reg2104,
                 reg2103,
                 forvar2102,
                 reg2101,
                 reg2100,
                 reg2099,
                 reg2098,
                 reg2097,
                 forvar2096,
                 reg2095,
                 reg2094,
                 forvar2093,
                 reg2092,
                 reg2091,
                 reg2090,
                 reg2089,
                 forvar2088,
                 reg2087,
                 reg2086,
                 reg2085,
                 reg2084,
                 reg2083,
                 forvar2082,
                 reg2081,
                 forvar2080,
                 forvar2079,
                 reg2078,
                 forvar2077,
                 reg2076,
                 reg2075,
                 reg2074,
                 forvar2073,
                 forvar2070,
                 reg2069,
                 reg2073,
                 reg2072,
                 reg2071,
                 reg2070,
                 forvar2069,
                 reg2068,
                 reg2067,
                 reg2063,
                 reg2056,
                 reg2066,
                 forvar2065,
                 reg2064,
                 forvar2063,
                 reg2062,
                 reg2061,
                 reg2060,
                 reg2059,
                 reg2058,
                 reg2057,
                 forvar2056,
                 forvar2055,
                 reg2054,
                 reg2053,
                 forvar2052,
                 reg2051,
                 reg2050,
                 reg2049,
                 reg2048,
                 reg2047,
                 reg2046,
                 reg2045,
                 reg2044,
                 forvar2043,
                 forvar2042,
                 forvar2041,
                 forvar2040,
                 wire2039,
                 wire2038,
                 wire2037,
                 wire2036,
                 reg2035,
                 reg2034,
                 reg2033,
                 forvar2032,
                 reg2031,
                 reg2030,
                 forvar2029,
                 forvar2028,
                 reg2027,
                 reg2026,
                 reg2025,
                 reg2024,
                 reg2023,
                 reg2022,
                 reg2021,
                 reg2020,
                 reg2019,
                 reg2018,
                 reg2017,
                 reg2016,
                 forvar2015,
                 reg2014,
                 reg2013,
                 reg2012,
                 reg2011,
                 forvar2010,
                 reg2009,
                 reg2008,
                 reg2007,
                 reg2006,
                 forvar2005,
                 forvar2004,
                 forvar2003,
                 reg2002,
                 reg2001,
                 reg2000,
                 reg1999,
                 reg1998,
                 forvar1997,
                 forvar1996,
                 forvar1995,
                 reg1982,
                 forvar1978,
                 reg1976,
                 reg1975,
                 forvar1972,
                 reg1970,
                 reg1968,
                 reg1967,
                 reg1987,
                 reg1994,
                 reg1993,
                 reg1992,
                 reg1991,
                 reg1990,
                 reg1989,
                 reg1988,
                 forvar1987,
                 reg1986,
                 reg1985,
                 reg1984,
                 reg1983,
                 forvar1982,
                 reg1981,
                 reg1980,
                 reg1979,
                 reg1978,
                 reg1977,
                 forvar1976,
                 forvar1975,
                 reg1974,
                 reg1973,
                 reg1972,
                 reg1971,
                 forvar1970,
                 reg1969,
                 forvar1968,
                 forvar1967,
                 forvar1966,
                 wire1965,
                 wire1964,
                 wire1963,
                 wire1962,
                 wire1961,
                 wire1960,
                 reg1886,
                 forvar1878,
                 forvar1877,
                 reg1931,
                 forvar1930,
                 reg1959,
                 reg1958,
                 reg1957,
                 forvar1956,
                 forvar1944,
                 reg1955,
                 reg1954,
                 reg1953,
                 reg1952,
                 reg1951,
                 reg1950,
                 reg1949,
                 reg1948,
                 reg1947,
                 reg1946,
                 reg1945,
                 reg1944,
                 reg1943,
                 reg1942,
                 reg1941,
                 forvar1940,
                 reg1939,
                 reg1938,
                 forvar1937,
                 forvar1936,
                 reg1935,
                 reg1934,
                 reg1933,
                 reg1932,
                 forvar1931,
                 reg1930,
                 reg1929,
                 forvar1928,
                 forvar1913,
                 reg1909,
                 forvar1906,
                 forvar1898,
                 reg1927,
                 reg1926,
                 forvar1925,
                 reg1924,
                 reg1919,
                 reg1923,
                 reg1922,
                 reg1921,
                 reg1920,
                 forvar1919,
                 reg1918,
                 forvar1917,
                 reg1916,
                 reg1915,
                 reg1914,
                 reg1913,
                 reg1912,
                 reg1911,
                 reg1910,
                 forvar1909,
                 reg1908,
                 reg1902,
                 reg1907,
                 reg1906,
                 reg1905,
                 reg1904,
                 reg1903,
                 forvar1902,
                 reg1901,
                 reg1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 reg1896,
                 forvar1895,
                 reg1894,
                 reg1893,
                 reg1892,
                 reg1891,
                 reg1890,
                 reg1889,
                 reg1888,
                 reg1887,
                 forvar1886,
                 reg1881,
                 forvar1879,
                 forvar1876,
                 forvar1875,
                 reg1874,
                 reg1885,
                 reg1884,
                 reg1883,
                 reg1882,
                 forvar1881,
                 reg1880,
                 reg1879,
                 reg1878,
                 reg1877,
                 reg1876,
                 reg1875,
                 forvar1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 reg1870,
                 reg1869,
                 reg1868,
                 forvar1867,
                 reg1867,
                 reg1866,
                 reg1865,
                 reg1864,
                 reg1863,
                 reg1859,
                 reg1857,
                 reg1862,
                 reg1861,
                 reg1860,
                 forvar1859,
                 reg1858,
                 forvar1857,
                 forvar1856,
                 forvar1855,
                 reg1854,
                 reg1853,
                 reg1852,
                 forvar1851,
                 reg1850,
                 forvar1849,
                 reg1848,
                 forvar1844,
                 reg1847,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1843,
                 forvar1842,
                 reg1841,
                 forvar1836,
                 forvar1832,
                 forvar1823,
                 forvar1816,
                 forvar1817,
                 forvar1838,
                 reg1840,
                 reg1839,
                 reg1838,
                 reg1837,
                 reg1836,
                 forvar1835,
                 forvar1830,
                 forvar1825,
                 reg1824,
                 reg1822,
                 forvar1821,
                 forvar1818,
                 forvar1814,
                 reg1834,
                 reg1833,
                 reg1832,
                 forvar1831,
                 reg1828,
                 forvar1826,
                 reg1831,
                 reg1830,
                 reg1829,
                 forvar1828,
                 reg1827,
                 reg1826,
                 reg1825,
                 forvar1824,
                 reg1823,
                 forvar1822,
                 reg1821,
                 reg1820,
                 reg1819,
                 reg1818,
                 reg1817,
                 reg1816,
                 reg1815,
                 reg1814,
                 wire1813,
                 wire1812,
                 wire1811,
                 wire1810,
                 wire1809,
                 (1'h0)};
  assign wire1809 = wire1808;
  assign wire1810 = (((wire1804 ?
                            (wire1806 ?
                                wire1805 : wire1806) : (wire1807 || (8'hb8))) ?
                        $unsigned($unsigned(wire1808)) : {$signed(wire1807)}) + $signed({(wire1806 ?
                            wire1808 : wire1808)}));
  assign wire1811 = {$signed(wire1808[(4'h8):(2'h2)])};
  assign wire1812 = ({(wire1811 <= wire1810)} ? $unsigned((8'hb0)) : wire1811);
  assign wire1813 = {{$signed((wire1807 ? wire1806 : (8'hae)))}};
  always
    @(posedge clk) begin
      if ($signed(wire1811[(4'h8):(2'h2)]))
        begin
          if ($signed(wire1812))
            begin
              if ((wire1812 <= $signed((wire1808[(4'h8):(3'h6)] ^~ ((8'ha5) ?
                  (8'h9c) : wire1808)))))
                begin
                  reg1814 <= wire1806[(3'h5):(2'h2)];
                  if (($signed($unsigned({wire1807})) ?
                      (($unsigned(wire1808) ?
                              wire1810[(3'h6):(1'h1)] : wire1809) ?
                          $unsigned(wire1808) : wire1804) : (8'had)))
                    begin
                      reg1815 <= (wire1806[(3'h5):(2'h2)] ~^ ({(wire1807 || wire1812)} != wire1808));
                      reg1816 <= ($signed(reg1814[(1'h0):(1'h0)]) <<< (^~{(^wire1811)}));
                      reg1817 <= $unsigned((wire1811 - ((wire1808 * (8'ha8)) ~^ {(8'hba)})));
                      reg1818 <= wire1806[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg1815 <= $signed($signed(($unsigned(wire1813) >>> $signed(reg1815))));
                      reg1816 <= $signed(wire1810);
                      reg1817 <= wire1811[(1'h1):(1'h0)];
                    end
                  if ($signed(wire1806))
                    begin
                      reg1819 <= ((^~(~|(wire1806 >>> reg1815))) | $signed(wire1813));
                      reg1820 <= wire1808;
                      reg1821 <= $signed($signed({(&reg1819)}));
                    end
                  else
                    begin
                      reg1819 <= reg1816[(1'h1):(1'h0)];
                      reg1820 <= {reg1816[(3'h4):(2'h3)]};
                      reg1821 <= (((~&wire1809) ^ wire1808[(4'h9):(2'h3)]) >>> (-{(wire1809 ^~ reg1821)}));
                    end
                end
              else
                begin
                  if ($signed((~|$unsigned((|(8'hb7))))))
                    begin
                      reg1814 <= wire1813;
                      reg1815 <= wire1805;
                      reg1816 <= (~^reg1818);
                      reg1817 <= $signed(((wire1811 <<< $signed(wire1806)) ?
                          reg1821 : reg1816[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg1814 <= (8'ha4);
                      reg1815 <= $unsigned(reg1820[(3'h6):(1'h0)]);
                      reg1816 <= wire1806[(2'h2):(1'h0)];
                      reg1817 <= $signed(wire1805);
                    end
                  if (wire1812)
                    begin
                      reg1818 <= {$signed(($unsigned(reg1815) ?
                              {reg1814} : (~^wire1808)))};
                      reg1819 <= ((wire1812 > (((8'hb2) ?
                          (8'hb2) : reg1819) >> (|wire1810))) <= $signed((~wire1812[(4'h9):(4'h9)])));
                    end
                  else
                    begin
                      reg1818 <= {(~^(~&$unsigned(reg1816)))};
                      reg1819 <= reg1820;
                      reg1820 <= reg1820[(3'h5):(1'h1)];
                      reg1821 <= $unsigned({(((8'had) < wire1812) ^~ $unsigned(reg1818))});
                    end
                  for (forvar1822 = (1'h0); (forvar1822 < (1'h0)); forvar1822 = (forvar1822 + (1'h1)))
                    begin
                      reg1823 <= wire1813[(2'h3):(2'h2)];
                    end
                end
              if ($unsigned($unsigned({(|(8'hb9))})))
                begin
                  for (forvar1824 = (1'h0); (forvar1824 < (2'h2)); forvar1824 = (forvar1824 + (1'h1)))
                    begin
                      reg1825 <= $unsigned(($unsigned(((8'h9c) ?
                          reg1814 : wire1804)) | wire1808));
                      reg1826 <= reg1816[(3'h4):(3'h4)];
                    end
                  reg1827 <= reg1816;
                  for (forvar1828 = (1'h0); (forvar1828 < (2'h2)); forvar1828 = (forvar1828 + (1'h1)))
                    begin
                      reg1829 <= (8'haa);
                    end
                  if ($signed(((8'hb7) | (~wire1811))))
                    begin
                      reg1830 <= {($signed((+reg1821)) ?
                              $unsigned($unsigned(reg1829)) : $signed((reg1818 | reg1819)))};
                      reg1831 <= $unsigned($signed($signed((+reg1821))));
                    end
                  else
                    begin
                      reg1830 <= {$unsigned($signed(forvar1828))};
                    end
                end
              else
                begin
                  for (forvar1824 = (1'h0); (forvar1824 < (1'h0)); forvar1824 = (forvar1824 + (1'h1)))
                    begin
                      reg1825 <= $signed($signed(((wire1807 >> reg1817) ?
                          forvar1824[(1'h0):(1'h0)] : {(8'hab)})));
                    end
                  for (forvar1826 = (1'h0); (forvar1826 < (2'h2)); forvar1826 = (forvar1826 + (1'h1)))
                    begin
                      reg1827 <= (reg1831 ?
                          ({reg1815[(2'h3):(2'h2)]} ?
                              reg1827[(1'h1):(1'h1)] : $unsigned({wire1812})) : wire1808);
                    end
                  if (reg1831[(3'h4):(1'h0)])
                    begin
                      reg1828 <= $unsigned($unsigned((&(reg1826 ?
                          (8'h9e) : wire1806))));
                      reg1829 <= reg1828[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1828 <= $signed(((8'hb5) & $signed({wire1811})));
                      reg1829 <= $signed(wire1806[(3'h6):(3'h5)]);
                      reg1830 <= {(~^$signed($signed(reg1821)))};
                    end
                  for (forvar1831 = (1'h0); (forvar1831 < (1'h0)); forvar1831 = (forvar1831 + (1'h1)))
                    begin
                      reg1832 <= ((~&(forvar1824[(2'h2):(1'h1)] ?
                              $signed(forvar1822) : forvar1831)) ?
                          (wire1804[(3'h5):(3'h5)] ?
                              reg1828[(2'h2):(2'h2)] : (~^(8'hb2))) : ((((8'hab) ?
                                  reg1821 : wire1810) ?
                              (reg1828 <= reg1821) : wire1804[(3'h6):(1'h0)]) | $signed({reg1825})));
                      reg1833 <= $unsigned((^~$signed({wire1804})));
                      reg1834 <= {reg1814[(4'h9):(3'h7)]};
                    end
                end
            end
          else
            begin
              for (forvar1814 = (1'h0); (forvar1814 < (1'h1)); forvar1814 = (forvar1814 + (1'h1)))
                begin
                  if ((($unsigned(reg1828[(2'h3):(2'h3)]) ^ $unsigned((^~reg1815))) ?
                      (reg1819[(2'h3):(2'h3)] ?
                          reg1819 : reg1831) : ($unsigned((reg1831 < reg1821)) ?
                          ((^~reg1834) ?
                              $unsigned((8'hab)) : ((8'hb4) <<< wire1808)) : wire1805)))
                    begin
                      reg1815 <= reg1819;
                      reg1816 <= wire1812[(1'h0):(1'h0)];
                      reg1817 <= (($signed($unsigned(wire1807)) || reg1823) ?
                          (forvar1814[(4'h8):(3'h7)] ^~ $unsigned({reg1816})) : $signed(($signed(wire1804) ^~ {reg1816})));
                    end
                  else
                    begin
                      reg1815 <= (+wire1808[(1'h0):(1'h0)]);
                      reg1816 <= ($signed($signed({reg1828})) ?
                          (~^((forvar1831 >>> wire1810) ?
                              reg1834[(4'hc):(1'h1)] : (wire1811 || reg1834))) : reg1826);
                    end
                  for (forvar1818 = (1'h0); (forvar1818 < (2'h3)); forvar1818 = (forvar1818 + (1'h1)))
                    begin
                      reg1819 <= ((&$unsigned((|wire1805))) & reg1818[(2'h3):(1'h1)]);
                      reg1820 <= reg1814;
                    end
                end
              for (forvar1821 = (1'h0); (forvar1821 < (2'h3)); forvar1821 = (forvar1821 + (1'h1)))
                begin
                  if (({$signed({wire1805})} != reg1833))
                    begin
                      reg1822 <= ({reg1823} + reg1817[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg1822 <= (wire1811 ? reg1831 : $unsigned(forvar1824));
                      reg1823 <= reg1834;
                      reg1824 <= {reg1817};
                    end
                end
              if ($unsigned((8'hb7)))
                begin
                  if ((^$signed((~(+forvar1822)))))
                    begin
                      reg1825 <= reg1825[(3'h5):(1'h1)];
                      reg1826 <= forvar1818[(4'hd):(1'h0)];
                      reg1827 <= (~^forvar1822);
                      reg1828 <= ($unsigned(({reg1820} < {reg1830})) != wire1808[(3'h7):(3'h5)]);
                    end
                  else
                    begin
                      reg1825 <= $signed(reg1828[(2'h3):(2'h3)]);
                      reg1826 <= ($signed((wire1813 ?
                              $signed((8'hb7)) : reg1831)) ?
                          (^wire1812[(3'h7):(2'h3)]) : (((reg1818 & reg1834) ?
                                  $unsigned(reg1823) : $signed(reg1834)) ?
                              (((8'h9d) != (8'hb5)) << (^wire1810)) : {(-forvar1826)}));
                      reg1827 <= reg1818;
                    end
                end
              else
                begin
                  for (forvar1825 = (1'h0); (forvar1825 < (2'h3)); forvar1825 = (forvar1825 + (1'h1)))
                    begin
                      reg1826 <= forvar1814;
                      reg1827 <= forvar1822;
                      reg1828 <= wire1805;
                      reg1829 <= reg1833[(2'h3):(1'h0)];
                    end
                  for (forvar1830 = (1'h0); (forvar1830 < (2'h2)); forvar1830 = (forvar1830 + (1'h1)))
                    begin
                      reg1831 <= ((((forvar1831 <= reg1832) ?
                              reg1830[(3'h4):(1'h0)] : $signed(forvar1818)) != $signed((wire1809 ?
                              wire1805 : reg1823))) ?
                          reg1817 : reg1826[(3'h5):(1'h0)]);
                      reg1832 <= reg1834[(3'h4):(2'h3)];
                      reg1833 <= $unsigned({forvar1830});
                      reg1834 <= {({forvar1828[(4'hb):(4'h9)]} ?
                              reg1825 : ($unsigned(reg1818) ?
                                  reg1831 : {reg1815}))};
                    end
                  for (forvar1835 = (1'h0); (forvar1835 < (1'h1)); forvar1835 = (forvar1835 + (1'h1)))
                    begin
                      reg1836 <= {reg1830[(1'h1):(1'h1)]};
                    end
                end
              if (reg1816[(3'h4):(2'h2)])
                begin
                  if (reg1829)
                    begin
                      reg1837 <= reg1827[(2'h3):(1'h1)];
                      reg1838 <= forvar1822;
                      reg1839 <= $unsigned(wire1811[(3'h6):(2'h3)]);
                      reg1840 <= forvar1818[(4'h8):(2'h3)];
                    end
                  else
                    begin
                      reg1837 <= ($signed({wire1807[(3'h4):(1'h1)]}) > {reg1820[(3'h7):(2'h2)]});
                    end
                end
              else
                begin
                  reg1837 <= forvar1822[(3'h7):(3'h5)];
                  for (forvar1838 = (1'h0); (forvar1838 < (1'h1)); forvar1838 = (forvar1838 + (1'h1)))
                    begin
                      reg1839 <= $signed(forvar1831);
                    end
                end
            end
        end
      else
        begin
          for (forvar1814 = (1'h0); (forvar1814 < (2'h3)); forvar1814 = (forvar1814 + (1'h1)))
            begin
              reg1815 <= ((^reg1821[(3'h6):(1'h1)]) >> $signed($signed((forvar1831 >> wire1807))));
              if (forvar1821[(4'hf):(4'hb)])
                begin
                  reg1816 <= forvar1838;
                  for (forvar1817 = (1'h0); (forvar1817 < (2'h2)); forvar1817 = (forvar1817 + (1'h1)))
                    begin
                      reg1818 <= (+wire1806);
                      reg1819 <= ({$signed($unsigned((8'ha1)))} ?
                          $signed((8'ha1)) : ((((8'hb1) ?
                              reg1819 : forvar1835) + {reg1839}) >= (8'haf)));
                    end
                  reg1820 <= wire1810;
                  reg1821 <= $signed($signed($signed((reg1823 ~^ reg1837))));
                end
              else
                begin
                  for (forvar1816 = (1'h0); (forvar1816 < (2'h3)); forvar1816 = (forvar1816 + (1'h1)))
                    begin
                      reg1817 <= (~&{($signed(wire1813) ?
                              $signed(reg1825) : (^~forvar1828))});
                      reg1818 <= ($signed($unsigned($unsigned(reg1815))) ?
                          ($signed($unsigned(reg1830)) ?
                              ({reg1820} <<< ((8'hb7) > forvar1828)) : reg1823[(3'h7):(3'h6)]) : wire1812);
                      reg1819 <= forvar1818[(3'h5):(2'h2)];
                    end
                  reg1820 <= $signed(reg1823);
                end
              reg1822 <= $signed(reg1839);
              for (forvar1823 = (1'h0); (forvar1823 < (2'h2)); forvar1823 = (forvar1823 + (1'h1)))
                begin
                  for (forvar1824 = (1'h0); (forvar1824 < (2'h3)); forvar1824 = (forvar1824 + (1'h1)))
                    begin
                      reg1825 <= wire1806;
                      reg1826 <= (8'ha5);
                      reg1827 <= $signed((~&forvar1824[(1'h1):(1'h1)]));
                    end
                  for (forvar1828 = (1'h0); (forvar1828 < (2'h2)); forvar1828 = (forvar1828 + (1'h1)))
                    begin
                      reg1829 <= ($unsigned($signed((wire1809 >> reg1828))) ?
                          $signed($signed((reg1821 && wire1811))) : reg1819[(2'h3):(2'h3)]);
                      reg1830 <= ($unsigned(reg1821[(3'h6):(2'h3)]) ?
                          (wire1812 ?
                              ((reg1829 ? reg1825 : forvar1814) ?
                                  $signed((8'ha8)) : forvar1831[(3'h6):(2'h3)]) : $unsigned(wire1807)) : $signed(forvar1831[(4'h9):(3'h7)]));
                      reg1831 <= {{(^forvar1814)}};
                    end
                  for (forvar1832 = (1'h0); (forvar1832 < (2'h2)); forvar1832 = (forvar1832 + (1'h1)))
                    begin
                      reg1833 <= $unsigned($unsigned(reg1824));
                      reg1834 <= (reg1833 ?
                          (wire1805[(4'h8):(1'h0)] & ($signed(reg1838) + (reg1827 ?
                              forvar1824 : (8'h9e)))) : {wire1806});
                    end
                end
            end
          for (forvar1835 = (1'h0); (forvar1835 < (2'h2)); forvar1835 = (forvar1835 + (1'h1)))
            begin
              for (forvar1836 = (1'h0); (forvar1836 < (1'h0)); forvar1836 = (forvar1836 + (1'h1)))
                begin
                  if (wire1811[(4'hb):(2'h2)])
                    begin
                      reg1837 <= (8'hb1);
                    end
                  else
                    begin
                      reg1837 <= ((8'ha2) ?
                          forvar1818[(4'hb):(4'hb)] : ({(forvar1814 + (8'hb2))} ^~ $signed({forvar1838})));
                    end
                  if ((8'hb9))
                    begin
                      reg1838 <= forvar1818[(3'h5):(2'h3)];
                      reg1839 <= (reg1830 * forvar1816);
                    end
                  else
                    begin
                      reg1838 <= forvar1821;
                      reg1839 <= ((8'h9c) != $unsigned($unsigned({reg1817})));
                      reg1840 <= (^(~&$unsigned(reg1840)));
                      reg1841 <= $unsigned({$signed($signed(reg1830))});
                    end
                end
              if (reg1829[(3'h4):(2'h2)])
                begin
                  for (forvar1842 = (1'h0); (forvar1842 < (2'h2)); forvar1842 = (forvar1842 + (1'h1)))
                    begin
                      reg1843 <= {$signed({$signed(reg1826)})};
                      reg1844 <= (((!((8'hb8) ? reg1815 : reg1843)) ?
                              (~|(reg1840 ?
                                  wire1810 : forvar1836)) : $unsigned((forvar1842 & (8'hb5)))) ?
                          {{(!reg1833)}} : ((((8'ha8) ~^ wire1804) ?
                                  (forvar1826 ? reg1823 : reg1826) : (reg1821 ?
                                      reg1839 : reg1822)) ?
                              reg1840 : (reg1816[(2'h2):(1'h1)] ~^ reg1839[(1'h0):(1'h0)])));
                      reg1845 <= $signed($unsigned($unsigned(reg1831[(3'h5):(1'h1)])));
                    end
                  if ((~&reg1832))
                    begin
                      reg1846 <= (8'hb5);
                    end
                  else
                    begin
                      reg1846 <= ((^~forvar1830[(1'h1):(1'h0)]) ?
                          forvar1832 : {$signed({reg1843})});
                    end
                  reg1847 <= {reg1824};
                end
              else
                begin
                  for (forvar1842 = (1'h0); (forvar1842 < (2'h3)); forvar1842 = (forvar1842 + (1'h1)))
                    begin
                      reg1843 <= reg1832[(4'hc):(3'h5)];
                    end
                  for (forvar1844 = (1'h0); (forvar1844 < (1'h1)); forvar1844 = (forvar1844 + (1'h1)))
                    begin
                      reg1845 <= (8'h9f);
                      reg1846 <= (!(reg1825[(2'h3):(1'h0)] ?
                          (reg1845 ^ forvar1821) : reg1840[(4'hd):(3'h5)]));
                      reg1847 <= wire1804;
                      reg1848 <= (reg1837[(1'h1):(1'h1)] <= wire1811);
                    end
                end
              for (forvar1849 = (1'h0); (forvar1849 < (1'h1)); forvar1849 = (forvar1849 + (1'h1)))
                begin
                  reg1850 <= $unsigned($unsigned(((+wire1812) ?
                      forvar1828 : $signed(reg1824))));
                  for (forvar1851 = (1'h0); (forvar1851 < (1'h0)); forvar1851 = (forvar1851 + (1'h1)))
                    begin
                      reg1852 <= {(~wire1807)};
                      reg1853 <= $signed(($unsigned({reg1816}) || wire1806));
                    end
                  reg1854 <= (reg1844[(4'ha):(1'h1)] ?
                      $unsigned(forvar1817) : (reg1833[(3'h5):(2'h2)] ?
                          {$signed(wire1810)} : reg1814[(3'h6):(1'h0)]));
                end
            end
        end
      for (forvar1855 = (1'h0); (forvar1855 < (2'h2)); forvar1855 = (forvar1855 + (1'h1)))
        begin
          for (forvar1856 = (1'h0); (forvar1856 < (2'h3)); forvar1856 = (forvar1856 + (1'h1)))
            begin
              if (forvar1831[(1'h1):(1'h0)])
                begin
                  for (forvar1857 = (1'h0); (forvar1857 < (1'h1)); forvar1857 = (forvar1857 + (1'h1)))
                    begin
                      reg1858 <= $signed($unsigned(($unsigned((8'ha6)) <<< (reg1816 >>> reg1822))));
                    end
                  for (forvar1859 = (1'h0); (forvar1859 < (2'h3)); forvar1859 = (forvar1859 + (1'h1)))
                    begin
                      reg1860 <= $unsigned(($unsigned({forvar1836}) ?
                          forvar1857[(1'h0):(1'h0)] : (^$signed(reg1819))));
                      reg1861 <= {(-reg1819[(3'h4):(2'h3)])};
                      reg1862 <= {{{wire1813[(2'h2):(1'h0)]}}};
                    end
                end
              else
                begin
                  if ((reg1841[(1'h1):(1'h1)] | reg1829))
                    begin
                      reg1857 <= $unsigned(forvar1835[(2'h3):(1'h0)]);
                      reg1858 <= $signed((((reg1843 ?
                          wire1806 : reg1822) && (wire1806 & reg1834)) >> reg1826));
                    end
                  else
                    begin
                      reg1857 <= $unsigned(wire1809);
                      reg1858 <= ((reg1834[(1'h1):(1'h0)] ?
                          $unsigned(reg1825[(4'hc):(3'h6)]) : ($unsigned(reg1828) + (8'hae))) >= (+reg1822[(1'h0):(1'h0)]));
                    end
                  reg1859 <= (+$signed(forvar1855[(2'h2):(1'h0)]));
                end
              if (((^$signed(reg1834[(4'ha):(4'h8)])) <= {$unsigned((^forvar1832))}))
                begin
                  reg1863 <= reg1841[(4'h8):(3'h4)];
                  if (reg1821[(4'hb):(1'h1)])
                    begin
                      reg1864 <= ($unsigned($unsigned($signed(reg1858))) ?
                          wire1805[(2'h3):(1'h0)] : {reg1823});
                      reg1865 <= wire1806[(1'h1):(1'h1)];
                      reg1866 <= ($unsigned(forvar1817[(3'h5):(3'h4)]) ?
                          ($signed((forvar1835 ?
                              (8'ha1) : reg1831)) > (^~(reg1857 ?
                              reg1825 : forvar1849))) : reg1818);
                      reg1867 <= $unsigned(forvar1824);
                    end
                  else
                    begin
                      reg1864 <= {(!$signed($unsigned(reg1836)))};
                    end
                end
              else
                begin
                  if (reg1818[(3'h6):(2'h3)])
                    begin
                      reg1863 <= (~|wire1812[(4'he):(4'h8)]);
                      reg1864 <= ($unsigned((reg1815 ^ $signed(reg1840))) ?
                          ((reg1857 >> (!wire1810)) ?
                              reg1815[(1'h1):(1'h1)] : $signed($signed((8'hb9)))) : (^reg1824[(1'h0):(1'h0)]));
                      reg1865 <= $signed($signed($signed(((8'hb8) ?
                          reg1826 : reg1854))));
                      reg1866 <= (-(~$unsigned((~reg1848))));
                    end
                  else
                    begin
                      reg1863 <= ((forvar1818[(3'h6):(3'h5)] < $unsigned((!(8'hb0)))) << wire1808[(1'h0):(1'h0)]);
                    end
                  for (forvar1867 = (1'h0); (forvar1867 < (1'h0)); forvar1867 = (forvar1867 + (1'h1)))
                    begin
                      reg1868 <= {((~&$unsigned(reg1858)) ?
                              $signed(((8'hb3) - wire1813)) : reg1846)};
                      reg1869 <= ($unsigned({reg1825[(4'hd):(4'hb)]}) ?
                          ($signed((wire1810 ? reg1865 : (8'haa))) ?
                              $unsigned((~^forvar1830)) : $unsigned((forvar1816 > forvar1836))) : $unsigned(((reg1815 ?
                              reg1853 : reg1858) << $signed(reg1847))));
                      reg1870 <= $signed($signed((reg1848[(1'h1):(1'h1)] ~^ $signed(reg1826))));
                    end
                  reg1871 <= reg1866[(3'h4):(1'h1)];
                  reg1872 <= reg1818;
                end
            end
        end
      reg1873 <= ((forvar1826[(4'h8):(3'h7)] ?
          $signed((!reg1844)) : (wire1805[(3'h6):(1'h0)] & {(8'ha7)})) == wire1810);
      if (reg1852)
        begin
          if ((8'ha6))
            begin
              if (forvar1821)
                begin
                  for (forvar1874 = (1'h0); (forvar1874 < (1'h1)); forvar1874 = (forvar1874 + (1'h1)))
                    begin
                      reg1875 <= (8'hb0);
                      reg1876 <= wire1810[(4'he):(4'h8)];
                    end
                  if (reg1834)
                    begin
                      reg1877 <= (&(^~{$signed(reg1870)}));
                      reg1878 <= $signed((&(~|{forvar1838})));
                    end
                  else
                    begin
                      reg1877 <= $unsigned(reg1831[(2'h2):(2'h2)]);
                      reg1878 <= reg1840[(3'h7):(1'h1)];
                      reg1879 <= {$signed(reg1819)};
                      reg1880 <= (!(wire1810[(4'hb):(1'h0)] ?
                          ((forvar1823 ?
                              forvar1859 : reg1876) | (^reg1826)) : reg1830));
                    end
                end
              else
                begin
                  for (forvar1874 = (1'h0); (forvar1874 < (2'h2)); forvar1874 = (forvar1874 + (1'h1)))
                    begin
                      reg1875 <= reg1825[(3'h6):(3'h5)];
                      reg1876 <= $signed($unsigned((((8'ha6) ?
                              reg1815 : reg1831) ?
                          reg1876[(2'h2):(1'h0)] : {reg1834})));
                      reg1877 <= ((reg1838[(3'h7):(2'h3)] >> reg1852[(2'h2):(1'h0)]) || (&($signed(reg1867) ?
                          (~reg1880) : $signed(reg1833))));
                      reg1878 <= forvar1838;
                    end
                end
              for (forvar1881 = (1'h0); (forvar1881 < (2'h3)); forvar1881 = (forvar1881 + (1'h1)))
                begin
                  if (reg1834)
                    begin
                      reg1882 <= reg1827[(1'h1):(1'h1)];
                      reg1883 <= (forvar1816[(4'ha):(1'h1)] ?
                          reg1875[(3'h4):(1'h1)] : (((-forvar1832) ^~ (~&wire1808)) ?
                              {(reg1872 >>> (8'hb7))} : $signed((forvar1816 ?
                                  reg1864 : reg1828))));
                      reg1884 <= $signed(reg1877);
                    end
                  else
                    begin
                      reg1882 <= $unsigned((forvar1818 ^~ {$unsigned(reg1822)}));
                      reg1883 <= $signed(((wire1807 ? forvar1838 : (-(8'hab))) ?
                          $unsigned((reg1827 ?
                              reg1883 : reg1857)) : ({forvar1816} && forvar1849[(3'h7):(2'h3)])));
                      reg1884 <= forvar1842;
                      reg1885 <= $unsigned($signed((~{reg1858})));
                    end
                end
            end
          else
            begin
              reg1874 <= (+{reg1865});
              for (forvar1875 = (1'h0); (forvar1875 < (2'h2)); forvar1875 = (forvar1875 + (1'h1)))
                begin
                  for (forvar1876 = (1'h0); (forvar1876 < (1'h0)); forvar1876 = (forvar1876 + (1'h1)))
                    begin
                      reg1877 <= $unsigned(((|reg1875[(2'h2):(2'h2)]) ?
                          $unsigned($signed(forvar1881)) : $signed((reg1879 >= reg1878))));
                    end
                  reg1878 <= {$signed($unsigned(forvar1875))};
                  for (forvar1879 = (1'h0); (forvar1879 < (1'h0)); forvar1879 = (forvar1879 + (1'h1)))
                    begin
                      reg1880 <= (forvar1817 ?
                          $unsigned(reg1836[(2'h3):(2'h2)]) : wire1813);
                    end
                  if (reg1822)
                    begin
                      reg1881 <= forvar1822[(3'h7):(1'h1)];
                      reg1882 <= $unsigned(({(|reg1883)} >> ((reg1861 & forvar1838) ?
                          (^~forvar1838) : (reg1876 ? reg1848 : forvar1867))));
                      reg1883 <= ({(+$unsigned(reg1880))} <= (&((~^(8'h9d)) ?
                          $unsigned(reg1863) : ((8'hac) | reg1865))));
                      reg1884 <= (-{$signed($unsigned(wire1804))});
                    end
                  else
                    begin
                      reg1881 <= $unsigned(reg1817[(3'h5):(1'h1)]);
                      reg1882 <= reg1834;
                      reg1883 <= ((reg1867[(3'h6):(3'h4)] << $unsigned(reg1877)) > (8'hb6));
                    end
                end
              reg1885 <= (~(((reg1871 ? forvar1855 : reg1845) ?
                      forvar1826 : (reg1885 + forvar1879)) ?
                  {forvar1831} : $signed(wire1812)));
              for (forvar1886 = (1'h0); (forvar1886 < (2'h2)); forvar1886 = (forvar1886 + (1'h1)))
                begin
                  if ($signed(($unsigned($unsigned(reg1837)) ?
                      (~|$unsigned((8'hba))) : (^~(8'h9e)))))
                    begin
                      reg1887 <= (($signed(reg1863) * (+(+reg1864))) ^~ ($signed({wire1806}) ?
                          $unsigned($unsigned(forvar1838)) : (^$signed((8'ha8)))));
                      reg1888 <= reg1846[(2'h2):(1'h1)];
                      reg1889 <= (reg1834 ?
                          forvar1838 : $unsigned($signed((reg1885 ?
                              wire1812 : reg1876))));
                    end
                  else
                    begin
                      reg1887 <= {$unsigned((+forvar1816[(3'h4):(3'h4)]))};
                      reg1888 <= $unsigned((forvar1825 >> $unsigned((^~(8'ha5)))));
                      reg1889 <= (forvar1844 == {forvar1824});
                      reg1890 <= ((reg1825[(4'h8):(3'h5)] ?
                          $unsigned((-reg1848)) : $unsigned((8'hb8))) | $unsigned($unsigned((8'ha4))));
                    end
                  if ($signed((^~$unsigned($signed(reg1837)))))
                    begin
                      reg1891 <= ((&(((8'h9d) * (8'hb3)) ?
                          reg1821 : (^~forvar1886))) >> (($unsigned((8'haa)) ?
                              reg1869[(4'ha):(2'h2)] : (^~(8'ha4))) ?
                          $signed(reg1838) : reg1824));
                      reg1892 <= reg1888;
                      reg1893 <= ($signed($signed((~&forvar1818))) ^ (&forvar1844));
                      reg1894 <= (($signed(reg1815) != $signed((reg1877 ?
                              reg1893 : reg1823))) ?
                          reg1868[(1'h0):(1'h0)] : reg1816[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1891 <= reg1873[(4'h8):(2'h3)];
                      reg1892 <= {((|reg1824[(3'h5):(3'h4)]) >> wire1804[(3'h4):(1'h1)])};
                      reg1893 <= reg1858[(2'h2):(1'h1)];
                      reg1894 <= (reg1860[(1'h0):(1'h0)] && (forvar1823[(2'h3):(1'h1)] ?
                          $signed($signed(reg1825)) : $signed((reg1819 * reg1885))));
                    end
                  for (forvar1895 = (1'h0); (forvar1895 < (1'h1)); forvar1895 = (forvar1895 + (1'h1)))
                    begin
                      reg1896 <= forvar1895[(1'h1):(1'h1)];
                      reg1897 <= (^$unsigned($signed($signed(reg1850))));
                    end
                end
            end
          if (reg1880)
            begin
              if (reg1893)
                begin
                  if ($signed(reg1819[(2'h2):(2'h2)]))
                    begin
                      reg1898 <= reg1828[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg1898 <= ((~^(^$unsigned((8'hb5)))) ?
                          reg1820 : (reg1826[(3'h6):(2'h2)] ?
                              $unsigned($unsigned(reg1837)) : $unsigned({reg1825})));
                    end
                  if ($unsigned($unsigned(forvar1814[(1'h1):(1'h1)])))
                    begin
                      reg1899 <= reg1816;
                      reg1900 <= ((&forvar1836) ?
                          reg1870 : (reg1819[(3'h5):(3'h5)] ?
                              (((8'ha4) ?
                                  reg1862 : reg1844) <<< (^~reg1854)) : forvar1823[(4'h9):(4'h8)]));
                      reg1901 <= $unsigned(((reg1893[(2'h2):(1'h0)] ?
                          (reg1824 && reg1889) : (reg1900 & reg1870)) >= (reg1837[(4'hc):(3'h6)] ~^ reg1837[(2'h3):(2'h3)])));
                    end
                  else
                    begin
                      reg1899 <= ($unsigned(forvar1832[(1'h1):(1'h0)]) & {({(8'ha9)} ?
                              (reg1868 ?
                                  forvar1823 : forvar1826) : (reg1862 ^~ reg1824))});
                    end
                  for (forvar1902 = (1'h0); (forvar1902 < (2'h3)); forvar1902 = (forvar1902 + (1'h1)))
                    begin
                      reg1903 <= forvar1867;
                      reg1904 <= (((|reg1823[(4'h9):(2'h3)]) ^ $unsigned((forvar1881 ?
                              reg1857 : reg1885))) ?
                          $unsigned((reg1890[(1'h0):(1'h0)] >= (reg1820 ?
                              (8'ha4) : forvar1879))) : $signed(($signed(forvar1902) ?
                              reg1899 : (forvar1875 ?
                                  forvar1828 : forvar1816))));
                      reg1905 <= $unsigned({({reg1863} ?
                              reg1869[(3'h7):(3'h7)] : (reg1871 ?
                                  reg1903 : reg1841))});
                    end
                  if (reg1894)
                    begin
                      reg1906 <= $signed((8'ha7));
                      reg1907 <= ($unsigned(($signed(reg1821) ?
                          reg1818[(3'h4):(2'h2)] : ((8'hae) ?
                              reg1843 : reg1819))) == {(^(~|reg1834))});
                    end
                  else
                    begin
                      reg1906 <= reg1873[(4'h9):(3'h5)];
                      reg1907 <= (reg1870 ?
                          wire1811 : $unsigned($unsigned(reg1846[(1'h1):(1'h0)])));
                    end
                end
              else
                begin
                  reg1898 <= $signed(reg1836[(2'h2):(1'h0)]);
                  if ((^$signed($signed(forvar1835))))
                    begin
                      reg1899 <= forvar1851[(4'h9):(3'h6)];
                    end
                  else
                    begin
                      reg1899 <= reg1838;
                      reg1900 <= wire1805[(1'h1):(1'h1)];
                      reg1901 <= {reg1818};
                    end
                  if ($signed({((8'hac) | $signed((8'h9d)))}))
                    begin
                      reg1902 <= {(forvar1842 ?
                              ($unsigned(reg1887) > $signed(reg1897)) : ((wire1804 ?
                                      forvar1828 : reg1825) ?
                                  (reg1836 & forvar1814) : reg1893[(2'h2):(1'h0)]))};
                    end
                  else
                    begin
                      reg1902 <= ($unsigned(forvar1874[(4'hd):(3'h4)]) ?
                          ($unsigned({reg1825}) >> reg1894) : ($signed($unsigned(reg1831)) != (~&$unsigned(reg1859))));
                    end
                end
              reg1908 <= $signed(reg1854);
              for (forvar1909 = (1'h0); (forvar1909 < (2'h2)); forvar1909 = (forvar1909 + (1'h1)))
                begin
                  if ({$signed($signed(wire1806[(1'h1):(1'h0)]))})
                    begin
                      reg1910 <= $unsigned($unsigned(forvar1835[(3'h7):(3'h5)]));
                    end
                  else
                    begin
                      reg1910 <= (((~&{reg1817}) && ($unsigned(forvar1875) ~^ $signed((8'ha8)))) ?
                          $unsigned((reg1872[(4'hb):(3'h7)] ?
                              reg1831 : forvar1879[(1'h1):(1'h1)])) : (|($unsigned((8'hb4)) + (reg1814 >= reg1840))));
                      reg1911 <= $unsigned((reg1822 ?
                          $signed(wire1807) : (-(reg1903 ?
                              (8'hb6) : forvar1874))));
                      reg1912 <= reg1852;
                    end
                  if ({$signed(($signed(forvar1822) * reg1910))})
                    begin
                      reg1913 <= (^~forvar1817);
                      reg1914 <= {reg1913[(2'h2):(2'h2)]};
                      reg1915 <= (reg1897 ?
                          $unsigned($signed((~|reg1852))) : (&((^~reg1868) >> forvar1830)));
                      reg1916 <= reg1911[(3'h7):(3'h4)];
                    end
                  else
                    begin
                      reg1913 <= $unsigned($signed((^(reg1913 ?
                          reg1874 : reg1854))));
                      reg1914 <= ((&$signed((~|reg1823))) && $signed((reg1846[(2'h2):(1'h1)] && (8'ha3))));
                    end
                  for (forvar1917 = (1'h0); (forvar1917 < (1'h0)); forvar1917 = (forvar1917 + (1'h1)))
                    begin
                      reg1918 <= $unsigned((+(reg1869[(3'h5):(2'h2)] ?
                          (8'ha8) : (forvar1856 ? reg1915 : reg1862))));
                    end
                end
              if (({reg1880[(1'h1):(1'h1)]} < (reg1820 ?
                  ((reg1833 ? reg1872 : reg1859) ?
                      reg1889[(1'h0):(1'h0)] : $unsigned(reg1823)) : $unsigned(reg1907))))
                begin
                  for (forvar1919 = (1'h0); (forvar1919 < (1'h0)); forvar1919 = (forvar1919 + (1'h1)))
                    begin
                      reg1920 <= (8'hae);
                      reg1921 <= (reg1906[(3'h4):(2'h2)] != $unsigned(($unsigned((8'ha5)) ?
                          $unsigned(reg1850) : ((8'ha2) ?
                              forvar1835 : reg1823))));
                      reg1922 <= (reg1857[(2'h2):(2'h2)] ?
                          {(-(reg1907 ? reg1881 : (8'haf)))} : {reg1921});
                      reg1923 <= {(~(reg1896 ?
                              (reg1875 ? wire1813 : reg1918) : {forvar1895}))};
                    end
                end
              else
                begin
                  if ($unsigned($signed($signed((reg1885 > (8'ha6))))))
                    begin
                      reg1919 <= $signed({$signed($signed(forvar1832))});
                      reg1920 <= reg1868[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg1919 <= (^~reg1860);
                    end
                  if ($unsigned(({(~|forvar1824)} ?
                      (!reg1817[(3'h4):(2'h3)]) : forvar1917[(3'h4):(1'h1)])))
                    begin
                      reg1921 <= $signed(($signed(forvar1821[(2'h3):(2'h3)]) ?
                          ((forvar1917 ? reg1877 : reg1854) ?
                              reg1880[(1'h1):(1'h0)] : $unsigned(forvar1823)) : (reg1864[(2'h2):(1'h1)] & $signed(reg1872))));
                      reg1922 <= (|reg1870);
                      reg1923 <= $signed(forvar1886);
                    end
                  else
                    begin
                      reg1921 <= (($unsigned(reg1880[(1'h1):(1'h0)]) == {forvar1875}) <<< $signed(reg1844));
                      reg1922 <= {$unsigned(forvar1828)};
                      reg1923 <= (reg1841 || reg1839[(3'h6):(1'h1)]);
                      reg1924 <= (($signed($signed(reg1899)) ~^ (-(reg1870 ?
                              reg1850 : (8'hb2)))) ?
                          (^reg1838[(4'hf):(1'h0)]) : ($unsigned(reg1858) < $unsigned((reg1876 >= reg1821))));
                    end
                  for (forvar1925 = (1'h0); (forvar1925 < (1'h1)); forvar1925 = (forvar1925 + (1'h1)))
                    begin
                      reg1926 <= ((~|reg1874) ?
                          (-$unsigned($signed((8'hb8)))) : reg1869);
                    end
                  reg1927 <= $signed($signed(reg1829[(3'h4):(2'h2)]));
                end
            end
          else
            begin
              for (forvar1898 = (1'h0); (forvar1898 < (2'h3)); forvar1898 = (forvar1898 + (1'h1)))
                begin
                  if (((reg1816 || forvar1823[(3'h5):(3'h5)]) ?
                      (reg1901 <= (-(reg1834 - reg1870))) : $signed($signed((reg1899 ?
                          reg1854 : forvar1824)))))
                    begin
                      reg1899 <= (($unsigned(wire1813) >= {$unsigned(reg1877)}) | $signed($unsigned((reg1871 ^ forvar1830))));
                    end
                  else
                    begin
                      reg1899 <= (!reg1902[(3'h4):(2'h2)]);
                    end
                  reg1900 <= $unsigned((((+(8'ha0)) ?
                          $unsigned(reg1820) : {reg1830}) ?
                      $signed((-forvar1822)) : $signed((8'hae))));
                end
              reg1901 <= (~^$unsigned((reg1828[(4'hb):(4'h9)] ?
                  reg1891 : ((8'ha3) ? reg1922 : reg1903))));
              for (forvar1902 = (1'h0); (forvar1902 < (1'h1)); forvar1902 = (forvar1902 + (1'h1)))
                begin
                  if (forvar1855[(2'h2):(2'h2)])
                    begin
                      reg1903 <= {(reg1827 ?
                              forvar1902[(3'h7):(2'h2)] : $unsigned((reg1880 | reg1902)))};
                      reg1904 <= $signed(reg1897[(2'h2):(2'h2)]);
                      reg1905 <= (^~forvar1875);
                    end
                  else
                    begin
                      reg1903 <= (-((~&(forvar1874 + wire1804)) ?
                          reg1845 : $signed({reg1857})));
                    end
                  for (forvar1906 = (1'h0); (forvar1906 < (1'h1)); forvar1906 = (forvar1906 + (1'h1)))
                    begin
                      reg1907 <= $unsigned($signed($signed(forvar1817)));
                      reg1908 <= $signed($signed((wire1805 ?
                          reg1891[(4'ha):(1'h1)] : $unsigned(forvar1842))));
                    end
                end
              if ($unsigned(((~$signed(reg1884)) || (^~reg1927))))
                begin
                  reg1909 <= reg1916;
                end
              else
                begin
                  if ($unsigned(reg1919[(4'hb):(1'h1)]))
                    begin
                      reg1909 <= reg1824[(1'h1):(1'h1)];
                      reg1910 <= $signed(($unsigned($signed(reg1864)) != $unsigned((forvar1835 || reg1833))));
                      reg1911 <= reg1926[(1'h0):(1'h0)];
                      reg1912 <= (^~$signed($unsigned($signed(reg1816))));
                    end
                  else
                    begin
                      reg1909 <= $signed($signed({(reg1846 ~^ reg1874)}));
                      reg1910 <= ((~|(-$signed(reg1912))) * (wire1807 << $unsigned($unsigned((8'hb3)))));
                    end
                  for (forvar1913 = (1'h0); (forvar1913 < (2'h2)); forvar1913 = (forvar1913 + (1'h1)))
                    begin
                      reg1914 <= {{reg1882}};
                      reg1915 <= (8'ha1);
                      reg1916 <= (~&forvar1832[(3'h6):(3'h6)]);
                    end
                end
            end
          if ((8'ha2))
            begin
              for (forvar1928 = (1'h0); (forvar1928 < (1'h0)); forvar1928 = (forvar1928 + (1'h1)))
                begin
                  if ((forvar1874[(1'h1):(1'h1)] ?
                      {$signed($signed(reg1911))} : reg1885))
                    begin
                      reg1929 <= reg1866[(2'h2):(1'h0)];
                      reg1930 <= (^($signed(reg1816) ?
                          ($unsigned(forvar1859) ?
                              (+forvar1844) : $signed((8'hb2))) : ((forvar1902 - (8'haf)) ?
                              reg1819 : forvar1881[(2'h2):(2'h2)])));
                    end
                  else
                    begin
                      reg1929 <= (&reg1927);
                      reg1930 <= reg1927;
                    end
                  for (forvar1931 = (1'h0); (forvar1931 < (1'h1)); forvar1931 = (forvar1931 + (1'h1)))
                    begin
                      reg1932 <= $unsigned((forvar1879[(1'h1):(1'h1)] > $signed((forvar1919 ?
                          (8'ha8) : forvar1818))));
                      reg1933 <= (8'h9c);
                      reg1934 <= $unsigned((reg1882 ?
                          (reg1868[(1'h1):(1'h0)] ?
                              (&wire1805) : $unsigned(forvar1902)) : {(8'hb4)}));
                      reg1935 <= reg1899;
                    end
                end
              for (forvar1936 = (1'h0); (forvar1936 < (2'h2)); forvar1936 = (forvar1936 + (1'h1)))
                begin
                  for (forvar1937 = (1'h0); (forvar1937 < (1'h0)); forvar1937 = (forvar1937 + (1'h1)))
                    begin
                      reg1938 <= $signed($signed({$signed(reg1865)}));
                      reg1939 <= wire1806[(3'h4):(1'h0)];
                    end
                  for (forvar1940 = (1'h0); (forvar1940 < (2'h3)); forvar1940 = (forvar1940 + (1'h1)))
                    begin
                      reg1941 <= $signed((forvar1844 ?
                          {(^(8'hb5))} : forvar1879));
                      reg1942 <= reg1833;
                    end
                  reg1943 <= $signed((~|reg1858[(3'h4):(1'h0)]));
                end
              if ({reg1843})
                begin
                  if ($signed((~reg1870)))
                    begin
                      reg1944 <= $unsigned(($signed(reg1871[(3'h6):(3'h4)]) > ({(8'ha8)} <<< (^reg1922))));
                      reg1945 <= {$unsigned($unsigned($unsigned(reg1922)))};
                      reg1946 <= $unsigned(($unsigned(forvar1823[(4'h9):(2'h3)]) & reg1837));
                      reg1947 <= {$signed($unsigned((reg1907 ?
                              wire1809 : forvar1867)))};
                    end
                  else
                    begin
                      reg1944 <= reg1915;
                    end
                  if ($signed($signed((~|$signed((8'hab))))))
                    begin
                      reg1948 <= ($unsigned(($unsigned(reg1899) ?
                          (forvar1818 ? reg1900 : (8'ha3)) : (reg1830 ?
                              reg1829 : reg1926))) & $signed((8'hb1)));
                      reg1949 <= {({reg1822[(3'h4):(2'h2)]} ?
                              {reg1919} : ({reg1938} ?
                                  (reg1938 ?
                                      reg1844 : reg1908) : $signed(wire1807)))};
                      reg1950 <= (reg1891[(2'h2):(1'h1)] ?
                          (reg1894[(3'h4):(3'h4)] ?
                              reg1920[(1'h1):(1'h0)] : (8'ha6)) : ((reg1898[(1'h0):(1'h0)] ^~ {forvar1906}) & (((8'hb7) >= (8'ha0)) ?
                              reg1853[(3'h7):(3'h5)] : reg1942)));
                      reg1951 <= (~(((8'hb8) + (8'hb8)) && $unsigned($signed(reg1839))));
                    end
                  else
                    begin
                      reg1948 <= (((reg1950[(1'h0):(1'h0)] ~^ reg1901) ?
                              ($unsigned((8'hae)) ?
                                  (reg1891 == reg1845) : $unsigned(forvar1886)) : reg1887[(2'h3):(1'h0)]) ?
                          ($signed((~^forvar1937)) != $unsigned({forvar1902})) : ({$unsigned(forvar1849)} ?
                              (wire1806[(2'h3):(1'h1)] ?
                                  (~forvar1818) : reg1875[(3'h4):(1'h0)]) : $unsigned(forvar1817[(2'h3):(2'h3)])));
                    end
                  if ((({{forvar1867}} ^ (reg1838 ?
                      (~^reg1898) : $signed(reg1898))) ^~ (-(~^$signed(reg1906)))))
                    begin
                      reg1952 <= (8'hba);
                      reg1953 <= (~(!($signed(reg1952) ?
                          (wire1806 ?
                              wire1805 : reg1879) : reg1952[(1'h1):(1'h1)])));
                      reg1954 <= ($signed((+$unsigned(reg1898))) ?
                          (($signed(wire1812) ?
                              {reg1834} : {(8'hb3)}) * (reg1823[(2'h2):(1'h0)] >= reg1904)) : (!reg1815[(1'h0):(1'h0)]));
                      reg1955 <= reg1830[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg1952 <= (reg1840 ?
                          {$signed((&wire1811))} : $signed($unsigned((reg1919 ?
                              reg1836 : wire1810))));
                      reg1953 <= $unsigned(forvar1842[(4'ha):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar1944 = (1'h0); (forvar1944 < (2'h3)); forvar1944 = (forvar1944 + (1'h1)))
                    begin
                      reg1945 <= ($signed((reg1867[(3'h7):(1'h1)] >>> (8'hb0))) + (((|forvar1830) > {forvar1814}) ?
                          ({(8'hb7)} ?
                              $signed(wire1806) : $unsigned(reg1930)) : $signed($unsigned((8'had)))));
                    end
                  reg1946 <= ((^reg1941[(3'h6):(3'h6)]) ?
                      (8'hb7) : (&{$unsigned((8'hb9))}));
                  reg1947 <= ({reg1846} ?
                      (~reg1951[(1'h1):(1'h1)]) : reg1871[(4'h9):(2'h2)]);
                end
              for (forvar1956 = (1'h0); (forvar1956 < (1'h1)); forvar1956 = (forvar1956 + (1'h1)))
                begin
                  if ((($signed((reg1829 ? forvar1835 : reg1904)) ?
                      $signed(reg1923) : (forvar1831 ?
                          $signed(reg1923) : (+reg1930))) | reg1823[(4'h8):(3'h7)]))
                    begin
                      reg1957 <= reg1941;
                      reg1958 <= reg1818;
                      reg1959 <= $signed($unsigned(reg1828[(4'ha):(3'h5)]));
                    end
                  else
                    begin
                      reg1957 <= {$unsigned($signed({forvar1821}))};
                      reg1958 <= (!$unsigned(((forvar1944 ?
                          reg1843 : (8'ha6)) ^~ (&reg1879))));
                      reg1959 <= {reg1831};
                    end
                end
            end
          else
            begin
              for (forvar1928 = (1'h0); (forvar1928 < (2'h2)); forvar1928 = (forvar1928 + (1'h1)))
                begin
                  reg1929 <= $signed($signed(($signed(reg1862) ?
                      forvar1928 : $signed((8'hb5)))));
                  for (forvar1930 = (1'h0); (forvar1930 < (1'h0)); forvar1930 = (forvar1930 + (1'h1)))
                    begin
                      reg1931 <= $signed(((reg1839[(1'h0):(1'h0)] ?
                              {reg1934} : (|(8'hb4))) ?
                          forvar1856[(1'h1):(1'h0)] : ($unsigned(reg1884) <= $signed(forvar1909))));
                      reg1932 <= (!($signed(forvar1830[(2'h2):(1'h0)]) || {(reg1841 - reg1860)}));
                      reg1933 <= forvar1814[(3'h6):(1'h0)];
                    end
                end
              reg1934 <= (8'h9c);
            end
        end
      else
        begin
          if ((8'hb6))
            begin
              if (reg1924[(2'h3):(2'h2)])
                begin
                  if (((forvar1849[(3'h7):(3'h5)] ?
                      $signed(((8'ha4) ^~ reg1864)) : reg1938[(3'h6):(1'h0)]) & ({(forvar1838 ?
                          forvar1857 : reg1839)} < ($unsigned(reg1939) ?
                      (wire1805 - reg1954) : $unsigned(reg1858)))))
                    begin
                      reg1874 <= ($signed($signed({forvar1828})) ?
                          (^~reg1869[(4'hd):(4'hd)]) : (!{(reg1893 ?
                                  reg1832 : reg1906)}));
                      reg1875 <= (8'hb4);
                      reg1876 <= (!($unsigned((~^forvar1913)) != ({forvar1913} ?
                          reg1823 : {reg1907})));
                    end
                  else
                    begin
                      reg1874 <= reg1946[(2'h3):(2'h2)];
                      reg1875 <= (reg1954 ?
                          $unsigned(((forvar1816 <= reg1844) ?
                              reg1911[(2'h2):(1'h0)] : (reg1873 ?
                                  reg1828 : reg1901))) : reg1930);
                      reg1876 <= reg1862[(3'h4):(3'h4)];
                      reg1877 <= forvar1906[(2'h3):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar1874 = (1'h0); (forvar1874 < (1'h0)); forvar1874 = (forvar1874 + (1'h1)))
                    begin
                      reg1875 <= $unsigned((|$signed(reg1929)));
                      reg1876 <= $signed((8'h9c));
                    end
                  for (forvar1877 = (1'h0); (forvar1877 < (1'h1)); forvar1877 = (forvar1877 + (1'h1)))
                    begin
                      reg1878 <= $signed(((wire1808[(3'h7):(1'h1)] ?
                          $unsigned(wire1806) : $signed(forvar1867)) == ($unsigned((8'ha0)) & $unsigned(reg1862))));
                    end
                end
              for (forvar1879 = (1'h0); (forvar1879 < (2'h3)); forvar1879 = (forvar1879 + (1'h1)))
                begin
                  reg1880 <= (^~(reg1826 ?
                      reg1945[(4'ha):(2'h3)] : $unsigned((reg1884 ?
                          reg1833 : wire1806))));
                  if ($unsigned($unsigned(({reg1848} ?
                      (reg1845 >>> reg1931) : (&wire1813)))))
                    begin
                      reg1881 <= (8'ha8);
                    end
                  else
                    begin
                      reg1881 <= reg1912;
                      reg1882 <= $signed((-reg1885));
                      reg1883 <= ((reg1938 == ($unsigned(reg1929) ^ (reg1843 * forvar1875))) ?
                          $unsigned(wire1804) : ($signed($unsigned(reg1866)) + ($unsigned(reg1955) ?
                              reg1834 : (~&reg1943))));
                      reg1884 <= reg1909[(3'h7):(3'h4)];
                    end
                end
            end
          else
            begin
              for (forvar1874 = (1'h0); (forvar1874 < (1'h1)); forvar1874 = (forvar1874 + (1'h1)))
                begin
                  for (forvar1875 = (1'h0); (forvar1875 < (2'h3)); forvar1875 = (forvar1875 + (1'h1)))
                    begin
                      reg1876 <= $signed(($signed(reg1920[(3'h7):(3'h5)]) >> $signed((forvar1940 ?
                          reg1832 : forvar1881))));
                    end
                end
              reg1877 <= $signed((~|$signed($unsigned((8'haa)))));
              if (((reg1836 ?
                      $unsigned($unsigned(reg1918)) : forvar1851[(3'h4):(1'h1)]) ?
                  reg1941 : $signed(forvar1855)))
                begin
                  for (forvar1878 = (1'h0); (forvar1878 < (2'h2)); forvar1878 = (forvar1878 + (1'h1)))
                    begin
                      reg1879 <= ((((reg1827 < reg1834) ?
                              forvar1828 : $signed(reg1821)) ?
                          $signed($signed((8'hac))) : $unsigned((reg1874 <= (8'hb1)))) - (~|forvar1822));
                      reg1880 <= $signed($signed(reg1892));
                    end
                  for (forvar1881 = (1'h0); (forvar1881 < (1'h1)); forvar1881 = (forvar1881 + (1'h1)))
                    begin
                      reg1882 <= (forvar1937 <<< reg1873[(4'h9):(4'h8)]);
                      reg1883 <= reg1931;
                      reg1884 <= (($unsigned($signed(forvar1874)) ^ $unsigned($unsigned(reg1829))) ?
                          (reg1880 ?
                              reg1908[(1'h1):(1'h1)] : reg1839) : (reg1952[(1'h0):(1'h0)] >>> (~&$unsigned((8'hb7)))));
                    end
                  reg1885 <= forvar1886[(1'h0):(1'h0)];
                  if ((~|(($signed((8'hb3)) <= forvar1835) >= {$unsigned(forvar1818)})))
                    begin
                      reg1886 <= $signed($unsigned((8'ha0)));
                    end
                  else
                    begin
                      reg1886 <= (8'hb9);
                      reg1887 <= reg1827;
                      reg1888 <= $signed($unsigned((~^{(8'ha9)})));
                    end
                end
              else
                begin
                  if ((reg1831[(3'h5):(2'h3)] ? (+(|{reg1890})) : reg1896))
                    begin
                      reg1878 <= ((8'h9f) * reg1892[(1'h1):(1'h1)]);
                      reg1879 <= reg1950[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1878 <= forvar1936;
                    end
                  if (reg1846[(1'h1):(1'h1)])
                    begin
                      reg1880 <= (reg1930[(2'h2):(2'h2)] * {$signed((+reg1948))});
                      reg1881 <= reg1958;
                    end
                  else
                    begin
                      reg1880 <= reg1930[(2'h2):(1'h0)];
                    end
                end
            end
        end
    end
  assign wire1960 = {(~&(~|$unsigned((8'ha2))))};
  assign wire1961 = (~&((^(|(8'ha3))) <= $unsigned($unsigned(forvar1824))));
  assign wire1962 = reg1874;
  assign wire1963 = (((reg1834 ?
                            $signed(reg1833) : ((8'hab) || reg1885)) == $unsigned({(8'ha7)})) ?
                        $unsigned(reg1887[(1'h0):(1'h0)]) : reg1915);
  assign wire1964 = (reg1872 + $unsigned($signed($signed(reg1926))));
  assign wire1965 = $unsigned((^$unsigned($unsigned(wire1806))));
  always
    @(posedge clk) begin
      for (forvar1966 = (1'h0); (forvar1966 < (1'h0)); forvar1966 = (forvar1966 + (1'h1)))
        begin
          if ($signed(reg1902[(3'h7):(2'h2)]))
            begin
              for (forvar1967 = (1'h0); (forvar1967 < (1'h1)); forvar1967 = (forvar1967 + (1'h1)))
                begin
                  for (forvar1968 = (1'h0); (forvar1968 < (1'h1)); forvar1968 = (forvar1968 + (1'h1)))
                    begin
                      reg1969 <= $signed(reg1820);
                    end
                  for (forvar1970 = (1'h0); (forvar1970 < (2'h3)); forvar1970 = (forvar1970 + (1'h1)))
                    begin
                      reg1971 <= (~&forvar1944[(2'h2):(2'h2)]);
                      reg1972 <= {(wire1963[(3'h5):(2'h3)] < {reg1840[(3'h7):(1'h0)]})};
                    end
                  if (($unsigned($signed({reg1820})) ?
                      (~&{$unsigned(reg1823)}) : $signed($signed($signed(forvar1830)))))
                    begin
                      reg1973 <= ($signed((((8'hb6) < reg1933) & (reg1885 >> reg1848))) ?
                          reg1844[(2'h2):(1'h0)] : $unsigned(reg1905[(4'h9):(2'h3)]));
                      reg1974 <= (reg1897 * $signed($signed(forvar1855)));
                    end
                  else
                    begin
                      reg1973 <= reg1947;
                      reg1974 <= $unsigned((&((reg1954 ^~ reg1837) || $unsigned((8'hb1)))));
                    end
                end
              for (forvar1975 = (1'h0); (forvar1975 < (2'h2)); forvar1975 = (forvar1975 + (1'h1)))
                begin
                  for (forvar1976 = (1'h0); (forvar1976 < (2'h3)); forvar1976 = (forvar1976 + (1'h1)))
                    begin
                      reg1977 <= $signed($signed(wire1960[(2'h2):(1'h1)]));
                    end
                  if (reg1858[(1'h1):(1'h0)])
                    begin
                      reg1978 <= (~reg1919[(3'h5):(3'h4)]);
                      reg1979 <= reg1874;
                      reg1980 <= $unsigned($signed(reg1857[(2'h2):(1'h0)]));
                      reg1981 <= $signed((8'h9e));
                    end
                  else
                    begin
                      reg1978 <= reg1843;
                      reg1979 <= wire1805[(3'h4):(2'h3)];
                      reg1980 <= ($unsigned((-{reg1916})) ~^ $unsigned(({reg1863} >= $unsigned(reg1933))));
                    end
                end
              if ((8'ha7))
                begin
                  for (forvar1982 = (1'h0); (forvar1982 < (2'h3)); forvar1982 = (forvar1982 + (1'h1)))
                    begin
                      reg1983 <= ((+(&$unsigned(forvar1917))) ?
                          $unsigned((~^(~&reg1899))) : (!(8'hba)));
                      reg1984 <= $unsigned((reg1823 ?
                          ((reg1914 ? (8'ha5) : reg1865) ?
                              wire1811 : (reg1840 ^ forvar1879)) : (^(reg1907 - reg1861))));
                      reg1985 <= $unsigned(((~reg1969[(4'he):(3'h7)]) ?
                          $unsigned((8'had)) : {{reg1952}}));
                      reg1986 <= $signed(($unsigned({reg1939}) <<< ((reg1933 ?
                          reg1903 : reg1979) * (!reg1897))));
                    end
                  for (forvar1987 = (1'h0); (forvar1987 < (1'h1)); forvar1987 = (forvar1987 + (1'h1)))
                    begin
                      reg1988 <= $unsigned(((^~$signed(forvar1825)) ?
                          forvar1830[(4'h8):(3'h5)] : (^~reg1863[(3'h4):(1'h1)])));
                      reg1989 <= (~|reg1911);
                      reg1990 <= $signed(reg1839);
                    end
                  if (({(reg1971 ?
                          forvar1956 : $unsigned(forvar1881))} == (8'hb6)))
                    begin
                      reg1991 <= (((&(reg1847 < reg1862)) ?
                              reg1883[(1'h0):(1'h0)] : ($unsigned(reg1945) ~^ (reg1926 * (8'hba)))) ?
                          ($signed($signed(reg1820)) ?
                              reg1950 : forvar1913) : reg1927);
                      reg1992 <= ((-(reg1863[(2'h2):(2'h2)] ?
                              $signed(reg1827) : reg1852[(1'h1):(1'h0)])) ?
                          $signed(reg1934[(2'h2):(1'h1)]) : $signed($unsigned((forvar1895 - reg1850))));
                      reg1993 <= (8'hb4);
                      reg1994 <= forvar1855;
                    end
                  else
                    begin
                      reg1991 <= $unsigned($signed(((reg1931 <<< reg1879) ~^ $signed(reg1977))));
                    end
                end
              else
                begin
                  for (forvar1982 = (1'h0); (forvar1982 < (1'h0)); forvar1982 = (forvar1982 + (1'h1)))
                    begin
                      reg1983 <= forvar1836[(3'h6):(3'h5)];
                      reg1984 <= reg1904[(2'h3):(2'h3)];
                      reg1985 <= reg1854[(1'h1):(1'h1)];
                      reg1986 <= reg1814[(4'h9):(4'h9)];
                    end
                  if ($unsigned((|reg1877)))
                    begin
                      reg1987 <= wire1804[(3'h4):(3'h4)];
                      reg1988 <= forvar1970[(4'ha):(2'h2)];
                    end
                  else
                    begin
                      reg1987 <= {$signed($signed((reg1916 * reg1893)))};
                      reg1988 <= (8'hae);
                    end
                end
            end
          else
            begin
              if (forvar1909)
                begin
                  reg1967 <= reg1969;
                  if ($signed($unsigned(((reg1902 ?
                      reg1921 : reg1883) >>> ((8'ha4) || (8'ha7))))))
                    begin
                      reg1968 <= {(~^reg1980[(4'h8):(3'h4)])};
                      reg1969 <= {{$unsigned($signed(wire1808))}};
                      reg1970 <= (~|($signed(reg1897[(2'h2):(1'h1)]) ?
                          ({reg1993} ?
                              (forvar1944 ?
                                  (8'hb3) : reg1911) : {(8'ha4)}) : (forvar1859 ^~ wire1960[(2'h2):(2'h2)])));
                      reg1971 <= $unsigned($unsigned({(wire1808 ?
                              (8'h9c) : reg1873)}));
                    end
                  else
                    begin
                      reg1968 <= (reg1864 << $signed(reg1974));
                      reg1969 <= $signed((forvar1849[(2'h3):(1'h0)] != ($unsigned(forvar1987) ?
                          forvar1879 : $signed(reg1991))));
                    end
                end
              else
                begin
                  for (forvar1967 = (1'h0); (forvar1967 < (2'h3)); forvar1967 = (forvar1967 + (1'h1)))
                    begin
                      reg1968 <= (($unsigned(reg1954) + $unsigned($signed(reg1968))) ?
                          reg1898 : $unsigned((8'h9e)));
                      reg1969 <= (!$signed($unsigned(reg1884)));
                      reg1970 <= (&(8'hb9));
                      reg1971 <= ((forvar1982 > {$signed((8'hb4))}) || (reg1986[(3'h6):(3'h4)] ?
                          ((reg1839 ? (8'haf) : reg1890) ~^ (reg1929 ?
                              reg1948 : (8'ha5))) : ($signed(reg1886) ^ (forvar1898 << reg1822))));
                    end
                  for (forvar1972 = (1'h0); (forvar1972 < (1'h1)); forvar1972 = (forvar1972 + (1'h1)))
                    begin
                      reg1973 <= (forvar1925 ?
                          (((^~forvar1881) ?
                              reg1886[(2'h3):(2'h2)] : reg1817) ^~ reg1909) : ($signed((reg1902 ?
                              (8'hb3) : forvar1902)) ^~ reg1875[(3'h6):(2'h2)]));
                      reg1974 <= $unsigned(reg1879[(4'h9):(4'h9)]);
                      reg1975 <= $signed(forvar1917[(1'h0):(1'h0)]);
                      reg1976 <= $unsigned($signed(reg1909[(4'h9):(4'h8)]));
                    end
                  reg1977 <= (^~$signed($unsigned((&reg1836))));
                  for (forvar1978 = (1'h0); (forvar1978 < (2'h2)); forvar1978 = (forvar1978 + (1'h1)))
                    begin
                      reg1979 <= {((^~$unsigned(forvar1849)) != ({reg1992} ?
                              (reg1991 ?
                                  wire1812 : (8'ha9)) : $signed((8'hae))))};
                      reg1980 <= $unsigned({(^~reg1881)});
                      reg1981 <= $signed(reg1975[(3'h4):(3'h4)]);
                      reg1982 <= $signed(reg1898);
                    end
                end
            end
          for (forvar1995 = (1'h0); (forvar1995 < (1'h1)); forvar1995 = (forvar1995 + (1'h1)))
            begin
              for (forvar1996 = (1'h0); (forvar1996 < (2'h3)); forvar1996 = (forvar1996 + (1'h1)))
                begin
                  for (forvar1997 = (1'h0); (forvar1997 < (2'h3)); forvar1997 = (forvar1997 + (1'h1)))
                    begin
                      reg1998 <= forvar1987[(4'hb):(1'h1)];
                    end
                  if ((^$unsigned($signed({forvar1877}))))
                    begin
                      reg1999 <= (~&($unsigned($signed(reg1980)) ?
                          reg1871[(3'h7):(2'h3)] : (reg1979 ?
                              $unsigned(forvar1909) : $signed(reg1992))));
                      reg2000 <= $unsigned(forvar1913[(1'h0):(1'h0)]);
                      reg2001 <= $unsigned($unsigned(reg1989));
                    end
                  else
                    begin
                      reg1999 <= ((8'h9c) ?
                          (~|reg1894[(3'h5):(3'h5)]) : $unsigned((^~reg1865[(1'h1):(1'h0)])));
                      reg2000 <= {$signed(((forvar1838 && reg1941) ?
                              reg1979[(1'h1):(1'h1)] : $unsigned(forvar1878)))};
                      reg2001 <= $signed(($signed($unsigned(reg1878)) << {(&reg1883)}));
                    end
                end
            end
          reg2002 <= (~(((reg1887 ?
                  reg1970 : forvar1855) + forvar1855[(1'h0):(1'h0)]) ?
              ($signed((8'haa)) ?
                  $unsigned(reg1859) : $signed(forvar1881)) : forvar1822));
          for (forvar2003 = (1'h0); (forvar2003 < (2'h2)); forvar2003 = (forvar2003 + (1'h1)))
            begin
              for (forvar2004 = (1'h0); (forvar2004 < (1'h1)); forvar2004 = (forvar2004 + (1'h1)))
                begin
                  for (forvar2005 = (1'h0); (forvar2005 < (1'h0)); forvar2005 = (forvar2005 + (1'h1)))
                    begin
                      reg2006 <= (~&reg1926[(2'h2):(2'h2)]);
                      reg2007 <= (~|forvar1940[(4'h8):(4'h8)]);
                      reg2008 <= reg1861[(3'h7):(3'h7)];
                      reg2009 <= reg1931;
                    end
                  for (forvar2010 = (1'h0); (forvar2010 < (2'h2)); forvar2010 = (forvar2010 + (1'h1)))
                    begin
                      reg2011 <= $unsigned((reg1837[(4'h9):(2'h3)] ?
                          $unsigned((reg1998 + reg1863)) : ($signed(reg1821) <<< wire1809)));
                      reg2012 <= (8'hb9);
                      reg2013 <= reg1972[(2'h2):(1'h1)];
                      reg2014 <= forvar1855[(2'h2):(1'h0)];
                    end
                  for (forvar2015 = (1'h0); (forvar2015 < (1'h1)); forvar2015 = (forvar2015 + (1'h1)))
                    begin
                      reg2016 <= ((forvar2004 - $signed($signed(reg1970))) >>> (+((^~reg1899) ?
                          (~forvar1878) : $signed(reg1827))));
                      reg2017 <= ($unsigned($signed(((8'had) <= forvar2010))) ?
                          forvar1982 : reg1838);
                      reg2018 <= reg1933[(1'h0):(1'h0)];
                      reg2019 <= (-$signed((^(-reg1863))));
                    end
                  if (($signed((forvar1940 ?
                      $unsigned(forvar1818) : (reg1901 ?
                          (8'hb8) : reg1903))) <= $unsigned(((+reg1837) ?
                      (8'ha7) : forvar2004))))
                    begin
                      reg2020 <= (forvar1830 ^~ forvar1817);
                      reg2021 <= $unsigned(($signed($unsigned(reg1931)) ?
                          $unsigned({reg1955}) : forvar1881[(2'h3):(2'h2)]));
                      reg2022 <= reg1872;
                    end
                  else
                    begin
                      reg2020 <= ($unsigned((~$unsigned(reg2011))) ?
                          (~|{$unsigned(forvar1976)}) : $unsigned((reg1886 & reg1932)));
                      reg2021 <= (^$unsigned(forvar1821[(4'hb):(4'hb)]));
                    end
                end
              reg2023 <= $unsigned(forvar1966);
              if ($signed($unsigned((8'hae))))
                begin
                  if ($signed(reg1929[(3'h5):(2'h3)]))
                    begin
                      reg2024 <= $unsigned((reg1939 ^ $unsigned((reg1860 ~^ reg1981))));
                      reg2025 <= (~^(^~((!forvar1877) ?
                          reg1818 : {forvar1818})));
                      reg2026 <= $signed($unsigned($unsigned($signed(wire1804))));
                    end
                  else
                    begin
                      reg2024 <= $signed($signed($signed($unsigned(reg1990))));
                      reg2025 <= reg1927;
                    end
                end
              else
                begin
                  if ({reg1974})
                    begin
                      reg2024 <= $unsigned((&$signed({(8'haa)})));
                      reg2025 <= $signed((-reg1881[(2'h3):(2'h2)]));
                    end
                  else
                    begin
                      reg2024 <= ({(8'hba)} ?
                          forvar1849 : {(!$unsigned(reg1915))});
                      reg2025 <= $signed({forvar1818[(3'h4):(1'h0)]});
                      reg2026 <= $unsigned($signed($unsigned($signed(reg1970))));
                      reg2027 <= reg1993;
                    end
                end
              for (forvar2028 = (1'h0); (forvar2028 < (2'h2)); forvar2028 = (forvar2028 + (1'h1)))
                begin
                  for (forvar2029 = (1'h0); (forvar2029 < (1'h1)); forvar2029 = (forvar2029 + (1'h1)))
                    begin
                      reg2030 <= reg1914[(1'h0):(1'h0)];
                      reg2031 <= (((wire1807[(1'h0):(1'h0)] != {reg1871}) ?
                          $unsigned(reg1927[(2'h2):(2'h2)]) : forvar1878) || $signed((reg1827[(1'h1):(1'h0)] ?
                          (|forvar1831) : $unsigned((8'h9d)))));
                    end
                  for (forvar2032 = (1'h0); (forvar2032 < (1'h0)); forvar2032 = (forvar2032 + (1'h1)))
                    begin
                      reg2033 <= ($signed(reg1952[(1'h0):(1'h0)]) & (((reg1893 != forvar1876) ?
                              $unsigned(forvar1849) : $signed(reg1972)) ?
                          forvar1817 : ($signed(reg1908) ?
                              $signed(reg1949) : (^reg1827))));
                      reg2034 <= reg1888;
                    end
                end
            end
        end
      reg2035 <= forvar1867[(2'h3):(2'h3)];
    end
  assign wire2036 = ((reg1826[(3'h5):(2'h3)] + (reg1953 >= (reg1927 ?
                        reg1908 : reg1843))) + {($signed(reg1848) ?
                            $unsigned(reg1919) : $signed((8'ha1)))});
  assign wire2037 = $unsigned(reg1817);
  assign wire2038 = (~&$unsigned($signed(forvar1855)));
  assign wire2039 = forvar1878[(4'h9):(1'h0)];
  always
    @(posedge clk) begin
      for (forvar2040 = (1'h0); (forvar2040 < (2'h2)); forvar2040 = (forvar2040 + (1'h1)))
        begin
          for (forvar2041 = (1'h0); (forvar2041 < (2'h3)); forvar2041 = (forvar2041 + (1'h1)))
            begin
              for (forvar2042 = (1'h0); (forvar2042 < (1'h0)); forvar2042 = (forvar2042 + (1'h1)))
                begin
                  for (forvar2043 = (1'h0); (forvar2043 < (1'h0)); forvar2043 = (forvar2043 + (1'h1)))
                    begin
                      reg2044 <= ($signed((~(reg1992 ?
                          wire1963 : reg2022))) * reg2014[(3'h6):(2'h3)]);
                      reg2045 <= reg1817;
                      reg2046 <= forvar1881[(1'h1):(1'h0)];
                    end
                  reg2047 <= $signed((^((+reg2026) << $unsigned(forvar1975))));
                  if (((^((reg1993 - reg1848) + $signed(wire1810))) > forvar1859[(2'h3):(1'h0)]))
                    begin
                      reg2048 <= {$unsigned($unsigned((reg1987 ?
                              (8'hb4) : reg1976)))};
                      reg2049 <= reg2006;
                      reg2050 <= $signed($unsigned(((reg1922 < reg2049) ^~ $unsigned(reg1871))));
                      reg2051 <= forvar1838;
                    end
                  else
                    begin
                      reg2048 <= (~&(reg1880 && (!$signed(forvar1995))));
                      reg2049 <= ($unsigned(forvar1849) ?
                          $signed(((forvar1823 <<< reg2002) & $unsigned(wire1965))) : reg1992);
                    end
                  for (forvar2052 = (1'h0); (forvar2052 < (1'h0)); forvar2052 = (forvar2052 + (1'h1)))
                    begin
                      reg2053 <= {{($signed(forvar1976) ?
                                  (forvar1881 ?
                                      reg1850 : forvar1919) : (~^reg1893))}};
                      reg2054 <= {reg1892};
                    end
                end
            end
          for (forvar2055 = (1'h0); (forvar2055 < (2'h3)); forvar2055 = (forvar2055 + (1'h1)))
            begin
              if ($signed(reg1929))
                begin
                  for (forvar2056 = (1'h0); (forvar2056 < (1'h1)); forvar2056 = (forvar2056 + (1'h1)))
                    begin
                      reg2057 <= reg1909[(1'h1):(1'h0)];
                      reg2058 <= (&$unsigned($unsigned(forvar2015[(2'h3):(2'h3)])));
                      reg2059 <= $unsigned($unsigned(forvar1972));
                      reg2060 <= reg1817[(2'h3):(2'h2)];
                    end
                  if ((!(reg1837[(3'h4):(2'h3)] ?
                      $unsigned($signed(reg1892)) : wire1810[(4'ha):(4'h8)])))
                    begin
                      reg2061 <= ({{{reg1955}}} ?
                          $signed({(reg1950 ?
                                  wire1807 : (8'h9e))}) : {(forvar1822 >> reg2020[(2'h2):(1'h1)])});
                      reg2062 <= ((reg1881[(4'hb):(4'h9)] ?
                          {reg1949} : reg1990) << reg1826);
                    end
                  else
                    begin
                      reg2061 <= ($unsigned($unsigned((forvar1996 ?
                          (8'ha1) : reg1831))) ^ (forvar1816 | $unsigned(reg1944[(1'h0):(1'h0)])));
                    end
                  for (forvar2063 = (1'h0); (forvar2063 < (1'h1)); forvar2063 = (forvar2063 + (1'h1)))
                    begin
                      reg2064 <= (reg1992 ?
                          ($signed((&reg1987)) >> reg1825[(4'hc):(4'hb)]) : (&($signed(forvar2028) ^~ (^~forvar2043))));
                    end
                  for (forvar2065 = (1'h0); (forvar2065 < (1'h1)); forvar2065 = (forvar2065 + (1'h1)))
                    begin
                      reg2066 <= {(reg2022 <<< reg1975)};
                    end
                end
              else
                begin
                  if (reg2006[(1'h1):(1'h0)])
                    begin
                      reg2056 <= $unsigned(($unsigned(forvar2004[(2'h3):(1'h1)]) ?
                          reg2066 : (-reg1859[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg2056 <= {reg1968[(4'hb):(1'h0)]};
                      reg2057 <= (~{((forvar1978 ?
                              reg1907 : reg1989) ^~ $unsigned((8'hb1)))});
                      reg2058 <= $unsigned(reg2011);
                      reg2059 <= wire1808[(3'h5):(1'h1)];
                    end
                  if (($signed($unsigned(((8'ha7) || reg1897))) ?
                      (~|(+$unsigned(reg1912))) : reg1906))
                    begin
                      reg2060 <= (~|({{forvar1826}} ?
                          ((reg1999 ?
                              (8'h9c) : reg1958) > (-reg1944)) : wire1811[(4'hc):(1'h1)]));
                      reg2061 <= ((((reg1871 ?
                              (8'ha7) : (8'hac)) ^ $signed((8'ha6))) >>> (~reg1901[(2'h2):(2'h2)])) ?
                          ($signed((~&(8'hab))) ?
                              ((reg1954 ? reg1892 : reg1944) ?
                                  (8'had) : $signed(reg1909)) : $unsigned($signed((8'ha4)))) : reg1947);
                      reg2062 <= $unsigned({reg1978});
                      reg2063 <= $unsigned($unsigned((&(reg1852 << reg1994))));
                    end
                  else
                    begin
                      reg2060 <= reg1833;
                    end
                end
              if ($signed((forvar2004 ?
                  ((-reg2001) ?
                      $unsigned(forvar1856) : $signed((8'haf))) : reg1880[(1'h0):(1'h0)])))
                begin
                  reg2067 <= reg2044;
                  reg2068 <= ($unsigned({(forvar2041 ?
                          reg2051 : forvar1970)}) << forvar1835[(1'h1):(1'h0)]);
                  for (forvar2069 = (1'h0); (forvar2069 < (1'h1)); forvar2069 = (forvar2069 + (1'h1)))
                    begin
                      reg2070 <= reg2025;
                      reg2071 <= (-((8'ha1) >= reg1979));
                      reg2072 <= reg1900[(2'h3):(1'h1)];
                      reg2073 <= $signed((+$unsigned((reg1852 > reg1872))));
                    end
                end
              else
                begin
                  if ((~&(reg1838[(3'h6):(2'h3)] + reg1922[(3'h4):(2'h3)])))
                    begin
                      reg2067 <= (~^reg2013[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2067 <= reg1993[(1'h1):(1'h1)];
                      reg2068 <= reg1846;
                      reg2069 <= (forvar1886[(1'h1):(1'h1)] ?
                          (!$unsigned({forvar2029})) : reg2024);
                    end
                  for (forvar2070 = (1'h0); (forvar2070 < (1'h1)); forvar2070 = (forvar2070 + (1'h1)))
                    begin
                      reg2071 <= (+(reg1834 ?
                          (reg1947 ~^ $signed(reg1881)) : reg1883));
                      reg2072 <= (reg1825 <<< (-((reg1990 ~^ reg1948) <= (reg1867 ?
                          (8'ha9) : reg1989))));
                    end
                  for (forvar2073 = (1'h0); (forvar2073 < (1'h1)); forvar2073 = (forvar2073 + (1'h1)))
                    begin
                      reg2074 <= (8'hb0);
                      reg2075 <= $unsigned(forvar1972[(4'hb):(3'h5)]);
                      reg2076 <= $signed(reg1884);
                    end
                end
            end
          for (forvar2077 = (1'h0); (forvar2077 < (1'h1)); forvar2077 = (forvar2077 + (1'h1)))
            begin
              reg2078 <= (((!(forvar1851 ?
                  forvar2004 : reg1827)) && (~&(reg1930 ~^ (8'hac)))) > (reg1904 ?
                  (^~reg2053) : reg1914[(2'h3):(2'h3)]));
            end
          for (forvar2079 = (1'h0); (forvar2079 < (2'h3)); forvar2079 = (forvar2079 + (1'h1)))
            begin
              for (forvar2080 = (1'h0); (forvar2080 < (2'h3)); forvar2080 = (forvar2080 + (1'h1)))
                begin
                  reg2081 <= reg1891[(4'h8):(3'h5)];
                  for (forvar2082 = (1'h0); (forvar2082 < (1'h1)); forvar2082 = (forvar2082 + (1'h1)))
                    begin
                      reg2083 <= {reg1871};
                    end
                  if (((~|reg1826[(2'h3):(2'h3)]) * reg1971))
                    begin
                      reg2084 <= (+$unsigned($unsigned(((8'hb8) ^~ reg2031))));
                      reg2085 <= (|($signed($signed((8'h9f))) >> $unsigned($unsigned(reg1952))));
                      reg2086 <= reg2017[(4'h8):(2'h3)];
                      reg2087 <= $unsigned($signed((reg2044[(3'h5):(3'h4)] ?
                          $unsigned((8'ha5)) : reg1840[(4'hb):(3'h5)])));
                    end
                  else
                    begin
                      reg2084 <= (reg1930 ?
                          $signed($unsigned((wire2037 | wire2036))) : reg2051[(2'h2):(1'h0)]);
                      reg2085 <= $signed({(forvar1917 ?
                              (reg1975 ? reg1894 : reg1822) : (^~reg1827))});
                    end
                  for (forvar2088 = (1'h0); (forvar2088 < (1'h1)); forvar2088 = (forvar2088 + (1'h1)))
                    begin
                      reg2089 <= wire1806;
                      reg2090 <= $signed({(~|(reg1970 ? reg2023 : reg1860))});
                      reg2091 <= $unsigned({(^~$signed(forvar1814))});
                      reg2092 <= ($unsigned(({reg1897} ?
                          (reg1972 >>> reg2019) : $signed(forvar2088))) ^ (~^(reg1819[(3'h6):(3'h4)] <<< (reg2057 ?
                          reg2018 : (8'ha7)))));
                    end
                end
              if ($unsigned(forvar1830[(4'ha):(2'h2)]))
                begin
                  for (forvar2093 = (1'h0); (forvar2093 < (2'h2)); forvar2093 = (forvar2093 + (1'h1)))
                    begin
                      reg2094 <= $signed(($signed((wire1804 ?
                              reg1983 : (8'hb5))) ?
                          forvar1906[(4'h9):(3'h6)] : (~&(wire2036 ?
                              (8'hba) : forvar1816))));
                      reg2095 <= (+(($signed(forvar1940) ?
                              (~|reg1894) : (forvar1828 ? reg1950 : wire1805)) ?
                          $signed((|reg1955)) : (reg2046[(2'h2):(2'h2)] && (|forvar1828))));
                    end
                  for (forvar2096 = (1'h0); (forvar2096 < (1'h1)); forvar2096 = (forvar2096 + (1'h1)))
                    begin
                      reg2097 <= (~&reg1955[(4'hd):(4'hd)]);
                      reg2098 <= $signed(((+{reg1982}) != ({(8'hb2)} ?
                          ((8'haa) != forvar1902) : wire1810)));
                      reg2099 <= $signed((~$unsigned((~&reg2095))));
                      reg2100 <= (reg1952 >= ((~^reg2011[(1'h0):(1'h0)]) ?
                          (~(|(8'haa))) : (forvar1928 == $signed(forvar2032))));
                    end
                  reg2101 <= (!$signed({reg1904}));
                  for (forvar2102 = (1'h0); (forvar2102 < (1'h1)); forvar2102 = (forvar2102 + (1'h1)))
                    begin
                      reg2103 <= {{reg1827[(2'h2):(1'h0)]}};
                      reg2104 <= ((8'hb6) * reg2048[(4'h8):(3'h5)]);
                      reg2105 <= wire1811;
                    end
                end
              else
                begin
                  if ($unsigned(($unsigned(reg2025) ?
                      $signed((8'hb6)) : $signed(forvar1940))))
                    begin
                      reg2093 <= (reg1931[(4'h9):(3'h6)] != reg1914[(1'h1):(1'h1)]);
                      reg2094 <= $unsigned($signed($signed((~|forvar1856))));
                    end
                  else
                    begin
                      reg2093 <= forvar1917;
                      reg2094 <= reg2095;
                    end
                end
            end
        end
      if (reg2007[(2'h2):(2'h2)])
        begin
          for (forvar2106 = (1'h0); (forvar2106 < (1'h0)); forvar2106 = (forvar2106 + (1'h1)))
            begin
              for (forvar2107 = (1'h0); (forvar2107 < (2'h3)); forvar2107 = (forvar2107 + (1'h1)))
                begin
                  reg2108 <= reg1902[(4'hc):(4'hb)];
                  for (forvar2109 = (1'h0); (forvar2109 < (2'h2)); forvar2109 = (forvar2109 + (1'h1)))
                    begin
                      reg2110 <= (~&(reg1926 ?
                          reg1830[(1'h1):(1'h1)] : $signed((forvar2010 ?
                              forvar2069 : reg2030))));
                      reg2111 <= (forvar1925 ~^ ({reg1950[(2'h2):(2'h2)]} ?
                          reg1860 : reg2062[(3'h6):(1'h1)]));
                      reg2112 <= (((~|{forvar2088}) ?
                              reg1826[(2'h2):(1'h1)] : $unsigned((forvar1956 ?
                                  (8'ha5) : reg1977))) ?
                          wire1812[(2'h2):(1'h0)] : (^~$unsigned(reg1819)));
                      reg2113 <= ((((~&reg1994) >> (reg1976 & forvar1824)) ~^ ($unsigned(reg1839) ?
                          (reg2045 ?
                              reg2050 : reg1845) : forvar2003[(2'h2):(1'h1)])) << ({(~reg1941)} <<< reg2054));
                    end
                  for (forvar2114 = (1'h0); (forvar2114 < (1'h1)); forvar2114 = (forvar2114 + (1'h1)))
                    begin
                      reg2115 <= reg1879;
                      reg2116 <= $unsigned($unsigned({reg2081[(3'h7):(3'h4)]}));
                      reg2117 <= $signed((($signed(reg1820) || reg1845[(1'h0):(1'h0)]) && $signed((reg2101 ?
                          reg2046 : reg2045))));
                    end
                  for (forvar2118 = (1'h0); (forvar2118 < (2'h2)); forvar2118 = (forvar2118 + (1'h1)))
                    begin
                      reg2119 <= $unsigned((^~$unsigned({reg1949})));
                      reg2120 <= $signed(((^~$unsigned(wire1813)) ?
                          (!((8'ha5) != reg1830)) : (reg1933[(1'h1):(1'h1)] ^~ $unsigned((8'haf)))));
                    end
                end
              for (forvar2121 = (1'h0); (forvar2121 < (1'h1)); forvar2121 = (forvar2121 + (1'h1)))
                begin
                  reg2122 <= $signed($unsigned(((reg2062 ?
                      reg2033 : (8'hac)) >= reg2067[(2'h3):(1'h1)])));
                  reg2123 <= $signed(reg1981[(2'h2):(1'h1)]);
                  for (forvar2124 = (1'h0); (forvar2124 < (2'h2)); forvar2124 = (forvar2124 + (1'h1)))
                    begin
                      reg2125 <= (~|$signed($signed($unsigned(forvar2003))));
                      reg2126 <= $unsigned($signed($signed((8'hab))));
                    end
                end
              for (forvar2127 = (1'h0); (forvar2127 < (1'h1)); forvar2127 = (forvar2127 + (1'h1)))
                begin
                  reg2128 <= $signed(reg2087);
                  reg2129 <= forvar1940[(1'h0):(1'h0)];
                  reg2130 <= reg2126;
                end
              reg2131 <= $signed(($unsigned($signed((8'ha4))) != forvar1972));
            end
          for (forvar2132 = (1'h0); (forvar2132 < (1'h1)); forvar2132 = (forvar2132 + (1'h1)))
            begin
              for (forvar2133 = (1'h0); (forvar2133 < (1'h0)); forvar2133 = (forvar2133 + (1'h1)))
                begin
                  reg2134 <= (wire2038 <= (~|((8'h9c) ?
                      $unsigned((8'ha9)) : (wire1810 ? reg1909 : reg2120))));
                  reg2135 <= (forvar2118 ?
                      ($unsigned((reg1908 <<< forvar2133)) + (forvar1995[(3'h6):(3'h4)] ?
                          (reg2131 ^~ reg2023) : {forvar2124})) : $unsigned(($unsigned((8'ha0)) ?
                          forvar1931 : forvar1855[(1'h1):(1'h0)])));
                  reg2136 <= (|forvar1851);
                  reg2137 <= (~|reg1922[(3'h7):(3'h7)]);
                end
            end
          for (forvar2138 = (1'h0); (forvar2138 < (1'h0)); forvar2138 = (forvar2138 + (1'h1)))
            begin
              if (($signed(($signed(forvar2138) || forvar1895[(2'h2):(1'h1)])) == (reg1909 ?
                  reg1978[(1'h0):(1'h0)] : ($unsigned(wire1962) >> (8'hac)))))
                begin
                  for (forvar2139 = (1'h0); (forvar2139 < (1'h0)); forvar2139 = (forvar2139 + (1'h1)))
                    begin
                      reg2140 <= $signed(({$unsigned(reg1973)} >> reg2108[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  reg2139 <= (+$unsigned(($signed((8'hb9)) ?
                      ((8'h9f) ? forvar2042 : forvar1886) : (reg2057 ?
                          reg1887 : reg2061))));
                  reg2140 <= forvar2096;
                end
              reg2141 <= forvar2070;
              for (forvar2142 = (1'h0); (forvar2142 < (2'h3)); forvar2142 = (forvar2142 + (1'h1)))
                begin
                  reg2143 <= (~&(reg2089[(1'h1):(1'h1)] || ({forvar1886} >>> $unsigned(reg2067))));
                  for (forvar2144 = (1'h0); (forvar2144 < (2'h3)); forvar2144 = (forvar2144 + (1'h1)))
                    begin
                      reg2145 <= $unsigned((({reg2140} ? {reg2075} : (8'h9f)) ?
                          (^~(reg2007 ?
                              reg1977 : forvar1902)) : (~^$signed(reg1916))));
                      reg2146 <= reg1939[(3'h7):(2'h2)];
                    end
                  if ((!(~$unsigned((reg1825 ? wire2038 : reg1931)))))
                    begin
                      reg2147 <= (^$signed(reg1942[(4'h9):(4'h8)]));
                      reg2148 <= $signed($signed(forvar1851[(3'h6):(3'h6)]));
                      reg2149 <= reg1876[(1'h0):(1'h0)];
                      reg2150 <= (((reg2068 - (reg2110 == reg2071)) <<< (!$signed(reg1836))) ?
                          $unsigned((~&$unsigned(reg2035))) : reg1892);
                    end
                  else
                    begin
                      reg2147 <= (~forvar1940[(4'hd):(3'h7)]);
                      reg2148 <= (&$signed(((^reg2150) ?
                          $unsigned(reg1885) : reg2116)));
                      reg2149 <= ($unsigned($signed({reg2104})) - ($unsigned(reg1983[(4'hd):(3'h4)]) > {$signed((8'hb3))}));
                      reg2150 <= ((reg1981 <<< {(-reg1948)}) == (8'ha0));
                    end
                  if (wire2036)
                    begin
                      reg2151 <= reg1844[(2'h2):(1'h0)];
                      reg2152 <= ((~&(|reg1870)) <<< $unsigned(reg2141));
                    end
                  else
                    begin
                      reg2151 <= (8'had);
                    end
                end
            end
        end
      else
        begin
          reg2106 <= $signed(reg1904[(3'h4):(1'h0)]);
          for (forvar2107 = (1'h0); (forvar2107 < (2'h2)); forvar2107 = (forvar2107 + (1'h1)))
            begin
              if ((~&wire1806))
                begin
                  for (forvar2108 = (1'h0); (forvar2108 < (2'h3)); forvar2108 = (forvar2108 + (1'h1)))
                    begin
                      reg2109 <= (&{{{forvar1997}}});
                    end
                  if ((~^$unsigned($signed(reg2139))))
                    begin
                      reg2110 <= (8'hb1);
                      reg2111 <= {reg1847};
                    end
                  else
                    begin
                      reg2110 <= $signed(forvar2056);
                      reg2111 <= $unsigned(reg1873[(4'h8):(3'h6)]);
                    end
                  reg2112 <= $unsigned((~|forvar1886));
                  for (forvar2113 = (1'h0); (forvar2113 < (1'h0)); forvar2113 = (forvar2113 + (1'h1)))
                    begin
                      reg2114 <= ($unsigned((|(reg1954 > reg1824))) && $unsigned({$unsigned(reg1834)}));
                      reg2115 <= reg1872;
                    end
                end
              else
                begin
                  if ({(($unsigned(reg1949) <<< $unsigned(reg2009)) >= $unsigned((~&reg1982)))})
                    begin
                      reg2108 <= $signed($unsigned(reg1815[(2'h3):(2'h2)]));
                      reg2109 <= (~reg1909[(2'h2):(1'h1)]);
                      reg2110 <= wire2038[(4'h8):(2'h3)];
                    end
                  else
                    begin
                      reg2108 <= ($unsigned(reg1820[(2'h3):(1'h0)]) >> $unsigned(((reg1920 ?
                          reg2076 : forvar2096) - (reg2056 ?
                          reg1887 : reg2113))));
                      reg2109 <= reg2031;
                      reg2110 <= (reg1845 ?
                          ({(~&reg1843)} ?
                              reg2051 : (reg1939 << (|reg2093))) : (reg1860 ?
                              (|reg2094[(2'h3):(1'h0)]) : {(wire1811 ?
                                      (8'ha8) : forvar2132)}));
                    end
                  for (forvar2111 = (1'h0); (forvar2111 < (2'h3)); forvar2111 = (forvar2111 + (1'h1)))
                    begin
                      reg2112 <= (($signed(reg2078) >> $signed(reg2048[(3'h7):(2'h2)])) ?
                          {{$unsigned((8'ha0))}} : (({(8'hb5)} ?
                              forvar2015 : $signed(reg1908)) << reg1922));
                      reg2113 <= $unsigned(reg2139);
                    end
                end
              for (forvar2116 = (1'h0); (forvar2116 < (2'h2)); forvar2116 = (forvar2116 + (1'h1)))
                begin
                  if ((^~$unsigned($signed((|forvar1816)))))
                    begin
                      reg2117 <= (forvar1842[(1'h1):(1'h0)] << (($signed(reg1959) ?
                          reg2071 : $signed(reg2047)) | $unsigned({reg2147})));
                      reg2118 <= ((reg2147[(1'h1):(1'h1)] ?
                              forvar2093 : reg2148) ?
                          {reg1857[(2'h2):(1'h1)]} : (&(wire2037[(4'h9):(3'h7)] >>> forvar1875)));
                      reg2119 <= $signed(($signed(reg2054[(1'h0):(1'h0)]) << ((reg1897 && reg1970) ?
                          (~&reg2021) : $unsigned(reg2024))));
                      reg2120 <= ((reg1832 | {(~&reg1908)}) ?
                          $unsigned(({forvar1857} ?
                              reg1873 : $signed(forvar2139))) : ((&$unsigned((8'hba))) ?
                              $signed((forvar1928 < reg2113)) : ((~&reg2008) ?
                                  forvar1987 : reg1817[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg2117 <= reg1958;
                    end
                  for (forvar2121 = (1'h0); (forvar2121 < (1'h1)); forvar2121 = (forvar2121 + (1'h1)))
                    begin
                      reg2122 <= reg1846[(1'h1):(1'h0)];
                      reg2123 <= (($unsigned(reg1991[(1'h0):(1'h0)]) ?
                              $unsigned($unsigned((8'hb9))) : ((reg2053 > reg2026) ?
                                  (reg2084 ? reg2051 : reg1923) : {reg2044})) ?
                          forvar2108 : (~|$signed(reg1986[(2'h3):(1'h1)])));
                    end
                  if (((forvar2142[(1'h0):(1'h0)] - $unsigned(reg1893)) & ($unsigned((forvar1987 ~^ reg1823)) <= ($unsigned(reg1887) ?
                      (~|forvar2070) : forvar2111[(1'h1):(1'h0)]))))
                    begin
                      reg2124 <= {(&$unsigned(((8'hb1) ?
                              forvar2096 : reg2075)))};
                      reg2125 <= $unsigned($signed((&(reg2099 ?
                          forvar2102 : reg1904))));
                    end
                  else
                    begin
                      reg2124 <= ((&(^$signed(reg1860))) || ((&(forvar2070 ^~ forvar2139)) != (reg1838[(3'h6):(3'h6)] & (forvar2096 >> reg1971))));
                      reg2125 <= (|((~|{forvar1821}) == {reg2072[(3'h4):(1'h1)]}));
                      reg2126 <= (reg1821[(4'hc):(3'h5)] ?
                          reg1893 : {reg1934[(1'h0):(1'h0)]});
                      reg2127 <= reg2139[(3'h6):(1'h1)];
                    end
                end
              for (forvar2128 = (1'h0); (forvar2128 < (2'h2)); forvar2128 = (forvar2128 + (1'h1)))
                begin
                  for (forvar2129 = (1'h0); (forvar2129 < (1'h0)); forvar2129 = (forvar2129 + (1'h1)))
                    begin
                      reg2130 <= $signed($signed({(forvar2139 == wire2037)}));
                      reg2131 <= reg2135;
                    end
                  if ((~&(({reg1821} || (reg1822 >= reg1845)) > $signed(reg2002[(1'h0):(1'h0)]))))
                    begin
                      reg2132 <= $unsigned((&(((8'ha4) ?
                          forvar2138 : reg2112) >> $unsigned(reg2140))));
                      reg2133 <= ({$unsigned(reg1988[(1'h0):(1'h0)])} ?
                          $unsigned((|wire1963)) : reg1867[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2132 <= (~&$unsigned({reg1867}));
                      reg2133 <= $unsigned(reg2008);
                    end
                  for (forvar2134 = (1'h0); (forvar2134 < (2'h3)); forvar2134 = (forvar2134 + (1'h1)))
                    begin
                      reg2135 <= (-$unsigned(((reg1899 ^~ reg1904) < reg1846[(2'h2):(1'h0)])));
                      reg2136 <= (($signed((reg1916 ?
                              reg2150 : reg1888)) * (~&$unsigned(reg2075))) ?
                          ($unsigned({reg1999}) ^ (reg2136[(3'h4):(1'h0)] > reg2017)) : $signed(($unsigned(reg2056) ~^ reg1976[(2'h3):(1'h0)])));
                      reg2137 <= forvar2138[(2'h2):(1'h1)];
                    end
                  for (forvar2138 = (1'h0); (forvar2138 < (1'h0)); forvar2138 = (forvar2138 + (1'h1)))
                    begin
                      reg2139 <= ((|(~^(reg1877 ?
                          reg2143 : (8'hb3)))) ^ $unsigned(forvar1825));
                      reg2140 <= reg2045;
                    end
                end
            end
        end
      reg2153 <= $signed((8'hb0));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2225
#(parameter param3109 = (~{((-(8'hac)) << ((8'h9f) ? (8'ha8) : (8'h9f)))}))
(y, clk, wire2229, wire2228, wire2227, wire2226);
  output wire [(32'h9d1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire2229;
  input wire signed [(3'h6):(1'h0)] wire2228;
  input wire [(4'hd):(1'h0)] wire2227;
  input wire [(4'ha):(1'h0)] wire2226;
  reg [(2'h3):(1'h0)] reg3108 = (1'h0);
  reg [(2'h3):(1'h0)] reg3107 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3078 = (1'h0);
  reg [(4'hb):(1'h0)] reg3081 = (1'h0);
  reg [(4'he):(1'h0)] forvar3094 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3088 = (1'h0);
  reg [(4'ha):(1'h0)] reg3084 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3083 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3082 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3080 = (1'h0);
  reg [(3'h7):(1'h0)] reg3106 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3105 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3104 = (1'h0);
  reg [(4'h8):(1'h0)] reg3103 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3102 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3101 = (1'h0);
  reg [(2'h3):(1'h0)] reg3100 = (1'h0);
  reg [(4'he):(1'h0)] reg3099 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3098 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3097 = (1'h0);
  reg [(4'hd):(1'h0)] reg3096 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3095 = (1'h0);
  reg [(4'he):(1'h0)] reg3094 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3093 = (1'h0);
  reg [(3'h6):(1'h0)] reg3092 = (1'h0);
  reg [(3'h7):(1'h0)] reg3091 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3090 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3089 = (1'h0);
  reg [(4'ha):(1'h0)] reg3088 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3087 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3086 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3085 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3084 = (1'h0);
  reg [(4'hd):(1'h0)] reg3083 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3082 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3081 = (1'h0);
  reg [(4'he):(1'h0)] reg3080 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3079 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3072 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3071 = (1'h0);
  reg [(2'h3):(1'h0)] reg3073 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3070 = (1'h0);
  reg [(3'h4):(1'h0)] reg3078 = (1'h0);
  reg [(2'h2):(1'h0)] reg3077 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3076 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3075 = (1'h0);
  reg [(5'h10):(1'h0)] reg3074 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3073 = (1'h0);
  reg [(4'hb):(1'h0)] reg3072 = (1'h0);
  reg [(4'hf):(1'h0)] reg3071 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3070 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3069 = (1'h0);
  reg [(4'hd):(1'h0)] reg3068 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3067 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3066 = (1'h0);
  reg [(2'h2):(1'h0)] reg3065 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3061 = (1'h0);
  reg [(3'h4):(1'h0)] reg3064 = (1'h0);
  reg [(4'hf):(1'h0)] reg3063 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3062 = (1'h0);
  reg [(4'hc):(1'h0)] reg3061 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3060 = (1'h0);
  reg [(2'h3):(1'h0)] reg3059 = (1'h0);
  reg [(4'h9):(1'h0)] reg3058 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3057 = (1'h0);
  reg [(4'hd):(1'h0)] reg3056 = (1'h0);
  reg [(3'h5):(1'h0)] reg3055 = (1'h0);
  reg [(4'hb):(1'h0)] reg3054 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3053 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3052 = (1'h0);
  reg [(4'he):(1'h0)] reg3051 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3050 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3049 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3048 = (1'h0);
  reg [(4'he):(1'h0)] forvar3047 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3046 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3045 = (1'h0);
  reg [(4'hd):(1'h0)] reg3044 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3043 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3042 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3041 = (1'h0);
  reg [(3'h7):(1'h0)] reg3040 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3039 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3038 = (1'h0);
  reg [(4'ha):(1'h0)] reg3037 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3036 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3035 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3034 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3029 = (1'h0);
  reg [(4'hc):(1'h0)] reg3028 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3026 = (1'h0);
  reg [(4'hf):(1'h0)] reg3024 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3023 = (1'h0);
  reg [(4'hf):(1'h0)] reg3033 = (1'h0);
  reg [(4'h8):(1'h0)] reg3032 = (1'h0);
  reg [(4'he):(1'h0)] reg3031 = (1'h0);
  reg [(4'h8):(1'h0)] reg3030 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3029 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3028 = (1'h0);
  reg [(4'hc):(1'h0)] reg3027 = (1'h0);
  reg [(4'ha):(1'h0)] reg3026 = (1'h0);
  reg [(3'h6):(1'h0)] reg3025 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3024 = (1'h0);
  reg [(4'hf):(1'h0)] reg3023 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3022 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3021 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire3020;
  wire signed [(4'hd):(1'h0)] wire3019;
  wire signed [(4'ha):(1'h0)] wire3018;
  wire signed [(4'hf):(1'h0)] wire3017;
  wire [(3'h4):(1'h0)] wire3016;
  wire signed [(4'hc):(1'h0)] wire3014;
  reg [(4'h9):(1'h0)] reg2352 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2351 = (1'h0);
  reg [(4'hd):(1'h0)] reg2350 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2347 = (1'h0);
  reg [(2'h2):(1'h0)] reg2344 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2339 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2335 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2334 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2332 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2366 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2365 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2364 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2363 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2362 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2361 = (1'h0);
  reg [(4'hf):(1'h0)] reg2360 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2359 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2357 = (1'h0);
  reg [(4'hc):(1'h0)] reg2356 = (1'h0);
  reg [(2'h3):(1'h0)] reg2355 = (1'h0);
  reg [(3'h7):(1'h0)] reg2354 = (1'h0);
  reg [(3'h4):(1'h0)] reg2353 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2352 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2351 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2350 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2349 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2348 = (1'h0);
  reg [(3'h7):(1'h0)] reg2347 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2346 = (1'h0);
  reg [(4'he):(1'h0)] reg2345 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2344 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2343 = (1'h0);
  reg [(3'h5):(1'h0)] reg2341 = (1'h0);
  reg [(4'h8):(1'h0)] reg2342 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2341 = (1'h0);
  reg [(4'ha):(1'h0)] reg2340 = (1'h0);
  reg [(3'h5):(1'h0)] reg2339 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2338 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2337 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2336 = (1'h0);
  reg [(3'h4):(1'h0)] reg2335 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2334 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2333 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2332 = (1'h0);
  reg [(4'ha):(1'h0)] reg2320 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2314 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2331 = (1'h0);
  reg [(4'he):(1'h0)] forvar2330 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2329 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2328 = (1'h0);
  reg [(4'ha):(1'h0)] reg2327 = (1'h0);
  reg [(2'h2):(1'h0)] reg2326 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2325 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2324 = (1'h0);
  reg [(2'h2):(1'h0)] reg2323 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2322 = (1'h0);
  reg [(4'hc):(1'h0)] reg2321 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2320 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2319 = (1'h0);
  reg [(4'ha):(1'h0)] reg2318 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2317 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2316 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2315 = (1'h0);
  reg [(5'h10):(1'h0)] reg2314 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2313 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2312 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2305 = (1'h0);
  reg [(4'hb):(1'h0)] reg2311 = (1'h0);
  reg [(4'he):(1'h0)] reg2310 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2309 = (1'h0);
  reg [(2'h3):(1'h0)] reg2308 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2302 = (1'h0);
  reg [(4'hd):(1'h0)] reg2301 = (1'h0);
  reg [(4'h8):(1'h0)] reg2307 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2306 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2305 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2304 = (1'h0);
  reg [(4'hd):(1'h0)] reg2303 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2302 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2301 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2300 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2253 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2257 = (1'h0);
  reg [(4'he):(1'h0)] forvar2249 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2248 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2296 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2291 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2290 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2299 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2298 = (1'h0);
  reg [(4'hd):(1'h0)] reg2297 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2296 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2295 = (1'h0);
  reg [(4'h9):(1'h0)] reg2294 = (1'h0);
  reg [(4'h8):(1'h0)] reg2293 = (1'h0);
  reg [(4'h8):(1'h0)] reg2292 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2291 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2290 = (1'h0);
  reg [(2'h2):(1'h0)] reg2289 = (1'h0);
  reg [(2'h2):(1'h0)] reg2288 = (1'h0);
  reg [(5'h10):(1'h0)] reg2287 = (1'h0);
  reg [(4'ha):(1'h0)] reg2286 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2285 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2282 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2281 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2277 = (1'h0);
  reg [(3'h6):(1'h0)] reg2284 = (1'h0);
  reg [(4'hf):(1'h0)] reg2283 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2282 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2281 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2280 = (1'h0);
  reg [(2'h2):(1'h0)] reg2279 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2278 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2277 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2276 = (1'h0);
  reg [(3'h6):(1'h0)] reg2275 = (1'h0);
  reg [(4'he):(1'h0)] reg2274 = (1'h0);
  reg [(4'hd):(1'h0)] reg2273 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2272 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2271 = (1'h0);
  reg [(3'h5):(1'h0)] reg2270 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2269 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2268 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2267 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2266 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2265 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2264 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2263 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2262 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2261 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2250 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2246 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2260 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2259 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2258 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2257 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2256 = (1'h0);
  reg [(4'ha):(1'h0)] reg2255 = (1'h0);
  reg [(4'hf):(1'h0)] reg2254 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2253 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2252 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2251 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2250 = (1'h0);
  reg [(2'h3):(1'h0)] reg2249 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2248 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2247 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2246 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2245 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2244 = (1'h0);
  reg [(2'h3):(1'h0)] reg2243 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2242 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2241 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2240 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2239 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2238 = (1'h0);
  reg [(2'h3):(1'h0)] reg2237 = (1'h0);
  reg [(2'h3):(1'h0)] reg2236 = (1'h0);
  reg [(3'h5):(1'h0)] reg2235 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2234 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2233 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2232 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2231 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2230 = (1'h0);
  assign y = {reg3108,
                 reg3107,
                 forvar3078,
                 reg3081,
                 forvar3094,
                 forvar3088,
                 reg3084,
                 forvar3083,
                 reg3082,
                 forvar3080,
                 reg3106,
                 reg3105,
                 forvar3104,
                 reg3103,
                 reg3102,
                 reg3101,
                 reg3100,
                 reg3099,
                 reg3098,
                 forvar3097,
                 reg3096,
                 reg3095,
                 reg3094,
                 reg3093,
                 reg3092,
                 reg3091,
                 reg3090,
                 forvar3089,
                 reg3088,
                 reg3087,
                 reg3086,
                 reg3085,
                 forvar3084,
                 reg3083,
                 forvar3082,
                 forvar3081,
                 reg3080,
                 reg3079,
                 forvar3072,
                 forvar3071,
                 reg3073,
                 reg3070,
                 reg3078,
                 reg3077,
                 reg3076,
                 reg3075,
                 reg3074,
                 forvar3073,
                 reg3072,
                 reg3071,
                 forvar3070,
                 reg3069,
                 reg3068,
                 reg3067,
                 forvar3066,
                 reg3065,
                 forvar3061,
                 reg3064,
                 reg3063,
                 reg3062,
                 reg3061,
                 reg3060,
                 reg3059,
                 reg3058,
                 reg3057,
                 reg3056,
                 reg3055,
                 reg3054,
                 reg3053,
                 reg3052,
                 reg3051,
                 reg3050,
                 forvar3049,
                 forvar3048,
                 forvar3047,
                 reg3046,
                 reg3045,
                 reg3044,
                 reg3043,
                 forvar3042,
                 reg3041,
                 reg3040,
                 reg3039,
                 forvar3038,
                 reg3037,
                 reg3036,
                 reg3035,
                 forvar3034,
                 forvar3029,
                 reg3028,
                 forvar3026,
                 reg3024,
                 forvar3023,
                 reg3033,
                 reg3032,
                 reg3031,
                 reg3030,
                 reg3029,
                 forvar3028,
                 reg3027,
                 reg3026,
                 reg3025,
                 forvar3024,
                 reg3023,
                 forvar3022,
                 reg3021,
                 wire3020,
                 wire3019,
                 wire3018,
                 wire3017,
                 wire3016,
                 wire3014,
                 reg2352,
                 reg2351,
                 reg2350,
                 forvar2347,
                 reg2344,
                 forvar2339,
                 forvar2335,
                 forvar2334,
                 reg2332,
                 reg2366,
                 reg2365,
                 reg2364,
                 reg2363,
                 reg2362,
                 reg2361,
                 reg2360,
                 reg2359,
                 reg2358,
                 reg2357,
                 reg2356,
                 reg2355,
                 reg2354,
                 reg2353,
                 forvar2352,
                 forvar2351,
                 forvar2350,
                 reg2349,
                 reg2348,
                 reg2347,
                 reg2346,
                 reg2345,
                 forvar2344,
                 reg2343,
                 reg2341,
                 reg2342,
                 forvar2341,
                 reg2340,
                 reg2339,
                 reg2338,
                 reg2337,
                 reg2336,
                 reg2335,
                 reg2334,
                 forvar2333,
                 forvar2332,
                 reg2320,
                 forvar2314,
                 reg2331,
                 forvar2330,
                 reg2329,
                 reg2328,
                 reg2327,
                 reg2326,
                 reg2325,
                 reg2324,
                 reg2323,
                 reg2322,
                 reg2321,
                 forvar2320,
                 forvar2319,
                 reg2318,
                 reg2317,
                 reg2316,
                 reg2315,
                 reg2314,
                 forvar2313,
                 reg2312,
                 reg2305,
                 reg2311,
                 reg2310,
                 reg2309,
                 reg2308,
                 forvar2302,
                 reg2301,
                 reg2307,
                 reg2306,
                 forvar2305,
                 reg2304,
                 reg2303,
                 reg2302,
                 forvar2301,
                 forvar2300,
                 reg2253,
                 reg2257,
                 forvar2249,
                 forvar2248,
                 reg2296,
                 reg2291,
                 forvar2290,
                 reg2299,
                 reg2298,
                 reg2297,
                 forvar2296,
                 reg2295,
                 reg2294,
                 reg2293,
                 reg2292,
                 forvar2291,
                 reg2290,
                 reg2289,
                 reg2288,
                 reg2287,
                 reg2286,
                 forvar2285,
                 reg2282,
                 forvar2281,
                 forvar2277,
                 reg2284,
                 reg2283,
                 forvar2282,
                 reg2281,
                 reg2280,
                 reg2279,
                 reg2278,
                 reg2277,
                 reg2276,
                 reg2275,
                 reg2274,
                 reg2273,
                 reg2272,
                 forvar2271,
                 reg2270,
                 reg2269,
                 reg2268,
                 reg2267,
                 forvar2266,
                 reg2265,
                 reg2264,
                 reg2263,
                 forvar2262,
                 forvar2261,
                 reg2250,
                 forvar2246,
                 reg2260,
                 reg2259,
                 reg2258,
                 forvar2257,
                 reg2256,
                 reg2255,
                 reg2254,
                 forvar2253,
                 reg2252,
                 reg2251,
                 forvar2250,
                 reg2249,
                 reg2248,
                 reg2247,
                 reg2246,
                 forvar2245,
                 reg2244,
                 reg2243,
                 reg2242,
                 forvar2241,
                 forvar2240,
                 reg2239,
                 reg2238,
                 reg2237,
                 reg2236,
                 reg2235,
                 reg2234,
                 forvar2233,
                 forvar2232,
                 forvar2231,
                 forvar2230,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar2230 = (1'h0); (forvar2230 < (1'h1)); forvar2230 = (forvar2230 + (1'h1)))
        begin
          for (forvar2231 = (1'h0); (forvar2231 < (1'h0)); forvar2231 = (forvar2231 + (1'h1)))
            begin
              for (forvar2232 = (1'h0); (forvar2232 < (2'h3)); forvar2232 = (forvar2232 + (1'h1)))
                begin
                  for (forvar2233 = (1'h0); (forvar2233 < (1'h0)); forvar2233 = (forvar2233 + (1'h1)))
                    begin
                      reg2234 <= ((~&forvar2233) ?
                          (&wire2226[(3'h4):(2'h3)]) : wire2228[(2'h2):(2'h2)]);
                    end
                  if (forvar2231[(2'h3):(1'h0)])
                    begin
                      reg2235 <= $signed(forvar2233);
                      reg2236 <= $unsigned(reg2234);
                    end
                  else
                    begin
                      reg2235 <= $unsigned(reg2235);
                      reg2236 <= (($unsigned((+wire2228)) ?
                              ((wire2229 >= reg2235) ?
                                  (^forvar2232) : $unsigned(wire2229)) : wire2227) ?
                          {forvar2230[(5'h10):(4'hd)]} : ({(~&wire2229)} && wire2228[(2'h3):(2'h2)]));
                      reg2237 <= $unsigned((reg2235[(2'h3):(2'h2)] ^ ((!(8'ha9)) ?
                          $signed(wire2227) : (8'hb8))));
                      reg2238 <= $signed(forvar2230);
                    end
                  reg2239 <= $unsigned(((+(reg2235 - (8'hb1))) ?
                      $unsigned($signed(forvar2231)) : wire2226[(4'h8):(3'h6)]));
                end
              for (forvar2240 = (1'h0); (forvar2240 < (1'h1)); forvar2240 = (forvar2240 + (1'h1)))
                begin
                  for (forvar2241 = (1'h0); (forvar2241 < (2'h2)); forvar2241 = (forvar2241 + (1'h1)))
                    begin
                      reg2242 <= wire2226[(3'h7):(2'h2)];
                      reg2243 <= $signed(reg2238[(2'h2):(2'h2)]);
                    end
                  reg2244 <= {(forvar2240 != (~|(forvar2233 ?
                          (8'h9d) : wire2228)))};
                end
            end
        end
      if ((!(~&{(reg2235 ? (8'hb7) : reg2243)})))
        begin
          if (({(reg2243[(2'h3):(2'h3)] ?
                      {reg2242} : wire2227[(4'hc):(1'h1)])} ?
              reg2244 : forvar2231[(1'h0):(1'h0)]))
            begin
              for (forvar2245 = (1'h0); (forvar2245 < (2'h2)); forvar2245 = (forvar2245 + (1'h1)))
                begin
                  if ((~forvar2240[(3'h5):(3'h5)]))
                    begin
                      reg2246 <= wire2228[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg2246 <= $unsigned({reg2234[(2'h2):(2'h2)]});
                      reg2247 <= $unsigned($signed($signed(((8'hac) - (8'ha2)))));
                      reg2248 <= {(reg2246 ?
                              reg2236[(1'h1):(1'h0)] : (&$unsigned(forvar2233)))};
                      reg2249 <= reg2248[(3'h4):(3'h4)];
                    end
                  for (forvar2250 = (1'h0); (forvar2250 < (2'h2)); forvar2250 = (forvar2250 + (1'h1)))
                    begin
                      reg2251 <= forvar2233[(3'h4):(1'h1)];
                      reg2252 <= $unsigned(wire2228);
                    end
                  for (forvar2253 = (1'h0); (forvar2253 < (2'h3)); forvar2253 = (forvar2253 + (1'h1)))
                    begin
                      reg2254 <= $signed((~|$unsigned((!reg2239))));
                      reg2255 <= wire2229[(3'h5):(1'h0)];
                      reg2256 <= (reg2251 ? wire2226 : reg2244);
                    end
                  for (forvar2257 = (1'h0); (forvar2257 < (2'h2)); forvar2257 = (forvar2257 + (1'h1)))
                    begin
                      reg2258 <= $signed($unsigned($signed((!reg2242))));
                      reg2259 <= $signed(wire2228);
                      reg2260 <= forvar2231;
                    end
                end
            end
          else
            begin
              for (forvar2245 = (1'h0); (forvar2245 < (1'h0)); forvar2245 = (forvar2245 + (1'h1)))
                begin
                  for (forvar2246 = (1'h0); (forvar2246 < (2'h2)); forvar2246 = (forvar2246 + (1'h1)))
                    begin
                      reg2247 <= $unsigned(($signed($unsigned(reg2259)) < (8'hac)));
                      reg2248 <= forvar2245[(4'ha):(3'h4)];
                      reg2249 <= $unsigned($unsigned($unsigned((+(8'ha7)))));
                    end
                  if (forvar2240)
                    begin
                      reg2250 <= (~&$unsigned(reg2259[(4'ha):(2'h3)]));
                    end
                  else
                    begin
                      reg2250 <= reg2249[(2'h2):(1'h1)];
                      reg2251 <= reg2234;
                      reg2252 <= {$signed($unsigned((reg2238 ?
                              reg2238 : reg2256)))};
                    end
                  for (forvar2253 = (1'h0); (forvar2253 < (1'h1)); forvar2253 = (forvar2253 + (1'h1)))
                    begin
                      reg2254 <= ($unsigned((~&(~^forvar2257))) & (forvar2232 ?
                          $unsigned((^forvar2246)) : $signed($signed((8'h9f)))));
                      reg2255 <= ((wire2226 != ((-wire2229) >= (wire2226 && wire2229))) < (8'haa));
                      reg2256 <= reg2258;
                    end
                  for (forvar2257 = (1'h0); (forvar2257 < (1'h0)); forvar2257 = (forvar2257 + (1'h1)))
                    begin
                      reg2258 <= ((!(|(reg2239 > reg2256))) + (~|({reg2246} >> reg2256)));
                      reg2259 <= forvar2240;
                      reg2260 <= reg2252[(3'h4):(3'h4)];
                    end
                end
              for (forvar2261 = (1'h0); (forvar2261 < (2'h3)); forvar2261 = (forvar2261 + (1'h1)))
                begin
                  for (forvar2262 = (1'h0); (forvar2262 < (1'h0)); forvar2262 = (forvar2262 + (1'h1)))
                    begin
                      reg2263 <= (~^reg2256[(4'h9):(3'h6)]);
                      reg2264 <= $signed({((wire2227 ? (8'h9e) : forvar2240) ?
                              reg2244[(4'h9):(4'h9)] : (reg2246 <= reg2247))});
                      reg2265 <= (8'hab);
                    end
                  for (forvar2266 = (1'h0); (forvar2266 < (1'h0)); forvar2266 = (forvar2266 + (1'h1)))
                    begin
                      reg2267 <= forvar2246[(4'hc):(1'h1)];
                      reg2268 <= reg2267;
                      reg2269 <= ((forvar2232 * (^~forvar2257)) * ($unsigned(reg2247) ?
                          $unsigned(reg2252[(2'h3):(1'h1)]) : forvar2245));
                      reg2270 <= ($unsigned((&(+(8'hb1)))) + wire2229);
                    end
                  for (forvar2271 = (1'h0); (forvar2271 < (1'h0)); forvar2271 = (forvar2271 + (1'h1)))
                    begin
                      reg2272 <= $unsigned({reg2270[(1'h1):(1'h1)]});
                      reg2273 <= forvar2253[(2'h2):(1'h0)];
                      reg2274 <= $unsigned($unsigned(((8'ha0) ^~ (~&forvar2261))));
                      reg2275 <= ((~^$unsigned((reg2260 ?
                              reg2259 : forvar2240))) ?
                          reg2239 : $signed($signed(forvar2245)));
                    end
                  reg2276 <= (~|$signed((8'ha2)));
                end
              if ({((~^(~&reg2268)) | ($unsigned(forvar2271) ?
                      reg2235[(3'h4):(1'h0)] : forvar2230))})
                begin
                  reg2277 <= reg2259[(4'hc):(2'h2)];
                  if ((((^~$signed((8'hb1))) * (~^(+reg2236))) & reg2236[(2'h2):(1'h0)]))
                    begin
                      reg2278 <= $signed((8'h9f));
                    end
                  else
                    begin
                      reg2278 <= (^~$signed((reg2243 * $unsigned(forvar2253))));
                    end
                  if (reg2273)
                    begin
                      reg2279 <= (((&wire2227) ?
                          reg2276[(4'h9):(3'h5)] : $signed({wire2229})) && reg2260);
                      reg2280 <= ($signed(reg2269) != wire2228);
                      reg2281 <= $signed($unsigned((-(reg2256 ?
                          wire2228 : reg2249))));
                    end
                  else
                    begin
                      reg2279 <= $signed(({(+forvar2245)} ?
                          reg2236 : $signed($unsigned((8'hb7)))));
                      reg2280 <= reg2259[(3'h4):(1'h1)];
                      reg2281 <= $signed(((^(reg2273 & reg2264)) ?
                          (~^(reg2276 ? reg2236 : reg2267)) : ((forvar2246 ?
                                  reg2236 : forvar2241) ?
                              {forvar2241} : (~forvar2253))));
                    end
                  for (forvar2282 = (1'h0); (forvar2282 < (2'h3)); forvar2282 = (forvar2282 + (1'h1)))
                    begin
                      reg2283 <= $signed((|($signed(reg2268) < reg2234)));
                      reg2284 <= (forvar2261 || forvar2230[(4'ha):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar2277 = (1'h0); (forvar2277 < (1'h1)); forvar2277 = (forvar2277 + (1'h1)))
                    begin
                      reg2278 <= {(~^(wire2226 ? {(8'h9d)} : forvar2253))};
                      reg2279 <= ((~forvar2246[(4'hc):(3'h5)]) >>> (^reg2234[(3'h5):(2'h2)]));
                    end
                  reg2280 <= (&reg2280);
                  for (forvar2281 = (1'h0); (forvar2281 < (2'h3)); forvar2281 = (forvar2281 + (1'h1)))
                    begin
                      reg2282 <= (8'ha0);
                    end
                end
            end
          for (forvar2285 = (1'h0); (forvar2285 < (1'h0)); forvar2285 = (forvar2285 + (1'h1)))
            begin
              reg2286 <= {($signed($unsigned(reg2265)) + (8'hb2))};
              if (($unsigned((-(reg2286 ? forvar2233 : reg2249))) ?
                  ($signed((&reg2277)) < reg2250[(2'h2):(1'h1)]) : (+$unsigned($signed(forvar2282)))))
                begin
                  if ((+reg2279[(2'h2):(1'h1)]))
                    begin
                      reg2287 <= wire2228[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2287 <= $signed(reg2269[(3'h6):(1'h1)]);
                      reg2288 <= $unsigned(({(reg2264 ? reg2234 : (8'ha1))} ?
                          reg2243 : (~^forvar2231)));
                    end
                  if (reg2234)
                    begin
                      reg2289 <= ((+$signed((forvar2246 ?
                          reg2286 : forvar2266))) ~^ (((forvar2257 ?
                          wire2226 : (8'h9e)) > $unsigned((8'h9c))) << $signed($signed(reg2259))));
                      reg2290 <= $signed((((forvar2240 * forvar2277) ?
                              wire2227 : (^(8'ha5))) ?
                          $unsigned(((8'h9e) == reg2275)) : $unsigned((forvar2241 ?
                              wire2228 : forvar2230))));
                    end
                  else
                    begin
                      reg2289 <= (reg2256[(2'h3):(2'h2)] ~^ reg2286);
                      reg2290 <= reg2276[(4'ha):(1'h1)];
                    end
                  for (forvar2291 = (1'h0); (forvar2291 < (1'h1)); forvar2291 = (forvar2291 + (1'h1)))
                    begin
                      reg2292 <= (8'ha8);
                      reg2293 <= (reg2272 ^~ $signed(reg2236[(2'h2):(1'h1)]));
                      reg2294 <= forvar2271[(3'h4):(2'h2)];
                      reg2295 <= reg2254[(4'h8):(1'h1)];
                    end
                  for (forvar2296 = (1'h0); (forvar2296 < (1'h0)); forvar2296 = (forvar2296 + (1'h1)))
                    begin
                      reg2297 <= (+$signed(($unsigned(reg2238) ?
                          reg2238 : $signed(reg2277))));
                      reg2298 <= {(|((forvar2285 - reg2284) | (^~reg2276)))};
                      reg2299 <= reg2297[(4'hd):(2'h2)];
                    end
                end
              else
                begin
                  if (reg2246)
                    begin
                      reg2287 <= reg2264[(1'h1):(1'h0)];
                      reg2288 <= $signed(reg2298[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg2287 <= ((8'hb9) >> (~^((reg2270 ?
                          reg2294 : wire2226) - reg2292[(2'h3):(1'h0)])));
                      reg2288 <= reg2252;
                      reg2289 <= wire2228[(2'h3):(2'h3)];
                    end
                  for (forvar2290 = (1'h0); (forvar2290 < (2'h3)); forvar2290 = (forvar2290 + (1'h1)))
                    begin
                      reg2291 <= ((({reg2294} ?
                          forvar2271 : reg2263[(3'h4):(3'h4)]) >>> forvar2285[(3'h6):(2'h3)]) < {($signed(wire2226) ^ $unsigned((8'ha7)))});
                      reg2292 <= reg2256;
                    end
                  if ((-reg2291))
                    begin
                      reg2293 <= {((|$signed(reg2284)) ^~ reg2288)};
                      reg2294 <= $unsigned(forvar2291);
                      reg2295 <= wire2226[(1'h0):(1'h0)];
                      reg2296 <= $unsigned(($signed($signed(reg2275)) < (+(reg2282 + reg2291))));
                    end
                  else
                    begin
                      reg2293 <= reg2263[(4'h9):(2'h3)];
                      reg2294 <= (reg2236 | (reg2280[(4'hd):(3'h6)] && ($signed(reg2299) <<< reg2256)));
                      reg2295 <= ((~reg2274) ? forvar2285 : forvar2285);
                    end
                  if ($signed((~^$unsigned((reg2235 | (8'ha9))))))
                    begin
                      reg2297 <= $signed({forvar2246[(3'h4):(1'h0)]});
                    end
                  else
                    begin
                      reg2297 <= $signed(reg2251[(3'h5):(2'h3)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar2245 = (1'h0); (forvar2245 < (2'h2)); forvar2245 = (forvar2245 + (1'h1)))
            begin
              reg2246 <= ({$unsigned(forvar2285)} ?
                  forvar2261 : reg2282[(3'h5):(1'h0)]);
              reg2247 <= $unsigned({((reg2250 ~^ reg2279) > (8'ha1))});
            end
          for (forvar2248 = (1'h0); (forvar2248 < (2'h2)); forvar2248 = (forvar2248 + (1'h1)))
            begin
              if ((^($unsigned(forvar2250[(1'h0):(1'h0)]) ?
                  (~^$unsigned(reg2242)) : $signed(reg2281[(1'h0):(1'h0)]))))
                begin
                  for (forvar2249 = (1'h0); (forvar2249 < (2'h2)); forvar2249 = (forvar2249 + (1'h1)))
                    begin
                      reg2250 <= reg2272;
                      reg2251 <= ((~$signed((forvar2277 ~^ forvar2266))) ?
                          $unsigned({$unsigned(reg2258)}) : (reg2259[(4'hd):(3'h6)] > $signed($signed(reg2291))));
                      reg2252 <= $signed(forvar2249);
                    end
                  for (forvar2253 = (1'h0); (forvar2253 < (1'h1)); forvar2253 = (forvar2253 + (1'h1)))
                    begin
                      reg2254 <= $unsigned(reg2267);
                      reg2255 <= $signed($unsigned(((!reg2239) & (reg2238 || reg2249))));
                      reg2256 <= (&(~^wire2226));
                    end
                  if ((($unsigned(forvar2249) ?
                          $unsigned((!forvar2296)) : reg2290) ?
                      forvar2291[(4'he):(4'hb)] : {wire2229}))
                    begin
                      reg2257 <= (-(forvar2231[(3'h4):(1'h1)] ?
                          reg2281[(2'h2):(2'h2)] : $unsigned((reg2272 < forvar2232))));
                    end
                  else
                    begin
                      reg2257 <= {reg2236[(1'h0):(1'h0)]};
                      reg2258 <= (~&($unsigned((|(8'ha6))) | ({wire2229} || (forvar2248 >> reg2298))));
                      reg2259 <= $signed(({$signed(reg2298)} ?
                          $unsigned(forvar2290[(3'h6):(3'h6)]) : reg2293));
                      reg2260 <= $unsigned($unsigned((~^(&reg2273))));
                    end
                end
              else
                begin
                  reg2249 <= $signed(reg2265);
                  if ((((reg2264 ^ reg2238) << reg2276) ?
                      (~reg2280[(2'h3):(1'h1)]) : (~&(-forvar2249[(2'h3):(2'h2)]))))
                    begin
                      reg2250 <= $unsigned(reg2284[(3'h6):(1'h1)]);
                      reg2251 <= $signed(($unsigned(forvar2245) ?
                          $unsigned((reg2290 ?
                              reg2264 : reg2290)) : $unsigned(reg2252)));
                      reg2252 <= (8'ha0);
                    end
                  else
                    begin
                      reg2250 <= forvar2249[(2'h3):(1'h1)];
                      reg2251 <= (~reg2251);
                      reg2252 <= (~$unsigned(reg2272[(1'h0):(1'h0)]));
                    end
                  if ({(~&($signed(reg2294) * reg2267))})
                    begin
                      reg2253 <= $unsigned((~|((reg2299 > reg2291) <<< (reg2237 <<< reg2275))));
                      reg2254 <= forvar2241[(1'h0):(1'h0)];
                      reg2255 <= (8'hb7);
                    end
                  else
                    begin
                      reg2253 <= $signed(wire2229[(2'h2):(1'h1)]);
                      reg2254 <= reg2291[(4'hd):(2'h2)];
                    end
                  if (($signed(((|forvar2230) == (forvar2291 <= reg2247))) ?
                      $unsigned($unsigned((reg2294 ?
                          forvar2291 : reg2260))) : $unsigned($signed($signed(reg2294)))))
                    begin
                      reg2256 <= $signed($unsigned(forvar2266[(1'h1):(1'h1)]));
                      reg2257 <= ((((!(8'ha7)) == {forvar2245}) == reg2246[(3'h7):(3'h7)]) << $unsigned(($signed(forvar2253) >= $signed(wire2229))));
                    end
                  else
                    begin
                      reg2256 <= ({(forvar2262 || (+reg2269))} ^ (-$unsigned({reg2249})));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2300 = (1'h0); (forvar2300 < (2'h2)); forvar2300 = (forvar2300 + (1'h1)))
        begin
          if ($signed(((reg2255 ?
              (reg2263 ? reg2287 : wire2227) : (~^(8'h9e))) * (8'hb1))))
            begin
              if ((&(reg2298[(3'h5):(3'h5)] - $unsigned(reg2254))))
                begin
                  for (forvar2301 = (1'h0); (forvar2301 < (1'h0)); forvar2301 = (forvar2301 + (1'h1)))
                    begin
                      reg2302 <= (reg2295 < ($unsigned((reg2249 ?
                          reg2292 : wire2226)) <= reg2280[(3'h7):(2'h2)]));
                      reg2303 <= ($signed(((wire2227 ?
                          forvar2241 : reg2276) > $unsigned(reg2278))) < reg2237);
                      reg2304 <= $unsigned(reg2295[(3'h5):(3'h5)]);
                    end
                  for (forvar2305 = (1'h0); (forvar2305 < (1'h0)); forvar2305 = (forvar2305 + (1'h1)))
                    begin
                      reg2306 <= forvar2246;
                      reg2307 <= reg2302[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  reg2301 <= ({(+(&(8'hb5)))} & $unsigned((!$signed(reg2276))));
                  for (forvar2302 = (1'h0); (forvar2302 < (1'h1)); forvar2302 = (forvar2302 + (1'h1)))
                    begin
                      reg2303 <= (({(forvar2233 ? forvar2248 : reg2237)} ?
                              {reg2281[(2'h2):(1'h1)]} : (reg2236 || $signed(reg2284))) ?
                          ($signed((~|(8'hb8))) ?
                              forvar2301[(3'h7):(2'h2)] : $unsigned($unsigned(forvar2253))) : reg2273);
                      reg2304 <= $signed((~&(-reg2243)));
                    end
                end
              if (reg2299)
                begin
                  if ($signed($signed($signed(forvar2240))))
                    begin
                      reg2308 <= reg2286;
                      reg2309 <= $signed((($unsigned((8'ha3)) ?
                          $unsigned((8'ha0)) : $unsigned(reg2243)) > ($unsigned((8'ha3)) ?
                          $signed(forvar2257) : $signed(reg2295))));
                      reg2310 <= reg2280;
                      reg2311 <= $signed($unsigned($signed(((8'h9d) ?
                          (8'hac) : forvar2290))));
                    end
                  else
                    begin
                      reg2308 <= {(|$signed(reg2283[(4'h8):(1'h0)]))};
                    end
                end
              else
                begin
                  if ((($signed((reg2253 ? (8'hb8) : forvar2233)) ?
                          reg2280[(4'hf):(1'h1)] : reg2299[(2'h3):(2'h2)]) ?
                      reg2236[(2'h2):(1'h0)] : $signed($unsigned($signed(forvar2245)))))
                    begin
                      reg2308 <= (!forvar2282[(1'h1):(1'h0)]);
                      reg2309 <= ((~((reg2238 <= (8'hb7)) ?
                          (~^forvar2232) : reg2290[(3'h7):(1'h1)])) != reg2247[(2'h3):(1'h0)]);
                      reg2310 <= (^~(({forvar2285} ?
                              reg2238[(2'h3):(1'h0)] : forvar2250[(1'h0):(1'h0)]) ?
                          (8'ha3) : forvar2271));
                      reg2311 <= ((reg2260 >> (8'ha1)) ~^ ({(reg2242 ?
                              reg2239 : forvar2232)} ^ $unsigned(reg2251)));
                    end
                  else
                    begin
                      reg2308 <= $signed({{$signed(reg2287)}});
                    end
                end
            end
          else
            begin
              if ((+$unsigned(forvar2305[(1'h0):(1'h0)])))
                begin
                  for (forvar2301 = (1'h0); (forvar2301 < (2'h2)); forvar2301 = (forvar2301 + (1'h1)))
                    begin
                      reg2302 <= reg2273[(4'hd):(4'h9)];
                      reg2303 <= ((((reg2269 >>> reg2252) ?
                              $signed(reg2293) : ((8'hb6) <<< (8'ha8))) ?
                          reg2267[(2'h2):(1'h0)] : reg2294) != (&forvar2290));
                      reg2304 <= $signed($signed($signed(reg2247[(4'ha):(3'h7)])));
                      reg2305 <= (reg2242[(1'h1):(1'h0)] ?
                          ({(!reg2307)} != $signed((reg2294 + forvar2253))) : ($signed((reg2251 >> reg2273)) - (reg2294 << $unsigned(reg2272))));
                    end
                end
              else
                begin
                  for (forvar2301 = (1'h0); (forvar2301 < (2'h3)); forvar2301 = (forvar2301 + (1'h1)))
                    begin
                      reg2302 <= $signed(forvar2266[(2'h2):(2'h2)]);
                      reg2303 <= ((forvar2245 <<< ((reg2237 <<< reg2247) ?
                              (-reg2253) : ((8'h9c) ? reg2265 : (8'hb6)))) ?
                          (!{{forvar2262}}) : {reg2268[(1'h1):(1'h1)]});
                      reg2304 <= reg2293[(1'h1):(1'h0)];
                    end
                  if ((((forvar2240[(3'h5):(1'h0)] * reg2287[(3'h5):(1'h1)]) ~^ reg2265[(1'h0):(1'h0)]) ~^ (forvar2248[(3'h4):(2'h3)] - wire2227[(4'hb):(3'h7)])))
                    begin
                      reg2305 <= {$signed(forvar2290)};
                      reg2306 <= ($unsigned(reg2280) & (^reg2292));
                      reg2307 <= (|(~|(!reg2281)));
                      reg2308 <= $signed(((|{forvar2300}) ?
                          {(reg2299 ? forvar2233 : reg2295)} : (~&reg2236)));
                    end
                  else
                    begin
                      reg2305 <= $signed(reg2238);
                      reg2306 <= forvar2230;
                    end
                  if (reg2247)
                    begin
                      reg2309 <= forvar2305;
                    end
                  else
                    begin
                      reg2309 <= $unsigned((($unsigned(reg2237) ?
                          $signed(reg2270) : (forvar2257 << reg2269)) & (8'h9c)));
                      reg2310 <= reg2295[(2'h2):(1'h0)];
                    end
                end
              reg2311 <= $unsigned({(~|$unsigned(reg2254))});
              reg2312 <= (8'hb3);
            end
          if ((~^(forvar2253 < ($signed(reg2243) - wire2228))))
            begin
              for (forvar2313 = (1'h0); (forvar2313 < (1'h0)); forvar2313 = (forvar2313 + (1'h1)))
                begin
                  reg2314 <= (^forvar2248);
                  if ({reg2295[(3'h7):(3'h6)]})
                    begin
                      reg2315 <= $unsigned($unsigned($signed(((8'ha2) ?
                          forvar2296 : reg2274))));
                      reg2316 <= reg2268;
                      reg2317 <= $unsigned((~^$unsigned($signed(reg2305))));
                      reg2318 <= (reg2268 ?
                          ({$signed(forvar2253)} ^ ((|forvar2300) && (reg2238 ?
                              reg2234 : forvar2241))) : ($signed(reg2234[(3'h4):(3'h4)]) << $signed(reg2238[(2'h3):(1'h1)])));
                    end
                  else
                    begin
                      reg2315 <= ({$signed($signed(reg2248))} >= reg2243);
                      reg2316 <= ($unsigned($unsigned((reg2247 ?
                              reg2274 : (8'haa)))) ?
                          {(^reg2308)} : $unsigned($unsigned($signed(wire2226))));
                      reg2317 <= $signed($unsigned((reg2248 ?
                          (8'haa) : ((8'ha2) ? forvar2249 : reg2238))));
                    end
                end
              for (forvar2319 = (1'h0); (forvar2319 < (1'h1)); forvar2319 = (forvar2319 + (1'h1)))
                begin
                  for (forvar2320 = (1'h0); (forvar2320 < (2'h2)); forvar2320 = (forvar2320 + (1'h1)))
                    begin
                      reg2321 <= (reg2239 + {reg2280});
                    end
                end
              if (forvar2320)
                begin
                  reg2322 <= ($unsigned(($unsigned(reg2307) ?
                      (reg2295 ? forvar2305 : forvar2302) : (reg2317 ?
                          (8'hb1) : reg2295))) * reg2302[(2'h2):(2'h2)]);
                  reg2323 <= forvar2320;
                end
              else
                begin
                  reg2322 <= (reg2307 ?
                      (reg2284[(2'h2):(2'h2)] <<< forvar2253) : (^(forvar2249[(4'h9):(3'h6)] ?
                          reg2265 : (~&reg2242))));
                  if (($signed((8'ha0)) ? (8'hb9) : wire2227[(3'h6):(3'h5)]))
                    begin
                      reg2323 <= {(~|$unsigned($unsigned(reg2312)))};
                      reg2324 <= (($signed((!(8'hb2))) || {(+reg2244)}) >>> {reg2235});
                      reg2325 <= $signed((reg2305 == reg2318[(3'h7):(2'h2)]));
                    end
                  else
                    begin
                      reg2323 <= $signed(forvar2231[(1'h0):(1'h0)]);
                      reg2324 <= $signed($unsigned({$signed((8'ha6))}));
                      reg2325 <= ($unsigned($unsigned((^reg2247))) ?
                          $unsigned(forvar2266) : (($unsigned((8'h9f)) ?
                                  $unsigned(reg2267) : $signed(wire2227)) ?
                              $unsigned(reg2248[(2'h2):(1'h0)]) : ((|reg2310) <= (forvar2240 ?
                                  forvar2241 : reg2252))));
                    end
                  if (reg2288[(1'h1):(1'h0)])
                    begin
                      reg2326 <= reg2252[(2'h2):(1'h1)];
                      reg2327 <= forvar2240;
                    end
                  else
                    begin
                      reg2326 <= ((&reg2312[(3'h5):(2'h2)]) ?
                          {$unsigned((forvar2240 ?
                                  (8'ha7) : forvar2301))} : (8'hb1));
                      reg2327 <= $unsigned((reg2267[(2'h2):(2'h2)] | reg2246[(3'h7):(1'h0)]));
                      reg2328 <= reg2238;
                      reg2329 <= (~&((+((8'ha0) | reg2297)) | (~&(reg2280 ?
                          forvar2296 : reg2328))));
                    end
                  for (forvar2330 = (1'h0); (forvar2330 < (2'h2)); forvar2330 = (forvar2330 + (1'h1)))
                    begin
                      reg2331 <= reg2315;
                    end
                end
            end
          else
            begin
              for (forvar2313 = (1'h0); (forvar2313 < (2'h2)); forvar2313 = (forvar2313 + (1'h1)))
                begin
                  for (forvar2314 = (1'h0); (forvar2314 < (1'h1)); forvar2314 = (forvar2314 + (1'h1)))
                    begin
                      reg2315 <= $unsigned(reg2277);
                    end
                  if (forvar2246[(2'h2):(1'h0)])
                    begin
                      reg2316 <= $unsigned((reg2248[(3'h7):(3'h4)] ?
                          (reg2327 >> {reg2298}) : {(~|forvar2302)}));
                      reg2317 <= (+(reg2246 << $signed($unsigned(forvar2245))));
                    end
                  else
                    begin
                      reg2316 <= reg2294[(3'h5):(1'h1)];
                      reg2317 <= ((((8'ha0) || $unsigned(wire2228)) < $signed((reg2263 ?
                          forvar2277 : (8'ha7)))) * (!{forvar2232[(2'h3):(2'h2)]}));
                      reg2318 <= (8'ha1);
                    end
                  for (forvar2319 = (1'h0); (forvar2319 < (1'h0)); forvar2319 = (forvar2319 + (1'h1)))
                    begin
                      reg2320 <= ($signed(reg2326) - forvar2330);
                      reg2321 <= reg2257[(1'h1):(1'h0)];
                      reg2322 <= reg2242[(1'h0):(1'h0)];
                    end
                end
              reg2323 <= (~(~reg2281));
            end
        end
      if ((~^({forvar2253[(3'h5):(1'h0)]} << reg2292[(3'h4):(2'h2)])))
        begin
          for (forvar2332 = (1'h0); (forvar2332 < (2'h2)); forvar2332 = (forvar2332 + (1'h1)))
            begin
              if ((|$unsigned(($unsigned(reg2267) ?
                  $signed((8'ha9)) : (8'hb0)))))
                begin
                  for (forvar2333 = (1'h0); (forvar2333 < (2'h3)); forvar2333 = (forvar2333 + (1'h1)))
                    begin
                      reg2334 <= $unsigned((reg2268 ?
                          reg2277[(3'h4):(2'h3)] : reg2322[(4'hb):(3'h5)]));
                      reg2335 <= (8'hac);
                      reg2336 <= $unsigned($signed($signed(reg2248[(1'h0):(1'h0)])));
                      reg2337 <= reg2238[(1'h0):(1'h0)];
                    end
                  if ((8'hb5))
                    begin
                      reg2338 <= ($unsigned($signed((!reg2282))) ~^ forvar2300);
                      reg2339 <= $signed((((~|forvar2296) ?
                              (~^forvar2257) : reg2317[(2'h2):(2'h2)]) ?
                          (+reg2323[(2'h2):(2'h2)]) : ((reg2257 * reg2259) ?
                              (^reg2259) : ((8'ha6) << reg2260))));
                    end
                  else
                    begin
                      reg2338 <= ({(((8'ha7) ? forvar2233 : forvar2233) ?
                                  reg2296 : (8'hb8))} ?
                          ($signed((reg2263 >> reg2238)) ?
                              reg2254[(2'h2):(1'h1)] : ($signed(reg2324) != reg2276[(4'h9):(1'h0)])) : ((forvar2231[(2'h3):(1'h0)] ~^ (&(8'hab))) ?
                              $signed((reg2338 >= forvar2271)) : reg2324[(1'h0):(1'h0)]));
                      reg2339 <= ((($unsigned(reg2247) ?
                          (-forvar2257) : $signed(reg2294)) > reg2236[(2'h2):(1'h0)]) >>> $signed($signed(reg2269)));
                      reg2340 <= forvar2320;
                    end
                  for (forvar2341 = (1'h0); (forvar2341 < (2'h3)); forvar2341 = (forvar2341 + (1'h1)))
                    begin
                      reg2342 <= $unsigned(reg2331);
                    end
                end
              else
                begin
                  for (forvar2333 = (1'h0); (forvar2333 < (2'h3)); forvar2333 = (forvar2333 + (1'h1)))
                    begin
                      reg2334 <= (^~(8'hac));
                    end
                  if ($unsigned($unsigned((^$signed(forvar2241)))))
                    begin
                      reg2335 <= $unsigned($unsigned(($signed((8'hb9)) ?
                          $signed(forvar2250) : reg2303)));
                      reg2336 <= $signed((($signed(reg2322) ?
                          (8'ha9) : ((8'h9f) ^ reg2234)) < (^{(8'h9c)})));
                      reg2337 <= reg2304[(2'h2):(1'h0)];
                      reg2338 <= (reg2253[(3'h5):(1'h1)] ?
                          $unsigned((+(reg2234 <= reg2301))) : (({reg2336} + $unsigned(reg2272)) ?
                              ($unsigned(forvar2261) ?
                                  $signed(forvar2245) : reg2252) : ($signed(forvar2233) ?
                                  {reg2340} : forvar2250[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg2335 <= forvar2290[(3'h6):(1'h1)];
                      reg2336 <= {forvar2233[(4'h9):(3'h4)]};
                    end
                  reg2339 <= (~|((~(reg2299 && reg2244)) ^ (8'hb1)));
                  if (forvar2300)
                    begin
                      reg2340 <= forvar2240[(1'h0):(1'h0)];
                      reg2341 <= reg2324[(1'h0):(1'h0)];
                      reg2342 <= ((((reg2317 ?
                                  reg2315 : reg2338) ^ $unsigned((8'hb1))) ?
                              ((|forvar2231) >= reg2258) : forvar2230) ?
                          $unsigned($signed($unsigned((8'hb0)))) : {($signed(reg2320) ?
                                  reg2237 : (reg2304 ? reg2318 : reg2259))});
                      reg2343 <= (reg2253 ?
                          (reg2291 ?
                              ({reg2247} ?
                                  wire2228 : (8'hb3)) : reg2303[(2'h2):(2'h2)]) : (8'ha8));
                    end
                  else
                    begin
                      reg2340 <= $signed($unsigned($signed((!reg2257))));
                      reg2341 <= (-(^reg2336));
                    end
                end
              for (forvar2344 = (1'h0); (forvar2344 < (1'h1)); forvar2344 = (forvar2344 + (1'h1)))
                begin
                  if ($unsigned((((reg2235 ^~ forvar2320) == $signed(reg2236)) ?
                      ((!reg2314) && reg2336) : $signed((+forvar2262)))))
                    begin
                      reg2345 <= (forvar2305[(1'h0):(1'h0)] ?
                          ((~$unsigned(reg2250)) ?
                              {((8'hae) ?
                                      forvar2313 : reg2305)} : {$unsigned(reg2248)}) : {($signed(forvar2319) ?
                                  $unsigned(forvar2232) : (forvar2333 ^~ reg2325))});
                      reg2346 <= reg2312;
                      reg2347 <= {($signed((~&reg2324)) ?
                              (+reg2343[(1'h1):(1'h0)]) : $signed((~|(8'hb4))))};
                    end
                  else
                    begin
                      reg2345 <= forvar2319;
                      reg2346 <= ($unsigned(wire2227[(1'h0):(1'h0)]) + ((reg2280[(4'ha):(4'h9)] ?
                          {reg2272} : $signed(forvar2271)) <= reg2316));
                      reg2347 <= ($signed(((~^wire2227) ?
                          forvar2241[(4'hc):(3'h7)] : forvar2257[(3'h6):(3'h4)])) - forvar2320[(3'h5):(3'h4)]);
                      reg2348 <= ((reg2267[(1'h1):(1'h1)] ?
                          (reg2238 ?
                              $unsigned(forvar2332) : (-reg2259)) : (|(reg2275 < forvar2341))) && reg2248[(2'h2):(2'h2)]);
                    end
                end
            end
          reg2349 <= wire2227;
          for (forvar2350 = (1'h0); (forvar2350 < (2'h2)); forvar2350 = (forvar2350 + (1'h1)))
            begin
              for (forvar2351 = (1'h0); (forvar2351 < (2'h3)); forvar2351 = (forvar2351 + (1'h1)))
                begin
                  for (forvar2352 = (1'h0); (forvar2352 < (2'h3)); forvar2352 = (forvar2352 + (1'h1)))
                    begin
                      reg2353 <= (~&(8'haf));
                      reg2354 <= {(~^{(reg2268 != forvar2233)})};
                      reg2355 <= (~&reg2299[(1'h1):(1'h0)]);
                      reg2356 <= reg2246;
                    end
                  if ($unsigned(reg2243))
                    begin
                      reg2357 <= forvar2314;
                      reg2358 <= ($signed(($signed(reg2336) * reg2310[(3'h7):(3'h6)])) ?
                          ((~&{reg2294}) ?
                              reg2270 : $unsigned($unsigned((8'h9f)))) : reg2341);
                    end
                  else
                    begin
                      reg2357 <= (reg2243 ^~ {$signed((8'h9d))});
                      reg2358 <= $signed($signed((|$unsigned(reg2278))));
                      reg2359 <= reg2314[(2'h3):(1'h0)];
                      reg2360 <= reg2237;
                    end
                end
              if ($unsigned($signed(reg2267[(1'h1):(1'h1)])))
                begin
                  reg2361 <= forvar2230;
                  if ((8'haa))
                    begin
                      reg2362 <= $unsigned((-wire2228[(3'h6):(3'h4)]));
                      reg2363 <= reg2248;
                    end
                  else
                    begin
                      reg2362 <= $signed($signed((((8'had) ?
                          reg2234 : reg2257) < {(8'hb2)})));
                      reg2363 <= (~|($signed(reg2302[(2'h2):(1'h1)]) + ({reg2253} | forvar2233)));
                    end
                end
              else
                begin
                  reg2361 <= $unsigned({(reg2264 << forvar2240)});
                  reg2362 <= reg2307[(2'h2):(1'h1)];
                  if ($unsigned({$signed((8'ha1))}))
                    begin
                      reg2363 <= ($unsigned($unsigned(((8'ha6) << reg2335))) == ((8'ha1) ^ (~&reg2353)));
                      reg2364 <= $signed(reg2325);
                      reg2365 <= ($unsigned($signed($unsigned(reg2346))) ?
                          (($unsigned(reg2342) ? (^~wire2226) : (|(8'hae))) ?
                              forvar2296 : (8'hb1)) : reg2327);
                      reg2366 <= (~|reg2268[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2363 <= (+(+$unsigned($unsigned(forvar2262))));
                      reg2364 <= (^~((^~(forvar2332 + forvar2240)) ?
                          $unsigned($unsigned(reg2339)) : forvar2285[(1'h1):(1'h1)]));
                      reg2365 <= ($signed(forvar2305[(1'h0):(1'h0)]) ?
                          $unsigned(forvar2282[(1'h0):(1'h0)]) : $signed(reg2356));
                      reg2366 <= {reg2327[(4'h8):(4'h8)]};
                    end
                end
            end
        end
      else
        begin
          reg2332 <= reg2253[(3'h6):(1'h0)];
          for (forvar2333 = (1'h0); (forvar2333 < (2'h2)); forvar2333 = (forvar2333 + (1'h1)))
            begin
              for (forvar2334 = (1'h0); (forvar2334 < (2'h3)); forvar2334 = (forvar2334 + (1'h1)))
                begin
                  for (forvar2335 = (1'h0); (forvar2335 < (2'h2)); forvar2335 = (forvar2335 + (1'h1)))
                    begin
                      reg2336 <= reg2276;
                      reg2337 <= {reg2263};
                      reg2338 <= ((&forvar2231[(1'h0):(1'h0)]) ?
                          (reg2295 ?
                              (^(-reg2334)) : (reg2284[(2'h3):(2'h2)] >>> $unsigned(reg2318))) : ((~|wire2226[(2'h2):(1'h1)]) && ($signed(reg2275) ?
                              $unsigned(forvar2335) : $signed(reg2249))));
                    end
                  for (forvar2339 = (1'h0); (forvar2339 < (1'h1)); forvar2339 = (forvar2339 + (1'h1)))
                    begin
                      reg2340 <= ((((forvar2351 ? reg2305 : forvar2351) ?
                              wire2226 : $unsigned((8'h9c))) * (~(^reg2250))) ?
                          (((8'hb9) ?
                              ((8'ha1) <<< reg2340) : $unsigned((8'ha5))) >>> (!wire2226[(2'h2):(1'h1)])) : $signed({reg2355[(2'h2):(1'h1)]}));
                      reg2341 <= (($unsigned(reg2365[(1'h1):(1'h0)]) != $unsigned($signed(reg2257))) != (^(^~((8'hb1) ?
                          (8'hb6) : reg2327))));
                      reg2342 <= ((reg2290 ?
                          (forvar2352[(2'h2):(1'h0)] ^~ $signed(reg2323)) : reg2254[(4'he):(4'h8)]) < $signed($unsigned(((8'hb6) ^~ reg2305))));
                    end
                  if ($signed($unsigned($unsigned((+(8'ha2))))))
                    begin
                      reg2343 <= {reg2363};
                      reg2344 <= (~forvar2290);
                      reg2345 <= (8'ha1);
                      reg2346 <= forvar2320;
                    end
                  else
                    begin
                      reg2343 <= $unsigned((^(reg2239[(4'h9):(3'h4)] ?
                          $signed(forvar2302) : (~^reg2297))));
                    end
                  for (forvar2347 = (1'h0); (forvar2347 < (2'h3)); forvar2347 = (forvar2347 + (1'h1)))
                    begin
                      reg2348 <= $signed(reg2365[(1'h0):(1'h0)]);
                      reg2349 <= $signed((^~forvar2352[(1'h1):(1'h1)]));
                      reg2350 <= $unsigned((|forvar2347));
                      reg2351 <= {$signed($unsigned(((8'had) <<< forvar2241)))};
                    end
                end
            end
          reg2352 <= ({((reg2307 == reg2264) ?
                  (-(8'ha2)) : $signed((8'ha2)))} & (!$signed(reg2234[(2'h3):(1'h0)])));
        end
    end
  module2367 modinst3015 (wire3014, clk, forvar2347, reg2287, reg2329, forvar2301);
  assign wire3016 = reg2252[(4'ha):(4'ha)];
  assign wire3017 = $signed(($unsigned((8'hb0)) ^~ $unsigned({reg2295})));
  assign wire3018 = (!reg2332);
  assign wire3019 = forvar2339[(3'h6):(2'h2)];
  assign wire3020 = wire3014;
  always
    @(posedge clk) begin
      if ($signed(wire3018))
        begin
          reg3021 <= $unsigned((reg2286 < $signed(reg2248)));
          for (forvar3022 = (1'h0); (forvar3022 < (1'h0)); forvar3022 = (forvar3022 + (1'h1)))
            begin
              if ({((8'ha3) << $unsigned((reg2321 < reg2249)))})
                begin
                  reg3023 <= $unsigned(reg2264);
                  for (forvar3024 = (1'h0); (forvar3024 < (1'h0)); forvar3024 = (forvar3024 + (1'h1)))
                    begin
                      reg3025 <= (reg2251 < (8'hb5));
                      reg3026 <= {$unsigned($unsigned((reg2290 ?
                              forvar2314 : reg2295)))};
                      reg3027 <= ((+(+forvar2335)) || reg2366);
                    end
                  for (forvar3028 = (1'h0); (forvar3028 < (1'h1)); forvar3028 = (forvar3028 + (1'h1)))
                    begin
                      reg3029 <= (^~((~|(reg2323 - reg2325)) <<< (~|reg2320[(2'h2):(2'h2)])));
                    end
                  if ((8'hba))
                    begin
                      reg3030 <= {$signed(($signed(reg2268) ?
                              {reg2358} : ((8'hb6) | forvar2320)))};
                      reg3031 <= $unsigned(({(wire3014 ?
                              (8'hb0) : (8'hb5))} << ((reg2359 && reg2274) & reg2277)));
                      reg3032 <= reg2335;
                      reg3033 <= ({(~&$signed(reg3032))} * forvar2313);
                    end
                  else
                    begin
                      reg3030 <= {wire3020[(3'h4):(2'h3)]};
                    end
                end
              else
                begin
                  for (forvar3023 = (1'h0); (forvar3023 < (1'h1)); forvar3023 = (forvar3023 + (1'h1)))
                    begin
                      reg3024 <= ({($signed(reg2276) | $unsigned(forvar2230))} ?
                          (^($unsigned(reg2243) ?
                              ((8'hb4) >>> reg2234) : (reg2237 & reg2314))) : $signed(((~^reg2360) ?
                              $signed(reg2284) : reg2249)));
                    end
                  reg3025 <= reg2332;
                  for (forvar3026 = (1'h0); (forvar3026 < (2'h2)); forvar3026 = (forvar3026 + (1'h1)))
                    begin
                      reg3027 <= {$signed($unsigned(forvar2291))};
                      reg3028 <= $unsigned((&(reg2351[(2'h2):(2'h2)] < reg2305)));
                    end
                  for (forvar3029 = (1'h0); (forvar3029 < (1'h1)); forvar3029 = (forvar3029 + (1'h1)))
                    begin
                      reg3030 <= $signed((|$unsigned($signed(reg2328))));
                    end
                end
              if ({reg2290})
                begin
                  for (forvar3034 = (1'h0); (forvar3034 < (1'h1)); forvar3034 = (forvar3034 + (1'h1)))
                    begin
                      reg3035 <= $signed(({$signed((8'haa))} <<< {$signed(reg2320)}));
                      reg3036 <= $unsigned((reg2323 ?
                          $signed((reg2243 ?
                              (8'hb5) : reg2250)) : (|reg2357[(4'hb):(4'hb)])));
                      reg3037 <= (~(^reg2249[(2'h2):(1'h0)]));
                    end
                  for (forvar3038 = (1'h0); (forvar3038 < (2'h2)); forvar3038 = (forvar3038 + (1'h1)))
                    begin
                      reg3039 <= reg2284;
                      reg3040 <= reg2339;
                      reg3041 <= $signed((({forvar3029} ?
                          forvar3023 : $signed(reg2305)) ~^ $unsigned((~forvar2266))));
                    end
                end
              else
                begin
                  for (forvar3034 = (1'h0); (forvar3034 < (2'h2)); forvar3034 = (forvar3034 + (1'h1)))
                    begin
                      reg3035 <= (forvar2233[(5'h10):(4'ha)] > reg2356[(4'h9):(4'h8)]);
                    end
                end
              for (forvar3042 = (1'h0); (forvar3042 < (1'h1)); forvar3042 = (forvar3042 + (1'h1)))
                begin
                  if ($unsigned({forvar2285}))
                    begin
                      reg3043 <= forvar2296[(3'h7):(2'h2)];
                    end
                  else
                    begin
                      reg3043 <= reg2349[(3'h5):(2'h3)];
                      reg3044 <= (+$signed($signed($unsigned(reg2270))));
                      reg3045 <= $unsigned((|(reg2358[(1'h0):(1'h0)] ?
                          $unsigned(reg2325) : (forvar2245 * reg2244))));
                      reg3046 <= {{{(8'hb2)}}};
                    end
                end
            end
          for (forvar3047 = (1'h0); (forvar3047 < (2'h3)); forvar3047 = (forvar3047 + (1'h1)))
            begin
              for (forvar3048 = (1'h0); (forvar3048 < (1'h0)); forvar3048 = (forvar3048 + (1'h1)))
                begin
                  for (forvar3049 = (1'h0); (forvar3049 < (2'h2)); forvar3049 = (forvar3049 + (1'h1)))
                    begin
                      reg3050 <= (^reg2275[(1'h1):(1'h0)]);
                      reg3051 <= (($signed((8'hb6)) * {(~^reg2303)}) ?
                          reg2317 : ($signed(reg3037[(4'h9):(1'h0)]) ?
                              ($signed(reg2283) ?
                                  $unsigned(forvar2290) : (reg2301 || (8'had))) : {$signed(wire3016)}));
                    end
                  if (((~^($unsigned(forvar2302) << (forvar3022 ?
                          reg3024 : reg2335))) ?
                      (-$signed({reg2260})) : ($signed(forvar3048) - (reg2274[(3'h6):(2'h2)] ?
                          reg2352[(3'h7):(2'h3)] : (8'ha4)))))
                    begin
                      reg3052 <= $signed(reg3035);
                      reg3053 <= (forvar2241 ?
                          reg2329[(4'h8):(3'h6)] : $signed($unsigned(reg2263)));
                      reg3054 <= {$unsigned((8'haa))};
                      reg3055 <= reg2272[(3'h7):(1'h0)];
                    end
                  else
                    begin
                      reg3052 <= reg2346[(2'h2):(1'h1)];
                      reg3053 <= $unsigned(forvar2344[(1'h0):(1'h0)]);
                    end
                  if (reg2316)
                    begin
                      reg3056 <= (forvar2271[(1'h0):(1'h0)] || (-($unsigned(reg2281) ?
                          $unsigned(reg2346) : (reg3029 ? reg2250 : (8'hb9)))));
                      reg3057 <= $unsigned($unsigned(reg2307));
                      reg3058 <= reg2343;
                    end
                  else
                    begin
                      reg3056 <= $unsigned(($signed(reg2292[(3'h4):(3'h4)]) ?
                          ((reg2299 ?
                              reg3056 : reg2306) << $unsigned(reg2282)) : ((reg2307 ^ reg2316) ?
                              (reg2243 ?
                                  reg2281 : reg2351) : $unsigned(reg2316))));
                      reg3057 <= ($unsigned((-((8'hb8) ? reg2346 : reg2332))) ?
                          ((-(reg2252 ?
                              (8'hb7) : reg3027)) * reg2316[(2'h2):(1'h1)]) : reg2360[(4'h9):(1'h1)]);
                      reg3058 <= forvar2301[(3'h4):(1'h0)];
                      reg3059 <= {reg2275[(3'h5):(3'h4)]};
                    end
                  reg3060 <= $unsigned(reg2292[(3'h6):(3'h5)]);
                end
              if ((reg2343 ~^ $signed($signed($unsigned(reg2342)))))
                begin
                  if (((8'hb3) && {(-reg2270[(1'h1):(1'h1)])}))
                    begin
                      reg3061 <= (^~({forvar3049} ?
                          forvar2250 : (~(~|reg3046))));
                    end
                  else
                    begin
                      reg3061 <= ({((reg3046 ?
                                  reg2237 : reg2350) - $signed(reg2280))} ?
                          (+forvar2250[(2'h3):(2'h2)]) : reg2339[(3'h4):(2'h3)]);
                      reg3062 <= $unsigned((|(^~forvar2332)));
                    end
                  reg3063 <= ((!$signed((forvar2347 ?
                      forvar2249 : reg2321))) && ($unsigned(reg2358[(1'h1):(1'h1)]) ?
                      reg2279 : (((8'h9d) <<< (8'hac)) >> forvar3038)));
                  reg3064 <= (^~(8'hac));
                end
              else
                begin
                  for (forvar3061 = (1'h0); (forvar3061 < (1'h1)); forvar3061 = (forvar3061 + (1'h1)))
                    begin
                      reg3062 <= (+$signed({reg3021}));
                      reg3063 <= {$unsigned({(!(8'hac))})};
                      reg3064 <= $unsigned(wire3016);
                      reg3065 <= $signed(($signed((&reg2305)) <<< $unsigned((&forvar2305))));
                    end
                  for (forvar3066 = (1'h0); (forvar3066 < (1'h1)); forvar3066 = (forvar3066 + (1'h1)))
                    begin
                      reg3067 <= ((($unsigned((8'ha9)) * reg2352[(4'h8):(1'h1)]) ?
                              (8'ha6) : $signed($unsigned(reg2337))) ?
                          $signed($signed(reg2280)) : $unsigned({$signed(reg2270)}));
                      reg3068 <= (^reg2235);
                    end
                end
              reg3069 <= ($unsigned((!((8'hac) > forvar2341))) ?
                  (~&reg2258[(3'h5):(1'h0)]) : $unsigned({reg2351[(3'h7):(3'h7)]}));
            end
        end
      else
        begin
          reg3021 <= reg2249[(1'h0):(1'h0)];
        end
      if (reg2336[(2'h2):(1'h0)])
        begin
          if ($unsigned(reg2317))
            begin
              if ((reg2323 >> reg2292[(2'h2):(1'h1)]))
                begin
                  for (forvar3070 = (1'h0); (forvar3070 < (2'h2)); forvar3070 = (forvar3070 + (1'h1)))
                    begin
                      reg3071 <= (!reg2314);
                      reg3072 <= reg3068[(3'h6):(2'h3)];
                    end
                  for (forvar3073 = (1'h0); (forvar3073 < (1'h0)); forvar3073 = (forvar3073 + (1'h1)))
                    begin
                      reg3074 <= $signed((forvar3024 ?
                          $unsigned((~reg2350)) : reg2298));
                    end
                  reg3075 <= $unsigned({{$signed(reg2251)}});
                  if ($signed($unsigned($signed({(8'ha0)}))))
                    begin
                      reg3076 <= {$unsigned($signed((&reg2283)))};
                      reg3077 <= $unsigned((8'hb7));
                      reg3078 <= forvar2233[(3'h7):(2'h2)];
                    end
                  else
                    begin
                      reg3076 <= $signed({$unsigned($signed((8'hb2)))});
                      reg3077 <= (reg2297[(3'h5):(1'h0)] || (wire3020[(2'h3):(1'h1)] ?
                          reg2358[(1'h0):(1'h0)] : (!(8'hba))));
                      reg3078 <= wire3020;
                    end
                end
              else
                begin
                  if (wire3018)
                    begin
                      reg3070 <= reg2356;
                      reg3071 <= $signed((((8'ha7) | $unsigned(reg2264)) * ({reg3078} * $signed(reg2329))));
                      reg3072 <= $signed((-(-{forvar2350})));
                      reg3073 <= forvar2240[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg3070 <= (^~($signed(reg3024[(3'h7):(1'h1)]) - ({reg2337} ?
                          $signed((8'h9e)) : (reg3078 ? reg2287 : reg2274))));
                      reg3071 <= forvar2319;
                      reg3072 <= reg3039[(2'h2):(2'h2)];
                    end
                end
            end
          else
            begin
              reg3070 <= $unsigned(forvar2233);
              for (forvar3071 = (1'h0); (forvar3071 < (2'h2)); forvar3071 = (forvar3071 + (1'h1)))
                begin
                  for (forvar3072 = (1'h0); (forvar3072 < (2'h2)); forvar3072 = (forvar3072 + (1'h1)))
                    begin
                      reg3073 <= $signed({(~^((8'hae) <<< reg3024))});
                    end
                  if ($signed(({$signed(reg3031)} && reg2248[(2'h2):(2'h2)])))
                    begin
                      reg3074 <= reg3029;
                      reg3075 <= reg2304[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3074 <= $unsigned(reg2297);
                    end
                  reg3076 <= (~(^~(|$signed(reg3036))));
                end
            end
          reg3079 <= $signed($unsigned(forvar3071[(2'h3):(1'h1)]));
          if (($signed(reg2366[(3'h4):(3'h4)]) ?
              $unsigned((reg2362[(4'hb):(4'hb)] ?
                  (reg2288 >> reg2355) : $signed(reg2269))) : {reg3075[(2'h2):(2'h2)]}))
            begin
              reg3080 <= reg2281;
              for (forvar3081 = (1'h0); (forvar3081 < (1'h0)); forvar3081 = (forvar3081 + (1'h1)))
                begin
                  for (forvar3082 = (1'h0); (forvar3082 < (1'h1)); forvar3082 = (forvar3082 + (1'h1)))
                    begin
                      reg3083 <= (-(-(!reg2290[(2'h3):(2'h2)])));
                    end
                  for (forvar3084 = (1'h0); (forvar3084 < (2'h2)); forvar3084 = (forvar3084 + (1'h1)))
                    begin
                      reg3085 <= (reg2301[(2'h2):(1'h0)] ?
                          ($signed((wire3018 - forvar2240)) ?
                              $signed((wire3018 ?
                                  (8'hb5) : forvar2277)) : forvar3038) : (~&reg2311));
                      reg3086 <= $unsigned(($unsigned((reg3070 > forvar2282)) <<< ({(8'ha3)} ?
                          (forvar3081 ^ reg2353) : (reg2291 >>> forvar3047))));
                      reg3087 <= reg2317[(3'h6):(3'h5)];
                      reg3088 <= (-(8'haf));
                    end
                  for (forvar3089 = (1'h0); (forvar3089 < (2'h2)); forvar3089 = (forvar3089 + (1'h1)))
                    begin
                      reg3090 <= $signed(((reg3061 ?
                              $signed(reg2263) : $unsigned(reg3064)) ?
                          $unsigned((reg2328 ?
                              reg2277 : forvar2334)) : $unsigned((^(8'hb2)))));
                      reg3091 <= reg3036[(3'h4):(1'h1)];
                      reg3092 <= ($unsigned(reg3056) ?
                          $unsigned(($unsigned(wire2227) ?
                              reg2354[(3'h6):(1'h0)] : forvar3024[(2'h2):(1'h1)])) : reg2341);
                    end
                  if ($unsigned({reg3087[(1'h0):(1'h0)]}))
                    begin
                      reg3093 <= {(({wire2226} ?
                                  (forvar2296 & forvar2334) : $unsigned(forvar2248)) ?
                              (^(forvar2291 ?
                                  (8'hb6) : reg2243)) : (reg3055[(2'h2):(2'h2)] ?
                                  {reg3076} : $signed(forvar2262)))};
                      reg3094 <= ((forvar2253 >>> $unsigned($signed((8'hb3)))) || $unsigned(reg3090));
                      reg3095 <= reg3087[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg3093 <= (($signed(reg2317[(2'h3):(1'h0)]) ?
                              reg2302 : ((forvar2344 ?
                                  forvar2250 : forvar2261) <<< forvar2233)) ?
                          reg2314[(2'h2):(1'h1)] : ((^~((8'h9d) <= forvar3024)) ?
                              $signed((reg2284 ?
                                  reg3093 : reg2350)) : (!(reg2282 | reg3072))));
                      reg3094 <= (~^reg3095[(1'h1):(1'h1)]);
                      reg3095 <= (((reg2242[(2'h3):(2'h2)] > $unsigned(reg3055)) + reg3040) ?
                          $unsigned(((reg2290 ? reg2347 : forvar3084) ?
                              reg3057 : {reg2320})) : $unsigned(reg2275[(1'h0):(1'h0)]));
                      reg3096 <= (reg2247 ?
                          $unsigned(((+reg2276) == (+reg2248))) : $unsigned(reg2280));
                    end
                end
              for (forvar3097 = (1'h0); (forvar3097 < (2'h3)); forvar3097 = (forvar3097 + (1'h1)))
                begin
                  if (reg2304)
                    begin
                      reg3098 <= $signed(((^(8'hb4)) ?
                          forvar2257[(4'h9):(2'h3)] : {(reg2236 ?
                                  wire3017 : reg3092)}));
                      reg3099 <= $signed(forvar2282[(3'h7):(1'h1)]);
                    end
                  else
                    begin
                      reg3098 <= forvar2245[(2'h2):(2'h2)];
                      reg3099 <= (+(reg2250 ^~ (~|(forvar2266 + reg2242))));
                    end
                  if (($unsigned($unsigned((reg3043 <= reg2252))) ?
                      (~$signed((^~reg3086))) : (reg2280[(4'hb):(3'h4)] + reg2326)))
                    begin
                      reg3100 <= ($unsigned((+(8'hb3))) + $signed($unsigned((~^(8'hb9)))));
                      reg3101 <= ($signed(($signed(reg2334) == $unsigned((8'ha3)))) * (((wire3016 ^ forvar2248) >> $signed(forvar3072)) * (~^$unsigned(reg3024))));
                      reg3102 <= $signed(((~^$signed(forvar2347)) ?
                          ($unsigned(forvar3022) > (|forvar2271)) : reg3050[(4'h9):(2'h2)]));
                      reg3103 <= $signed({((forvar2352 ? (8'hb7) : reg3045) ?
                              forvar3034[(4'he):(4'he)] : (reg3045 ^ reg3073))});
                    end
                  else
                    begin
                      reg3100 <= ($unsigned((~^$unsigned((8'ha1)))) ?
                          ((^~reg2288) == (reg3087[(3'h4):(3'h4)] ^ ((8'hb9) != reg3035))) : (8'h9d));
                      reg3101 <= ($signed((|(reg2312 >= forvar2249))) <= (((reg2263 ?
                              reg2326 : reg3027) ?
                          $unsigned(reg3051) : wire3019) | (&reg2341)));
                      reg3102 <= (~(reg3036 ?
                          {wire3018[(1'h1):(1'h0)]} : reg3040[(3'h5):(1'h1)]));
                    end
                  for (forvar3104 = (1'h0); (forvar3104 < (1'h0)); forvar3104 = (forvar3104 + (1'h1)))
                    begin
                      reg3105 <= $unsigned((~^$unsigned($signed(reg2350))));
                      reg3106 <= (((8'ha3) ?
                              $unsigned((reg3091 > (8'ha0))) : (forvar2344[(2'h2):(2'h2)] ?
                                  (8'hb8) : (reg2354 ? reg2323 : reg3071))) ?
                          $signed($unsigned({reg2272})) : (~&(reg3079[(1'h1):(1'h1)] ?
                              (reg3032 ? reg2332 : wire3017) : (reg3026 ?
                                  (8'h9c) : forvar2305))));
                    end
                end
            end
          else
            begin
              for (forvar3080 = (1'h0); (forvar3080 < (1'h0)); forvar3080 = (forvar3080 + (1'h1)))
                begin
                  for (forvar3081 = (1'h0); (forvar3081 < (2'h3)); forvar3081 = (forvar3081 + (1'h1)))
                    begin
                      reg3082 <= reg2314[(4'h9):(4'h9)];
                    end
                end
              for (forvar3083 = (1'h0); (forvar3083 < (1'h1)); forvar3083 = (forvar3083 + (1'h1)))
                begin
                  if ({(~^$signed(reg3074))})
                    begin
                      reg3084 <= (($unsigned(reg3077[(1'h1):(1'h1)]) << forvar2248) ?
                          (!$unsigned($unsigned(reg3055))) : (!reg2349[(1'h1):(1'h1)]));
                      reg3085 <= reg2361;
                      reg3086 <= reg2352[(2'h2):(1'h1)];
                      reg3087 <= reg2278;
                    end
                  else
                    begin
                      reg3084 <= $signed(((~&((8'h9f) ?
                          reg3041 : reg3063)) <= (8'ha8)));
                    end
                end
              for (forvar3088 = (1'h0); (forvar3088 < (1'h1)); forvar3088 = (forvar3088 + (1'h1)))
                begin
                  for (forvar3089 = (1'h0); (forvar3089 < (1'h1)); forvar3089 = (forvar3089 + (1'h1)))
                    begin
                      reg3090 <= (&forvar2248);
                      reg3091 <= (reg2237 ?
                          $signed($signed((~reg2246))) : reg2344);
                      reg3092 <= $signed((reg2352[(2'h3):(2'h3)] ?
                          {reg2298} : {$unsigned(reg2297)}));
                      reg3093 <= reg3050[(2'h2):(1'h0)];
                    end
                  for (forvar3094 = (1'h0); (forvar3094 < (2'h2)); forvar3094 = (forvar3094 + (1'h1)))
                    begin
                      reg3095 <= ((+$unsigned($unsigned(reg2264))) ?
                          reg2341 : (^reg2362[(3'h7):(3'h5)]));
                    end
                end
            end
        end
      else
        begin
          if (reg2239)
            begin
              reg3070 <= (8'hb8);
              for (forvar3071 = (1'h0); (forvar3071 < (1'h0)); forvar3071 = (forvar3071 + (1'h1)))
                begin
                  reg3072 <= reg2238;
                  for (forvar3073 = (1'h0); (forvar3073 < (2'h3)); forvar3073 = (forvar3073 + (1'h1)))
                    begin
                      reg3074 <= ($signed($signed((^reg2304))) ?
                          $signed(reg2289) : {reg2268[(2'h2):(1'h1)]});
                      reg3075 <= $signed((forvar2341 * reg3078[(1'h0):(1'h0)]));
                      reg3076 <= reg2327;
                    end
                end
            end
          else
            begin
              if (($unsigned(forvar3049) & (!(8'h9f))))
                begin
                  for (forvar3070 = (1'h0); (forvar3070 < (2'h2)); forvar3070 = (forvar3070 + (1'h1)))
                    begin
                      reg3071 <= (-$unsigned(reg3069));
                    end
                  reg3072 <= $unsigned((~^(8'haf)));
                  for (forvar3073 = (1'h0); (forvar3073 < (1'h1)); forvar3073 = (forvar3073 + (1'h1)))
                    begin
                      reg3074 <= reg2257;
                      reg3075 <= (~|$unsigned(forvar3048));
                      reg3076 <= $signed((((reg2295 ?
                          reg2243 : forvar2314) | reg2356) && reg2288));
                      reg3077 <= reg2276[(2'h3):(1'h0)];
                    end
                  if ($unsigned((((reg2236 != reg2263) ?
                          (reg2281 ?
                              reg2296 : wire3018) : $signed(forvar2262)) ?
                      $unsigned((^~reg3086)) : reg2269[(1'h0):(1'h0)])))
                    begin
                      reg3078 <= {$signed($signed((reg3052 ?
                              reg2297 : forvar2352)))};
                      reg3079 <= {forvar2253[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg3078 <= $unsigned(reg3028);
                      reg3079 <= (^($signed((8'hb7)) == (8'hb4)));
                      reg3080 <= (^((!$signed(reg2294)) ?
                          reg2310[(4'hd):(1'h1)] : reg2349));
                      reg3081 <= {reg3025};
                    end
                end
              else
                begin
                  if ((+(&{$signed(reg2273)})))
                    begin
                      reg3070 <= (^$unsigned({(forvar2290 ?
                              forvar3029 : forvar3094)}));
                      reg3071 <= reg2275;
                    end
                  else
                    begin
                      reg3070 <= $signed((reg3062 < (((8'ha6) << wire3016) ?
                          reg2292 : (reg2258 | reg2363))));
                      reg3071 <= {$signed(((wire2229 ^~ reg2263) ?
                              {reg2237} : (reg3079 ? reg2327 : (8'hb2))))};
                    end
                  for (forvar3072 = (1'h0); (forvar3072 < (1'h0)); forvar3072 = (forvar3072 + (1'h1)))
                    begin
                      reg3073 <= $unsigned((~{(forvar2253 ~^ forvar2347)}));
                    end
                  if ($unsigned((reg2362 > {{reg2287}})))
                    begin
                      reg3074 <= ($signed($unsigned($signed(wire2226))) != {(^~$signed(reg2350))});
                      reg3075 <= forvar2245;
                      reg3076 <= ((~^((reg2243 ?
                          wire2227 : reg2357) > (8'ha1))) ^~ ((reg2320[(3'h7):(1'h1)] ?
                              (reg3055 ? (8'hb4) : (8'h9d)) : (reg2256 ?
                                  reg2362 : reg3090)) ?
                          reg2311[(4'hb):(1'h0)] : reg2304));
                    end
                  else
                    begin
                      reg3074 <= (&{((|reg3085) ?
                              (reg3057 <<< wire2228) : $signed(reg3065))});
                      reg3075 <= $signed((reg3024 >= $signed($signed((8'ha1)))));
                      reg3076 <= ($signed((8'haa)) ?
                          ({{reg2295}} ?
                              reg3095 : $signed($unsigned(wire3014))) : (+(~|(reg2287 && forvar2296))));
                      reg3077 <= ($unsigned($signed($unsigned(reg2325))) ?
                          reg2343 : $unsigned(forvar3023));
                    end
                  for (forvar3078 = (1'h0); (forvar3078 < (1'h1)); forvar3078 = (forvar3078 + (1'h1)))
                    begin
                      reg3079 <= (forvar2262 ?
                          $unsigned($unsigned((reg2349 ?
                              reg2265 : reg2345))) : ({$signed(reg2315)} | {$unsigned(reg2301)}));
                      reg3080 <= forvar2230;
                      reg3081 <= ((|reg2284[(1'h0):(1'h0)]) ?
                          ((+reg3043) ?
                              ((8'hb7) || forvar3024) : forvar2240) : (&reg2355));
                    end
                end
            end
        end
      reg3107 <= ((~^((~|reg2322) ? {wire3019} : (8'hb6))) ?
          $signed((8'haa)) : reg3060[(3'h7):(2'h2)]);
      reg3108 <= reg3041;
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2367  (y, clk, wire2371, wire2370, wire2369, wire2368);
  output wire [(32'h1a47):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire2371;
  input wire [(3'h7):(1'h0)] wire2370;
  input wire [(3'h4):(1'h0)] wire2369;
  input wire [(4'hf):(1'h0)] wire2368;
  reg [(4'he):(1'h0)] reg3010 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3013 = (1'h0);
  reg [(4'h9):(1'h0)] reg3012 = (1'h0);
  reg [(4'he):(1'h0)] reg3011 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3010 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3009 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3008 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3007 = (1'h0);
  reg [(4'he):(1'h0)] reg3006 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3005 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3004 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3003 = (1'h0);
  reg [(2'h3):(1'h0)] reg3002 = (1'h0);
  reg [(4'h8):(1'h0)] reg3001 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3000 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2999 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2997 = (1'h0);
  reg [(4'h9):(1'h0)] reg2991 = (1'h0);
  reg [(4'he):(1'h0)] reg2990 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2987 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2986 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2983 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2980 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2979 = (1'h0);
  reg [(4'hc):(1'h0)] reg2973 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2971 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2961 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2968 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2967 = (1'h0);
  reg [(3'h5):(1'h0)] reg2965 = (1'h0);
  reg [(4'hd):(1'h0)] reg2963 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2957 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2995 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2998 = (1'h0);
  reg [(4'hc):(1'h0)] reg2997 = (1'h0);
  reg [(3'h7):(1'h0)] reg2996 = (1'h0);
  reg [(5'h10):(1'h0)] reg2995 = (1'h0);
  reg [(4'h9):(1'h0)] reg2994 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2993 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2992 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2991 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2990 = (1'h0);
  reg [(3'h7):(1'h0)] reg2989 = (1'h0);
  reg [(4'h8):(1'h0)] reg2988 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2987 = (1'h0);
  reg [(2'h2):(1'h0)] reg2986 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2985 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2984 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2983 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2982 = (1'h0);
  reg [(4'he):(1'h0)] forvar2981 = (1'h0);
  reg [(4'hd):(1'h0)] reg2980 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2979 = (1'h0);
  reg [(3'h5):(1'h0)] reg2978 = (1'h0);
  reg [(3'h6):(1'h0)] reg2977 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2976 = (1'h0);
  reg [(3'h6):(1'h0)] reg2975 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2974 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2973 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2972 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2971 = (1'h0);
  reg [(4'h8):(1'h0)] reg2970 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2969 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2968 = (1'h0);
  reg [(4'h8):(1'h0)] reg2967 = (1'h0);
  reg [(5'h10):(1'h0)] reg2956 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2966 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2965 = (1'h0);
  reg [(3'h4):(1'h0)] reg2964 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2963 = (1'h0);
  reg [(3'h6):(1'h0)] reg2962 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2961 = (1'h0);
  reg [(3'h5):(1'h0)] reg2960 = (1'h0);
  reg [(4'hc):(1'h0)] reg2959 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2958 = (1'h0);
  reg [(4'h8):(1'h0)] reg2957 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2956 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2955 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2954 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2945 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2953 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2952 = (1'h0);
  reg [(4'h8):(1'h0)] reg2951 = (1'h0);
  reg [(4'hc):(1'h0)] reg2950 = (1'h0);
  reg [(3'h7):(1'h0)] reg2949 = (1'h0);
  reg [(4'hb):(1'h0)] reg2948 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2947 = (1'h0);
  reg [(2'h3):(1'h0)] reg2946 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2945 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2944 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2943 = (1'h0);
  reg [(3'h4):(1'h0)] reg2942 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2941 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2940 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2939 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2938 = (1'h0);
  reg [(3'h5):(1'h0)] reg2937 = (1'h0);
  reg [(4'he):(1'h0)] reg2936 = (1'h0);
  reg [(4'he):(1'h0)] reg2935 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2934 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2933 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2932 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2931 = (1'h0);
  reg [(2'h3):(1'h0)] reg2930 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2929 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2928 = (1'h0);
  reg [(2'h3):(1'h0)] reg2927 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2926 = (1'h0);
  reg [(4'ha):(1'h0)] reg2925 = (1'h0);
  reg [(3'h5):(1'h0)] reg2924 = (1'h0);
  reg [(3'h5):(1'h0)] reg2923 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2922 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2921 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2920 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2919 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2918 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2882 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2891 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2885 = (1'h0);
  reg [(3'h5):(1'h0)] reg2876 = (1'h0);
  reg [(4'h8):(1'h0)] reg2917 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2904 = (1'h0);
  reg [(4'h9):(1'h0)] reg2916 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2915 = (1'h0);
  reg [(3'h7):(1'h0)] reg2914 = (1'h0);
  reg [(4'ha):(1'h0)] reg2913 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2912 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2911 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2910 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2909 = (1'h0);
  reg [(3'h7):(1'h0)] reg2908 = (1'h0);
  reg [(4'hf):(1'h0)] reg2907 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2906 = (1'h0);
  reg [(4'hc):(1'h0)] reg2905 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2904 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2903 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2902 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2901 = (1'h0);
  reg [(4'he):(1'h0)] forvar2897 = (1'h0);
  reg [(4'he):(1'h0)] reg2896 = (1'h0);
  reg [(3'h5):(1'h0)] reg2894 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2893 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2900 = (1'h0);
  reg [(4'hd):(1'h0)] reg2899 = (1'h0);
  reg [(4'h9):(1'h0)] reg2898 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2897 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2896 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2895 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2894 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2893 = (1'h0);
  reg [(3'h5):(1'h0)] reg2892 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2891 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2888 = (1'h0);
  reg [(4'hb):(1'h0)] reg2883 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2881 = (1'h0);
  reg [(4'h8):(1'h0)] reg2880 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2890 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2889 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2888 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2887 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2886 = (1'h0);
  reg [(4'hf):(1'h0)] reg2885 = (1'h0);
  reg [(4'ha):(1'h0)] reg2884 = (1'h0);
  reg [(4'he):(1'h0)] forvar2883 = (1'h0);
  reg [(3'h5):(1'h0)] reg2882 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2881 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2880 = (1'h0);
  reg [(4'hb):(1'h0)] reg2879 = (1'h0);
  reg [(5'h10):(1'h0)] reg2878 = (1'h0);
  reg [(2'h2):(1'h0)] reg2877 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2876 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2875 = (1'h0);
  wire [(4'hd):(1'h0)] wire2874;
  reg signed [(4'hb):(1'h0)] reg2873 = (1'h0);
  reg [(2'h2):(1'h0)] reg2864 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2872 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2871 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2870 = (1'h0);
  reg [(2'h3):(1'h0)] reg2869 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2868 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2867 = (1'h0);
  reg [(4'he):(1'h0)] reg2866 = (1'h0);
  reg [(4'hc):(1'h0)] reg2865 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2864 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2861 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2860 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2856 = (1'h0);
  reg [(4'hc):(1'h0)] reg2863 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2862 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2861 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2860 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2859 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2858 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2857 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2856 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2855 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2833 = (1'h0);
  reg [(3'h4):(1'h0)] reg2831 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2828 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2854 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2853 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2852 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2851 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2850 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2849 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2848 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2847 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2846 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2845 = (1'h0);
  reg [(5'h10):(1'h0)] reg2844 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2843 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2842 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2841 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2840 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2839 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2838 = (1'h0);
  reg [(3'h5):(1'h0)] reg2837 = (1'h0);
  reg [(3'h6):(1'h0)] reg2836 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2835 = (1'h0);
  reg [(3'h7):(1'h0)] reg2834 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2833 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2832 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2831 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2830 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2829 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2828 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2827 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2826 = (1'h0);
  wire [(3'h5):(1'h0)] wire2825;
  reg [(4'hc):(1'h0)] reg2824 = (1'h0);
  reg [(4'hd):(1'h0)] reg2823 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2822 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2821 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2820 = (1'h0);
  reg [(4'ha):(1'h0)] reg2819 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2818 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2817 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2816 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2815 = (1'h0);
  reg [(4'hf):(1'h0)] reg2814 = (1'h0);
  reg [(4'he):(1'h0)] forvar2813 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2812 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2811 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2810 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2809 = (1'h0);
  reg [(4'h9):(1'h0)] reg2808 = (1'h0);
  reg [(4'hb):(1'h0)] reg2807 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2806 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2805 = (1'h0);
  reg [(2'h3):(1'h0)] reg2804 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2803 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2802 = (1'h0);
  reg [(4'hb):(1'h0)] reg2801 = (1'h0);
  reg [(3'h7):(1'h0)] reg2800 = (1'h0);
  reg [(4'hb):(1'h0)] reg2799 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2798 = (1'h0);
  reg [(4'he):(1'h0)] forvar2797 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2796 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2795 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2794 = (1'h0);
  reg [(4'hf):(1'h0)] reg2793 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2792 = (1'h0);
  reg [(4'hf):(1'h0)] reg2791 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2790 = (1'h0);
  reg [(3'h5):(1'h0)] reg2789 = (1'h0);
  reg [(4'hb):(1'h0)] reg2788 = (1'h0);
  reg [(3'h5):(1'h0)] reg2787 = (1'h0);
  reg [(4'hf):(1'h0)] reg2786 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2785 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2784 = (1'h0);
  reg [(4'h9):(1'h0)] reg2783 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2782 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2781 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2775 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2780 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2779 = (1'h0);
  reg [(4'h8):(1'h0)] reg2778 = (1'h0);
  reg [(2'h3):(1'h0)] reg2777 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2776 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2775 = (1'h0);
  reg [(3'h4):(1'h0)] reg2774 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2773 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2772 = (1'h0);
  reg [(3'h4):(1'h0)] reg2771 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2770 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2769 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2768 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2767 = (1'h0);
  reg [(4'h8):(1'h0)] reg2766 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2765 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2764 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2763 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2762 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2761 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2757 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2760 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2759 = (1'h0);
  reg [(4'h9):(1'h0)] reg2758 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2757 = (1'h0);
  reg [(3'h7):(1'h0)] reg2756 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2755 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2754 = (1'h0);
  reg [(4'h9):(1'h0)] reg2753 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2752 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2751 = (1'h0);
  reg [(4'hd):(1'h0)] reg2741 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2739 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2737 = (1'h0);
  reg [(3'h5):(1'h0)] reg2750 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2749 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2748 = (1'h0);
  reg [(5'h10):(1'h0)] reg2747 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2746 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2744 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2745 = (1'h0);
  reg [(3'h5):(1'h0)] reg2744 = (1'h0);
  reg [(4'hd):(1'h0)] reg2743 = (1'h0);
  reg [(2'h3):(1'h0)] reg2742 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2741 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2740 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2739 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2738 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2737 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2736 = (1'h0);
  reg [(3'h4):(1'h0)] reg2735 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2734 = (1'h0);
  reg [(2'h3):(1'h0)] reg2733 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2732 = (1'h0);
  reg [(4'hc):(1'h0)] reg2731 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2730 = (1'h0);
  reg [(4'ha):(1'h0)] reg2729 = (1'h0);
  reg [(2'h3):(1'h0)] reg2728 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2727 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2726 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2725 = (1'h0);
  reg [(4'h8):(1'h0)] reg2724 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2723 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2722 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2721 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2720 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2719 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2718 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2717 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2703 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2702 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2714 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2711 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2710 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2717 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2716 = (1'h0);
  reg [(4'h9):(1'h0)] reg2715 = (1'h0);
  reg [(3'h4):(1'h0)] reg2714 = (1'h0);
  reg [(4'hc):(1'h0)] reg2713 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2712 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2711 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2709 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2708 = (1'h0);
  reg [(4'hd):(1'h0)] reg2710 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2709 = (1'h0);
  reg [(4'h8):(1'h0)] reg2708 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2707 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2706 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2705 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2704 = (1'h0);
  reg [(4'hb):(1'h0)] reg2701 = (1'h0);
  reg [(4'hb):(1'h0)] reg2703 = (1'h0);
  reg [(3'h5):(1'h0)] reg2702 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2701 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2700 = (1'h0);
  reg [(4'h8):(1'h0)] reg2699 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2698 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2697 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2696 = (1'h0);
  reg [(4'hb):(1'h0)] reg2695 = (1'h0);
  reg [(5'h10):(1'h0)] reg2694 = (1'h0);
  reg [(4'h8):(1'h0)] reg2693 = (1'h0);
  reg [(4'he):(1'h0)] reg2692 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2691 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2690 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2689 = (1'h0);
  reg [(4'h9):(1'h0)] reg2688 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2687 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2686 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2685 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2684 = (1'h0);
  reg [(4'h9):(1'h0)] reg2683 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2682 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2681 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2681 = (1'h0);
  reg [(2'h3):(1'h0)] reg2680 = (1'h0);
  reg [(2'h2):(1'h0)] reg2679 = (1'h0);
  reg [(2'h3):(1'h0)] reg2678 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2677 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2676 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2675 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2674 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2673 = (1'h0);
  reg [(4'hb):(1'h0)] reg2672 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2670 = (1'h0);
  reg [(3'h7):(1'h0)] reg2671 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2670 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2668 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2664 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2663 = (1'h0);
  reg [(4'h9):(1'h0)] reg2662 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2669 = (1'h0);
  reg [(3'h4):(1'h0)] reg2668 = (1'h0);
  reg [(3'h5):(1'h0)] reg2667 = (1'h0);
  reg [(5'h10):(1'h0)] reg2666 = (1'h0);
  reg [(3'h6):(1'h0)] reg2665 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2664 = (1'h0);
  reg [(3'h6):(1'h0)] reg2663 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2662 = (1'h0);
  reg [(4'he):(1'h0)] reg2661 = (1'h0);
  reg [(4'hb):(1'h0)] reg2660 = (1'h0);
  reg [(2'h3):(1'h0)] reg2659 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2658 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2657 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2656 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2655 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2654 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2653 = (1'h0);
  reg [(4'h8):(1'h0)] reg2652 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2651 = (1'h0);
  reg [(3'h4):(1'h0)] reg2650 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2649 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2648 = (1'h0);
  reg [(4'hb):(1'h0)] reg2647 = (1'h0);
  reg [(4'ha):(1'h0)] reg2646 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2645 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2644 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2643 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2642 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2641 = (1'h0);
  reg [(5'h10):(1'h0)] reg2640 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2639 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2638 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2637 = (1'h0);
  reg [(3'h5):(1'h0)] reg2636 = (1'h0);
  reg [(5'h10):(1'h0)] reg2635 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2634 = (1'h0);
  reg [(3'h7):(1'h0)] reg2633 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2632 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2631 = (1'h0);
  reg [(3'h5):(1'h0)] reg2630 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2629 = (1'h0);
  reg [(4'he):(1'h0)] reg2628 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2627 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2626 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2625 = (1'h0);
  reg [(4'hb):(1'h0)] reg2624 = (1'h0);
  reg [(4'h9):(1'h0)] reg2620 = (1'h0);
  reg [(3'h7):(1'h0)] reg2615 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2613 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2611 = (1'h0);
  reg [(4'h9):(1'h0)] reg2610 = (1'h0);
  reg [(2'h2):(1'h0)] reg2609 = (1'h0);
  reg [(5'h10):(1'h0)] reg2623 = (1'h0);
  reg [(3'h7):(1'h0)] reg2622 = (1'h0);
  reg [(3'h5):(1'h0)] reg2621 = (1'h0);
  reg [(4'he):(1'h0)] forvar2620 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2619 = (1'h0);
  reg [(3'h6):(1'h0)] reg2618 = (1'h0);
  reg [(4'hb):(1'h0)] reg2617 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2616 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2615 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2614 = (1'h0);
  reg [(4'h8):(1'h0)] reg2613 = (1'h0);
  reg [(5'h10):(1'h0)] reg2612 = (1'h0);
  reg [(3'h7):(1'h0)] reg2611 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2610 = (1'h0);
  reg [(4'he):(1'h0)] forvar2609 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2608 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2550 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2607 = (1'h0);
  reg [(4'hb):(1'h0)] reg2606 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2605 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2604 = (1'h0);
  reg [(5'h10):(1'h0)] reg2603 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2602 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2601 = (1'h0);
  reg [(4'ha):(1'h0)] reg2600 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2599 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2598 = (1'h0);
  reg [(4'he):(1'h0)] reg2597 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2596 = (1'h0);
  reg [(4'hc):(1'h0)] reg2595 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2594 = (1'h0);
  reg [(4'hb):(1'h0)] reg2593 = (1'h0);
  reg [(4'hf):(1'h0)] reg2592 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2591 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2590 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2586 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2579 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2589 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2588 = (1'h0);
  reg [(3'h4):(1'h0)] reg2587 = (1'h0);
  reg [(4'hd):(1'h0)] reg2586 = (1'h0);
  reg [(3'h5):(1'h0)] reg2585 = (1'h0);
  reg [(3'h6):(1'h0)] reg2584 = (1'h0);
  reg [(2'h3):(1'h0)] reg2583 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2582 = (1'h0);
  reg [(4'h8):(1'h0)] reg2581 = (1'h0);
  reg [(4'hf):(1'h0)] reg2580 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2579 = (1'h0);
  reg [(4'hb):(1'h0)] reg2578 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2577 = (1'h0);
  reg [(2'h3):(1'h0)] reg2576 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2575 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2574 = (1'h0);
  reg [(5'h10):(1'h0)] reg2573 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2572 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2571 = (1'h0);
  reg [(4'ha):(1'h0)] reg2570 = (1'h0);
  reg [(4'h9):(1'h0)] reg2569 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2568 = (1'h0);
  reg [(4'hb):(1'h0)] reg2567 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2566 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2565 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2564 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2563 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2562 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2561 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2560 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2559 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2558 = (1'h0);
  reg [(4'hc):(1'h0)] reg2554 = (1'h0);
  reg [(5'h10):(1'h0)] reg2557 = (1'h0);
  reg [(4'h9):(1'h0)] reg2556 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2555 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2553 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2552 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2551 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2550 = (1'h0);
  reg [(2'h3):(1'h0)] reg2549 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2548 = (1'h0);
  reg [(4'hb):(1'h0)] reg2547 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire2546;
  wire [(4'ha):(1'h0)] wire2545;
  wire signed [(4'hf):(1'h0)] wire2544;
  wire [(4'h8):(1'h0)] wire2543;
  reg signed [(3'h5):(1'h0)] reg2542 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2541 = (1'h0);
  reg [(4'hc):(1'h0)] reg2540 = (1'h0);
  reg [(3'h4):(1'h0)] reg2539 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2538 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2537 = (1'h0);
  reg [(4'hc):(1'h0)] reg2536 = (1'h0);
  reg [(4'hc):(1'h0)] reg2535 = (1'h0);
  reg [(3'h6):(1'h0)] reg2534 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2533 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2530 = (1'h0);
  reg [(4'h8):(1'h0)] reg2529 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2527 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2532 = (1'h0);
  reg [(2'h2):(1'h0)] reg2531 = (1'h0);
  reg [(3'h5):(1'h0)] reg2530 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2529 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2528 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2527 = (1'h0);
  reg [(3'h7):(1'h0)] reg2526 = (1'h0);
  reg [(4'h9):(1'h0)] reg2525 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2520 = (1'h0);
  reg [(2'h2):(1'h0)] reg2519 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2524 = (1'h0);
  reg [(4'hd):(1'h0)] reg2523 = (1'h0);
  reg [(4'hb):(1'h0)] reg2522 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2521 = (1'h0);
  reg [(3'h7):(1'h0)] reg2520 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2519 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2518 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2517 = (1'h0);
  reg [(4'he):(1'h0)] reg2516 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2515 = (1'h0);
  reg [(4'h9):(1'h0)] reg2511 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2508 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2514 = (1'h0);
  reg [(3'h7):(1'h0)] reg2513 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2512 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2511 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2510 = (1'h0);
  reg [(4'h8):(1'h0)] reg2509 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2508 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2507 = (1'h0);
  reg [(2'h2):(1'h0)] reg2506 = (1'h0);
  reg [(4'he):(1'h0)] reg2505 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2504 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2503 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2502 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2501 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2500 = (1'h0);
  reg [(3'h4):(1'h0)] reg2499 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2498 = (1'h0);
  reg [(4'ha):(1'h0)] reg2497 = (1'h0);
  reg [(4'h8):(1'h0)] reg2496 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2495 = (1'h0);
  reg [(3'h5):(1'h0)] reg2494 = (1'h0);
  reg [(3'h7):(1'h0)] reg2493 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2492 = (1'h0);
  reg [(4'ha):(1'h0)] reg2491 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2490 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2489 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2488 = (1'h0);
  reg [(4'h8):(1'h0)] reg2487 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2486 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2485 = (1'h0);
  reg [(2'h2):(1'h0)] reg2484 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2483 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2482 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2481 = (1'h0);
  reg [(4'he):(1'h0)] reg2480 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2479 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2478 = (1'h0);
  reg [(4'he):(1'h0)] reg2477 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2476 = (1'h0);
  reg [(4'hb):(1'h0)] reg2475 = (1'h0);
  reg [(5'h10):(1'h0)] reg2474 = (1'h0);
  reg [(4'he):(1'h0)] forvar2473 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2472 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2471 = (1'h0);
  reg [(2'h2):(1'h0)] reg2470 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2469 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2468 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2467 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2466 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2465 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2464 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2463 = (1'h0);
  reg [(3'h6):(1'h0)] reg2462 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2448 = (1'h0);
  reg [(4'he):(1'h0)] reg2445 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2461 = (1'h0);
  reg [(4'h8):(1'h0)] reg2460 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2459 = (1'h0);
  reg [(3'h5):(1'h0)] reg2458 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2457 = (1'h0);
  reg [(4'he):(1'h0)] forvar2452 = (1'h0);
  reg [(4'hf):(1'h0)] reg2450 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2449 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2446 = (1'h0);
  reg [(4'h8):(1'h0)] reg2456 = (1'h0);
  reg [(4'ha):(1'h0)] reg2455 = (1'h0);
  reg [(3'h5):(1'h0)] reg2454 = (1'h0);
  reg [(4'ha):(1'h0)] reg2453 = (1'h0);
  reg [(4'hd):(1'h0)] reg2452 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2451 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2450 = (1'h0);
  reg [(4'hd):(1'h0)] reg2449 = (1'h0);
  reg [(3'h7):(1'h0)] reg2448 = (1'h0);
  reg [(3'h5):(1'h0)] reg2447 = (1'h0);
  reg [(3'h5):(1'h0)] reg2446 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2445 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2387 = (1'h0);
  reg [(3'h7):(1'h0)] reg2379 = (1'h0);
  reg [(4'hb):(1'h0)] reg2377 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2397 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2394 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2389 = (1'h0);
  reg [(2'h3):(1'h0)] reg2386 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2385 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2382 = (1'h0);
  reg [(4'hb):(1'h0)] reg2378 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2428 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2422 = (1'h0);
  reg [(3'h6):(1'h0)] reg2444 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2443 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2442 = (1'h0);
  reg [(4'h9):(1'h0)] reg2441 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2440 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2439 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2438 = (1'h0);
  reg [(5'h10):(1'h0)] reg2434 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2433 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2437 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2436 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2435 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2434 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2433 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2432 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2431 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2430 = (1'h0);
  reg [(4'h9):(1'h0)] reg2429 = (1'h0);
  reg [(4'h9):(1'h0)] reg2428 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2427 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2423 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2420 = (1'h0);
  reg [(4'hd):(1'h0)] reg2426 = (1'h0);
  reg [(4'hb):(1'h0)] reg2425 = (1'h0);
  reg [(4'he):(1'h0)] reg2424 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2423 = (1'h0);
  reg [(4'he):(1'h0)] reg2422 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2421 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2420 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2398 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2419 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2418 = (1'h0);
  reg [(2'h2):(1'h0)] reg2416 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2415 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2413 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2417 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2416 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2415 = (1'h0);
  reg [(3'h5):(1'h0)] reg2414 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2413 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2408 = (1'h0);
  reg [(3'h6):(1'h0)] reg2407 = (1'h0);
  reg [(3'h4):(1'h0)] reg2412 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2411 = (1'h0);
  reg [(2'h3):(1'h0)] reg2410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2409 = (1'h0);
  reg [(4'hb):(1'h0)] reg2408 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2407 = (1'h0);
  reg [(4'hb):(1'h0)] reg2406 = (1'h0);
  reg [(4'hc):(1'h0)] reg2405 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2404 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2403 = (1'h0);
  reg [(4'hb):(1'h0)] reg2402 = (1'h0);
  reg [(4'he):(1'h0)] reg2401 = (1'h0);
  reg [(2'h3):(1'h0)] reg2400 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2399 = (1'h0);
  reg [(4'he):(1'h0)] forvar2398 = (1'h0);
  reg [(4'hb):(1'h0)] reg2397 = (1'h0);
  reg [(4'ha):(1'h0)] reg2396 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2395 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2391 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2388 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2394 = (1'h0);
  reg [(4'hb):(1'h0)] reg2393 = (1'h0);
  reg [(5'h10):(1'h0)] reg2392 = (1'h0);
  reg [(5'h10):(1'h0)] reg2391 = (1'h0);
  reg [(2'h2):(1'h0)] reg2390 = (1'h0);
  reg [(5'h10):(1'h0)] reg2389 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2388 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2384 = (1'h0);
  reg [(3'h7):(1'h0)] reg2383 = (1'h0);
  reg [(5'h10):(1'h0)] reg2387 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2386 = (1'h0);
  reg [(3'h7):(1'h0)] reg2385 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2384 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2383 = (1'h0);
  reg [(4'h9):(1'h0)] reg2382 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2381 = (1'h0);
  reg [(3'h7):(1'h0)] reg2380 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2379 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2378 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2377 = (1'h0);
  wire [(4'hc):(1'h0)] wire2376;
  wire [(4'hb):(1'h0)] wire2375;
  wire [(3'h4):(1'h0)] wire2374;
  wire [(4'he):(1'h0)] wire2373;
  wire signed [(4'hd):(1'h0)] wire2372;
  assign y = {reg3010,
                 reg3013,
                 reg3012,
                 reg3011,
                 forvar3010,
                 reg3009,
                 reg3008,
                 reg3007,
                 reg3006,
                 reg3005,
                 reg3004,
                 reg3003,
                 reg3002,
                 reg3001,
                 reg3000,
                 reg2999,
                 forvar2997,
                 reg2991,
                 reg2990,
                 forvar2987,
                 forvar2986,
                 reg2983,
                 forvar2980,
                 reg2979,
                 reg2973,
                 forvar2971,
                 forvar2961,
                 reg2968,
                 forvar2967,
                 reg2965,
                 reg2963,
                 forvar2957,
                 forvar2995,
                 reg2998,
                 reg2997,
                 reg2996,
                 reg2995,
                 reg2994,
                 reg2993,
                 reg2992,
                 forvar2991,
                 forvar2990,
                 reg2989,
                 reg2988,
                 reg2987,
                 reg2986,
                 reg2985,
                 forvar2984,
                 forvar2983,
                 reg2982,
                 forvar2981,
                 reg2980,
                 forvar2979,
                 reg2978,
                 reg2977,
                 reg2976,
                 reg2975,
                 forvar2974,
                 forvar2973,
                 forvar2972,
                 reg2971,
                 reg2970,
                 reg2969,
                 forvar2968,
                 reg2967,
                 reg2956,
                 reg2966,
                 forvar2965,
                 reg2964,
                 forvar2963,
                 reg2962,
                 reg2961,
                 reg2960,
                 reg2959,
                 reg2958,
                 reg2957,
                 forvar2956,
                 forvar2955,
                 reg2954,
                 reg2945,
                 reg2953,
                 reg2952,
                 reg2951,
                 reg2950,
                 reg2949,
                 reg2948,
                 reg2947,
                 reg2946,
                 forvar2945,
                 reg2944,
                 forvar2943,
                 reg2942,
                 reg2941,
                 forvar2940,
                 forvar2939,
                 reg2938,
                 reg2937,
                 reg2936,
                 reg2935,
                 forvar2934,
                 forvar2933,
                 forvar2932,
                 reg2931,
                 reg2930,
                 forvar2929,
                 reg2928,
                 reg2927,
                 forvar2926,
                 reg2925,
                 reg2924,
                 reg2923,
                 reg2922,
                 forvar2921,
                 forvar2920,
                 forvar2919,
                 forvar2918,
                 forvar2882,
                 forvar2891,
                 forvar2885,
                 reg2876,
                 reg2917,
                 reg2904,
                 reg2916,
                 reg2915,
                 reg2914,
                 reg2913,
                 reg2912,
                 reg2911,
                 reg2910,
                 forvar2909,
                 reg2908,
                 reg2907,
                 reg2906,
                 reg2905,
                 forvar2904,
                 reg2903,
                 forvar2902,
                 reg2901,
                 forvar2897,
                 reg2896,
                 reg2894,
                 forvar2893,
                 reg2900,
                 reg2899,
                 reg2898,
                 reg2897,
                 forvar2896,
                 reg2895,
                 forvar2894,
                 reg2893,
                 reg2892,
                 reg2891,
                 reg2888,
                 reg2883,
                 forvar2881,
                 reg2880,
                 reg2890,
                 reg2889,
                 forvar2888,
                 reg2887,
                 reg2886,
                 reg2885,
                 reg2884,
                 forvar2883,
                 reg2882,
                 reg2881,
                 forvar2880,
                 reg2879,
                 reg2878,
                 reg2877,
                 forvar2876,
                 forvar2875,
                 wire2874,
                 reg2873,
                 reg2864,
                 reg2872,
                 reg2871,
                 reg2870,
                 reg2869,
                 forvar2868,
                 reg2867,
                 reg2866,
                 reg2865,
                 forvar2864,
                 reg2861,
                 forvar2860,
                 reg2856,
                 reg2863,
                 reg2862,
                 forvar2861,
                 reg2860,
                 reg2859,
                 reg2858,
                 reg2857,
                 forvar2856,
                 forvar2855,
                 reg2833,
                 reg2831,
                 reg2828,
                 reg2854,
                 reg2853,
                 reg2852,
                 forvar2851,
                 reg2850,
                 forvar2849,
                 reg2848,
                 reg2847,
                 forvar2846,
                 forvar2845,
                 reg2844,
                 reg2843,
                 reg2842,
                 reg2841,
                 reg2840,
                 forvar2839,
                 forvar2838,
                 reg2837,
                 reg2836,
                 reg2835,
                 reg2834,
                 forvar2833,
                 reg2832,
                 forvar2831,
                 reg2830,
                 reg2829,
                 forvar2828,
                 forvar2827,
                 reg2826,
                 wire2825,
                 reg2824,
                 reg2823,
                 forvar2822,
                 reg2821,
                 reg2820,
                 reg2819,
                 reg2818,
                 forvar2817,
                 reg2816,
                 reg2815,
                 reg2814,
                 forvar2813,
                 reg2812,
                 forvar2811,
                 forvar2810,
                 reg2809,
                 reg2808,
                 reg2807,
                 reg2806,
                 forvar2805,
                 reg2804,
                 reg2803,
                 forvar2802,
                 reg2801,
                 reg2800,
                 reg2799,
                 reg2798,
                 forvar2797,
                 reg2796,
                 reg2795,
                 reg2794,
                 reg2793,
                 forvar2792,
                 reg2791,
                 reg2790,
                 reg2789,
                 reg2788,
                 reg2787,
                 reg2786,
                 reg2785,
                 forvar2784,
                 reg2783,
                 forvar2782,
                 forvar2781,
                 reg2775,
                 reg2780,
                 reg2779,
                 reg2778,
                 reg2777,
                 reg2776,
                 forvar2775,
                 reg2774,
                 reg2773,
                 reg2772,
                 reg2771,
                 reg2770,
                 reg2769,
                 reg2768,
                 forvar2767,
                 reg2766,
                 reg2765,
                 reg2764,
                 forvar2763,
                 reg2762,
                 reg2761,
                 reg2757,
                 reg2760,
                 reg2759,
                 reg2758,
                 forvar2757,
                 reg2756,
                 reg2755,
                 forvar2754,
                 reg2753,
                 forvar2752,
                 forvar2751,
                 reg2741,
                 reg2739,
                 forvar2737,
                 reg2750,
                 forvar2749,
                 reg2748,
                 reg2747,
                 reg2746,
                 forvar2744,
                 reg2745,
                 reg2744,
                 reg2743,
                 reg2742,
                 forvar2741,
                 reg2740,
                 forvar2739,
                 forvar2738,
                 reg2737,
                 reg2736,
                 reg2735,
                 reg2734,
                 reg2733,
                 reg2732,
                 reg2731,
                 forvar2730,
                 reg2729,
                 reg2728,
                 reg2727,
                 reg2726,
                 forvar2725,
                 reg2724,
                 reg2723,
                 reg2722,
                 reg2721,
                 forvar2720,
                 forvar2719,
                 reg2718,
                 forvar2717,
                 forvar2703,
                 forvar2702,
                 forvar2714,
                 reg2711,
                 forvar2710,
                 reg2717,
                 reg2716,
                 reg2715,
                 reg2714,
                 reg2713,
                 reg2712,
                 forvar2711,
                 reg2709,
                 forvar2708,
                 reg2710,
                 forvar2709,
                 reg2708,
                 reg2707,
                 reg2706,
                 reg2705,
                 reg2704,
                 reg2701,
                 reg2703,
                 reg2702,
                 forvar2701,
                 reg2700,
                 reg2699,
                 reg2698,
                 reg2697,
                 forvar2696,
                 reg2695,
                 reg2694,
                 reg2693,
                 reg2692,
                 forvar2691,
                 forvar2690,
                 reg2689,
                 reg2688,
                 reg2687,
                 reg2686,
                 reg2685,
                 reg2684,
                 reg2683,
                 reg2682,
                 forvar2681,
                 reg2681,
                 reg2680,
                 reg2679,
                 reg2678,
                 forvar2677,
                 reg2676,
                 forvar2675,
                 forvar2674,
                 reg2673,
                 reg2672,
                 forvar2670,
                 reg2671,
                 reg2670,
                 forvar2668,
                 reg2664,
                 forvar2663,
                 reg2662,
                 reg2669,
                 reg2668,
                 reg2667,
                 reg2666,
                 reg2665,
                 forvar2664,
                 reg2663,
                 forvar2662,
                 reg2661,
                 reg2660,
                 reg2659,
                 reg2658,
                 reg2657,
                 forvar2656,
                 forvar2655,
                 reg2654,
                 reg2653,
                 reg2652,
                 reg2651,
                 reg2650,
                 forvar2649,
                 forvar2648,
                 reg2647,
                 reg2646,
                 reg2645,
                 reg2644,
                 forvar2643,
                 forvar2642,
                 forvar2641,
                 reg2640,
                 reg2639,
                 forvar2638,
                 reg2637,
                 reg2636,
                 reg2635,
                 reg2634,
                 reg2633,
                 reg2632,
                 forvar2631,
                 reg2630,
                 reg2629,
                 reg2628,
                 reg2627,
                 forvar2626,
                 forvar2625,
                 reg2624,
                 reg2620,
                 reg2615,
                 forvar2613,
                 forvar2611,
                 reg2610,
                 reg2609,
                 reg2623,
                 reg2622,
                 reg2621,
                 forvar2620,
                 reg2619,
                 reg2618,
                 reg2617,
                 reg2616,
                 forvar2615,
                 reg2614,
                 reg2613,
                 reg2612,
                 reg2611,
                 forvar2610,
                 forvar2609,
                 forvar2608,
                 reg2550,
                 reg2607,
                 reg2606,
                 reg2605,
                 reg2604,
                 reg2603,
                 reg2602,
                 reg2601,
                 reg2600,
                 forvar2599,
                 reg2598,
                 reg2597,
                 forvar2596,
                 reg2595,
                 reg2594,
                 reg2593,
                 reg2592,
                 forvar2591,
                 reg2590,
                 forvar2586,
                 forvar2579,
                 reg2589,
                 reg2588,
                 reg2587,
                 reg2586,
                 reg2585,
                 reg2584,
                 reg2583,
                 reg2582,
                 reg2581,
                 reg2580,
                 reg2579,
                 reg2578,
                 reg2577,
                 reg2576,
                 forvar2575,
                 forvar2574,
                 reg2573,
                 reg2572,
                 forvar2571,
                 reg2570,
                 reg2569,
                 reg2568,
                 reg2567,
                 reg2566,
                 forvar2565,
                 reg2564,
                 reg2563,
                 reg2562,
                 reg2561,
                 forvar2560,
                 reg2559,
                 forvar2558,
                 reg2554,
                 reg2557,
                 reg2556,
                 reg2555,
                 forvar2554,
                 reg2553,
                 reg2552,
                 forvar2551,
                 forvar2550,
                 reg2549,
                 forvar2548,
                 reg2547,
                 wire2546,
                 wire2545,
                 wire2544,
                 wire2543,
                 reg2542,
                 forvar2541,
                 reg2540,
                 reg2539,
                 reg2538,
                 reg2537,
                 reg2536,
                 reg2535,
                 reg2534,
                 reg2533,
                 forvar2530,
                 reg2529,
                 reg2527,
                 reg2532,
                 reg2531,
                 reg2530,
                 forvar2529,
                 reg2528,
                 forvar2527,
                 reg2526,
                 reg2525,
                 forvar2520,
                 reg2519,
                 reg2524,
                 reg2523,
                 reg2522,
                 reg2521,
                 reg2520,
                 forvar2519,
                 forvar2518,
                 reg2517,
                 reg2516,
                 forvar2515,
                 reg2511,
                 forvar2508,
                 reg2514,
                 reg2513,
                 reg2512,
                 forvar2511,
                 reg2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 reg2506,
                 reg2505,
                 reg2504,
                 forvar2503,
                 forvar2502,
                 forvar2501,
                 forvar2500,
                 reg2499,
                 reg2498,
                 reg2497,
                 reg2496,
                 reg2495,
                 reg2494,
                 reg2493,
                 forvar2492,
                 reg2491,
                 reg2490,
                 reg2489,
                 reg2488,
                 reg2487,
                 forvar2486,
                 forvar2485,
                 reg2484,
                 reg2483,
                 forvar2482,
                 reg2481,
                 reg2480,
                 reg2479,
                 reg2478,
                 reg2477,
                 reg2476,
                 reg2475,
                 reg2474,
                 forvar2473,
                 forvar2472,
                 reg2471,
                 reg2470,
                 reg2469,
                 reg2468,
                 reg2467,
                 reg2466,
                 forvar2465,
                 reg2464,
                 reg2463,
                 reg2462,
                 forvar2448,
                 reg2445,
                 reg2461,
                 reg2460,
                 reg2459,
                 reg2458,
                 forvar2457,
                 forvar2452,
                 reg2450,
                 forvar2449,
                 forvar2446,
                 reg2456,
                 reg2455,
                 reg2454,
                 reg2453,
                 reg2452,
                 reg2451,
                 forvar2450,
                 reg2449,
                 reg2448,
                 reg2447,
                 reg2446,
                 forvar2445,
                 forvar2387,
                 reg2379,
                 reg2377,
                 forvar2397,
                 forvar2394,
                 forvar2389,
                 reg2386,
                 forvar2385,
                 forvar2382,
                 reg2378,
                 forvar2428,
                 forvar2422,
                 reg2444,
                 forvar2443,
                 reg2442,
                 reg2441,
                 reg2440,
                 reg2439,
                 forvar2438,
                 reg2434,
                 forvar2433,
                 reg2437,
                 reg2436,
                 reg2435,
                 forvar2434,
                 reg2433,
                 reg2432,
                 reg2431,
                 reg2430,
                 reg2429,
                 reg2428,
                 reg2427,
                 reg2423,
                 forvar2420,
                 reg2426,
                 reg2425,
                 reg2424,
                 forvar2423,
                 reg2422,
                 reg2421,
                 reg2420,
                 reg2398,
                 reg2419,
                 forvar2418,
                 reg2416,
                 forvar2415,
                 forvar2413,
                 reg2417,
                 forvar2416,
                 reg2415,
                 reg2414,
                 reg2413,
                 forvar2408,
                 reg2407,
                 reg2412,
                 reg2411,
                 reg2410,
                 reg2409,
                 reg2408,
                 forvar2407,
                 reg2406,
                 reg2405,
                 reg2404,
                 reg2403,
                 reg2402,
                 reg2401,
                 reg2400,
                 reg2399,
                 forvar2398,
                 reg2397,
                 reg2396,
                 reg2395,
                 forvar2391,
                 reg2388,
                 reg2394,
                 reg2393,
                 reg2392,
                 reg2391,
                 reg2390,
                 reg2389,
                 forvar2388,
                 forvar2384,
                 reg2383,
                 reg2387,
                 forvar2386,
                 reg2385,
                 reg2384,
                 forvar2383,
                 reg2382,
                 reg2381,
                 reg2380,
                 forvar2379,
                 forvar2378,
                 forvar2377,
                 wire2376,
                 wire2375,
                 wire2374,
                 wire2373,
                 wire2372,
                 (1'h0)};
  assign wire2372 = (^~wire2369);
  assign wire2373 = (^(wire2372 <<< (!(~&wire2370))));
  assign wire2374 = wire2371[(1'h0):(1'h0)];
  assign wire2375 = ((-(+$signed(wire2371))) ?
                        $signed($unsigned(((8'ha8) && wire2372))) : $unsigned(($signed(wire2368) ?
                            $signed((8'ha9)) : wire2373)));
  assign wire2376 = $signed(($signed((wire2370 ? wire2372 : (8'ha4))) ?
                        {(wire2374 ?
                                (8'h9d) : wire2371)} : (~|(wire2371 >>> wire2370))));
  always
    @(posedge clk) begin
      if ((($unsigned(wire2376) ?
          {(wire2372 ? wire2371 : wire2368)} : ((wire2373 ?
              wire2368 : wire2376) == $unsigned((8'ha7)))) <<< (^$signed($unsigned(wire2370)))))
        begin
          for (forvar2377 = (1'h0); (forvar2377 < (2'h3)); forvar2377 = (forvar2377 + (1'h1)))
            begin
              for (forvar2378 = (1'h0); (forvar2378 < (1'h0)); forvar2378 = (forvar2378 + (1'h1)))
                begin
                  for (forvar2379 = (1'h0); (forvar2379 < (2'h3)); forvar2379 = (forvar2379 + (1'h1)))
                    begin
                      reg2380 <= wire2370;
                      reg2381 <= ($unsigned($unsigned(wire2369)) ^~ (-((wire2368 != wire2373) ?
                          forvar2379 : (wire2368 << reg2380))));
                      reg2382 <= wire2372[(3'h7):(3'h6)];
                    end
                end
              if ((|wire2376[(1'h1):(1'h0)]))
                begin
                  for (forvar2383 = (1'h0); (forvar2383 < (1'h0)); forvar2383 = (forvar2383 + (1'h1)))
                    begin
                      reg2384 <= wire2373;
                      reg2385 <= (+reg2382);
                    end
                  for (forvar2386 = (1'h0); (forvar2386 < (1'h0)); forvar2386 = (forvar2386 + (1'h1)))
                    begin
                      reg2387 <= $signed((!($unsigned((8'ha6)) ^~ (wire2376 ?
                          reg2385 : (8'ha0)))));
                    end
                end
              else
                begin
                  if ({(+$unsigned($unsigned(forvar2386)))})
                    begin
                      reg2383 <= {$unsigned($unsigned(wire2375[(1'h1):(1'h0)]))};
                    end
                  else
                    begin
                      reg2383 <= (^~(((reg2385 ~^ reg2385) ?
                          (~wire2376) : $signed(wire2374)) >> (~^reg2384[(4'he):(4'hd)])));
                    end
                  for (forvar2384 = (1'h0); (forvar2384 < (2'h2)); forvar2384 = (forvar2384 + (1'h1)))
                    begin
                      reg2385 <= $signed($signed((wire2373 * $unsigned((8'hb5)))));
                    end
                end
              if ((~&($unsigned($signed((8'hab))) & forvar2384)))
                begin
                  for (forvar2388 = (1'h0); (forvar2388 < (2'h3)); forvar2388 = (forvar2388 + (1'h1)))
                    begin
                      reg2389 <= ((~((wire2372 ?
                          (8'h9e) : reg2387) <<< (|reg2382))) + $unsigned(($signed(wire2375) ?
                          forvar2377[(1'h1):(1'h1)] : {forvar2378})));
                      reg2390 <= (((^(wire2369 ?
                          forvar2388 : wire2372)) > wire2369[(3'h4):(3'h4)]) <= forvar2378);
                      reg2391 <= {{(forvar2377 < forvar2377[(1'h0):(1'h0)])}};
                      reg2392 <= (|{({reg2384} ?
                              (reg2381 + reg2384) : ((8'hb8) <<< forvar2386))});
                    end
                  if ($signed((^$signed(forvar2386[(1'h1):(1'h0)]))))
                    begin
                      reg2393 <= $unsigned(((reg2391[(3'h4):(3'h4)] | $unsigned(forvar2383)) - (reg2381[(3'h7):(2'h2)] ?
                          (wire2376 <<< (8'h9f)) : {reg2390})));
                      reg2394 <= $signed($unsigned(((forvar2386 || reg2389) >>> (wire2375 ?
                          (8'ha1) : wire2376))));
                    end
                  else
                    begin
                      reg2393 <= (|wire2370);
                    end
                end
              else
                begin
                  if ($unsigned($signed($signed($unsigned(forvar2378)))))
                    begin
                      reg2388 <= $unsigned({((reg2384 >>> wire2375) == (reg2393 ^ (8'hb3)))});
                    end
                  else
                    begin
                      reg2388 <= $signed($signed($signed((^reg2387))));
                      reg2389 <= reg2383[(3'h5):(3'h4)];
                      reg2390 <= (wire2372[(3'h7):(3'h5)] & $signed($unsigned($unsigned(reg2388))));
                    end
                  for (forvar2391 = (1'h0); (forvar2391 < (1'h1)); forvar2391 = (forvar2391 + (1'h1)))
                    begin
                      reg2392 <= forvar2379;
                    end
                  reg2393 <= (-{(-wire2369[(2'h2):(1'h0)])});
                  if ($signed(reg2381))
                    begin
                      reg2394 <= (~&(reg2392 && $signed((reg2384 >> reg2384))));
                      reg2395 <= $unsigned(((~&{wire2368}) < $signed((~|reg2391))));
                      reg2396 <= $signed(reg2392);
                    end
                  else
                    begin
                      reg2394 <= $unsigned(($signed({reg2387}) != (|(reg2382 == reg2389))));
                    end
                end
              reg2397 <= forvar2384;
            end
          if ({{({(8'ha2)} ? (~|wire2374) : (forvar2383 <<< reg2387))}})
            begin
              for (forvar2398 = (1'h0); (forvar2398 < (2'h3)); forvar2398 = (forvar2398 + (1'h1)))
                begin
                  reg2399 <= (8'ha4);
                  if ((~&$signed($unsigned(reg2388[(3'h7):(1'h0)]))))
                    begin
                      reg2400 <= wire2374[(3'h4):(1'h1)];
                      reg2401 <= (!reg2397[(3'h5):(2'h3)]);
                      reg2402 <= (~^$signed(forvar2383[(1'h0):(1'h0)]));
                      reg2403 <= (reg2384 >>> {$unsigned(reg2397[(3'h7):(1'h1)])});
                    end
                  else
                    begin
                      reg2400 <= ($signed(reg2381) ~^ reg2380[(1'h0):(1'h0)]);
                      reg2401 <= $unsigned((^~($unsigned(wire2373) ?
                          $signed(wire2369) : $signed(reg2387))));
                      reg2402 <= ((reg2382[(3'h5):(3'h5)] ?
                          wire2376 : forvar2378[(1'h0):(1'h0)]) < ($unsigned($signed((8'ha5))) ?
                          reg2387[(5'h10):(4'ha)] : reg2391[(4'hb):(3'h5)]));
                      reg2403 <= forvar2377[(1'h0):(1'h0)];
                    end
                end
              if (($signed(((reg2382 ? reg2401 : forvar2378) ?
                      (~^reg2399) : forvar2391[(3'h4):(1'h1)])) ?
                  (reg2402[(2'h3):(2'h2)] ?
                      $signed(((8'hb1) == wire2372)) : (reg2400[(2'h3):(2'h3)] || $unsigned(wire2374))) : $signed(({forvar2398} * $signed(reg2385)))))
                begin
                  if (($signed((-(forvar2377 >> reg2393))) ?
                      $signed((|$signed(wire2371))) : $unsigned((reg2380[(3'h5):(3'h5)] >>> $unsigned(forvar2386)))))
                    begin
                      reg2404 <= (8'h9e);
                      reg2405 <= reg2384[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg2404 <= (reg2400 ?
                          $signed(forvar2379) : (forvar2377[(1'h1):(1'h1)] >> (^wire2369)));
                      reg2405 <= $unsigned($unsigned(reg2392[(3'h6):(1'h1)]));
                      reg2406 <= $signed($signed(reg2388[(3'h6):(3'h5)]));
                    end
                  for (forvar2407 = (1'h0); (forvar2407 < (2'h3)); forvar2407 = (forvar2407 + (1'h1)))
                    begin
                      reg2408 <= ({((~|reg2396) ?
                              ((8'hba) == reg2382) : $signed(forvar2386))} | (wire2373 ?
                          $unsigned({forvar2384}) : reg2396[(4'h9):(1'h1)]));
                      reg2409 <= reg2390[(1'h0):(1'h0)];
                    end
                  if (reg2401)
                    begin
                      reg2410 <= reg2403;
                      reg2411 <= $unsigned($unsigned(($unsigned(forvar2386) ^ ((8'hba) ?
                          wire2375 : forvar2388))));
                      reg2412 <= (^$unsigned($signed(reg2393)));
                    end
                  else
                    begin
                      reg2410 <= ($unsigned(forvar2407) ?
                          reg2396 : wire2368[(3'h6):(1'h1)]);
                    end
                end
              else
                begin
                  if (forvar2377[(3'h5):(3'h5)])
                    begin
                      reg2404 <= forvar2407[(2'h2):(1'h0)];
                      reg2405 <= (~&$unsigned(((forvar2388 ?
                              reg2388 : forvar2378) ?
                          $signed(forvar2391) : forvar2377)));
                      reg2406 <= $signed(wire2370);
                      reg2407 <= $signed($unsigned(forvar2407[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg2404 <= $signed((((&reg2383) ?
                          reg2394[(2'h2):(1'h0)] : ((8'hb2) ?
                              wire2368 : reg2393)) != (reg2392 ?
                          reg2394[(2'h2):(2'h2)] : $unsigned((8'h9d)))));
                      reg2405 <= (forvar2384[(1'h1):(1'h0)] ?
                          $signed(((^forvar2384) ?
                              {reg2382} : ((8'hb3) >>> (8'hab)))) : ({(forvar2383 && wire2374)} + ($signed((8'hb5)) - forvar2407)));
                      reg2406 <= $signed(wire2371);
                    end
                  for (forvar2408 = (1'h0); (forvar2408 < (1'h0)); forvar2408 = (forvar2408 + (1'h1)))
                    begin
                      reg2409 <= $unsigned($unsigned((8'hb4)));
                    end
                end
              if ($signed($unsigned({{wire2369}})))
                begin
                  if ($signed((!({forvar2407} ?
                      $unsigned(reg2401) : (reg2390 ? forvar2407 : reg2380)))))
                    begin
                      reg2413 <= wire2376[(3'h7):(3'h5)];
                    end
                  else
                    begin
                      reg2413 <= $signed((-(reg2392[(4'hc):(3'h6)] ?
                          wire2376[(3'h6):(2'h2)] : $unsigned(wire2374))));
                      reg2414 <= ((reg2389 ?
                              (reg2401[(4'hc):(4'h8)] < wire2372) : $unsigned($unsigned(reg2396))) ?
                          (reg2404[(1'h0):(1'h0)] ?
                              {(~|reg2404)} : $signed({(8'h9e)})) : reg2388);
                      reg2415 <= $signed((reg2405 ?
                          $unsigned((forvar2398 ?
                              forvar2407 : (8'hb7))) : reg2411));
                    end
                  for (forvar2416 = (1'h0); (forvar2416 < (1'h1)); forvar2416 = (forvar2416 + (1'h1)))
                    begin
                      reg2417 <= ($unsigned((|(reg2402 ? reg2399 : (8'hb5)))) ?
                          (!$signed((reg2387 ?
                              wire2372 : reg2405))) : (((^forvar2377) ?
                              $signed(forvar2377) : (reg2388 <= wire2368)) <= (reg2397 <= (reg2381 ?
                              (8'hae) : forvar2398))));
                    end
                end
              else
                begin
                  for (forvar2413 = (1'h0); (forvar2413 < (2'h2)); forvar2413 = (forvar2413 + (1'h1)))
                    begin
                      reg2414 <= $signed(reg2417[(2'h2):(1'h1)]);
                    end
                  for (forvar2415 = (1'h0); (forvar2415 < (2'h3)); forvar2415 = (forvar2415 + (1'h1)))
                    begin
                      reg2416 <= $unsigned($signed(((forvar2407 != reg2411) << $unsigned(wire2368))));
                      reg2417 <= $signed(forvar2413);
                    end
                  for (forvar2418 = (1'h0); (forvar2418 < (1'h1)); forvar2418 = (forvar2418 + (1'h1)))
                    begin
                      reg2419 <= {forvar2407[(2'h2):(1'h1)]};
                    end
                end
            end
          else
            begin
              reg2398 <= (|{$signed((forvar2415 ^~ forvar2378))});
            end
          if (reg2413[(1'h1):(1'h0)])
            begin
              if (((-$unsigned((&(8'h9c)))) ?
                  (&$signed({reg2406})) : $signed({$signed(reg2382)})))
                begin
                  if ((~|((~&(-(8'ha6))) ?
                      $signed(reg2385[(3'h6):(3'h5)]) : ((!reg2415) ?
                          ((8'h9e) ? reg2390 : (8'ha0)) : {reg2388}))))
                    begin
                      reg2420 <= (+$signed($unsigned(reg2394[(3'h7):(3'h7)])));
                      reg2421 <= reg2405[(2'h3):(1'h0)];
                      reg2422 <= (((&(reg2382 <<< reg2383)) * reg2414) + $unsigned((forvar2416 ?
                          reg2404 : forvar2398[(4'hb):(4'h8)])));
                    end
                  else
                    begin
                      reg2420 <= (reg2400 ^~ wire2371[(2'h2):(1'h0)]);
                    end
                  for (forvar2423 = (1'h0); (forvar2423 < (2'h2)); forvar2423 = (forvar2423 + (1'h1)))
                    begin
                      reg2424 <= forvar2415[(4'h8):(1'h0)];
                      reg2425 <= forvar2398[(3'h6):(3'h4)];
                      reg2426 <= reg2408[(2'h3):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar2420 = (1'h0); (forvar2420 < (2'h3)); forvar2420 = (forvar2420 + (1'h1)))
                    begin
                      reg2421 <= (~^($signed((~&reg2419)) ?
                          $signed((reg2381 >= wire2374)) : $unsigned((reg2380 ^ reg2426))));
                      reg2422 <= ($signed(($signed(reg2391) > forvar2398[(1'h1):(1'h0)])) ?
                          (reg2408 ?
                              $unsigned(wire2371[(3'h5):(1'h0)]) : wire2370) : (+forvar2386[(4'ha):(3'h4)]));
                      reg2423 <= (wire2374 ?
                          (reg2392 != $unsigned((reg2409 <= (8'ha6)))) : reg2380);
                      reg2424 <= ($signed((forvar2391[(2'h3):(1'h0)] ^ forvar2377[(3'h4):(1'h1)])) >> ({wire2376[(4'ha):(4'h8)]} ?
                          reg2402 : (forvar2378[(1'h0):(1'h0)] ?
                              (wire2376 ^ reg2402) : $signed((8'h9e)))));
                    end
                  if ($signed(((~reg2383[(3'h6):(1'h0)]) ?
                      wire2371 : (wire2374[(3'h4):(2'h2)] | reg2394[(3'h7):(3'h6)]))))
                    begin
                      reg2425 <= (($unsigned($unsigned(reg2397)) != ($signed(reg2396) ~^ (reg2392 ?
                              (8'ha7) : forvar2407))) ?
                          $unsigned((&forvar2388[(3'h7):(3'h7)])) : (^~(~&$unsigned(forvar2408))));
                      reg2426 <= $signed(forvar2377[(1'h1):(1'h0)]);
                      reg2427 <= ((reg2423[(1'h1):(1'h0)] << reg2383) ?
                          $unsigned(($signed(forvar2388) <= $signed(reg2409))) : ($unsigned($unsigned(wire2372)) | ((wire2369 ^ wire2373) ?
                              $signed(reg2416) : ((8'h9e) ?
                                  (8'ha7) : reg2384))));
                    end
                  else
                    begin
                      reg2425 <= {$signed($signed({reg2415}))};
                      reg2426 <= $unsigned(reg2409[(2'h2):(1'h1)]);
                      reg2427 <= {($signed((reg2427 ^~ reg2397)) ~^ $signed(reg2391[(1'h0):(1'h0)]))};
                    end
                  reg2428 <= reg2383;
                  reg2429 <= $signed(forvar2386);
                end
              if ((((^reg2391) <<< (forvar2408 ~^ {reg2401})) << reg2396))
                begin
                  if (forvar2383[(1'h1):(1'h0)])
                    begin
                      reg2430 <= {(+reg2390)};
                      reg2431 <= (!(((^reg2389) ?
                          $unsigned(wire2371) : (-(8'hac))) * (~|$signed(reg2404))));
                      reg2432 <= (reg2413 ?
                          (forvar2407 <= ($signed(forvar2383) >> {wire2371})) : (|((wire2373 ?
                                  reg2428 : reg2393) ?
                              reg2411 : reg2412[(3'h4):(3'h4)])));
                      reg2433 <= (-forvar2383);
                    end
                  else
                    begin
                      reg2430 <= (|reg2409[(1'h0):(1'h0)]);
                      reg2431 <= reg2409;
                      reg2432 <= forvar2377[(2'h3):(1'h0)];
                    end
                  for (forvar2434 = (1'h0); (forvar2434 < (1'h1)); forvar2434 = (forvar2434 + (1'h1)))
                    begin
                      reg2435 <= (({reg2417} - $unsigned(reg2413[(1'h1):(1'h1)])) && forvar2434[(1'h0):(1'h0)]);
                    end
                  if (((8'ha2) >>> forvar2418[(1'h1):(1'h1)]))
                    begin
                      reg2436 <= $signed((((8'ha2) ?
                          ((8'haf) && reg2399) : (reg2405 & reg2426)) == $unsigned({reg2382})));
                      reg2437 <= reg2403;
                    end
                  else
                    begin
                      reg2436 <= $unsigned($signed((-(reg2432 ?
                          forvar2434 : forvar2420))));
                      reg2437 <= $unsigned((($unsigned(reg2406) ?
                          $unsigned(forvar2420) : (reg2431 << reg2392)) <<< $signed($signed(wire2369))));
                    end
                end
              else
                begin
                  if ({{($unsigned(forvar2415) | (8'hb6))}})
                    begin
                      reg2430 <= ($unsigned((~&{reg2396})) ?
                          (^((reg2421 ?
                              forvar2416 : forvar2378) ~^ {reg2421})) : ((forvar2407[(2'h2):(1'h1)] ?
                                  (reg2399 ?
                                      reg2425 : (8'hba)) : $unsigned(reg2394)) ?
                              forvar2383[(1'h0):(1'h0)] : wire2375));
                      reg2431 <= ($unsigned($signed((~&reg2399))) & forvar2413[(4'h9):(1'h0)]);
                      reg2432 <= $unsigned(reg2420);
                    end
                  else
                    begin
                      reg2430 <= (({reg2407} ?
                          (+$signed(reg2419)) : $signed(reg2407)) ~^ wire2374);
                      reg2431 <= $signed((^~((8'h9f) ?
                          (forvar2398 ? reg2403 : forvar2407) : reg2429)));
                      reg2432 <= ((wire2374[(1'h0):(1'h0)] ?
                          $unsigned($signed((8'ha2))) : ((reg2436 ?
                                  reg2437 : reg2402) ?
                              reg2407 : (forvar2418 ~^ reg2381))) ~^ (~^{(reg2409 << reg2437)}));
                    end
                  for (forvar2433 = (1'h0); (forvar2433 < (2'h2)); forvar2433 = (forvar2433 + (1'h1)))
                    begin
                      reg2434 <= (~&(^~(wire2371 ?
                          $signed((8'ha9)) : (reg2435 == reg2381))));
                      reg2435 <= $unsigned(reg2417);
                      reg2436 <= (!((forvar2418[(2'h2):(1'h0)] << $unsigned(reg2405)) - (^~reg2437[(2'h3):(2'h3)])));
                      reg2437 <= wire2375;
                    end
                  for (forvar2438 = (1'h0); (forvar2438 < (2'h3)); forvar2438 = (forvar2438 + (1'h1)))
                    begin
                      reg2439 <= reg2409[(2'h2):(1'h0)];
                      reg2440 <= reg2416[(2'h2):(1'h1)];
                      reg2441 <= reg2381[(3'h5):(3'h5)];
                      reg2442 <= $unsigned(((^{reg2404}) >> (~(~reg2428))));
                    end
                  for (forvar2443 = (1'h0); (forvar2443 < (2'h3)); forvar2443 = (forvar2443 + (1'h1)))
                    begin
                      reg2444 <= {reg2413};
                    end
                end
            end
          else
            begin
              if ($signed((8'haa)))
                begin
                  for (forvar2420 = (1'h0); (forvar2420 < (2'h3)); forvar2420 = (forvar2420 + (1'h1)))
                    begin
                      reg2421 <= ((wire2371 == {$signed(forvar2408)}) + (!reg2422));
                    end
                  for (forvar2422 = (1'h0); (forvar2422 < (1'h0)); forvar2422 = (forvar2422 + (1'h1)))
                    begin
                      reg2423 <= reg2384[(5'h10):(2'h2)];
                    end
                end
              else
                begin
                  reg2420 <= $unsigned(reg2426);
                  reg2421 <= reg2410[(2'h2):(1'h0)];
                  for (forvar2422 = (1'h0); (forvar2422 < (1'h1)); forvar2422 = (forvar2422 + (1'h1)))
                    begin
                      reg2423 <= reg2411[(4'hb):(3'h5)];
                      reg2424 <= ({((reg2444 ?
                              reg2400 : forvar2416) == reg2437)} * (($unsigned(reg2384) > reg2414[(3'h4):(2'h2)]) ?
                          reg2394 : ((!forvar2377) <= $signed((8'h9e)))));
                    end
                  if (((~|(8'h9e)) | (!(~^(8'ha1)))))
                    begin
                      reg2425 <= ($signed((^wire2374[(1'h0):(1'h0)])) != ((reg2388[(3'h6):(2'h3)] > (reg2414 ?
                          reg2419 : wire2374)) >= reg2405[(4'ha):(1'h0)]));
                    end
                  else
                    begin
                      reg2425 <= $unsigned(forvar2413[(4'hd):(4'hb)]);
                      reg2426 <= reg2419[(3'h7):(1'h0)];
                      reg2427 <= (~|(&(&reg2408)));
                    end
                end
              for (forvar2428 = (1'h0); (forvar2428 < (2'h3)); forvar2428 = (forvar2428 + (1'h1)))
                begin
                  if (($signed($signed(reg2430)) ?
                      (forvar2443 ?
                          forvar2416 : $unsigned($signed(wire2375))) : (reg2400 ?
                          reg2403 : $unsigned((reg2380 < forvar2384)))))
                    begin
                      reg2429 <= ($unsigned((8'ha8)) != $unsigned(($unsigned(reg2429) <<< (reg2411 << (8'hac)))));
                      reg2430 <= ((reg2435 ?
                              $signed((~reg2387)) : ((forvar2438 >= (8'hb7)) >> (+reg2400))) ?
                          wire2376[(3'h7):(2'h3)] : (8'h9d));
                    end
                  else
                    begin
                      reg2429 <= ((+($signed(reg2433) >= $signed(wire2375))) << reg2406[(4'ha):(3'h6)]);
                    end
                end
            end
        end
      else
        begin
          if (reg2406)
            begin
              for (forvar2377 = (1'h0); (forvar2377 < (1'h1)); forvar2377 = (forvar2377 + (1'h1)))
                begin
                  reg2378 <= (~|forvar2378);
                  for (forvar2379 = (1'h0); (forvar2379 < (2'h2)); forvar2379 = (forvar2379 + (1'h1)))
                    begin
                      reg2380 <= ((8'hab) ?
                          (forvar2418[(1'h0):(1'h0)] ?
                              ((reg2402 ? forvar2434 : forvar2413) ?
                                  wire2373[(4'hc):(4'h9)] : (forvar2416 ?
                                      wire2368 : reg2382)) : wire2371) : $signed((~|(^~reg2388))));
                      reg2381 <= {(^reg2433[(3'h7):(2'h2)])};
                    end
                end
              if ((8'ha9))
                begin
                  reg2382 <= reg2440;
                  reg2383 <= $unsigned(($unsigned((forvar2434 << reg2439)) & $unsigned(reg2416[(2'h2):(2'h2)])));
                end
              else
                begin
                  for (forvar2382 = (1'h0); (forvar2382 < (2'h3)); forvar2382 = (forvar2382 + (1'h1)))
                    begin
                      reg2383 <= (!(8'hb6));
                      reg2384 <= $signed($signed(reg2425[(4'hb):(4'ha)]));
                    end
                  for (forvar2385 = (1'h0); (forvar2385 < (2'h3)); forvar2385 = (forvar2385 + (1'h1)))
                    begin
                      reg2386 <= $unsigned($signed(reg2382[(2'h2):(1'h0)]));
                      reg2387 <= (($unsigned($unsigned(forvar2407)) ?
                          (^~(~forvar2418)) : (+reg2410[(1'h0):(1'h0)])) ^~ ((8'ha8) ?
                          (8'hab) : (+(reg2405 > reg2383))));
                      reg2388 <= reg2391[(4'ha):(4'ha)];
                    end
                  for (forvar2389 = (1'h0); (forvar2389 < (2'h2)); forvar2389 = (forvar2389 + (1'h1)))
                    begin
                      reg2390 <= forvar2428[(1'h0):(1'h0)];
                    end
                end
              for (forvar2391 = (1'h0); (forvar2391 < (1'h1)); forvar2391 = (forvar2391 + (1'h1)))
                begin
                  if ($signed({$unsigned(((8'hb4) ? reg2408 : reg2420))}))
                    begin
                      reg2392 <= ({$signed(reg2410[(2'h2):(1'h1)])} ?
                          (reg2384[(4'hd):(3'h5)] != ((8'haf) ?
                              $unsigned(reg2410) : forvar2433)) : (~&$unsigned(reg2440)));
                    end
                  else
                    begin
                      reg2392 <= $signed(($unsigned({reg2415}) ?
                          {reg2435} : (reg2399 ?
                              (~reg2398) : reg2383[(3'h4):(2'h2)])));
                      reg2393 <= $unsigned(forvar2408[(1'h0):(1'h0)]);
                    end
                  for (forvar2394 = (1'h0); (forvar2394 < (2'h2)); forvar2394 = (forvar2394 + (1'h1)))
                    begin
                      reg2395 <= ((^~reg2414) ?
                          {$unsigned((reg2392 ?
                                  (8'ha6) : reg2395))} : (((reg2435 ~^ (8'hb5)) ?
                                  $unsigned(forvar2385) : $signed((8'h9f))) ?
                              reg2411[(3'h4):(1'h0)] : {reg2426[(1'h0):(1'h0)]}));
                      reg2396 <= forvar2443[(4'h8):(2'h2)];
                    end
                end
              for (forvar2397 = (1'h0); (forvar2397 < (2'h3)); forvar2397 = (forvar2397 + (1'h1)))
                begin
                  if (reg2440[(4'hd):(3'h6)])
                    begin
                      reg2398 <= {(^~($unsigned(reg2394) + {forvar2389}))};
                      reg2399 <= wire2374[(1'h0):(1'h0)];
                      reg2400 <= $signed(forvar2434[(1'h0):(1'h0)]);
                      reg2401 <= ($unsigned((forvar2422[(3'h6):(2'h3)] * (8'ha1))) == reg2384[(5'h10):(4'h8)]);
                    end
                  else
                    begin
                      reg2398 <= $unsigned((-{reg2383}));
                    end
                end
            end
          else
            begin
              if ({reg2404})
                begin
                  if (((~{(reg2432 ? reg2407 : reg2444)}) | $unsigned(reg2391)))
                    begin
                      reg2377 <= {(((reg2381 - reg2437) != (reg2401 * forvar2391)) ?
                              forvar2443 : ((reg2411 ^ reg2440) ?
                                  (8'ha7) : $signed(wire2368)))};
                      reg2378 <= $unsigned((({forvar2433} != reg2399) ^ (~|reg2393[(3'h7):(2'h2)])));
                    end
                  else
                    begin
                      reg2377 <= (^(8'ha0));
                      reg2378 <= (~(~&wire2372));
                    end
                  if (((forvar2377[(2'h2):(2'h2)] ^ wire2372[(4'h9):(3'h6)]) ^~ (+forvar2408[(2'h2):(2'h2)])))
                    begin
                      reg2379 <= reg2440[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg2379 <= $signed(reg2423);
                      reg2380 <= (^~$signed({(~^forvar2398)}));
                      reg2381 <= $signed((reg2415 ?
                          ($signed(forvar2397) << (reg2390 ^~ forvar2443)) : $signed($signed((8'had)))));
                      reg2382 <= ({$unsigned((forvar2388 + reg2389))} <<< (~&reg2379[(3'h5):(1'h0)]));
                    end
                  if ((~&reg2435[(2'h3):(1'h0)]))
                    begin
                      reg2383 <= (&($unsigned($signed(reg2403)) ?
                          reg2429 : {(reg2378 * wire2369)}));
                      reg2384 <= wire2370[(1'h0):(1'h0)];
                      reg2385 <= $signed(($signed($signed(reg2395)) >>> (~^$unsigned(forvar2416))));
                      reg2386 <= (+((~^(forvar2407 ?
                          forvar2397 : reg2405)) ~^ reg2415));
                    end
                  else
                    begin
                      reg2383 <= $signed(forvar2416[(2'h3):(2'h2)]);
                      reg2384 <= (&($signed((~|wire2373)) ~^ ($unsigned(reg2428) ?
                          (reg2424 ? (8'ha2) : reg2407) : $signed(reg2423))));
                    end
                  for (forvar2387 = (1'h0); (forvar2387 < (2'h3)); forvar2387 = (forvar2387 + (1'h1)))
                    begin
                      reg2388 <= $unsigned({$unsigned(reg2387[(4'he):(3'h6)])});
                      reg2389 <= (+$signed($unsigned($unsigned((8'hb3)))));
                      reg2390 <= $unsigned((8'ha9));
                      reg2391 <= (^$signed(((reg2410 ^~ (8'hb6)) ?
                          ((8'haf) ?
                              reg2428 : forvar2389) : $unsigned(forvar2423))));
                    end
                end
              else
                begin
                  reg2377 <= (forvar2433 ^~ $signed(forvar2389));
                  reg2378 <= (~&{forvar2397[(3'h4):(2'h2)]});
                  if ($signed($signed($signed(reg2427))))
                    begin
                      reg2379 <= $signed((reg2412[(3'h4):(2'h2)] || reg2428[(2'h3):(1'h0)]));
                      reg2380 <= (forvar2398 < $signed(({forvar2428} ?
                          $signed(reg2433) : wire2376)));
                      reg2381 <= (|$signed(forvar2378[(3'h4):(2'h3)]));
                      reg2382 <= ($signed((8'haa)) ?
                          reg2400[(2'h2):(2'h2)] : $unsigned(forvar2408));
                    end
                  else
                    begin
                      reg2379 <= (|($signed(reg2412[(2'h2):(1'h1)]) ?
                          forvar2438[(1'h0):(1'h0)] : {$signed(reg2381)}));
                      reg2380 <= reg2403;
                      reg2381 <= $unsigned((!forvar2418));
                      reg2382 <= reg2425;
                    end
                  if ((((-(^~reg2410)) ?
                      {(wire2376 && forvar2420)} : {forvar2415}) ^ ((+(wire2370 ?
                          reg2442 : (8'ha8))) ?
                      $signed((forvar2434 ?
                          reg2392 : reg2423)) : ($signed(reg2403) >= {reg2410}))))
                    begin
                      reg2383 <= (8'hb7);
                      reg2384 <= {{(|reg2442[(1'h1):(1'h0)])}};
                      reg2385 <= ($signed(((reg2385 ?
                          (8'hae) : forvar2434) >= reg2384)) ~^ (~^(~^(reg2422 - reg2428))));
                      reg2386 <= ({$signed((~&reg2423))} | forvar2387[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg2383 <= $signed($signed($unsigned($signed(reg2403))));
                      reg2384 <= (!$unsigned(reg2410));
                    end
                end
            end
          reg2402 <= ($signed(wire2371[(3'h4):(3'h4)]) ? wire2368 : reg2423);
        end
      if ({(!($signed(forvar2382) && reg2417[(2'h3):(2'h3)]))})
        begin
          if (reg2390)
            begin
              if ($signed($unsigned((8'hb7))))
                begin
                  for (forvar2445 = (1'h0); (forvar2445 < (2'h2)); forvar2445 = (forvar2445 + (1'h1)))
                    begin
                      reg2446 <= $unsigned((((|forvar2388) ?
                              forvar2377 : forvar2433) ?
                          (~&reg2441) : {$signed(reg2444)}));
                      reg2447 <= (|forvar2415[(4'hd):(4'h8)]);
                      reg2448 <= (~^(~^reg2396));
                      reg2449 <= forvar2433[(2'h3):(2'h2)];
                    end
                  for (forvar2450 = (1'h0); (forvar2450 < (2'h3)); forvar2450 = (forvar2450 + (1'h1)))
                    begin
                      reg2451 <= reg2395;
                      reg2452 <= (~&{reg2434});
                      reg2453 <= forvar2420;
                    end
                  if ($signed(forvar2391[(1'h1):(1'h0)]))
                    begin
                      reg2454 <= {forvar2388};
                      reg2455 <= ({reg2426} * (&reg2377[(1'h0):(1'h0)]));
                      reg2456 <= reg2451;
                    end
                  else
                    begin
                      reg2454 <= (reg2405[(3'h4):(1'h0)] * reg2453);
                      reg2455 <= $signed((forvar2387[(1'h1):(1'h0)] <= forvar2413[(4'hd):(4'hc)]));
                    end
                end
              else
                begin
                  for (forvar2445 = (1'h0); (forvar2445 < (1'h1)); forvar2445 = (forvar2445 + (1'h1)))
                    begin
                      reg2446 <= ($unsigned($unsigned(forvar2416)) ?
                          $unsigned($unsigned((-forvar2388))) : wire2375[(1'h1):(1'h0)]);
                      reg2447 <= reg2422;
                      reg2448 <= reg2423;
                      reg2449 <= $unsigned((($signed((8'hb8)) ?
                              ((8'hb2) <= reg2454) : (reg2411 ?
                                  forvar2383 : reg2417)) ?
                          reg2387[(5'h10):(4'he)] : reg2455));
                    end
                end
            end
          else
            begin
              for (forvar2445 = (1'h0); (forvar2445 < (1'h1)); forvar2445 = (forvar2445 + (1'h1)))
                begin
                  for (forvar2446 = (1'h0); (forvar2446 < (2'h2)); forvar2446 = (forvar2446 + (1'h1)))
                    begin
                      reg2447 <= ((&$signed((reg2393 ? wire2374 : wire2369))) ?
                          $unsigned(($signed(reg2378) + (^(8'hba)))) : (reg2392 | (~|$unsigned((8'hb4)))));
                      reg2448 <= (~$unsigned((~&(reg2442 ?
                          reg2408 : forvar2450))));
                    end
                  for (forvar2449 = (1'h0); (forvar2449 < (2'h2)); forvar2449 = (forvar2449 + (1'h1)))
                    begin
                      reg2450 <= reg2421[(1'h0):(1'h0)];
                      reg2451 <= (&$unsigned(((8'hb2) ?
                          (reg2450 ~^ reg2454) : ((8'ha0) ?
                              (8'ha1) : forvar2434))));
                    end
                  for (forvar2452 = (1'h0); (forvar2452 < (2'h2)); forvar2452 = (forvar2452 + (1'h1)))
                    begin
                      reg2453 <= (|$signed($unsigned((wire2373 <<< wire2375))));
                      reg2454 <= ($signed((&(forvar2443 ? reg2408 : reg2441))) ?
                          $unsigned(reg2434[(1'h1):(1'h1)]) : reg2407);
                      reg2455 <= (($unsigned({reg2412}) ?
                              ({reg2388} ?
                                  reg2455[(3'h7):(3'h6)] : $unsigned(forvar2386)) : reg2377[(3'h6):(3'h4)]) ?
                          $signed(reg2408[(2'h2):(2'h2)]) : (($signed((8'haa)) ^~ {(8'ha4)}) ?
                              reg2455 : $signed($signed(forvar2388))));
                      reg2456 <= reg2423[(1'h0):(1'h0)];
                    end
                  for (forvar2457 = (1'h0); (forvar2457 < (2'h3)); forvar2457 = (forvar2457 + (1'h1)))
                    begin
                      reg2458 <= reg2411;
                      reg2459 <= {reg2403};
                      reg2460 <= ($unsigned(({reg2387} || $unsigned(reg2424))) - (+{reg2381}));
                      reg2461 <= {reg2449};
                    end
                end
            end
        end
      else
        begin
          if (reg2456)
            begin
              reg2445 <= (reg2377 ?
                  (reg2397[(2'h2):(2'h2)] <= (8'hb4)) : $signed(forvar2428[(3'h5):(2'h3)]));
            end
          else
            begin
              if ($unsigned(reg2437))
                begin
                  for (forvar2445 = (1'h0); (forvar2445 < (1'h1)); forvar2445 = (forvar2445 + (1'h1)))
                    begin
                      reg2446 <= (+reg2421[(1'h1):(1'h0)]);
                      reg2447 <= reg2458[(3'h5):(3'h5)];
                    end
                  for (forvar2448 = (1'h0); (forvar2448 < (2'h2)); forvar2448 = (forvar2448 + (1'h1)))
                    begin
                      reg2449 <= ($unsigned((&$signed(wire2373))) ?
                          ((forvar2388 == wire2368[(3'h7):(3'h6)]) ?
                              reg2453[(4'h8):(1'h1)] : $signed((reg2400 <<< (8'hba)))) : $signed(((reg2380 <<< forvar2445) != $signed(reg2450))));
                      reg2450 <= reg2426;
                      reg2451 <= (^((!(&reg2387)) ?
                          (~|$signed(reg2414)) : $unsigned(forvar2388[(4'h8):(2'h2)])));
                    end
                  for (forvar2452 = (1'h0); (forvar2452 < (2'h2)); forvar2452 = (forvar2452 + (1'h1)))
                    begin
                      reg2453 <= (forvar2385 && $signed((|$signed(reg2413))));
                      reg2454 <= (reg2390[(1'h1):(1'h0)] ?
                          ((~(+reg2390)) | reg2422) : forvar2398);
                      reg2455 <= $signed(reg2396);
                    end
                  reg2456 <= ((((-reg2382) ?
                          (wire2368 ? (8'h9e) : (8'hb7)) : ((8'ha7) ?
                              wire2374 : reg2430)) ^ ((wire2371 ^~ reg2432) >>> (forvar2397 <= reg2430))) ?
                      $signed($signed({reg2382})) : $unsigned($signed((forvar2438 | (8'ha2)))));
                end
              else
                begin
                  if ($signed({(!(~|wire2376))}))
                    begin
                      reg2445 <= $unsigned(forvar2434[(4'he):(3'h4)]);
                      reg2446 <= wire2369;
                      reg2447 <= reg2446;
                    end
                  else
                    begin
                      reg2445 <= forvar2457;
                    end
                  if (((^(+(~&(8'ha4)))) <<< reg2408))
                    begin
                      reg2448 <= $unsigned(((reg2437 ?
                          (reg2404 >= reg2442) : (~^wire2370)) | (wire2369 * $unsigned(reg2401))));
                    end
                  else
                    begin
                      reg2448 <= $unsigned((((!reg2409) ?
                          $signed(reg2404) : (reg2400 >>> reg2451)) || reg2429[(3'h6):(3'h6)]));
                      reg2449 <= $signed($signed($signed((wire2369 >>> forvar2387))));
                    end
                  if (($unsigned(reg2456[(3'h6):(3'h5)]) ?
                      {((reg2430 <= reg2381) >>> (forvar2449 ?
                              reg2403 : (8'hb6)))} : (reg2427 ?
                          ($signed(reg2446) << (reg2407 ^~ reg2416)) : $signed($unsigned(forvar2422)))))
                    begin
                      reg2450 <= forvar2379;
                      reg2451 <= (reg2459[(1'h0):(1'h0)] || $signed(forvar2385[(2'h2):(2'h2)]));
                      reg2452 <= ($unsigned({(8'haa)}) ?
                          ($unsigned($unsigned(reg2392)) - {(forvar2378 <= forvar2384)}) : (!(-(reg2387 ^ reg2444))));
                      reg2453 <= {(&((reg2423 ? forvar2384 : reg2432) ?
                              {wire2374} : (forvar2387 ? reg2434 : reg2452)))};
                    end
                  else
                    begin
                      reg2450 <= reg2380;
                    end
                  reg2454 <= $unsigned(((-(~&reg2449)) + $unsigned(reg2378[(4'hb):(4'hb)])));
                end
              for (forvar2457 = (1'h0); (forvar2457 < (2'h2)); forvar2457 = (forvar2457 + (1'h1)))
                begin
                  if ((reg2454[(1'h1):(1'h0)] == ($unsigned((wire2373 ?
                      (8'hb5) : reg2380)) != $signed(((8'ha4) ?
                      reg2455 : forvar2407)))))
                    begin
                      reg2458 <= ((+reg2453[(1'h1):(1'h0)]) ?
                          {$unsigned(forvar2385)} : (8'ha9));
                      reg2459 <= (+(^{$signed((8'ha4))}));
                      reg2460 <= $unsigned($signed(forvar2386));
                      reg2461 <= (($signed((reg2422 >> reg2381)) >= ($signed(reg2392) != wire2372[(3'h7):(1'h0)])) ?
                          $signed((~|(+(8'haa)))) : (reg2423 + {(reg2434 <= reg2415)}));
                    end
                  else
                    begin
                      reg2458 <= ($signed({((8'haf) ?
                              forvar2387 : reg2422)}) < forvar2423[(2'h2):(2'h2)]);
                      reg2459 <= forvar2378;
                      reg2460 <= reg2456;
                    end
                  if ((forvar2418[(1'h1):(1'h1)] | (reg2395[(1'h1):(1'h1)] ?
                      $unsigned(reg2430) : (wire2373 || (wire2370 || reg2404)))))
                    begin
                      reg2462 <= (!(($unsigned(reg2404) ?
                              (reg2387 && forvar2383) : (reg2380 ?
                                  reg2442 : forvar2443)) ?
                          ($unsigned(wire2374) ?
                              (^~reg2422) : reg2382[(3'h4):(1'h0)]) : (reg2392 - $signed(reg2420))));
                      reg2463 <= (~|$unsigned($signed($signed(reg2447))));
                      reg2464 <= $unsigned((^(8'had)));
                    end
                  else
                    begin
                      reg2462 <= {(((forvar2416 ?
                              reg2448 : reg2458) != reg2435[(1'h0):(1'h0)]) + ((-reg2435) ?
                              forvar2386 : (reg2388 ? reg2420 : reg2409)))};
                      reg2463 <= reg2381;
                    end
                  for (forvar2465 = (1'h0); (forvar2465 < (2'h2)); forvar2465 = (forvar2465 + (1'h1)))
                    begin
                      reg2466 <= $unsigned(wire2376);
                      reg2467 <= (reg2448 ?
                          ((~(reg2434 | reg2428)) != ((&reg2426) ?
                              {reg2392} : (reg2393 ?
                                  forvar2434 : reg2431))) : reg2383[(2'h3):(1'h1)]);
                    end
                  if (reg2432)
                    begin
                      reg2468 <= reg2406[(1'h0):(1'h0)];
                      reg2469 <= {$signed((|(reg2421 ^~ forvar2452)))};
                      reg2470 <= {($signed($signed(forvar2423)) ^~ wire2374[(2'h3):(1'h0)])};
                    end
                  else
                    begin
                      reg2468 <= reg2426;
                      reg2469 <= reg2422[(1'h0):(1'h0)];
                      reg2470 <= reg2388;
                      reg2471 <= (~^$unsigned(reg2403[(3'h4):(2'h2)]));
                    end
                end
              for (forvar2472 = (1'h0); (forvar2472 < (1'h0)); forvar2472 = (forvar2472 + (1'h1)))
                begin
                  for (forvar2473 = (1'h0); (forvar2473 < (2'h3)); forvar2473 = (forvar2473 + (1'h1)))
                    begin
                      reg2474 <= $signed($unsigned($signed({reg2444})));
                      reg2475 <= (^~(reg2415 * reg2417));
                      reg2476 <= $signed(forvar2379[(3'h5):(2'h2)]);
                      reg2477 <= forvar2386[(3'h5):(3'h5)];
                    end
                  if ((forvar2377[(2'h3):(1'h1)] >>> wire2371))
                    begin
                      reg2478 <= forvar2382;
                      reg2479 <= ((!(forvar2398 & $unsigned(forvar2449))) << $signed($signed($unsigned(reg2381))));
                      reg2480 <= forvar2449;
                    end
                  else
                    begin
                      reg2478 <= (&wire2374[(2'h2):(2'h2)]);
                    end
                end
              reg2481 <= forvar2433;
            end
          for (forvar2482 = (1'h0); (forvar2482 < (2'h3)); forvar2482 = (forvar2482 + (1'h1)))
            begin
              reg2483 <= wire2373[(4'ha):(4'ha)];
              reg2484 <= ($unsigned(((^forvar2418) == wire2372)) ?
                  {$signed($unsigned(forvar2389))} : ({forvar2472[(3'h6):(3'h5)]} ?
                      wire2369[(1'h1):(1'h0)] : $unsigned(((8'ha2) != reg2448))));
              for (forvar2485 = (1'h0); (forvar2485 < (1'h1)); forvar2485 = (forvar2485 + (1'h1)))
                begin
                  for (forvar2486 = (1'h0); (forvar2486 < (2'h2)); forvar2486 = (forvar2486 + (1'h1)))
                    begin
                      reg2487 <= forvar2394;
                    end
                  if ({$unsigned((8'had))})
                    begin
                      reg2488 <= $signed($signed($signed((reg2476 - forvar2378))));
                      reg2489 <= (^~({(~reg2388)} & $signed((reg2422 ?
                          forvar2397 : reg2450))));
                      reg2490 <= (+({reg2466} ?
                          $unsigned(reg2403) : (~^$unsigned(forvar2387))));
                      reg2491 <= reg2442;
                    end
                  else
                    begin
                      reg2488 <= (~&(reg2478[(4'he):(4'he)] ^~ $signed(reg2428[(1'h0):(1'h0)])));
                      reg2489 <= reg2463[(3'h6):(3'h4)];
                    end
                  for (forvar2492 = (1'h0); (forvar2492 < (1'h0)); forvar2492 = (forvar2492 + (1'h1)))
                    begin
                      reg2493 <= $signed({reg2479[(2'h2):(1'h0)]});
                      reg2494 <= $unsigned($signed((!reg2419[(3'h4):(3'h4)])));
                      reg2495 <= reg2439;
                    end
                  if ({reg2495})
                    begin
                      reg2496 <= (reg2403 ?
                          (8'hac) : (reg2463[(1'h0):(1'h0)] ?
                              reg2459 : ($unsigned(reg2493) * reg2462)));
                    end
                  else
                    begin
                      reg2496 <= $unsigned($unsigned(((-reg2470) ?
                          (forvar2438 <= reg2467) : $signed(forvar2387))));
                      reg2497 <= $unsigned($signed(((forvar2485 ?
                          forvar2415 : (8'ha8)) && (wire2373 & reg2474))));
                    end
                end
              reg2498 <= (|$signed(forvar2472[(3'h7):(3'h6)]));
            end
          reg2499 <= reg2393[(4'ha):(4'h9)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar2500 = (1'h0); (forvar2500 < (2'h3)); forvar2500 = (forvar2500 + (1'h1)))
        begin
          for (forvar2501 = (1'h0); (forvar2501 < (1'h1)); forvar2501 = (forvar2501 + (1'h1)))
            begin
              for (forvar2502 = (1'h0); (forvar2502 < (2'h2)); forvar2502 = (forvar2502 + (1'h1)))
                begin
                  for (forvar2503 = (1'h0); (forvar2503 < (2'h3)); forvar2503 = (forvar2503 + (1'h1)))
                    begin
                      reg2504 <= {(|$signed({(8'hae)}))};
                      reg2505 <= $unsigned($signed((^~reg2495)));
                      reg2506 <= (^{$signed($unsigned((8'ha2)))});
                    end
                end
              reg2507 <= $signed(forvar2457[(3'h6):(2'h3)]);
              if ($unsigned(reg2469[(3'h4):(3'h4)]))
                begin
                  if ($signed(({{(8'ha2)}} ?
                      (forvar2492[(4'hc):(4'ha)] <= (forvar2408 > reg2467)) : $unsigned($signed((8'ha2))))))
                    begin
                      reg2508 <= ({(^~(reg2404 != reg2460))} ?
                          forvar2383 : reg2468[(3'h7):(2'h3)]);
                      reg2509 <= $unsigned(((reg2381[(3'h7):(3'h5)] ?
                              $signed(reg2385) : (reg2481 >= reg2422)) ?
                          (+$signed(forvar2386)) : (((8'hb0) ?
                                  reg2497 : reg2430) ?
                              reg2412 : reg2490)));
                      reg2510 <= (forvar2485[(3'h6):(3'h4)] ?
                          reg2506 : (~^reg2390[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2508 <= reg2441[(3'h4):(2'h3)];
                    end
                  for (forvar2511 = (1'h0); (forvar2511 < (2'h2)); forvar2511 = (forvar2511 + (1'h1)))
                    begin
                      reg2512 <= forvar2511;
                      reg2513 <= (reg2414[(1'h0):(1'h0)] ~^ ((~^(~^reg2387)) == $unsigned((|reg2493))));
                      reg2514 <= (&(reg2419[(2'h2):(1'h1)] ?
                          (reg2432 == reg2495[(3'h5):(2'h2)]) : {reg2450[(3'h4):(2'h3)]}));
                    end
                end
              else
                begin
                  for (forvar2508 = (1'h0); (forvar2508 < (2'h2)); forvar2508 = (forvar2508 + (1'h1)))
                    begin
                      reg2509 <= ((-$unsigned((8'hb9))) ?
                          reg2483 : forvar2438[(3'h4):(1'h1)]);
                      reg2510 <= (^~$signed($unsigned((reg2474 ?
                          (8'hab) : reg2403))));
                      reg2511 <= reg2432[(1'h1):(1'h1)];
                      reg2512 <= $unsigned(reg2474[(2'h3):(2'h2)]);
                    end
                end
              for (forvar2515 = (1'h0); (forvar2515 < (1'h1)); forvar2515 = (forvar2515 + (1'h1)))
                begin
                  if ((reg2451 >>> forvar2450[(1'h1):(1'h1)]))
                    begin
                      reg2516 <= reg2379;
                      reg2517 <= $unsigned(reg2377);
                    end
                  else
                    begin
                      reg2516 <= $signed(wire2374);
                    end
                end
            end
        end
      for (forvar2518 = (1'h0); (forvar2518 < (1'h1)); forvar2518 = (forvar2518 + (1'h1)))
        begin
          if ({(~&{$signed((8'hae))})})
            begin
              for (forvar2519 = (1'h0); (forvar2519 < (1'h0)); forvar2519 = (forvar2519 + (1'h1)))
                begin
                  reg2520 <= $unsigned($unsigned(forvar2433));
                  if ((^$signed(reg2505)))
                    begin
                      reg2521 <= {forvar2511};
                    end
                  else
                    begin
                      reg2521 <= {({(~&forvar2397)} ^ (8'ha3))};
                      reg2522 <= $unsigned((!($signed((8'ha5)) > reg2408)));
                      reg2523 <= {$signed(({reg2411} ?
                              $unsigned(reg2452) : reg2469[(1'h0):(1'h0)]))};
                      reg2524 <= {{reg2403[(3'h5):(3'h5)]}};
                    end
                end
            end
          else
            begin
              reg2519 <= (8'ha9);
              for (forvar2520 = (1'h0); (forvar2520 < (2'h3)); forvar2520 = (forvar2520 + (1'h1)))
                begin
                  if ($signed(($unsigned({reg2453}) ?
                      wire2370[(1'h1):(1'h0)] : $signed(reg2387[(3'h7):(2'h2)]))))
                    begin
                      reg2521 <= reg2460[(3'h5):(3'h5)];
                      reg2522 <= ((!(~&reg2499[(2'h3):(2'h2)])) ?
                          (^~reg2471) : (|({(8'ha0)} != {(8'hb6)})));
                      reg2523 <= $unsigned($unsigned(reg2389[(3'h6):(1'h0)]));
                      reg2524 <= (((|reg2442) != $unsigned(((8'ha4) ?
                              (8'h9d) : reg2426))) ?
                          {forvar2519} : ((reg2424[(4'hc):(1'h0)] || (&reg2436)) || reg2463));
                    end
                  else
                    begin
                      reg2521 <= reg2398[(3'h4):(2'h3)];
                    end
                end
              if ((|reg2523[(3'h4):(1'h1)]))
                begin
                  reg2525 <= $unsigned(reg2383[(1'h1):(1'h0)]);
                  if ({((-forvar2383) ~^ (8'h9d))})
                    begin
                      reg2526 <= (~|$unsigned((((8'h9c) ?
                          wire2374 : reg2387) ^ (reg2424 ?
                          (8'ha6) : reg2399))));
                    end
                  else
                    begin
                      reg2526 <= (reg2430[(1'h1):(1'h0)] ?
                          $signed(($unsigned(forvar2503) != {(8'ha7)})) : ((((8'had) + (8'h9e)) ?
                              (forvar2388 ?
                                  forvar2391 : reg2525) : (~&reg2521)) == ((&forvar2389) ?
                              (reg2441 ? (8'hb1) : reg2412) : (-(8'hb4)))));
                    end
                end
              else
                begin
                  reg2525 <= $signed($unsigned(forvar2382[(1'h1):(1'h1)]));
                end
              if (reg2406)
                begin
                  for (forvar2527 = (1'h0); (forvar2527 < (2'h2)); forvar2527 = (forvar2527 + (1'h1)))
                    begin
                      reg2528 <= (reg2523 + $signed({reg2394[(3'h5):(1'h0)]}));
                    end
                  for (forvar2529 = (1'h0); (forvar2529 < (2'h2)); forvar2529 = (forvar2529 + (1'h1)))
                    begin
                      reg2530 <= {$unsigned(forvar2529)};
                      reg2531 <= ($signed(((forvar2420 >> reg2456) ?
                              (^(8'ha3)) : {forvar2383})) ?
                          $unsigned(reg2442[(4'h9):(3'h4)]) : reg2393[(3'h7):(3'h7)]);
                    end
                  reg2532 <= ((8'ha2) ?
                      {$unsigned($unsigned((8'ha8)))} : reg2526[(3'h5):(2'h2)]);
                end
              else
                begin
                  if ($unsigned(reg2511))
                    begin
                      reg2527 <= (-reg2514);
                      reg2528 <= ($signed(reg2386[(1'h0):(1'h0)]) ?
                          forvar2501[(1'h0):(1'h0)] : $signed(reg2514[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2527 <= (~(^~reg2377[(3'h7):(1'h0)]));
                      reg2528 <= (($signed(reg2525[(1'h0):(1'h0)]) ?
                              ({reg2424} ?
                                  (!forvar2394) : {forvar2434}) : (~(forvar2450 ?
                                  forvar2520 : (8'h9d)))) ?
                          (reg2509[(2'h2):(1'h1)] != reg2462) : forvar2443);
                      reg2529 <= $unsigned($unsigned((|$unsigned(reg2487))));
                    end
                  for (forvar2530 = (1'h0); (forvar2530 < (2'h3)); forvar2530 = (forvar2530 + (1'h1)))
                    begin
                      reg2531 <= (+(&$signed({forvar2485})));
                      reg2532 <= forvar2457;
                      reg2533 <= forvar2385[(4'hc):(4'hc)];
                    end
                  if (reg2422)
                    begin
                      reg2534 <= $signed($unsigned(forvar2501));
                      reg2535 <= (reg2428[(2'h2):(1'h1)] >> $unsigned($unsigned((^~reg2466))));
                      reg2536 <= {(8'hb7)};
                    end
                  else
                    begin
                      reg2534 <= (!$unsigned(wire2374));
                      reg2535 <= (~^(($signed(forvar2518) ^ (reg2396 ?
                              (8'hb1) : (8'haf))) ?
                          forvar2413 : reg2392[(2'h2):(1'h0)]));
                      reg2536 <= $signed(({(forvar2518 ^ reg2449)} ^ (~|forvar2416)));
                    end
                  if ($signed(((!(|reg2449)) ?
                      {(reg2399 >> reg2447)} : $unsigned($unsigned(reg2405)))))
                    begin
                      reg2537 <= reg2469;
                      reg2538 <= $signed($unsigned((reg2469[(3'h6):(2'h3)] ?
                          $signed(reg2477) : (forvar2492 ?
                              reg2458 : forvar2384))));
                    end
                  else
                    begin
                      reg2537 <= (forvar2450[(3'h5):(2'h3)] >>> reg2532[(1'h1):(1'h0)]);
                      reg2538 <= $signed(($unsigned((reg2468 ?
                              (8'hb9) : reg2416)) ?
                          (((8'hb0) != (8'hb5)) ?
                              reg2408 : (reg2436 ?
                                  reg2527 : reg2394)) : reg2378[(4'h9):(1'h0)]));
                      reg2539 <= reg2402[(2'h3):(2'h3)];
                      reg2540 <= forvar2492[(4'hc):(3'h6)];
                    end
                end
            end
        end
      for (forvar2541 = (1'h0); (forvar2541 < (1'h0)); forvar2541 = (forvar2541 + (1'h1)))
        begin
          reg2542 <= {$unsigned(((~(8'ha4)) ? {reg2404} : $signed(reg2439)))};
        end
    end
  assign wire2543 = (&((reg2452[(4'hd):(4'h8)] ?
                        (forvar2452 ^~ reg2527) : (reg2483 == forvar2379)) >= reg2410[(1'h1):(1'h1)]));
  assign wire2544 = $signed(($unsigned($unsigned(forvar2508)) > {wire2543}));
  assign wire2545 = reg2517;
  assign wire2546 = forvar2450;
  always
    @(posedge clk) begin
      reg2547 <= $unsigned({$signed($signed(reg2397))});
      for (forvar2548 = (1'h0); (forvar2548 < (1'h0)); forvar2548 = (forvar2548 + (1'h1)))
        begin
          reg2549 <= {$unsigned(forvar2389)};
        end
      if ($signed(reg2479[(2'h3):(1'h0)]))
        begin
          for (forvar2550 = (1'h0); (forvar2550 < (1'h0)); forvar2550 = (forvar2550 + (1'h1)))
            begin
              if ($signed($unsigned($signed(reg2542[(2'h3):(2'h2)]))))
                begin
                  for (forvar2551 = (1'h0); (forvar2551 < (2'h3)); forvar2551 = (forvar2551 + (1'h1)))
                    begin
                      reg2552 <= $unsigned(((reg2510 ?
                              (forvar2527 & reg2427) : {reg2445}) ?
                          ((8'h9e) ?
                              reg2433[(2'h2):(1'h0)] : (^(8'hb3))) : ((reg2514 ?
                              reg2480 : reg2542) + (reg2439 <<< forvar2508))));
                      reg2553 <= reg2397;
                    end
                  for (forvar2554 = (1'h0); (forvar2554 < (2'h3)); forvar2554 = (forvar2554 + (1'h1)))
                    begin
                      reg2555 <= ((8'hb0) + reg2412);
                    end
                  if (($unsigned(reg2434) != $signed($unsigned($signed(forvar2500)))))
                    begin
                      reg2556 <= reg2487;
                      reg2557 <= $unsigned(reg2505[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg2556 <= reg2455;
                    end
                end
              else
                begin
                  for (forvar2551 = (1'h0); (forvar2551 < (1'h1)); forvar2551 = (forvar2551 + (1'h1)))
                    begin
                      reg2552 <= forvar2434[(1'h0):(1'h0)];
                    end
                  if ($unsigned($unsigned({$signed(forvar2511)})))
                    begin
                      reg2553 <= forvar2377;
                      reg2554 <= reg2496;
                      reg2555 <= ((reg2381[(3'h5):(2'h3)] ~^ reg2419[(1'h0):(1'h0)]) ?
                          reg2380 : {{$signed(reg2397)}});
                    end
                  else
                    begin
                      reg2553 <= ((reg2426 ?
                              reg2538[(4'hd):(4'hc)] : ($signed(forvar2386) ?
                                  (reg2382 && wire2369) : $unsigned((8'haa)))) ?
                          $signed({(8'hb8)}) : reg2549[(1'h1):(1'h1)]);
                      reg2554 <= reg2390[(2'h2):(1'h0)];
                    end
                  if (reg2534[(3'h4):(1'h0)])
                    begin
                      reg2556 <= $unsigned((((|forvar2383) | $signed(reg2412)) ?
                          (reg2509 == {reg2462}) : $unsigned($signed(reg2407))));
                      reg2557 <= $unsigned($unsigned(reg2479[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg2556 <= forvar2527;
                      reg2557 <= forvar2472[(3'h6):(1'h1)];
                    end
                  for (forvar2558 = (1'h0); (forvar2558 < (1'h1)); forvar2558 = (forvar2558 + (1'h1)))
                    begin
                      reg2559 <= wire2375;
                    end
                end
              for (forvar2560 = (1'h0); (forvar2560 < (2'h3)); forvar2560 = (forvar2560 + (1'h1)))
                begin
                  if ((8'h9f))
                    begin
                      reg2561 <= {(-$signed({reg2519}))};
                    end
                  else
                    begin
                      reg2561 <= reg2525[(2'h3):(1'h0)];
                    end
                  if (reg2424)
                    begin
                      reg2562 <= reg2414;
                      reg2563 <= $unsigned($signed((reg2405[(1'h0):(1'h0)] != reg2435[(3'h6):(1'h0)])));
                      reg2564 <= reg2494;
                    end
                  else
                    begin
                      reg2562 <= reg2506[(1'h1):(1'h0)];
                      reg2563 <= $unsigned((^~reg2456));
                    end
                  for (forvar2565 = (1'h0); (forvar2565 < (1'h1)); forvar2565 = (forvar2565 + (1'h1)))
                    begin
                      reg2566 <= $signed($unsigned(reg2506[(2'h2):(1'h1)]));
                      reg2567 <= $signed(reg2488);
                      reg2568 <= ($unsigned({$signed(reg2552)}) ?
                          {$unsigned($unsigned(forvar2434))} : reg2397[(1'h0):(1'h0)]);
                      reg2569 <= (^$unsigned(forvar2560));
                    end
                  reg2570 <= ((^(reg2414[(2'h2):(1'h1)] || reg2505)) >>> ((reg2526[(1'h1):(1'h1)] & $unsigned(reg2481)) || ({(8'ha9)} ?
                      $unsigned(wire2374) : (~(8'hb0)))));
                end
              for (forvar2571 = (1'h0); (forvar2571 < (1'h0)); forvar2571 = (forvar2571 + (1'h1)))
                begin
                  if (((~$signed((reg2509 || forvar2501))) ?
                      $unsigned(reg2481[(3'h4):(2'h2)]) : (&(-reg2379[(1'h0):(1'h0)]))))
                    begin
                      reg2572 <= ($signed($signed((reg2489 < reg2437))) * (+reg2470[(2'h2):(1'h0)]));
                      reg2573 <= reg2563;
                    end
                  else
                    begin
                      reg2572 <= ((({forvar2445} ?
                              reg2407 : forvar2550[(3'h6):(3'h4)]) ^ $unsigned(reg2508[(4'hb):(3'h6)])) ?
                          reg2563[(1'h0):(1'h0)] : reg2411[(4'he):(1'h0)]);
                    end
                end
            end
          for (forvar2574 = (1'h0); (forvar2574 < (2'h3)); forvar2574 = (forvar2574 + (1'h1)))
            begin
              for (forvar2575 = (1'h0); (forvar2575 < (1'h1)); forvar2575 = (forvar2575 + (1'h1)))
                begin
                  reg2576 <= (~reg2386);
                  if (((8'ha9) ^~ $unsigned($signed((~^forvar2420)))))
                    begin
                      reg2577 <= ($unsigned(reg2470[(1'h1):(1'h0)]) ?
                          $signed(((reg2380 ?
                              reg2400 : reg2562) * forvar2386[(4'hd):(4'hd)])) : forvar2422);
                      reg2578 <= $unsigned(reg2495[(3'h7):(3'h4)]);
                    end
                  else
                    begin
                      reg2577 <= ($unsigned(((~reg2459) | forvar2500[(3'h4):(2'h2)])) ?
                          (8'ha0) : {reg2396});
                      reg2578 <= (~|($signed((reg2447 ?
                          reg2547 : wire2546)) ^ forvar2438[(4'h9):(4'h9)]));
                    end
                end
            end
          if (reg2497[(3'h7):(2'h2)])
            begin
              if (reg2529[(3'h7):(1'h0)])
                begin
                  if ((|(reg2540 ~^ $signed((reg2525 <= forvar2554)))))
                    begin
                      reg2579 <= (8'h9c);
                      reg2580 <= ((^(reg2381[(3'h4):(1'h1)] ^ ((8'hb1) & reg2520))) ?
                          forvar2433 : ((&$signed(forvar2515)) != reg2382[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg2579 <= ($unsigned(reg2554[(3'h7):(3'h5)]) ?
                          reg2567 : (+(^~reg2520)));
                      reg2580 <= ($signed($signed(reg2495)) ?
                          {(~|(+reg2400))} : forvar2448[(1'h0):(1'h0)]);
                      reg2581 <= {reg2453[(1'h1):(1'h0)]};
                    end
                  reg2582 <= forvar2565;
                  if ((+reg2425))
                    begin
                      reg2583 <= $signed((~$signed($signed(reg2384))));
                      reg2584 <= forvar2473[(2'h3):(2'h2)];
                      reg2585 <= reg2540;
                    end
                  else
                    begin
                      reg2583 <= ($signed((8'hb2)) ?
                          $unsigned((forvar2550 ^~ forvar2389)) : $unsigned($unsigned((forvar2450 > reg2553))));
                    end
                  if ($signed(wire2372))
                    begin
                      reg2586 <= ($signed(forvar2415[(4'h8):(3'h4)]) * (8'ha9));
                      reg2587 <= $unsigned(reg2554[(4'hc):(4'hc)]);
                      reg2588 <= (((8'hae) ?
                              $signed((forvar2575 ^~ forvar2388)) : (reg2404 >>> $signed(wire2372))) ?
                          $signed(((&(8'hb2)) - (wire2543 == (8'hb5)))) : {$unsigned((-forvar2501))});
                      reg2589 <= forvar2445[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg2586 <= ((!(~$unsigned(forvar2519))) ?
                          forvar2391 : ({$signed(reg2429)} ?
                              (!(forvar2428 ?
                                  reg2463 : (8'hb4))) : $signed((~&(8'haa)))));
                      reg2587 <= reg2579[(2'h3):(2'h2)];
                      reg2588 <= ($unsigned((reg2585 ?
                          forvar2398 : $unsigned((8'had)))) != (-((reg2388 | (8'ha4)) ?
                          $signed(reg2537) : {reg2393})));
                      reg2589 <= ((reg2395 << (reg2525 ?
                              ((8'hab) ?
                                  wire2546 : reg2495) : reg2449[(4'hb):(3'h5)])) ?
                          (reg2417[(2'h2):(2'h2)] ?
                              $unsigned((forvar2575 - (8'ha2))) : $signed(forvar2558[(2'h3):(2'h3)])) : wire2372);
                    end
                end
              else
                begin
                  reg2579 <= reg2580;
                  if (reg2426[(3'h5):(2'h2)])
                    begin
                      reg2580 <= $unsigned(($signed(reg2433) ?
                          reg2456 : (&{reg2383})));
                      reg2581 <= {(reg2408 && ($unsigned(reg2536) ?
                              (forvar2508 <<< reg2400) : (reg2584 ?
                                  reg2422 : reg2542)))};
                      reg2582 <= (~reg2416[(1'h0):(1'h0)]);
                      reg2583 <= (|forvar2389[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg2580 <= (~^reg2509);
                      reg2581 <= (((^$unsigned(reg2384)) ?
                          reg2495[(3'h6):(3'h6)] : reg2399[(1'h1):(1'h0)]) * $signed(((|forvar2433) ?
                          ((8'hb7) ? reg2437 : forvar2560) : (8'ha9))));
                      reg2582 <= reg2377;
                      reg2583 <= (~^reg2379);
                    end
                  reg2584 <= (~^(8'ha1));
                end
            end
          else
            begin
              for (forvar2579 = (1'h0); (forvar2579 < (1'h0)); forvar2579 = (forvar2579 + (1'h1)))
                begin
                  if ((^~$signed(reg2432[(1'h0):(1'h0)])))
                    begin
                      reg2580 <= reg2475;
                      reg2581 <= $unsigned($signed($unsigned($signed(reg2449))));
                      reg2582 <= $unsigned((reg2529[(3'h4):(1'h0)] ?
                          (forvar2445 ?
                              ((8'h9f) ^ reg2406) : ((8'hba) + reg2409)) : reg2377[(1'h1):(1'h0)]));
                      reg2583 <= {$signed((((8'ha2) ? reg2580 : forvar2443) ?
                              (reg2559 ? reg2466 : forvar2486) : reg2488))};
                    end
                  else
                    begin
                      reg2580 <= ($unsigned((((8'haf) ?
                          forvar2416 : reg2430) >>> $signed(reg2582))) >>> ($signed((!reg2383)) + (~^$unsigned(reg2528))));
                      reg2581 <= reg2408[(4'hb):(4'h9)];
                      reg2582 <= ((~^reg2380) ?
                          $unsigned(reg2494[(3'h5):(3'h5)]) : (~^((reg2581 ^ (8'h9e)) ?
                              reg2476[(3'h4):(2'h3)] : $unsigned(reg2549))));
                      reg2583 <= (~^reg2586[(4'hc):(2'h3)]);
                    end
                  if ((((~^(reg2542 ? reg2483 : reg2407)) ?
                          $unsigned($unsigned(forvar2457)) : forvar2420[(1'h0):(1'h0)]) ?
                      reg2556[(2'h2):(1'h0)] : (!wire2543)))
                    begin
                      reg2584 <= (($signed($signed(reg2564)) ?
                          ((reg2521 ? (8'ha5) : forvar2541) ?
                              reg2378 : (reg2579 ?
                                  (8'hb1) : (8'ha4))) : reg2578) ~^ {{$signed((8'hb0))}});
                      reg2585 <= (&reg2509);
                    end
                  else
                    begin
                      reg2584 <= forvar2415[(4'hd):(3'h5)];
                      reg2585 <= (|$unsigned($unsigned((&reg2563))));
                    end
                  for (forvar2586 = (1'h0); (forvar2586 < (2'h3)); forvar2586 = (forvar2586 + (1'h1)))
                    begin
                      reg2587 <= ((|{$unsigned((8'hb2))}) ?
                          (wire2373 ?
                              (8'ha4) : reg2534) : (forvar2377 + reg2391));
                      reg2588 <= $signed({(|$signed(reg2404))});
                      reg2589 <= $signed($unsigned(((forvar2383 > (8'hba)) ^~ $signed(reg2416))));
                      reg2590 <= {{reg2586}};
                    end
                  for (forvar2591 = (1'h0); (forvar2591 < (2'h2)); forvar2591 = (forvar2591 + (1'h1)))
                    begin
                      reg2592 <= $signed($unsigned((^(reg2566 * forvar2422))));
                      reg2593 <= (8'hb2);
                      reg2594 <= ($unsigned(((reg2511 ?
                              reg2559 : reg2442) < $signed(reg2527))) ?
                          {reg2464} : (($signed(reg2524) ?
                                  {forvar2565} : (wire2543 >= reg2446)) ?
                              ($signed(reg2593) ?
                                  (forvar2397 < reg2426) : $unsigned(reg2423)) : (&$unsigned((8'ha1)))));
                      reg2595 <= (!$unsigned(((reg2516 & reg2517) ?
                          (8'hb0) : (reg2522 <<< reg2578))));
                    end
                end
              for (forvar2596 = (1'h0); (forvar2596 < (2'h2)); forvar2596 = (forvar2596 + (1'h1)))
                begin
                  if (reg2478[(1'h0):(1'h0)])
                    begin
                      reg2597 <= reg2505;
                      reg2598 <= $signed({(reg2389[(2'h2):(1'h1)] ~^ $signed(reg2470))});
                    end
                  else
                    begin
                      reg2597 <= ((^reg2408[(4'hb):(3'h6)]) >= (((8'ha7) << (forvar2511 >> reg2507)) ?
                          {reg2561} : $unsigned($unsigned((8'hac)))));
                      reg2598 <= reg2398;
                    end
                  for (forvar2599 = (1'h0); (forvar2599 < (2'h2)); forvar2599 = (forvar2599 + (1'h1)))
                    begin
                      reg2600 <= $signed((({forvar2397} ?
                              $unsigned(forvar2511) : (reg2493 ?
                                  (8'hae) : (8'haa))) ?
                          (~&{(8'hb2)}) : $unsigned((wire2371 ?
                              reg2491 : (8'hb4)))));
                      reg2601 <= $signed($unsigned(reg2564[(2'h3):(2'h3)]));
                      reg2602 <= ($unsigned($unsigned(reg2600[(4'h9):(2'h2)])) <= $signed(forvar2423));
                      reg2603 <= $signed(((!$signed(reg2434)) >> $unsigned((reg2563 > reg2408))));
                    end
                  if ($signed($unsigned(((reg2409 >= reg2533) || reg2471[(4'h8):(1'h1)]))))
                    begin
                      reg2604 <= (^reg2526[(1'h1):(1'h0)]);
                      reg2605 <= {(^~((-reg2405) >>> (reg2434 ?
                              reg2424 : forvar2438)))};
                    end
                  else
                    begin
                      reg2604 <= {reg2470};
                      reg2605 <= forvar2541[(4'h9):(3'h7)];
                    end
                end
              reg2606 <= forvar2434[(2'h2):(1'h0)];
              reg2607 <= reg2454;
            end
        end
      else
        begin
          reg2550 <= ($unsigned($unsigned(reg2423[(4'h8):(3'h5)])) ?
              {reg2521} : $unsigned({$unsigned(forvar2501)}));
        end
    end
  always
    @(posedge clk) begin
      if (forvar2501[(2'h2):(1'h1)])
        begin
          for (forvar2608 = (1'h0); (forvar2608 < (1'h0)); forvar2608 = (forvar2608 + (1'h1)))
            begin
              for (forvar2609 = (1'h0); (forvar2609 < (1'h0)); forvar2609 = (forvar2609 + (1'h1)))
                begin
                  for (forvar2610 = (1'h0); (forvar2610 < (2'h3)); forvar2610 = (forvar2610 + (1'h1)))
                    begin
                      reg2611 <= $unsigned($unsigned((forvar2378[(1'h1):(1'h1)] ?
                          $signed((8'haa)) : $unsigned(reg2420))));
                      reg2612 <= (-$signed(({reg2514} ? {reg2605} : reg2455)));
                      reg2613 <= reg2612[(4'hf):(4'hc)];
                    end
                  reg2614 <= {reg2387};
                  for (forvar2615 = (1'h0); (forvar2615 < (1'h1)); forvar2615 = (forvar2615 + (1'h1)))
                    begin
                      reg2616 <= $signed($signed(((reg2428 ?
                              reg2553 : (8'ha3)) ?
                          {reg2586} : reg2414[(2'h2):(1'h0)])));
                      reg2617 <= (forvar2438[(3'h7):(1'h0)] ?
                          reg2395[(1'h0):(1'h0)] : (+((~|(8'hb3)) ?
                              forvar2541[(1'h0):(1'h0)] : ((8'hb0) && (8'hb6)))));
                      reg2618 <= (^(8'hb4));
                      reg2619 <= {(reg2450 > (-wire2545[(2'h2):(1'h1)]))};
                    end
                  for (forvar2620 = (1'h0); (forvar2620 < (1'h1)); forvar2620 = (forvar2620 + (1'h1)))
                    begin
                      reg2621 <= $signed({reg2440[(3'h4):(1'h0)]});
                      reg2622 <= $signed($signed((8'hba)));
                      reg2623 <= reg2397[(1'h1):(1'h0)];
                    end
                end
            end
        end
      else
        begin
          if (({($unsigned(reg2514) ^ $signed(reg2550))} ?
              reg2556[(3'h5):(3'h5)] : reg2417))
            begin
              if ((($unsigned((^~reg2525)) ?
                      ({reg2388} == reg2498[(3'h4):(2'h3)]) : $unsigned((|reg2450))) ?
                  $signed($signed(reg2402[(2'h2):(2'h2)])) : ($unsigned((forvar2449 > forvar2520)) || (~(~|(8'hb9))))))
                begin
                  for (forvar2608 = (1'h0); (forvar2608 < (2'h3)); forvar2608 = (forvar2608 + (1'h1)))
                    begin
                      reg2609 <= forvar2378[(3'h5):(2'h2)];
                    end
                  reg2610 <= (~|reg2526);
                  for (forvar2611 = (1'h0); (forvar2611 < (2'h2)); forvar2611 = (forvar2611 + (1'h1)))
                    begin
                      reg2612 <= $signed((8'hac));
                      reg2613 <= (reg2393 ?
                          reg2477[(2'h3):(1'h1)] : $signed(forvar2391[(3'h4):(3'h4)]));
                    end
                end
              else
                begin
                  for (forvar2608 = (1'h0); (forvar2608 < (1'h1)); forvar2608 = (forvar2608 + (1'h1)))
                    begin
                      reg2609 <= reg2554;
                      reg2610 <= reg2419;
                      reg2611 <= $signed({((8'ha4) ^ (8'ha5))});
                      reg2612 <= $unsigned({((!forvar2620) ?
                              (reg2469 ? reg2483 : (8'ha9)) : {reg2436})});
                    end
                  for (forvar2613 = (1'h0); (forvar2613 < (1'h1)); forvar2613 = (forvar2613 + (1'h1)))
                    begin
                      reg2614 <= (forvar2397[(4'hb):(3'h4)] ?
                          reg2440 : forvar2377[(2'h3):(2'h2)]);
                      reg2615 <= reg2401;
                      reg2616 <= reg2445[(4'ha):(2'h2)];
                      reg2617 <= (~(~^reg2456));
                    end
                end
            end
          else
            begin
              for (forvar2608 = (1'h0); (forvar2608 < (2'h2)); forvar2608 = (forvar2608 + (1'h1)))
                begin
                  if (($unsigned(reg2459[(3'h6):(2'h3)]) * wire2543[(3'h5):(3'h5)]))
                    begin
                      reg2609 <= ({$unsigned(reg2553[(4'ha):(3'h4)])} ?
                          $unsigned({$signed(reg2562)}) : reg2487);
                      reg2610 <= (^(($signed((8'ha2)) ?
                              $unsigned(reg2461) : (forvar2398 ?
                                  forvar2446 : forvar2384)) ?
                          $unsigned((reg2623 * wire2376)) : wire2370));
                      reg2611 <= forvar2511[(4'ha):(1'h0)];
                    end
                  else
                    begin
                      reg2609 <= $signed(reg2597);
                      reg2610 <= reg2388[(3'h6):(1'h0)];
                      reg2611 <= $signed($signed(forvar2591));
                      reg2612 <= reg2425;
                    end
                end
              for (forvar2613 = (1'h0); (forvar2613 < (2'h2)); forvar2613 = (forvar2613 + (1'h1)))
                begin
                  if ($signed(reg2594))
                    begin
                      reg2614 <= (~|$unsigned({$unsigned(forvar2398)}));
                    end
                  else
                    begin
                      reg2614 <= {(reg2378[(1'h1):(1'h0)] ?
                              (~reg2440[(4'hb):(3'h7)]) : $unsigned(((8'hac) ?
                                  reg2550 : reg2401)))};
                      reg2615 <= $unsigned(($signed(reg2387[(3'h7):(3'h6)]) ?
                          (|((8'hb8) ? reg2419 : forvar2486)) : {reg2456}));
                      reg2616 <= $signed((forvar2473[(1'h0):(1'h0)] | $signed(reg2381[(3'h5):(1'h1)])));
                    end
                  if ($signed(reg2381))
                    begin
                      reg2617 <= ((forvar2416 >> (forvar2407[(1'h1):(1'h0)] ?
                              reg2623 : reg2383[(2'h2):(2'h2)])) ?
                          (reg2463 && reg2533) : reg2382[(2'h2):(1'h0)]);
                      reg2618 <= $unsigned((&$unsigned($signed(reg2617))));
                      reg2619 <= $unsigned((8'haf));
                      reg2620 <= reg2613;
                    end
                  else
                    begin
                      reg2617 <= $unsigned(reg2533[(3'h4):(1'h0)]);
                      reg2618 <= forvar2586;
                    end
                  reg2621 <= reg2614;
                  if (($unsigned((~&(reg2580 ? forvar2530 : (8'h9d)))) ?
                      (reg2477[(1'h1):(1'h1)] ?
                          (^~forvar2379[(3'h4):(1'h1)]) : forvar2472[(2'h3):(2'h3)]) : (!($signed(reg2411) ?
                          $unsigned(forvar2377) : ((8'ha4) * (8'hb4))))))
                    begin
                      reg2622 <= (($signed($signed(reg2420)) * ((forvar2611 <= reg2517) ?
                          (reg2526 ?
                              forvar2452 : reg2604) : {reg2484})) | reg2433);
                      reg2623 <= {(+$unsigned({reg2384}))};
                    end
                  else
                    begin
                      reg2622 <= reg2510;
                      reg2623 <= ($signed(reg2389) ^~ ({(reg2405 ?
                                  forvar2378 : reg2467)} ?
                          $unsigned($unsigned((8'ha4))) : reg2484));
                      reg2624 <= reg2559[(1'h0):(1'h0)];
                    end
                end
              for (forvar2625 = (1'h0); (forvar2625 < (2'h2)); forvar2625 = (forvar2625 + (1'h1)))
                begin
                  for (forvar2626 = (1'h0); (forvar2626 < (1'h0)); forvar2626 = (forvar2626 + (1'h1)))
                    begin
                      reg2627 <= wire2545;
                      reg2628 <= forvar2515[(3'h5):(3'h5)];
                      reg2629 <= ((8'hab) | $unsigned({$signed((8'ha0))}));
                      reg2630 <= (8'hb3);
                    end
                  for (forvar2631 = (1'h0); (forvar2631 < (1'h0)); forvar2631 = (forvar2631 + (1'h1)))
                    begin
                      reg2632 <= ((+$unsigned((forvar2386 ?
                              (8'ha2) : reg2542))) ?
                          (reg2462[(3'h4):(1'h1)] ?
                              reg2535[(3'h7):(2'h3)] : reg2614) : (reg2620[(3'h4):(3'h4)] ?
                              $signed(((8'ha7) + reg2532)) : reg2564[(2'h3):(1'h0)]));
                      reg2633 <= reg2552;
                    end
                  if ((~reg2407[(3'h5):(3'h5)]))
                    begin
                      reg2634 <= (^~forvar2511[(3'h7):(1'h0)]);
                    end
                  else
                    begin
                      reg2634 <= (~^$unsigned(((forvar2382 ?
                              (8'haa) : reg2427) ?
                          (reg2447 ?
                              reg2522 : reg2407) : $signed(forvar2579))));
                      reg2635 <= (forvar2550 << reg2398);
                      reg2636 <= reg2568;
                      reg2637 <= $signed(reg2627);
                    end
                  for (forvar2638 = (1'h0); (forvar2638 < (1'h1)); forvar2638 = (forvar2638 + (1'h1)))
                    begin
                      reg2639 <= forvar2379[(3'h5):(2'h2)];
                      reg2640 <= {$signed(wire2372[(3'h7):(3'h7)])};
                    end
                end
            end
          for (forvar2641 = (1'h0); (forvar2641 < (2'h3)); forvar2641 = (forvar2641 + (1'h1)))
            begin
              for (forvar2642 = (1'h0); (forvar2642 < (2'h2)); forvar2642 = (forvar2642 + (1'h1)))
                begin
                  for (forvar2643 = (1'h0); (forvar2643 < (2'h2)); forvar2643 = (forvar2643 + (1'h1)))
                    begin
                      reg2644 <= ((reg2404[(4'h8):(2'h2)] ?
                              $unsigned((8'ha0)) : (^(forvar2465 <<< reg2623))) ?
                          wire2546[(3'h4):(1'h1)] : {((~|forvar2642) | wire2368)});
                    end
                  if ((~reg2617[(3'h7):(3'h7)]))
                    begin
                      reg2645 <= reg2428;
                      reg2646 <= reg2506;
                      reg2647 <= ((~reg2564[(2'h3):(1'h0)]) ^ (8'hae));
                    end
                  else
                    begin
                      reg2645 <= ((!$unsigned((!reg2490))) != (+($signed(wire2545) ?
                          forvar2611[(2'h2):(2'h2)] : $signed(forvar2641))));
                    end
                end
              for (forvar2648 = (1'h0); (forvar2648 < (1'h0)); forvar2648 = (forvar2648 + (1'h1)))
                begin
                  for (forvar2649 = (1'h0); (forvar2649 < (2'h2)); forvar2649 = (forvar2649 + (1'h1)))
                    begin
                      reg2650 <= ((+$unsigned((reg2611 == forvar2502))) >> (forvar2434 || $unsigned(wire2546)));
                      reg2651 <= ($signed(reg2411) ?
                          $signed(((reg2566 ? (8'h9d) : reg2436) ?
                              wire2543[(3'h7):(3'h5)] : {(8'hb9)})) : forvar2642[(4'hb):(3'h4)]);
                      reg2652 <= $unsigned($unsigned((reg2624 ?
                          forvar2586 : (~|reg2509))));
                      reg2653 <= ({reg2424} ?
                          $signed(reg2390) : (($unsigned(reg2632) ?
                              reg2605[(2'h2):(1'h1)] : {reg2590}) == reg2432[(1'h1):(1'h1)]));
                    end
                  reg2654 <= $unsigned((($unsigned(reg2650) >= $unsigned(reg2611)) ?
                      $signed($signed(forvar2500)) : forvar2379[(3'h4):(1'h0)]));
                end
              for (forvar2655 = (1'h0); (forvar2655 < (2'h3)); forvar2655 = (forvar2655 + (1'h1)))
                begin
                  for (forvar2656 = (1'h0); (forvar2656 < (1'h1)); forvar2656 = (forvar2656 + (1'h1)))
                    begin
                      reg2657 <= reg2397[(3'h7):(1'h0)];
                      reg2658 <= {$signed($unsigned((reg2414 ?
                              reg2445 : forvar2434)))};
                      reg2659 <= forvar2413;
                      reg2660 <= $unsigned((($unsigned(reg2637) ?
                              reg2526 : (~&reg2483)) ?
                          $signed($unsigned((8'ha6))) : $unsigned(reg2654[(1'h1):(1'h0)])));
                    end
                  reg2661 <= (reg2469 << forvar2502[(1'h0):(1'h0)]);
                end
            end
          if ($unsigned(reg2444))
            begin
              for (forvar2662 = (1'h0); (forvar2662 < (2'h3)); forvar2662 = (forvar2662 + (1'h1)))
                begin
                  reg2663 <= wire2376;
                  for (forvar2664 = (1'h0); (forvar2664 < (2'h2)); forvar2664 = (forvar2664 + (1'h1)))
                    begin
                      reg2665 <= reg2531;
                      reg2666 <= ($unsigned(($signed((8'ha2)) ?
                          $signed(reg2585) : $unsigned((8'ha5)))) && ((reg2470[(1'h0):(1'h0)] ?
                          (forvar2662 <<< reg2632) : $signed(reg2553)) == (!reg2451[(4'h8):(3'h7)])));
                      reg2667 <= $signed((~&$unsigned(reg2528[(3'h4):(2'h3)])));
                    end
                  if ($signed((($unsigned(reg2579) || {reg2554}) && (8'hb6))))
                    begin
                      reg2668 <= {$unsigned($unsigned(reg2380[(3'h5):(3'h5)]))};
                    end
                  else
                    begin
                      reg2668 <= (-reg2629);
                      reg2669 <= (($signed($unsigned(reg2517)) >> reg2557) ?
                          ((~&$unsigned(reg2615)) ?
                              $unsigned((reg2517 ?
                                  reg2445 : reg2632)) : $signed(reg2421)) : reg2542);
                    end
                end
            end
          else
            begin
              if ((8'had))
                begin
                  reg2662 <= $signed($signed(forvar2560[(3'h4):(1'h0)]));
                  for (forvar2663 = (1'h0); (forvar2663 < (1'h1)); forvar2663 = (forvar2663 + (1'h1)))
                    begin
                      reg2664 <= $signed((8'ha0));
                      reg2665 <= (8'hb2);
                      reg2666 <= $unsigned($signed(((reg2667 == reg2610) == (forvar2551 ?
                          forvar2502 : reg2401))));
                    end
                  reg2667 <= (8'hb2);
                  for (forvar2668 = (1'h0); (forvar2668 < (1'h1)); forvar2668 = (forvar2668 + (1'h1)))
                    begin
                      reg2669 <= $unsigned($unsigned((^~(reg2663 ~^ (8'hab)))));
                      reg2670 <= (~|(($unsigned((8'hb3)) ?
                              forvar2384 : $signed((8'ha3))) ?
                          {(forvar2383 ?
                                  (8'h9e) : (8'had))} : $unsigned($unsigned(forvar2449))));
                      reg2671 <= (8'ha5);
                    end
                end
              else
                begin
                  for (forvar2662 = (1'h0); (forvar2662 < (2'h3)); forvar2662 = (forvar2662 + (1'h1)))
                    begin
                      reg2663 <= $unsigned((((8'haf) ^ $unsigned((8'hb0))) ?
                          forvar2388[(2'h2):(2'h2)] : {(|reg2477)}));
                      reg2664 <= reg2505;
                      reg2665 <= (~$signed(($unsigned((8'haa)) << $unsigned(reg2487))));
                    end
                  if ({reg2437})
                    begin
                      reg2666 <= (reg2667 ^ reg2448[(3'h5):(2'h3)]);
                    end
                  else
                    begin
                      reg2666 <= $signed(((-(reg2435 >>> reg2380)) + (8'haf)));
                      reg2667 <= forvar2643[(3'h7):(2'h3)];
                      reg2668 <= $unsigned($unsigned(((reg2392 ?
                              (8'hac) : reg2477) ?
                          $signed(reg2657) : (+forvar2515))));
                      reg2669 <= $unsigned(reg2391[(3'h6):(2'h3)]);
                    end
                  for (forvar2670 = (1'h0); (forvar2670 < (1'h0)); forvar2670 = (forvar2670 + (1'h1)))
                    begin
                      reg2671 <= (forvar2541 ^~ ($signed(reg2523[(4'h9):(2'h2)]) ?
                          forvar2613 : (8'ha0)));
                    end
                  if (forvar2620)
                    begin
                      reg2672 <= forvar2649;
                    end
                  else
                    begin
                      reg2672 <= $unsigned($unsigned(reg2385[(1'h1):(1'h1)]));
                      reg2673 <= forvar2448[(2'h3):(2'h2)];
                    end
                end
              for (forvar2674 = (1'h0); (forvar2674 < (1'h0)); forvar2674 = (forvar2674 + (1'h1)))
                begin
                  for (forvar2675 = (1'h0); (forvar2675 < (2'h2)); forvar2675 = (forvar2675 + (1'h1)))
                    begin
                      reg2676 <= $signed(reg2409);
                    end
                end
              if ((~|$signed(((&reg2421) << (^~reg2640)))))
                begin
                  for (forvar2677 = (1'h0); (forvar2677 < (2'h2)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= ($unsigned($unsigned($unsigned(reg2657))) ?
                          {($signed(reg2612) ?
                                  reg2605[(1'h0):(1'h0)] : (wire2368 ?
                                      reg2564 : forvar2558))} : reg2394[(3'h6):(3'h5)]);
                      reg2679 <= ($signed({$signed(reg2388)}) <<< reg2484);
                      reg2680 <= forvar2615[(3'h7):(2'h3)];
                      reg2681 <= (($signed(reg2440) <= (reg2397 * $signed(reg2530))) ?
                          {forvar2398[(4'h8):(1'h0)]} : forvar2452);
                    end
                end
              else
                begin
                  for (forvar2677 = (1'h0); (forvar2677 < (2'h2)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= ({{(&reg2396)}} * (((reg2406 & reg2428) ?
                              reg2583[(2'h3):(1'h0)] : wire2545) ?
                          (-(&reg2586)) : $signed({forvar2530})));
                      reg2679 <= $signed((!$unsigned($unsigned(reg2408))));
                      reg2680 <= reg2673;
                    end
                  for (forvar2681 = (1'h0); (forvar2681 < (1'h1)); forvar2681 = (forvar2681 + (1'h1)))
                    begin
                      reg2682 <= {(^reg2615[(2'h2):(1'h1)])};
                      reg2683 <= (reg2598[(4'h9):(4'h8)] <<< (($unsigned((8'hab)) <<< reg2441) + {$signed(reg2602)}));
                      reg2684 <= (~^(8'hab));
                      reg2685 <= reg2439;
                    end
                  reg2686 <= ($signed(forvar2518[(2'h2):(1'h0)]) > reg2437[(3'h5):(1'h1)]);
                  if (($unsigned((|$unsigned(reg2624))) + (-reg2671[(3'h4):(2'h2)])))
                    begin
                      reg2687 <= $signed($unsigned($unsigned($signed(reg2603))));
                    end
                  else
                    begin
                      reg2687 <= $signed($signed((~&$signed(reg2568))));
                      reg2688 <= (~^($signed((reg2429 | (8'hb7))) ?
                          ($unsigned(reg2624) ?
                              (reg2597 + forvar2508) : $unsigned(reg2522)) : ((reg2600 <<< wire2372) ?
                              {reg2380} : (forvar2675 ?
                                  forvar2448 : reg2585))));
                      reg2689 <= {$signed($signed((reg2463 * (8'ha0))))};
                    end
                end
              for (forvar2690 = (1'h0); (forvar2690 < (1'h1)); forvar2690 = (forvar2690 + (1'h1)))
                begin
                  for (forvar2691 = (1'h0); (forvar2691 < (2'h3)); forvar2691 = (forvar2691 + (1'h1)))
                    begin
                      reg2692 <= (($signed((wire2543 ?
                          reg2526 : (8'ha4))) | $unsigned(reg2496[(2'h2):(1'h1)])) > ((~^forvar2518) ?
                          $unsigned((reg2387 < reg2507)) : {reg2532[(3'h5):(3'h5)]}));
                      reg2693 <= $unsigned((($signed(reg2449) ?
                          (forvar2579 * reg2535) : (reg2542 ?
                              (8'hb0) : reg2605)) <<< $unsigned((^(8'h9c)))));
                      reg2694 <= (forvar2418 ~^ ($signed($signed(reg2516)) <= $signed(((8'hb8) ?
                          reg2555 : (8'ha2)))));
                      reg2695 <= reg2667;
                    end
                  for (forvar2696 = (1'h0); (forvar2696 < (2'h2)); forvar2696 = (forvar2696 + (1'h1)))
                    begin
                      reg2697 <= ($signed($unsigned((reg2587 ?
                          reg2669 : (8'ha2)))) > (&(~&(forvar2663 * reg2416))));
                      reg2698 <= $signed(((reg2459[(3'h7):(2'h3)] | reg2426) ?
                          (~&{wire2370}) : reg2685));
                      reg2699 <= (-$unsigned(({forvar2382} ?
                          (~reg2614) : $signed(reg2634))));
                      reg2700 <= (reg2519 && ({$signed(wire2376)} < {(reg2556 ?
                              reg2550 : reg2395)}));
                    end
                end
            end
        end
      if (forvar2407[(1'h0):(1'h0)])
        begin
          if (((8'hb0) ?
              $signed(reg2448) : ($signed(reg2427) ?
                  ($signed(reg2669) ?
                      $unsigned(forvar2389) : forvar2656) : $unsigned(reg2659))))
            begin
              if ({$signed($signed((reg2617 && reg2445)))})
                begin
                  for (forvar2701 = (1'h0); (forvar2701 < (2'h3)); forvar2701 = (forvar2701 + (1'h1)))
                    begin
                      reg2702 <= reg2660[(4'h8):(2'h3)];
                      reg2703 <= $signed((~$unsigned((&(8'hac)))));
                    end
                end
              else
                begin
                  reg2701 <= {forvar2656[(2'h2):(2'h2)]};
                  reg2702 <= $unsigned(reg2390[(1'h0):(1'h0)]);
                  if ((($unsigned(((8'ha0) - reg2637)) * forvar2656) || $unsigned($unsigned(reg2621[(2'h2):(2'h2)]))))
                    begin
                      reg2703 <= {reg2602};
                      reg2704 <= $unsigned($unsigned($signed(forvar2677)));
                      reg2705 <= (8'hb9);
                      reg2706 <= reg2540[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg2703 <= $signed(forvar2677);
                    end
                  reg2707 <= ((((-forvar2388) >>> $unsigned(wire2374)) & reg2425[(1'h0):(1'h0)]) ^~ reg2701[(4'h8):(3'h7)]);
                end
              if (reg2471[(3'h5):(2'h2)])
                begin
                  reg2708 <= $signed(reg2668[(1'h1):(1'h1)]);
                  for (forvar2709 = (1'h0); (forvar2709 < (1'h0)); forvar2709 = (forvar2709 + (1'h1)))
                    begin
                      reg2710 <= ($unsigned($unsigned((^~reg2469))) & ((reg2681[(3'h7):(2'h2)] ?
                          reg2508[(4'ha):(3'h6)] : (!reg2688)) & $unsigned(reg2491[(2'h3):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar2708 = (1'h0); (forvar2708 < (2'h2)); forvar2708 = (forvar2708 + (1'h1)))
                    begin
                      reg2709 <= reg2555[(1'h1):(1'h0)];
                      reg2710 <= {(~^$signed(reg2540))};
                    end
                  for (forvar2711 = (1'h0); (forvar2711 < (1'h0)); forvar2711 = (forvar2711 + (1'h1)))
                    begin
                      reg2712 <= $unsigned($signed({forvar2486}));
                      reg2713 <= ($unsigned($unsigned(reg2489[(2'h2):(1'h0)])) || $unsigned({$signed(reg2699)}));
                      reg2714 <= {reg2637[(3'h5):(1'h1)]};
                    end
                  if (reg2619[(4'hb):(1'h0)])
                    begin
                      reg2715 <= reg2416;
                    end
                  else
                    begin
                      reg2715 <= $signed(forvar2394);
                      reg2716 <= forvar2620[(4'h8):(4'h8)];
                    end
                end
              reg2717 <= reg2387;
            end
          else
            begin
              if ($signed($signed((~^(&reg2487)))))
                begin
                  if (reg2379[(2'h2):(2'h2)])
                    begin
                      reg2701 <= reg2628;
                      reg2702 <= (reg2610 >= ({{wire2375}} ?
                          $signed((reg2597 <<< (8'ha7))) : $unsigned($signed((8'ha2)))));
                      reg2703 <= $signed({(~&$signed(forvar2662))});
                      reg2704 <= forvar2472;
                    end
                  else
                    begin
                      reg2701 <= $unsigned((~|((reg2479 || reg2618) ?
                          forvar2625 : reg2510)));
                      reg2702 <= reg2521[(1'h0):(1'h0)];
                      reg2703 <= reg2539[(2'h3):(1'h0)];
                      reg2704 <= $signed((((~reg2645) ?
                          (^reg2509) : $signed(forvar2696)) >> $unsigned((-reg2666))));
                    end
                  reg2705 <= reg2698;
                  if ((reg2377[(4'h9):(1'h0)] ?
                      ((~&(~&forvar2674)) * (reg2630 & reg2583[(2'h2):(2'h2)])) : $signed({((8'hb3) ?
                              reg2409 : reg2555)})))
                    begin
                      reg2706 <= reg2429[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg2706 <= ($unsigned($signed((forvar2520 ?
                          reg2554 : reg2509))) || (8'ha0));
                      reg2707 <= (($unsigned((forvar2708 ? reg2507 : reg2582)) ?
                          {reg2661} : $signed($signed((8'h9c)))) || {(!$unsigned((8'hb2)))});
                      reg2708 <= $unsigned(reg2505[(4'h9):(4'h9)]);
                      reg2709 <= $signed((reg2553[(4'h9):(3'h4)] ?
                          ($signed(forvar2625) + reg2527) : reg2704));
                    end
                end
              else
                begin
                  if (({((+reg2611) ?
                              reg2695[(3'h6):(1'h0)] : $signed(reg2428))} ?
                      forvar2550[(2'h3):(1'h0)] : reg2509[(3'h6):(3'h5)]))
                    begin
                      reg2701 <= reg2598;
                      reg2702 <= $signed($unsigned(reg2389[(4'hc):(1'h0)]));
                      reg2703 <= forvar2382;
                      reg2704 <= reg2491;
                    end
                  else
                    begin
                      reg2701 <= $signed($signed($signed(reg2593[(3'h4):(2'h2)])));
                    end
                end
              for (forvar2710 = (1'h0); (forvar2710 < (1'h0)); forvar2710 = (forvar2710 + (1'h1)))
                begin
                  if ($unsigned($unsigned((~reg2681))))
                    begin
                      reg2711 <= reg2602[(4'h9):(4'h9)];
                      reg2712 <= $signed(((!$signed(reg2709)) ?
                          reg2609 : ($signed(forvar2438) ?
                              $unsigned(forvar2391) : $signed(forvar2626))));
                    end
                  else
                    begin
                      reg2711 <= (-$unsigned((~reg2636[(3'h5):(2'h2)])));
                      reg2712 <= (8'hba);
                      reg2713 <= $signed((reg2683[(2'h3):(2'h2)] && (&(!(8'hb4)))));
                    end
                  for (forvar2714 = (1'h0); (forvar2714 < (1'h0)); forvar2714 = (forvar2714 + (1'h1)))
                    begin
                      reg2715 <= (~^((|reg2592) <= reg2542[(2'h3):(1'h0)]));
                      reg2716 <= $unsigned($unsigned(reg2670));
                      reg2717 <= (($unsigned((reg2496 <= reg2523)) ?
                          (~&((8'ha4) ^ reg2698)) : (forvar2449[(1'h1):(1'h0)] ?
                              $unsigned((8'ha4)) : $signed(wire2546))) << {{reg2386}});
                    end
                end
            end
        end
      else
        begin
          for (forvar2701 = (1'h0); (forvar2701 < (1'h0)); forvar2701 = (forvar2701 + (1'h1)))
            begin
              for (forvar2702 = (1'h0); (forvar2702 < (1'h1)); forvar2702 = (forvar2702 + (1'h1)))
                begin
                  for (forvar2703 = (1'h0); (forvar2703 < (2'h3)); forvar2703 = (forvar2703 + (1'h1)))
                    begin
                      reg2704 <= $signed($signed($unsigned({forvar2518})));
                      reg2705 <= $signed((~|($signed(forvar2385) ?
                          {(8'hb7)} : (reg2670 - forvar2530))));
                    end
                  if (reg2650[(1'h0):(1'h0)])
                    begin
                      reg2706 <= reg2706[(4'hd):(2'h3)];
                      reg2707 <= (~&(forvar2452[(2'h3):(2'h2)] >>> reg2646[(1'h0):(1'h0)]));
                      reg2708 <= $signed(reg2669[(4'hb):(4'h9)]);
                    end
                  else
                    begin
                      reg2706 <= ((+wire2371[(2'h2):(2'h2)]) ?
                          $signed((^~$signed(reg2414))) : ($signed($signed(reg2633)) ^ ($signed(reg2514) ?
                              (forvar2571 ?
                                  forvar2631 : (8'ha2)) : $signed(reg2617))));
                      reg2707 <= {$unsigned(((reg2459 ?
                              forvar2638 : reg2577) && wire2543))};
                      reg2708 <= forvar2541[(4'h9):(1'h0)];
                      reg2709 <= reg2555[(1'h0):(1'h0)];
                    end
                end
              for (forvar2710 = (1'h0); (forvar2710 < (2'h3)); forvar2710 = (forvar2710 + (1'h1)))
                begin
                  reg2711 <= (8'haf);
                  reg2712 <= ($unsigned((reg2695[(4'h8):(2'h2)] ?
                      (&reg2539) : (8'ha2))) == ($unsigned($signed(forvar2391)) ?
                      (~^forvar2541[(3'h5):(1'h1)]) : (~(8'h9e))));
                  if ((reg2601 ?
                      (~^(forvar2465 ~^ (forvar2433 && reg2483))) : (|reg2542[(3'h4):(3'h4)])))
                    begin
                      reg2713 <= ((~$unsigned((reg2525 ? reg2708 : reg2406))) ?
                          ((8'hb4) != $unsigned((forvar2452 ?
                              reg2469 : reg2566))) : wire2374[(2'h2):(1'h0)]);
                      reg2714 <= forvar2415;
                      reg2715 <= {(forvar2485[(3'h4):(1'h0)] ?
                              (8'ha9) : (wire2544 ?
                                  reg2587 : $signed(reg2537)))};
                      reg2716 <= (~|forvar2391);
                    end
                  else
                    begin
                      reg2713 <= {(~((~^(8'hb4)) ? (&reg2563) : {reg2454}))};
                      reg2714 <= $unsigned(reg2699);
                    end
                  for (forvar2717 = (1'h0); (forvar2717 < (2'h2)); forvar2717 = (forvar2717 + (1'h1)))
                    begin
                      reg2718 <= {reg2669[(4'h9):(1'h0)]};
                    end
                end
              for (forvar2719 = (1'h0); (forvar2719 < (1'h1)); forvar2719 = (forvar2719 + (1'h1)))
                begin
                  for (forvar2720 = (1'h0); (forvar2720 < (2'h3)); forvar2720 = (forvar2720 + (1'h1)))
                    begin
                      reg2721 <= forvar2648[(4'hd):(4'hd)];
                    end
                  if (wire2368[(4'hf):(4'hd)])
                    begin
                      reg2722 <= reg2487;
                      reg2723 <= reg2410;
                      reg2724 <= reg2477[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2722 <= {$unsigned((~reg2394[(3'h5):(1'h1)]))};
                      reg2723 <= $unsigned(forvar2385);
                    end
                  for (forvar2725 = (1'h0); (forvar2725 < (2'h3)); forvar2725 = (forvar2725 + (1'h1)))
                    begin
                      reg2726 <= reg2693[(2'h3):(2'h2)];
                      reg2727 <= reg2383[(2'h3):(2'h3)];
                      reg2728 <= $signed((reg2568[(3'h5):(3'h5)] ?
                          ((~forvar2674) ?
                              (+(8'ha1)) : (reg2561 << (8'h9f))) : ((forvar2664 ~^ (8'hb9)) ?
                              (reg2407 == reg2471) : (reg2490 <<< reg2602))));
                      reg2729 <= ({$signed((~reg2682))} ?
                          reg2379 : reg2387[(1'h0):(1'h0)]);
                    end
                end
              for (forvar2730 = (1'h0); (forvar2730 < (1'h1)); forvar2730 = (forvar2730 + (1'h1)))
                begin
                  reg2731 <= wire2375;
                  reg2732 <= forvar2408[(2'h2):(1'h0)];
                  if ((~^reg2383[(3'h5):(2'h2)]))
                    begin
                      reg2733 <= {((reg2692 == $signed(forvar2675)) ?
                              $signed(wire2371[(3'h4):(1'h0)]) : ($unsigned((8'hae)) | {wire2373}))};
                      reg2734 <= reg2426[(2'h2):(1'h0)];
                      reg2735 <= forvar2407;
                      reg2736 <= reg2528[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg2733 <= $signed($signed(forvar2691));
                    end
                end
            end
          if (reg2426[(1'h0):(1'h0)])
            begin
              reg2737 <= {{((reg2396 << reg2639) ?
                          reg2534[(1'h0):(1'h0)] : $unsigned(reg2661))}};
              for (forvar2738 = (1'h0); (forvar2738 < (2'h3)); forvar2738 = (forvar2738 + (1'h1)))
                begin
                  for (forvar2739 = (1'h0); (forvar2739 < (2'h3)); forvar2739 = (forvar2739 + (1'h1)))
                    begin
                      reg2740 <= (-((~reg2512[(3'h5):(3'h4)]) ?
                          ((^reg2470) ?
                              $signed(reg2453) : ((8'hb3) & (8'ha9))) : $signed($unsigned(reg2672))));
                    end
                  for (forvar2741 = (1'h0); (forvar2741 < (1'h0)); forvar2741 = (forvar2741 + (1'h1)))
                    begin
                      reg2742 <= ({((-reg2549) ?
                              (8'h9c) : (^reg2621))} < ($signed($signed(reg2661)) ?
                          (reg2629 & (!(8'hba))) : ((8'ha9) != ((8'ha2) > forvar2500))));
                    end
                  reg2743 <= $unsigned({forvar2739});
                end
              if ((((^~$unsigned((8'ha2))) | forvar2620) ?
                  reg2524[(2'h3):(1'h0)] : $unsigned(({reg2589} <= $signed(reg2535)))))
                begin
                  if (reg2511)
                    begin
                      reg2744 <= $signed(reg2553);
                      reg2745 <= (+$signed(forvar2599[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg2744 <= ((|reg2519[(2'h2):(1'h1)]) ?
                          ({reg2444} ?
                              (reg2469[(3'h4):(1'h0)] ?
                                  (reg2678 ?
                                      reg2614 : forvar2709) : {reg2718}) : ($unsigned(forvar2739) ^~ (reg2699 != reg2550))) : $signed($unsigned($unsigned(reg2744))));
                      reg2745 <= {($unsigned($signed(reg2590)) >> reg2701[(2'h3):(1'h0)])};
                    end
                end
              else
                begin
                  for (forvar2744 = (1'h0); (forvar2744 < (1'h0)); forvar2744 = (forvar2744 + (1'h1)))
                    begin
                      reg2745 <= $signed(($unsigned((-forvar2388)) ?
                          reg2452 : $signed($signed((8'ha2)))));
                      reg2746 <= ($unsigned(({reg2573} | $signed(reg2446))) ^~ reg2535);
                      reg2747 <= reg2529;
                      reg2748 <= (|(8'h9c));
                    end
                  for (forvar2749 = (1'h0); (forvar2749 < (2'h3)); forvar2749 = (forvar2749 + (1'h1)))
                    begin
                      reg2750 <= reg2702;
                    end
                end
            end
          else
            begin
              for (forvar2737 = (1'h0); (forvar2737 < (2'h2)); forvar2737 = (forvar2737 + (1'h1)))
                begin
                  for (forvar2738 = (1'h0); (forvar2738 < (1'h1)); forvar2738 = (forvar2738 + (1'h1)))
                    begin
                      reg2739 <= (!($unsigned(forvar2551) ?
                          (forvar2418[(2'h2):(1'h0)] ?
                              (reg2619 ?
                                  reg2448 : (8'h9e)) : reg2576) : forvar2675[(2'h3):(2'h2)]));
                      reg2740 <= $signed($unsigned($unsigned(reg2497[(2'h3):(2'h3)])));
                      reg2741 <= $signed($unsigned(((reg2453 ^ forvar2663) ?
                          (reg2459 ? forvar2386 : forvar2445) : (^reg2701))));
                      reg2742 <= {reg2668[(2'h3):(1'h1)]};
                    end
                  reg2743 <= reg2512;
                  reg2744 <= $signed(forvar2418[(1'h0):(1'h0)]);
                end
            end
        end
      for (forvar2751 = (1'h0); (forvar2751 < (2'h3)); forvar2751 = (forvar2751 + (1'h1)))
        begin
          for (forvar2752 = (1'h0); (forvar2752 < (2'h3)); forvar2752 = (forvar2752 + (1'h1)))
            begin
              reg2753 <= ($unsigned($unsigned(forvar2501)) > ($signed((reg2710 ~^ forvar2508)) ?
                  reg2669[(3'h6):(3'h4)] : ((&reg2688) >> ((8'hb0) ?
                      forvar2449 : wire2545))));
            end
          for (forvar2754 = (1'h0); (forvar2754 < (2'h2)); forvar2754 = (forvar2754 + (1'h1)))
            begin
              if (reg2579)
                begin
                  if ((8'hb7))
                    begin
                      reg2755 <= forvar2446[(3'h7):(2'h2)];
                      reg2756 <= {{forvar2388}};
                    end
                  else
                    begin
                      reg2755 <= (~forvar2668);
                    end
                  for (forvar2757 = (1'h0); (forvar2757 < (2'h3)); forvar2757 = (forvar2757 + (1'h1)))
                    begin
                      reg2758 <= (8'h9f);
                      reg2759 <= $signed((~|(8'hb9)));
                      reg2760 <= ((~$signed((&(8'hb4)))) ?
                          {forvar2500[(2'h2):(1'h1)]} : $signed($unsigned({reg2562})));
                    end
                end
              else
                begin
                  if ($signed($unsigned(reg2451[(4'hb):(3'h5)])))
                    begin
                      reg2755 <= (reg2412[(3'h4):(3'h4)] || ((~&$unsigned((8'hb3))) ?
                          ((reg2600 ? reg2676 : reg2399) ?
                              reg2383[(3'h4):(2'h2)] : reg2432[(2'h2):(1'h0)]) : (reg2623 ?
                              $signed(reg2672) : reg2520[(1'h0):(1'h0)])));
                      reg2756 <= (!((8'haa) << $signed($unsigned(forvar2389))));
                    end
                  else
                    begin
                      reg2755 <= reg2586[(1'h0):(1'h0)];
                      reg2756 <= $signed((^~$signed(reg2721[(2'h3):(1'h0)])));
                      reg2757 <= (|reg2564[(2'h2):(2'h2)]);
                      reg2758 <= reg2535[(3'h7):(2'h3)];
                    end
                  reg2759 <= {$unsigned((8'ha7))};
                  if (reg2412)
                    begin
                      reg2760 <= $signed(reg2713[(4'ha):(4'ha)]);
                      reg2761 <= (8'hae);
                      reg2762 <= wire2545;
                    end
                  else
                    begin
                      reg2760 <= $unsigned((~($signed((8'h9d)) + (+(8'hb8)))));
                      reg2761 <= (^$unsigned(($unsigned(reg2739) + (forvar2615 < reg2744))));
                      reg2762 <= {$unsigned($signed((+reg2616)))};
                    end
                end
              for (forvar2763 = (1'h0); (forvar2763 < (2'h3)); forvar2763 = (forvar2763 + (1'h1)))
                begin
                  reg2764 <= $unsigned((|reg2621));
                  if ((~&(~&$signed(((8'hb9) ? reg2531 : (8'hb7))))))
                    begin
                      reg2765 <= (reg2756 ?
                          reg2416[(2'h2):(1'h0)] : (-($signed(reg2682) ?
                              $unsigned(reg2427) : $unsigned(forvar2387))));
                      reg2766 <= reg2420[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2765 <= $unsigned((reg2710[(4'ha):(3'h5)] ?
                          forvar2575 : (forvar2625[(4'hc):(2'h2)] << {forvar2554})));
                      reg2766 <= $unsigned(forvar2565[(3'h4):(2'h2)]);
                    end
                  for (forvar2767 = (1'h0); (forvar2767 < (2'h3)); forvar2767 = (forvar2767 + (1'h1)))
                    begin
                      reg2768 <= (reg2662 ? reg2423 : $unsigned((8'hb6)));
                      reg2769 <= reg2514[(2'h3):(2'h3)];
                      reg2770 <= reg2488;
                      reg2771 <= wire2374[(3'h4):(3'h4)];
                    end
                  if ($signed({$signed($signed(forvar2378))}))
                    begin
                      reg2772 <= $signed(reg2620[(4'h8):(4'h8)]);
                      reg2773 <= (^$signed({(+reg2664)}));
                      reg2774 <= ($unsigned(((~reg2704) * (reg2593 ?
                          reg2612 : forvar2560))) > {$signed($signed(reg2422))});
                    end
                  else
                    begin
                      reg2772 <= ($unsigned($unsigned((reg2466 <<< reg2451))) + (($signed(forvar2502) >> $signed(reg2456)) ^ (^$unsigned(forvar2413))));
                      reg2773 <= $unsigned((($signed(reg2423) <= (reg2400 - forvar2749)) ?
                          reg2671 : $signed($signed(reg2597))));
                      reg2774 <= (($signed(((8'h9d) * reg2535)) ?
                          (~|{reg2744}) : {(reg2433 ?
                                  reg2640 : (8'hb0))}) + ((^~forvar2677[(1'h0):(1'h0)]) & $unsigned((8'ha5))));
                    end
                end
              if ($signed({$signed(reg2721[(4'hd):(4'hc)])}))
                begin
                  for (forvar2775 = (1'h0); (forvar2775 < (1'h1)); forvar2775 = (forvar2775 + (1'h1)))
                    begin
                      reg2776 <= (^~(forvar2420[(1'h1):(1'h0)] >>> (-(8'hb2))));
                    end
                  if ($unsigned(({{reg2705}} && (^$unsigned(reg2705)))))
                    begin
                      reg2777 <= reg2512[(1'h1):(1'h0)];
                      reg2778 <= $signed($unsigned($unsigned($signed(reg2406))));
                      reg2779 <= ($signed((&$signed(wire2368))) >>> $unsigned({(reg2557 > reg2616)}));
                      reg2780 <= $signed(reg2639);
                    end
                  else
                    begin
                      reg2777 <= reg2408;
                      reg2778 <= {reg2744[(2'h2):(2'h2)]};
                      reg2779 <= $signed((forvar2690 ?
                          (^~(forvar2591 ?
                              forvar2457 : forvar2465)) : (|reg2542[(1'h0):(1'h0)])));
                      reg2780 <= forvar2575[(3'h7):(3'h4)];
                    end
                end
              else
                begin
                  reg2775 <= $unsigned(reg2393);
                end
            end
          for (forvar2781 = (1'h0); (forvar2781 < (1'h0)); forvar2781 = (forvar2781 + (1'h1)))
            begin
              if (((($unsigned((8'hb2)) ?
                      reg2464[(1'h1):(1'h0)] : (forvar2579 <= (8'hb0))) ?
                  (-$unsigned(reg2693)) : reg2505[(1'h1):(1'h1)]) ^~ $signed($unsigned((reg2387 + forvar2550)))))
                begin
                  for (forvar2782 = (1'h0); (forvar2782 < (1'h1)); forvar2782 = (forvar2782 + (1'h1)))
                    begin
                      reg2783 <= (reg2477 ?
                          ($unsigned($unsigned(reg2671)) > (8'ha2)) : reg2529[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar2782 = (1'h0); (forvar2782 < (1'h0)); forvar2782 = (forvar2782 + (1'h1)))
                    begin
                      reg2783 <= forvar2472;
                    end
                  for (forvar2784 = (1'h0); (forvar2784 < (1'h0)); forvar2784 = (forvar2784 + (1'h1)))
                    begin
                      reg2785 <= $unsigned((8'hab));
                      reg2786 <= $unsigned((reg2529[(1'h0):(1'h0)] ?
                          (forvar2720[(4'hd):(2'h2)] ?
                              (reg2562 - forvar2609) : (forvar2515 ?
                                  reg2534 : reg2603)) : reg2616));
                      reg2787 <= $unsigned((reg2405 ?
                          {{forvar2473}} : reg2496[(3'h4):(2'h2)]));
                    end
                  if (forvar2378)
                    begin
                      reg2788 <= ((reg2745[(1'h1):(1'h1)] && (reg2718 < (~|reg2658))) != ($unsigned(reg2768[(2'h2):(2'h2)]) ?
                          forvar2530[(1'h0):(1'h0)] : $unsigned((8'ha3))));
                      reg2789 <= reg2663[(1'h1):(1'h0)];
                      reg2790 <= ((((reg2536 ? forvar2397 : reg2478) ?
                          ((8'hb6) ?
                              reg2622 : forvar2668) : (reg2755 && reg2584)) << ($unsigned(reg2583) ?
                          {reg2681} : (reg2460 ?
                              forvar2422 : reg2483))) - reg2427[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg2788 <= (reg2683[(2'h2):(2'h2)] ?
                          $unsigned($unsigned((!forvar2751))) : reg2452[(4'hb):(3'h4)]);
                      reg2789 <= ($signed(((reg2440 ?
                          forvar2670 : forvar2501) >= (forvar2613 >= (8'hb1)))) - {reg2733[(2'h3):(2'h2)]});
                      reg2790 <= forvar2625;
                    end
                  reg2791 <= (^$signed((reg2597[(4'hb):(3'h7)] >> (8'hb0))));
                end
              for (forvar2792 = (1'h0); (forvar2792 < (2'h2)); forvar2792 = (forvar2792 + (1'h1)))
                begin
                  if ({$unsigned($unsigned($signed(reg2470)))})
                    begin
                      reg2793 <= (8'h9e);
                    end
                  else
                    begin
                      reg2793 <= reg2572[(4'ha):(2'h2)];
                      reg2794 <= ($unsigned($signed({reg2621})) >>> $signed(($signed((8'ha0)) >> (reg2609 ?
                          reg2671 : reg2587))));
                      reg2795 <= $signed({reg2668});
                    end
                  reg2796 <= $unsigned((^~reg2721));
                end
              if (((|wire2368[(1'h1):(1'h1)]) ^~ {(^(reg2480 > (8'ha6)))}))
                begin
                  for (forvar2797 = (1'h0); (forvar2797 < (2'h2)); forvar2797 = (forvar2797 + (1'h1)))
                    begin
                      reg2798 <= {(wire2374 | $signed((reg2391 || reg2724)))};
                      reg2799 <= $signed($unsigned((-reg2616)));
                    end
                end
              else
                begin
                  for (forvar2797 = (1'h0); (forvar2797 < (2'h3)); forvar2797 = (forvar2797 + (1'h1)))
                    begin
                      reg2798 <= $signed(reg2403);
                      reg2799 <= ((+(reg2755[(2'h2):(2'h2)] ?
                          (reg2692 ~^ reg2570) : reg2604[(3'h5):(2'h2)])) ~^ ((^reg2601[(1'h0):(1'h0)]) <= (~|((8'hb3) ?
                          forvar2664 : reg2506))));
                      reg2800 <= (+(($signed((8'hac)) ?
                              (reg2524 ?
                                  forvar2388 : reg2519) : (reg2454 - reg2497)) ?
                          reg2610[(1'h0):(1'h0)] : ((~&forvar2503) << ((8'ha4) >> reg2707))));
                    end
                  reg2801 <= (^~(~&reg2429[(2'h2):(1'h0)]));
                  for (forvar2802 = (1'h0); (forvar2802 < (2'h3)); forvar2802 = (forvar2802 + (1'h1)))
                    begin
                      reg2803 <= {reg2602[(4'h8):(3'h7)]};
                      reg2804 <= ((reg2536 == ($unsigned(reg2699) ?
                              (~^reg2412) : forvar2677[(2'h3):(1'h1)])) ?
                          $signed(reg2381[(3'h4):(2'h3)]) : $signed($signed($signed(reg2612))));
                    end
                  for (forvar2805 = (1'h0); (forvar2805 < (2'h2)); forvar2805 = (forvar2805 + (1'h1)))
                    begin
                      reg2806 <= {reg2758[(1'h1):(1'h0)]};
                      reg2807 <= reg2612[(1'h0):(1'h0)];
                      reg2808 <= $signed($unsigned(((reg2390 ?
                          reg2480 : reg2727) <= reg2423[(1'h1):(1'h1)])));
                      reg2809 <= $signed((-(^reg2552[(2'h3):(1'h1)])));
                    end
                end
              for (forvar2810 = (1'h0); (forvar2810 < (1'h1)); forvar2810 = (forvar2810 + (1'h1)))
                begin
                  for (forvar2811 = (1'h0); (forvar2811 < (1'h1)); forvar2811 = (forvar2811 + (1'h1)))
                    begin
                      reg2812 <= reg2714[(2'h2):(1'h1)];
                    end
                  for (forvar2813 = (1'h0); (forvar2813 < (2'h2)); forvar2813 = (forvar2813 + (1'h1)))
                    begin
                      reg2814 <= forvar2717;
                      reg2815 <= ($signed(forvar2385[(2'h3):(2'h3)]) ?
                          $signed(reg2547[(3'h4):(1'h0)]) : reg2387[(3'h5):(1'h1)]);
                      reg2816 <= (($unsigned(((8'hb3) ? reg2385 : forvar2642)) ?
                          (reg2479[(3'h4):(2'h2)] ?
                              {reg2475} : reg2639[(2'h2):(1'h1)]) : reg2406[(2'h3):(1'h0)]) == $unsigned(($signed(reg2390) ?
                          reg2721[(4'h8):(4'h8)] : reg2556[(1'h0):(1'h0)])));
                    end
                  for (forvar2817 = (1'h0); (forvar2817 < (1'h0)); forvar2817 = (forvar2817 + (1'h1)))
                    begin
                      reg2818 <= $signed($unsigned($unsigned($unsigned((8'ha1)))));
                      reg2819 <= $unsigned($signed(forvar2591[(4'h8):(2'h2)]));
                      reg2820 <= {reg2549};
                      reg2821 <= forvar2668;
                    end
                  for (forvar2822 = (1'h0); (forvar2822 < (1'h0)); forvar2822 = (forvar2822 + (1'h1)))
                    begin
                      reg2823 <= {(~forvar2388)};
                      reg2824 <= forvar2730[(4'h9):(3'h6)];
                    end
                end
            end
        end
    end
  assign wire2825 = ($signed(reg2436) ?
                        $unsigned(forvar2418[(1'h0):(1'h0)]) : ($signed($signed(reg2475)) ?
                            ((reg2552 ? forvar2382 : reg2567) <= (reg2666 ?
                                forvar2670 : reg2607)) : forvar2423[(2'h2):(1'h0)]));
  always
    @(posedge clk) begin
      reg2826 <= reg2388[(1'h0):(1'h0)];
      for (forvar2827 = (1'h0); (forvar2827 < (2'h3)); forvar2827 = (forvar2827 + (1'h1)))
        begin
          if (($signed($unsigned(reg2731)) * forvar2656[(4'hb):(2'h2)]))
            begin
              for (forvar2828 = (1'h0); (forvar2828 < (1'h1)); forvar2828 = (forvar2828 + (1'h1)))
                begin
                  if (((forvar2642[(3'h6):(3'h4)] ?
                          forvar2554 : (forvar2541[(1'h1):(1'h1)] ?
                              (reg2398 ?
                                  (8'hb6) : reg2723) : forvar2389[(3'h6):(1'h1)])) ?
                      forvar2518[(1'h1):(1'h1)] : {{$signed(reg2557)}}))
                    begin
                      reg2829 <= $unsigned(({$unsigned(reg2451)} ?
                          $unsigned((reg2384 >>> reg2427)) : $unsigned($unsigned(reg2378))));
                      reg2830 <= ($signed($unsigned($signed((8'ha9)))) ?
                          reg2508 : forvar2613);
                    end
                  else
                    begin
                      reg2829 <= (!($unsigned((~|reg2718)) ~^ (^(reg2532 ?
                          forvar2822 : reg2496))));
                      reg2830 <= (|reg2396);
                    end
                  for (forvar2831 = (1'h0); (forvar2831 < (2'h2)); forvar2831 = (forvar2831 + (1'h1)))
                    begin
                      reg2832 <= (reg2724 ?
                          (((forvar2420 || forvar2642) ?
                              (-forvar2763) : (8'ha2)) | (^~(reg2567 || reg2496))) : forvar2725[(3'h4):(2'h2)]);
                    end
                  for (forvar2833 = (1'h0); (forvar2833 < (2'h3)); forvar2833 = (forvar2833 + (1'h1)))
                    begin
                      reg2834 <= (8'h9d);
                      reg2835 <= (~reg2718);
                      reg2836 <= $signed(reg2804);
                    end
                  reg2837 <= (+reg2496[(2'h2):(2'h2)]);
                end
              for (forvar2838 = (1'h0); (forvar2838 < (1'h1)); forvar2838 = (forvar2838 + (1'h1)))
                begin
                  for (forvar2839 = (1'h0); (forvar2839 < (1'h0)); forvar2839 = (forvar2839 + (1'h1)))
                    begin
                      reg2840 <= ($signed(reg2693) ?
                          reg2627 : $unsigned(reg2796[(3'h7):(3'h6)]));
                      reg2841 <= $unsigned((|(|((8'ha1) ? (8'hb6) : reg2530))));
                      reg2842 <= forvar2548[(4'ha):(3'h6)];
                    end
                  if (reg2623)
                    begin
                      reg2843 <= ($unsigned(({reg2498} | $signed(reg2771))) ?
                          reg2427 : reg2708[(1'h0):(1'h0)]);
                      reg2844 <= {((|(reg2684 ? reg2439 : forvar2518)) ?
                              $signed((~forvar2407)) : reg2654)};
                    end
                  else
                    begin
                      reg2843 <= (((!$unsigned(reg2785)) ?
                              $signed((^(8'had))) : $unsigned((~^reg2576))) ?
                          $unsigned(reg2680[(1'h0):(1'h0)]) : $signed($signed((reg2771 <<< forvar2754))));
                      reg2844 <= ($signed((+$unsigned((8'h9e)))) & reg2814[(3'h7):(2'h2)]);
                    end
                end
              for (forvar2845 = (1'h0); (forvar2845 < (1'h0)); forvar2845 = (forvar2845 + (1'h1)))
                begin
                  for (forvar2846 = (1'h0); (forvar2846 < (2'h2)); forvar2846 = (forvar2846 + (1'h1)))
                    begin
                      reg2847 <= $unsigned(($unsigned(forvar2717) ?
                          $unsigned(reg2692[(4'hb):(1'h1)]) : $unsigned($signed((8'hb2)))));
                      reg2848 <= $signed({(forvar2620[(2'h3):(2'h2)] ?
                              reg2651[(2'h3):(2'h3)] : reg2819)});
                    end
                  for (forvar2849 = (1'h0); (forvar2849 < (2'h2)); forvar2849 = (forvar2849 + (1'h1)))
                    begin
                      reg2850 <= ($unsigned($signed(wire2372)) ?
                          ($unsigned((reg2798 & (8'hba))) ?
                              {$unsigned((8'hb7))} : ((^(8'ha6)) ^ reg2829[(4'hb):(2'h3)])) : ((!(forvar2408 == reg2753)) ?
                              ($unsigned(forvar2591) || reg2630[(3'h5):(2'h2)]) : forvar2565));
                    end
                  for (forvar2851 = (1'h0); (forvar2851 < (1'h0)); forvar2851 = (forvar2851 + (1'h1)))
                    begin
                      reg2852 <= ($signed({$signed(forvar2702)}) ?
                          (~reg2620) : (($signed(reg2609) ?
                              $unsigned(reg2808) : reg2570[(4'h8):(3'h6)]) ^~ $unsigned((8'ha0))));
                      reg2853 <= {forvar2485};
                      reg2854 <= $unsigned(wire2546[(3'h7):(3'h4)]);
                    end
                end
            end
          else
            begin
              if ($unsigned((|reg2657[(4'h8):(1'h1)])))
                begin
                  if ((reg2816[(1'h1):(1'h0)] ?
                      reg2617 : {$unsigned($unsigned(forvar2418))}))
                    begin
                      reg2828 <= (($unsigned($signed(forvar2473)) ?
                              (reg2528[(4'ha):(3'h7)] - reg2540[(3'h5):(1'h1)]) : ($signed(reg2487) ?
                                  (~&reg2843) : (reg2790 > forvar2379))) ?
                          $signed(reg2847) : {(~$signed(reg2533))});
                    end
                  else
                    begin
                      reg2828 <= $unsigned($signed(($unsigned(reg2629) ?
                          $unsigned(reg2676) : (reg2414 ~^ reg2430))));
                      reg2829 <= $signed((&reg2746[(2'h2):(2'h2)]));
                    end
                  if ((^($signed((reg2786 ? (8'hb8) : forvar2394)) ?
                      {reg2588} : $unsigned($unsigned(forvar2811)))))
                    begin
                      reg2830 <= $signed(reg2801[(3'h6):(3'h4)]);
                      reg2831 <= reg2744;
                      reg2832 <= $signed({$signed($signed(reg2539))});
                    end
                  else
                    begin
                      reg2830 <= {{{(forvar2548 && reg2420)}}};
                      reg2831 <= $unsigned(({{forvar2805}} ?
                          {(forvar2664 ?
                                  forvar2415 : forvar2391)} : ({reg2570} ?
                              reg2786 : $signed(reg2392))));
                      reg2832 <= ((~(^$signed((8'ha1)))) || $unsigned(forvar2379[(2'h3):(1'h0)]));
                    end
                  if ({$unsigned(($signed((8'hae)) << reg2449[(4'hd):(3'h5)]))})
                    begin
                      reg2833 <= ((reg2440[(3'h5):(2'h2)] ?
                          $signed((reg2722 ^ reg2490)) : (~|$signed(reg2384))) <<< (&(~&$unsigned(reg2598))));
                    end
                  else
                    begin
                      reg2833 <= $unsigned({$unsigned(forvar2638)});
                      reg2834 <= (~(~|(|(^reg2576))));
                      reg2835 <= ((-$signed($signed(forvar2558))) ?
                          (^~$unsigned($unsigned(reg2549))) : {({reg2743} ?
                                  reg2837[(1'h1):(1'h1)] : {reg2395})});
                      reg2836 <= $signed(reg2412);
                    end
                end
              else
                begin
                  for (forvar2828 = (1'h0); (forvar2828 < (1'h0)); forvar2828 = (forvar2828 + (1'h1)))
                    begin
                      reg2829 <= (reg2497[(4'h9):(3'h6)] ?
                          (^~(&{reg2577})) : $unsigned(forvar2599));
                    end
                end
            end
          if ((~forvar2611[(3'h5):(1'h0)]))
            begin
              for (forvar2855 = (1'h0); (forvar2855 < (2'h3)); forvar2855 = (forvar2855 + (1'h1)))
                begin
                  for (forvar2856 = (1'h0); (forvar2856 < (1'h1)); forvar2856 = (forvar2856 + (1'h1)))
                    begin
                      reg2857 <= reg2570[(2'h3):(2'h2)];
                      reg2858 <= reg2513;
                      reg2859 <= reg2731;
                      reg2860 <= (^reg2522[(4'h8):(3'h6)]);
                    end
                  for (forvar2861 = (1'h0); (forvar2861 < (2'h3)); forvar2861 = (forvar2861 + (1'h1)))
                    begin
                      reg2862 <= reg2466;
                      reg2863 <= $signed((~&$signed((&reg2835))));
                    end
                end
            end
          else
            begin
              for (forvar2855 = (1'h0); (forvar2855 < (1'h0)); forvar2855 = (forvar2855 + (1'h1)))
                begin
                  reg2856 <= {(~&(forvar2413 ~^ $signed(reg2460)))};
                  reg2857 <= (8'hb1);
                  if ($signed($signed((^~$unsigned((8'hb7))))))
                    begin
                      reg2858 <= forvar2503[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg2858 <= ($unsigned(reg2460[(2'h2):(1'h1)]) ?
                          $signed(((reg2506 >> reg2673) || $signed((8'ha0)))) : (($unsigned(reg2511) >>> (^reg2383)) ^~ $signed($unsigned(reg2844))));
                      reg2859 <= $unsigned({{reg2481}});
                    end
                end
              if ((~^(!{$signed(reg2525)})))
                begin
                  for (forvar2860 = (1'h0); (forvar2860 < (1'h0)); forvar2860 = (forvar2860 + (1'h1)))
                    begin
                      reg2861 <= reg2777;
                      reg2862 <= ((^~(^~$unsigned(reg2759))) ?
                          $unsigned((reg2402 >= $signed(reg2463))) : (forvar2626[(4'h9):(2'h2)] ?
                              (|$signed(reg2422)) : $signed({reg2517})));
                    end
                  reg2863 <= $signed(reg2523);
                  for (forvar2864 = (1'h0); (forvar2864 < (2'h3)); forvar2864 = (forvar2864 + (1'h1)))
                    begin
                      reg2865 <= ((((~|forvar2596) ?
                          (forvar2519 ^ reg2766) : forvar2701[(2'h2):(1'h1)]) ^~ (reg2681 >> (reg2829 ?
                          reg2580 : reg2402))) <= $unsigned($unsigned($unsigned(reg2759))));
                      reg2866 <= reg2841[(4'h8):(1'h0)];
                      reg2867 <= $unsigned(($unsigned((reg2397 ?
                          reg2746 : forvar2828)) >> reg2446[(1'h0):(1'h0)]));
                    end
                  for (forvar2868 = (1'h0); (forvar2868 < (2'h2)); forvar2868 = (forvar2868 + (1'h1)))
                    begin
                      reg2869 <= reg2504;
                      reg2870 <= ($unsigned($unsigned((reg2776 < reg2637))) ?
                          $unsigned(reg2863[(3'h7):(1'h1)]) : ($signed($unsigned(reg2659)) ?
                              (!(8'had)) : reg2709));
                      reg2871 <= {reg2780[(3'h4):(2'h2)]};
                      reg2872 <= (&reg2710);
                    end
                end
              else
                begin
                  if (forvar2596)
                    begin
                      reg2860 <= (8'hb5);
                    end
                  else
                    begin
                      reg2860 <= (reg2865[(4'ha):(2'h3)] - reg2697);
                    end
                  if ((reg2452 - ($signed(((8'ha3) > reg2833)) ?
                      (+(reg2837 ? (8'hb0) : reg2787)) : forvar2781)))
                    begin
                      reg2861 <= $unsigned($unsigned(((reg2700 ?
                              forvar2448 : forvar2452) ?
                          $signed(reg2577) : reg2762[(3'h4):(2'h3)])));
                      reg2862 <= {{(-(wire2543 >>> reg2708))}};
                      reg2863 <= $signed(($signed($signed((8'ha6))) != $unsigned((-reg2441))));
                      reg2864 <= (+reg2401[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg2861 <= (8'hb3);
                      reg2862 <= ((reg2676 ?
                          forvar2613 : {$signed((8'haf))}) > $unsigned(((reg2491 >>> (8'ha3)) ^~ {forvar2805})));
                    end
                end
              reg2873 <= forvar2767[(3'h7):(3'h7)];
            end
        end
    end
  assign wire2874 = reg2410;
  always
    @(posedge clk) begin
      if ($unsigned((8'haf)))
        begin
          for (forvar2875 = (1'h0); (forvar2875 < (1'h0)); forvar2875 = (forvar2875 + (1'h1)))
            begin
              if (((~&$signed((reg2408 != forvar2574))) ?
                  reg2579 : $signed({{reg2436}})))
                begin
                  for (forvar2876 = (1'h0); (forvar2876 < (2'h3)); forvar2876 = (forvar2876 + (1'h1)))
                    begin
                      reg2877 <= forvar2702[(1'h1):(1'h0)];
                      reg2878 <= $signed((forvar2433 ?
                          ((^reg2742) ?
                              (reg2440 >= forvar2500) : $signed(wire2545)) : forvar2450[(4'ha):(4'h8)]));
                      reg2879 <= reg2816[(1'h0):(1'h0)];
                    end
                  for (forvar2880 = (1'h0); (forvar2880 < (2'h2)); forvar2880 = (forvar2880 + (1'h1)))
                    begin
                      reg2881 <= (reg2510 ?
                          $unsigned((!((8'hb4) > (8'hb6)))) : (reg2721[(3'h5):(1'h0)] <= $signed((reg2553 ?
                              reg2640 : forvar2792))));
                      reg2882 <= (8'hb0);
                    end
                  for (forvar2883 = (1'h0); (forvar2883 < (2'h3)); forvar2883 = (forvar2883 + (1'h1)))
                    begin
                      reg2884 <= reg2800;
                      reg2885 <= ((!($unsigned((8'hb4)) ?
                              reg2581 : forvar2784[(4'ha):(2'h3)])) ?
                          (+((reg2600 <= reg2508) ?
                              {forvar2416} : ((8'hb4) ~^ reg2710))) : $signed({((8'hae) ?
                                  reg2645 : reg2729)}));
                      reg2886 <= ((({forvar2413} - (^~reg2525)) != (+$unsigned((8'hab)))) ^~ $unsigned({(~&forvar2656)}));
                      reg2887 <= forvar2560[(2'h2):(1'h0)];
                    end
                  for (forvar2888 = (1'h0); (forvar2888 < (1'h1)); forvar2888 = (forvar2888 + (1'h1)))
                    begin
                      reg2889 <= (|$signed((^$unsigned(reg2757))));
                      reg2890 <= forvar2710;
                    end
                end
              else
                begin
                  for (forvar2876 = (1'h0); (forvar2876 < (2'h3)); forvar2876 = (forvar2876 + (1'h1)))
                    begin
                      reg2877 <= reg2778[(1'h1):(1'h1)];
                      reg2878 <= ($signed((|(^forvar2711))) ?
                          $signed(((&reg2669) ^ (^forvar2738))) : reg2771[(2'h2):(1'h0)]);
                      reg2879 <= ((reg2861 ?
                              ($unsigned((8'ha7)) ^ $signed((8'hb4))) : ((-(8'hb6)) ?
                                  forvar2856[(3'h7):(3'h5)] : $signed((8'ha7)))) ?
                          reg2475[(2'h2):(1'h1)] : wire2376);
                      reg2880 <= $signed($unsigned({(8'h9d)}));
                    end
                  for (forvar2881 = (1'h0); (forvar2881 < (2'h2)); forvar2881 = (forvar2881 + (1'h1)))
                    begin
                      reg2882 <= (($unsigned((~forvar2465)) ?
                              (reg2873 ?
                                  $unsigned(wire2374) : {forvar2738}) : ((|reg2713) || (reg2576 ?
                                  (8'had) : reg2632))) ?
                          ((~|$unsigned((8'hb4))) ?
                              reg2668 : (((8'hb8) ?
                                  wire2544 : forvar2846) - forvar2501)) : {reg2388});
                      reg2883 <= $unsigned($unsigned(reg2828));
                      reg2884 <= {reg2647[(3'h7):(3'h5)]};
                    end
                  if ((forvar2754 ?
                      (~reg2783[(1'h1):(1'h1)]) : (~|((reg2863 ?
                              reg2758 : reg2693) ?
                          (8'hae) : $unsigned(forvar2554)))))
                    begin
                      reg2885 <= ($signed(((forvar2529 ?
                              reg2553 : forvar2674) || reg2400)) ?
                          $unsigned((reg2549[(1'h0):(1'h0)] ?
                              forvar2554 : {reg2507})) : (reg2821[(2'h3):(2'h2)] ?
                              reg2636 : (~|reg2819[(3'h7):(2'h3)])));
                      reg2886 <= (forvar2611 ?
                          (reg2510 ~^ $signed($unsigned((8'hb5)))) : (-reg2441[(2'h3):(2'h3)]));
                      reg2887 <= $unsigned(($signed(reg2644) ?
                          $unsigned((~|reg2710)) : $unsigned((reg2889 >= forvar2714))));
                      reg2888 <= reg2401;
                    end
                  else
                    begin
                      reg2885 <= reg2622;
                    end
                  if (reg2382[(3'h6):(1'h0)])
                    begin
                      reg2889 <= reg2604[(2'h2):(1'h0)];
                      reg2890 <= reg2411[(4'he):(4'ha)];
                      reg2891 <= (|(~&((~^forvar2579) & $signed(reg2389))));
                      reg2892 <= $unsigned((((+reg2509) ?
                          (^(8'h9c)) : forvar2875[(1'h0):(1'h0)]) + (+(~|reg2427))));
                    end
                  else
                    begin
                      reg2889 <= {({$signed(forvar2752)} ?
                              (((8'ha2) < reg2536) ?
                                  $signed(reg2882) : $signed((8'hb5))) : $unsigned(reg2578))};
                      reg2890 <= ($unsigned((~^reg2440[(4'hd):(2'h2)])) ?
                          reg2505 : $signed($unsigned($unsigned(forvar2415))));
                    end
                end
              if ($signed($signed(({reg2389} ?
                  $unsigned(forvar2389) : (reg2794 ? reg2723 : reg2389)))))
                begin
                  reg2893 <= {$signed(($signed((8'h9c)) ?
                          (^reg2589) : {reg2889}))};
                  for (forvar2894 = (1'h0); (forvar2894 < (2'h2)); forvar2894 = (forvar2894 + (1'h1)))
                    begin
                      reg2895 <= ($signed(((^~(8'hac)) ?
                              reg2521 : forvar2579)) ?
                          $unsigned(reg2688) : (~|((~^reg2840) ?
                              (&reg2853) : (reg2718 || (8'ha8)))));
                    end
                  for (forvar2896 = (1'h0); (forvar2896 < (2'h3)); forvar2896 = (forvar2896 + (1'h1)))
                    begin
                      reg2897 <= $signed(forvar2565[(4'hc):(4'h8)]);
                      reg2898 <= $signed($unsigned(reg2746));
                      reg2899 <= reg2521[(1'h0):(1'h0)];
                      reg2900 <= $unsigned((((reg2379 - (8'hb5)) <= (~^reg2430)) <<< ($signed(forvar2828) ?
                          (8'hb0) : reg2380[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  for (forvar2893 = (1'h0); (forvar2893 < (1'h0)); forvar2893 = (forvar2893 + (1'h1)))
                    begin
                      reg2894 <= $signed((~^(reg2461[(1'h1):(1'h1)] ?
                          $unsigned(reg2415) : $signed(forvar2856))));
                      reg2895 <= $signed(({{forvar2422}} > $signed(reg2477[(3'h5):(2'h2)])));
                      reg2896 <= forvar2674;
                    end
                  for (forvar2897 = (1'h0); (forvar2897 < (2'h3)); forvar2897 = (forvar2897 + (1'h1)))
                    begin
                      reg2898 <= (~&reg2882[(2'h3):(1'h0)]);
                      reg2899 <= {(reg2773[(2'h2):(1'h0)] ^~ (&(reg2895 * reg2768)))};
                      reg2900 <= forvar2664[(1'h1):(1'h1)];
                      reg2901 <= {$unsigned(reg2419)};
                    end
                  for (forvar2902 = (1'h0); (forvar2902 < (2'h2)); forvar2902 = (forvar2902 + (1'h1)))
                    begin
                      reg2903 <= $unsigned((({reg2816} >>> reg2791[(4'hf):(4'he)]) ?
                          $signed($signed((8'had))) : $unsigned(reg2708[(3'h4):(2'h2)])));
                    end
                end
              if ({(+reg2898)})
                begin
                  for (forvar2904 = (1'h0); (forvar2904 < (2'h3)); forvar2904 = (forvar2904 + (1'h1)))
                    begin
                      reg2905 <= $unsigned((forvar2418 ?
                          ({forvar2473} ?
                              (reg2644 ?
                                  forvar2382 : (8'ha6)) : {(8'hb6)}) : $unsigned(reg2471[(1'h0):(1'h0)])));
                      reg2906 <= $unsigned(reg2398);
                      reg2907 <= (reg2521 ?
                          $signed(reg2753) : (forvar2397 << $unsigned((+reg2440))));
                      reg2908 <= ((((^forvar2383) >= {reg2898}) >= {reg2441[(2'h2):(2'h2)]}) * (-{$signed(reg2736)}));
                    end
                  for (forvar2909 = (1'h0); (forvar2909 < (1'h1)); forvar2909 = (forvar2909 + (1'h1)))
                    begin
                      reg2910 <= reg2529[(3'h5):(1'h1)];
                      reg2911 <= (~|$unsigned(forvar2626[(1'h0):(1'h0)]));
                      reg2912 <= reg2895[(3'h4):(3'h4)];
                    end
                  if ((|((reg2434[(4'h9):(2'h2)] ?
                      (reg2480 >= reg2606) : forvar2398) == $signed(forvar2416[(3'h4):(2'h2)]))))
                    begin
                      reg2913 <= (($signed(reg2464) + $signed($signed(forvar2520))) >>> (8'ha3));
                    end
                  else
                    begin
                      reg2913 <= reg2568[(1'h0):(1'h0)];
                      reg2914 <= $signed($unsigned(reg2721[(1'h1):(1'h0)]));
                      reg2915 <= {forvar2881};
                      reg2916 <= (({(reg2624 < reg2681)} * forvar2511[(3'h7):(2'h3)]) ?
                          $signed(reg2683) : ({$signed(reg2381)} ?
                              {$unsigned(reg2403)} : forvar2883[(4'hd):(4'hb)]));
                    end
                end
              else
                begin
                  if ((~^(8'ha0)))
                    begin
                      reg2904 <= reg2658;
                      reg2905 <= $unsigned($signed((8'h9c)));
                      reg2906 <= ((forvar2754 ?
                          reg2890[(3'h4):(2'h2)] : forvar2822) >>> ($unsigned($unsigned(reg2870)) ?
                          (8'ha9) : ($signed((8'haf)) & $unsigned((8'haa)))));
                      reg2907 <= (8'hba);
                    end
                  else
                    begin
                      reg2904 <= $unsigned(((8'haf) ? (8'hb2) : reg2411));
                      reg2905 <= (-((~&reg2416) ?
                          reg2684[(3'h6):(2'h2)] : reg2647[(4'h9):(2'h2)]));
                      reg2906 <= reg2612[(1'h0):(1'h0)];
                      reg2907 <= $unsigned((^~$signed($signed(reg2383))));
                    end
                end
            end
          reg2917 <= (($signed($signed(reg2906)) ?
                  (reg2463 ?
                      $signed(reg2517) : ((8'h9d) | reg2761)) : ((-reg2786) >> reg2778)) ?
              {(|((8'hab) >= reg2859))} : $signed(forvar2511));
        end
      else
        begin
          if (reg2383)
            begin
              for (forvar2875 = (1'h0); (forvar2875 < (2'h2)); forvar2875 = (forvar2875 + (1'h1)))
                begin
                  if ((forvar2708 ? forvar2508 : reg2665))
                    begin
                      reg2876 <= reg2476[(4'hc):(4'hc)];
                    end
                  else
                    begin
                      reg2876 <= ($unsigned(reg2713) ?
                          reg2861[(4'hf):(3'h4)] : $signed($unsigned((8'hb2))));
                      reg2877 <= $unsigned((!((~&reg2886) & (reg2568 == (8'hb3)))));
                      reg2878 <= ($signed((~^{reg2824})) >> (-(reg2561 ?
                          $signed(forvar2457) : reg2384)));
                    end
                  reg2879 <= $signed({(|$signed(forvar2709))});
                  for (forvar2880 = (1'h0); (forvar2880 < (2'h3)); forvar2880 = (forvar2880 + (1'h1)))
                    begin
                      reg2881 <= reg2622;
                    end
                  if (forvar2822[(3'h4):(1'h1)])
                    begin
                      reg2882 <= forvar2703[(4'ha):(1'h0)];
                      reg2883 <= reg2761[(2'h3):(2'h3)];
                      reg2884 <= $unsigned($signed((((8'h9e) ?
                              reg2604 : reg2820) ?
                          reg2633 : reg2460)));
                    end
                  else
                    begin
                      reg2882 <= reg2475;
                      reg2883 <= {$signed((reg2689 ?
                              (forvar2388 ?
                                  reg2884 : forvar2662) : $signed(forvar2571)))};
                    end
                end
              for (forvar2885 = (1'h0); (forvar2885 < (2'h2)); forvar2885 = (forvar2885 + (1'h1)))
                begin
                  if (($unsigned($unsigned(reg2844)) * $signed(reg2382)))
                    begin
                      reg2886 <= (~&((forvar2782[(1'h1):(1'h1)] ?
                              ((8'ha5) ?
                                  reg2870 : forvar2792) : ((8'hac) ^~ forvar2875)) ?
                          ($unsigned(reg2460) ?
                              reg2671[(1'h1):(1'h0)] : $signed(forvar2501)) : reg2400));
                      reg2887 <= $signed((forvar2717[(3'h5):(1'h1)] ?
                          ($signed(reg2718) >>> reg2569[(3'h5):(3'h4)]) : (~{forvar2482})));
                    end
                  else
                    begin
                      reg2886 <= $signed((!{(forvar2492 ? reg2449 : (8'hba))}));
                      reg2887 <= ({reg2678} ?
                          $signed((^~{forvar2503})) : ({(reg2435 <<< reg2734)} ^~ (~|(reg2907 ?
                              forvar2596 : forvar2452))));
                      reg2888 <= (reg2466[(3'h6):(3'h5)] ?
                          {((!reg2379) ?
                                  (reg2831 > reg2766) : (8'hae))} : forvar2529[(2'h2):(1'h1)]);
                      reg2889 <= reg2519;
                    end
                  reg2890 <= ((reg2512 ? reg2437 : reg2807[(2'h2):(2'h2)]) ?
                      $unsigned($signed((reg2569 == (8'ha8)))) : (~|(reg2750[(3'h4):(2'h3)] ?
                          $unsigned(reg2709) : $signed(reg2858))));
                  for (forvar2891 = (1'h0); (forvar2891 < (1'h0)); forvar2891 = (forvar2891 + (1'h1)))
                    begin
                      reg2892 <= ((($signed(forvar2875) ?
                          $signed((8'h9f)) : $signed(reg2821)) >> $signed({forvar2643})) >= $unsigned(($unsigned(reg2681) << ((8'haa) ?
                          reg2391 : reg2508))));
                    end
                  for (forvar2893 = (1'h0); (forvar2893 < (2'h2)); forvar2893 = (forvar2893 + (1'h1)))
                    begin
                      reg2894 <= reg2914;
                      reg2895 <= (forvar2625[(3'h7):(3'h7)] ?
                          $signed(reg2798) : $signed((~(reg2487 & (8'h9c)))));
                      reg2896 <= $unsigned((~^{{reg2699}}));
                    end
                end
            end
          else
            begin
              for (forvar2875 = (1'h0); (forvar2875 < (1'h0)); forvar2875 = (forvar2875 + (1'h1)))
                begin
                  for (forvar2876 = (1'h0); (forvar2876 < (2'h2)); forvar2876 = (forvar2876 + (1'h1)))
                    begin
                      reg2877 <= ((|reg2676) >>> reg2533);
                      reg2878 <= reg2793;
                      reg2879 <= (-(^$unsigned((forvar2751 ~^ reg2406))));
                    end
                  reg2880 <= ($signed((8'hb4)) * reg2847[(4'he):(4'h8)]);
                end
              for (forvar2881 = (1'h0); (forvar2881 < (1'h0)); forvar2881 = (forvar2881 + (1'h1)))
                begin
                  for (forvar2882 = (1'h0); (forvar2882 < (2'h3)); forvar2882 = (forvar2882 + (1'h1)))
                    begin
                      reg2883 <= (~|(8'ha8));
                      reg2884 <= forvar2413[(4'ha):(3'h5)];
                      reg2885 <= ((+(^(reg2431 && forvar2503))) | (!{((8'hb8) && reg2892)}));
                      reg2886 <= ((8'hb6) ?
                          forvar2485[(1'h1):(1'h1)] : (^$unsigned((~forvar2385))));
                    end
                  if ({$signed($signed((~^reg2679)))})
                    begin
                      reg2887 <= (~^(($unsigned(reg2736) == forvar2881) != forvar2861[(2'h2):(1'h0)]));
                      reg2888 <= $signed((($unsigned(reg2444) >> reg2458[(3'h4):(1'h0)]) ?
                          $signed((reg2439 ?
                              forvar2709 : reg2635)) : reg2470[(1'h1):(1'h1)]));
                      reg2889 <= (({$unsigned(reg2636)} ?
                              $signed((reg2619 ?
                                  reg2453 : (8'ha3))) : (^$signed(reg2491))) ?
                          {$signed(reg2387[(4'h8):(3'h5)])} : reg2686[(1'h1):(1'h1)]);
                      reg2890 <= forvar2882;
                    end
                  else
                    begin
                      reg2887 <= $unsigned((8'hb0));
                    end
                end
            end
        end
      for (forvar2918 = (1'h0); (forvar2918 < (1'h0)); forvar2918 = (forvar2918 + (1'h1)))
        begin
          for (forvar2919 = (1'h0); (forvar2919 < (2'h2)); forvar2919 = (forvar2919 + (1'h1)))
            begin
              for (forvar2920 = (1'h0); (forvar2920 < (2'h3)); forvar2920 = (forvar2920 + (1'h1)))
                begin
                  for (forvar2921 = (1'h0); (forvar2921 < (1'h0)); forvar2921 = (forvar2921 + (1'h1)))
                    begin
                      reg2922 <= forvar2529;
                      reg2923 <= ($unsigned(reg2852[(1'h1):(1'h0)]) == $unsigned(($signed(reg2734) ?
                          (forvar2554 ? reg2862 : reg2632) : reg2632)));
                      reg2924 <= ((^forvar2519) << {((reg2417 ?
                                  (8'ha3) : reg2800) ?
                              (forvar2919 ?
                                  forvar2560 : reg2864) : (~forvar2893))});
                    end
                  reg2925 <= (~|(forvar2625[(4'hd):(4'h8)] ?
                      (+(forvar2641 & reg2441)) : (reg2425 << (-reg2613))));
                  for (forvar2926 = (1'h0); (forvar2926 < (2'h2)); forvar2926 = (forvar2926 + (1'h1)))
                    begin
                      reg2927 <= reg2462;
                      reg2928 <= $signed(((8'hb0) <<< {(forvar2377 >> forvar2861)}));
                    end
                  for (forvar2929 = (1'h0); (forvar2929 < (1'h0)); forvar2929 = (forvar2929 + (1'h1)))
                    begin
                      reg2930 <= (reg2787[(3'h5):(2'h3)] ?
                          {$signed($unsigned(forvar2415))} : (reg2508 | reg2870));
                      reg2931 <= reg2804[(2'h2):(2'h2)];
                    end
                end
            end
          for (forvar2932 = (1'h0); (forvar2932 < (1'h0)); forvar2932 = (forvar2932 + (1'h1)))
            begin
              for (forvar2933 = (1'h0); (forvar2933 < (1'h1)); forvar2933 = (forvar2933 + (1'h1)))
                begin
                  for (forvar2934 = (1'h0); (forvar2934 < (2'h2)); forvar2934 = (forvar2934 + (1'h1)))
                    begin
                      reg2935 <= $signed($unsigned($signed(wire2370)));
                      reg2936 <= {($unsigned($unsigned(reg2390)) ?
                              $unsigned($signed(reg2393)) : {{reg2889}})};
                      reg2937 <= reg2406;
                    end
                  reg2938 <= $unsigned(reg2529);
                end
              for (forvar2939 = (1'h0); (forvar2939 < (1'h1)); forvar2939 = (forvar2939 + (1'h1)))
                begin
                  for (forvar2940 = (1'h0); (forvar2940 < (2'h2)); forvar2940 = (forvar2940 + (1'h1)))
                    begin
                      reg2941 <= reg2592[(4'h8):(3'h7)];
                      reg2942 <= (~$unsigned((8'hb1)));
                    end
                  for (forvar2943 = (1'h0); (forvar2943 < (2'h2)); forvar2943 = (forvar2943 + (1'h1)))
                    begin
                      reg2944 <= (^reg2776[(3'h6):(1'h0)]);
                    end
                end
            end
          if ($unsigned(reg2645[(3'h7):(1'h1)]))
            begin
              if ($unsigned($signed(((&reg2523) ^~ $unsigned(reg2663)))))
                begin
                  for (forvar2945 = (1'h0); (forvar2945 < (1'h0)); forvar2945 = (forvar2945 + (1'h1)))
                    begin
                      reg2946 <= ((($signed(reg2478) ?
                              reg2941[(3'h6):(1'h0)] : (wire2545 >> reg2878)) ?
                          (!$unsigned(reg2679)) : (reg2711 ?
                              forvar2710[(3'h4):(1'h1)] : reg2837)) & $unsigned($signed(reg2862[(1'h1):(1'h0)])));
                      reg2947 <= (~&forvar2416[(3'h5):(1'h1)]);
                      reg2948 <= forvar2655[(4'hd):(4'hd)];
                    end
                  reg2949 <= ($signed((!{reg2520})) ?
                      $unsigned(reg2403[(3'h5):(1'h0)]) : (({reg2764} ?
                              $unsigned(reg2561) : {reg2384}) ?
                          $signed((reg2740 != forvar2754)) : reg2880[(3'h7):(3'h4)]));
                  if ((^~{$signed($signed(reg2528))}))
                    begin
                      reg2950 <= ($unsigned($unsigned((reg2621 ?
                              reg2685 : forvar2434))) ?
                          ((reg2531[(1'h1):(1'h1)] ?
                                  reg2448[(2'h2):(1'h0)] : $unsigned(forvar2394)) ?
                              $unsigned({reg2700}) : reg2676) : reg2916);
                    end
                  else
                    begin
                      reg2950 <= (~|({$unsigned(forvar2415)} + reg2700[(2'h3):(1'h0)]));
                      reg2951 <= (reg2598 != (8'ha0));
                      reg2952 <= ((reg2628 ?
                          ({(8'ha3)} ?
                              reg2910 : (forvar2851 << reg2542)) : ($signed((8'ha3)) < (wire2874 | reg2378))) >> ($unsigned((reg2583 ?
                              (8'h9d) : reg2732)) ?
                          $unsigned($signed((8'ha9))) : {reg2938}));
                      reg2953 <= reg2775[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar2945 = (1'h0); (forvar2945 < (1'h0)); forvar2945 = (forvar2945 + (1'h1)))
                    begin
                      reg2946 <= ($unsigned((!(+forvar2448))) ?
                          $unsigned($signed(reg2498[(3'h6):(1'h1)])) : $signed($signed((reg2467 >>> reg2867))));
                      reg2947 <= $unsigned((^~reg2481[(1'h1):(1'h1)]));
                    end
                end
            end
          else
            begin
              reg2945 <= (reg2390[(2'h2):(2'h2)] ?
                  $signed(reg2456[(4'h8):(3'h6)]) : reg2609);
              reg2946 <= reg2722;
            end
        end
      reg2954 <= ({reg2778[(1'h0):(1'h0)]} ?
          {((~^forvar2448) >= $unsigned(reg2685))} : $unsigned(({reg2728} || (~&reg2685))));
      if ({$signed($signed((+reg2916)))})
        begin
          for (forvar2955 = (1'h0); (forvar2955 < (1'h0)); forvar2955 = (forvar2955 + (1'h1)))
            begin
              if ($signed(((reg2911 >>> reg2741) != (wire2369 & ((8'ha2) & forvar2885)))))
                begin
                  for (forvar2956 = (1'h0); (forvar2956 < (1'h0)); forvar2956 = (forvar2956 + (1'h1)))
                    begin
                      reg2957 <= $signed($unsigned($unsigned((~(8'hba)))));
                      reg2958 <= $signed(reg2394[(4'h8):(3'h7)]);
                    end
                  if ((!reg2665))
                    begin
                      reg2959 <= reg2740[(3'h7):(3'h4)];
                      reg2960 <= (reg2883[(3'h6):(1'h0)] ?
                          (~|$signed($unsigned((8'hb0)))) : (~reg2947));
                      reg2961 <= $signed(reg2463[(1'h1):(1'h1)]);
                      reg2962 <= $signed(forvar2625[(4'hc):(3'h5)]);
                    end
                  else
                    begin
                      reg2959 <= {(reg2742 ? reg2566 : reg2439[(1'h1):(1'h1)])};
                    end
                  for (forvar2963 = (1'h0); (forvar2963 < (2'h2)); forvar2963 = (forvar2963 + (1'h1)))
                    begin
                      reg2964 <= ((8'ha3) | ($unsigned($unsigned(forvar2797)) << (8'h9d)));
                    end
                  for (forvar2965 = (1'h0); (forvar2965 < (2'h2)); forvar2965 = (forvar2965 + (1'h1)))
                    begin
                      reg2966 <= ((|{{reg2517}}) == (|$unsigned({reg2907})));
                    end
                end
              else
                begin
                  if ($unsigned({((!reg2779) ?
                          (reg2442 ? (8'ha7) : reg2948) : (8'ha4))}))
                    begin
                      reg2956 <= ($unsigned(reg2627) ^ (!($signed(reg2382) & reg2387[(1'h1):(1'h1)])));
                      reg2957 <= (($unsigned($signed((8'hb8))) ?
                          (((8'h9d) ^ forvar2797) ?
                              reg2964 : $signed(reg2723)) : forvar2574) ~^ forvar2775[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg2956 <= reg2892[(2'h3):(2'h2)];
                      reg2957 <= ($unsigned(reg2452[(2'h2):(1'h1)]) ?
                          $signed($signed($unsigned(reg2664))) : (|{forvar2465}));
                    end
                  reg2958 <= $signed(reg2689[(1'h1):(1'h0)]);
                  if (forvar2433[(3'h6):(1'h1)])
                    begin
                      reg2959 <= (&(^(8'hb2)));
                      reg2960 <= (~|$unsigned((((8'ha3) ?
                          reg2658 : reg2603) || {(8'ha3)})));
                      reg2961 <= ($signed($unsigned(reg2646)) ?
                          (~&($signed(forvar2730) - (~reg2595))) : forvar2450);
                    end
                  else
                    begin
                      reg2959 <= ((~reg2521) ^~ $signed(reg2786));
                      reg2960 <= (~&reg2829);
                    end
                end
              reg2967 <= $unsigned((reg2403[(2'h2):(1'h0)] ?
                  forvar2448 : (^~reg2836)));
              for (forvar2968 = (1'h0); (forvar2968 < (1'h0)); forvar2968 = (forvar2968 + (1'h1)))
                begin
                  reg2969 <= $unsigned(reg2561);
                  reg2970 <= ($signed((^(reg2794 - reg2404))) << $unsigned((-$signed(reg2686))));
                end
            end
          reg2971 <= $unsigned((forvar2855 ?
              ($signed(reg2602) >>> (reg2441 ? (8'hb8) : reg2724)) : reg2669));
          for (forvar2972 = (1'h0); (forvar2972 < (2'h2)); forvar2972 = (forvar2972 + (1'h1)))
            begin
              for (forvar2973 = (1'h0); (forvar2973 < (1'h1)); forvar2973 = (forvar2973 + (1'h1)))
                begin
                  for (forvar2974 = (1'h0); (forvar2974 < (1'h0)); forvar2974 = (forvar2974 + (1'h1)))
                    begin
                      reg2975 <= (reg2410[(1'h0):(1'h0)] ?
                          reg2832[(4'ha):(3'h7)] : ($unsigned({forvar2383}) == $unsigned((&forvar2741))));
                      reg2976 <= (~|$unsigned(forvar2394));
                      reg2977 <= reg2481;
                      reg2978 <= (reg2732[(2'h2):(1'h0)] ?
                          (+(^~(reg2841 ? reg2382 : (8'hb6)))) : (reg2807 ?
                              reg2589[(2'h3):(2'h3)] : (~|forvar2620)));
                    end
                  for (forvar2979 = (1'h0); (forvar2979 < (1'h0)); forvar2979 = (forvar2979 + (1'h1)))
                    begin
                      reg2980 <= ($signed(((reg2615 && reg2687) ?
                              forvar2648[(3'h6):(2'h3)] : $signed(forvar2527))) ?
                          reg2461[(2'h2):(2'h2)] : (^~(&{reg2441})));
                    end
                  for (forvar2981 = (1'h0); (forvar2981 < (2'h2)); forvar2981 = (forvar2981 + (1'h1)))
                    begin
                      reg2982 <= {$signed($unsigned((forvar2445 ?
                              forvar2730 : forvar2894)))};
                    end
                end
              for (forvar2983 = (1'h0); (forvar2983 < (2'h3)); forvar2983 = (forvar2983 + (1'h1)))
                begin
                  for (forvar2984 = (1'h0); (forvar2984 < (2'h3)); forvar2984 = (forvar2984 + (1'h1)))
                    begin
                      reg2985 <= reg2391;
                      reg2986 <= {$unsigned(($unsigned(reg2688) ?
                              (reg2428 ?
                                  forvar2415 : forvar2560) : $signed(reg2850)))};
                      reg2987 <= $signed((8'hb7));
                    end
                  if ($signed((-reg2395[(1'h1):(1'h0)])))
                    begin
                      reg2988 <= (($signed((8'haf)) ?
                              $signed(forvar2575[(3'h5):(2'h3)]) : (^reg2402)) ?
                          $signed((+$signed(reg2678))) : {(reg2853[(2'h2):(1'h1)] ?
                                  {reg2563} : (reg2779 < forvar2620))});
                      reg2989 <= (^~(~&$unsigned({reg2891})));
                    end
                  else
                    begin
                      reg2988 <= (&(((|reg2679) ?
                              (forvar2670 ? reg2888 : reg2789) : reg2942) ?
                          ((forvar2638 || reg2470) ?
                              (reg2951 == reg2894) : (reg2714 ?
                                  reg2451 : reg2531)) : $unsigned($signed(reg2916))));
                      reg2989 <= (reg2731[(4'h8):(4'h8)] - $signed((|forvar2691)));
                    end
                end
              for (forvar2990 = (1'h0); (forvar2990 < (2'h2)); forvar2990 = (forvar2990 + (1'h1)))
                begin
                  for (forvar2991 = (1'h0); (forvar2991 < (2'h2)); forvar2991 = (forvar2991 + (1'h1)))
                    begin
                      reg2992 <= ($unsigned((8'ha6)) ?
                          $unsigned(($signed((8'hb9)) == (reg2773 ?
                              reg2441 : reg2881))) : (^(reg2953 & (reg2666 ?
                              (8'hb0) : reg2709))));
                      reg2993 <= (+reg2448);
                      reg2994 <= (!reg2837);
                    end
                end
              if (reg2454)
                begin
                  reg2995 <= {($unsigned(((8'ha9) ? reg2931 : reg2739)) ?
                          reg2694[(3'h7):(3'h7)] : reg2697[(2'h3):(2'h2)])};
                  if (reg2538)
                    begin
                      reg2996 <= ((!(~(8'hb8))) ~^ reg2514[(3'h5):(1'h1)]);
                      reg2997 <= {$signed($unsigned({reg2967}))};
                      reg2998 <= reg2682;
                    end
                  else
                    begin
                      reg2996 <= (^~reg2605[(2'h2):(1'h1)]);
                      reg2997 <= (($signed({reg2899}) == (forvar2739 ?
                          reg2447[(3'h4):(2'h3)] : reg2722[(4'h8):(1'h0)])) != $unsigned(((reg2636 ?
                              reg2858 : reg2455) ?
                          (~|reg2609) : reg2727)));
                      reg2998 <= $signed($unsigned($signed(((8'hb9) ^ reg2904))));
                    end
                end
              else
                begin
                  for (forvar2995 = (1'h0); (forvar2995 < (1'h0)); forvar2995 = (forvar2995 + (1'h1)))
                    begin
                      reg2996 <= $unsigned(reg2734);
                    end
                end
            end
        end
      else
        begin
          if (({reg2422} ?
              {$signed(reg2431[(2'h2):(2'h2)])} : (~(^~{reg2581}))))
            begin
              for (forvar2955 = (1'h0); (forvar2955 < (2'h3)); forvar2955 = (forvar2955 + (1'h1)))
                begin
                  reg2956 <= ($unsigned(reg2867) ^ $unsigned(reg2714[(1'h0):(1'h0)]));
                  for (forvar2957 = (1'h0); (forvar2957 < (2'h2)); forvar2957 = (forvar2957 + (1'h1)))
                    begin
                      reg2958 <= $unsigned(wire2825[(1'h1):(1'h0)]);
                      reg2959 <= ((reg2997 ?
                              ((forvar2875 ? forvar2893 : forvar2662) ?
                                  $unsigned(reg2653) : (forvar2631 ?
                                      (8'hb0) : forvar2615)) : (+(-forvar2656))) ?
                          ($unsigned({reg2445}) ?
                              forvar2902 : reg2906) : ($signed(forvar2757) ^~ reg2841));
                      reg2960 <= reg2510[(4'h9):(3'h5)];
                    end
                end
              if (reg2879)
                begin
                  if ($unsigned((^($signed(forvar2965) ?
                      reg2837 : (forvar2921 ? reg2993 : reg2833)))))
                    begin
                      reg2961 <= ((^~$signed({forvar2939})) ?
                          reg2478[(4'h8):(3'h6)] : forvar2737[(2'h2):(1'h1)]);
                      reg2962 <= ((^~reg2956[(3'h5):(2'h2)]) & {$unsigned({reg2998})});
                      reg2963 <= {reg2799[(2'h2):(1'h0)]};
                    end
                  else
                    begin
                      reg2961 <= $signed(reg2858);
                      reg2962 <= reg2533[(3'h5):(2'h2)];
                    end
                  if (reg2841)
                    begin
                      reg2964 <= (forvar2472[(3'h7):(2'h2)] ?
                          $signed(reg2538) : ({reg2534} ?
                              reg2901 : $unsigned({forvar2891})));
                      reg2965 <= (forvar2608[(3'h6):(3'h5)] <<< reg2899);
                      reg2966 <= $unsigned((forvar2452[(3'h7):(2'h3)] ~^ (|(forvar2880 & forvar2894))));
                    end
                  else
                    begin
                      reg2964 <= $signed((&(((8'ha0) ? reg2758 : (8'ha8)) ?
                          $unsigned(reg2622) : forvar2921[(2'h3):(2'h3)])));
                      reg2965 <= $signed(reg2594);
                      reg2966 <= reg2736[(1'h0):(1'h0)];
                    end
                  for (forvar2967 = (1'h0); (forvar2967 < (2'h2)); forvar2967 = (forvar2967 + (1'h1)))
                    begin
                      reg2968 <= ((8'hac) - {(~reg2474[(1'h1):(1'h1)])});
                    end
                  if ((reg2819 | forvar2991[(1'h0):(1'h0)]))
                    begin
                      reg2969 <= $unsigned((!(~^{(8'haa)})));
                    end
                  else
                    begin
                      reg2969 <= $unsigned(({{forvar2445}} == {$unsigned(forvar2663)}));
                      reg2970 <= (reg2618 >= $unsigned($signed($unsigned(reg2624))));
                    end
                end
              else
                begin
                  for (forvar2961 = (1'h0); (forvar2961 < (2'h3)); forvar2961 = (forvar2961 + (1'h1)))
                    begin
                      reg2962 <= ((+($unsigned(reg2477) <= $unsigned(reg2487))) ?
                          $signed(reg2954[(3'h5):(3'h4)]) : {reg2953});
                      reg2963 <= forvar2784[(4'h9):(3'h7)];
                      reg2964 <= $signed(reg2580[(1'h1):(1'h1)]);
                      reg2965 <= $unsigned($unsigned(reg2966[(1'h1):(1'h1)]));
                    end
                end
              for (forvar2971 = (1'h0); (forvar2971 < (2'h3)); forvar2971 = (forvar2971 + (1'h1)))
                begin
                  for (forvar2972 = (1'h0); (forvar2972 < (1'h1)); forvar2972 = (forvar2972 + (1'h1)))
                    begin
                      reg2973 <= {{{((8'hb8) ? reg2987 : forvar2920)}}};
                    end
                  for (forvar2974 = (1'h0); (forvar2974 < (1'h0)); forvar2974 = (forvar2974 + (1'h1)))
                    begin
                      reg2975 <= reg2853;
                    end
                  if ({$unsigned({reg2997})})
                    begin
                      reg2976 <= (forvar2610 ?
                          forvar2717[(2'h2):(1'h1)] : reg2526[(3'h7):(3'h7)]);
                    end
                  else
                    begin
                      reg2976 <= $unsigned(reg2597);
                      reg2977 <= $signed((&((!(8'hb4)) < $signed(reg2964))));
                      reg2978 <= forvar2990;
                      reg2979 <= {((reg2678[(2'h2):(2'h2)] - (forvar2861 ?
                              reg2774 : reg2676)) - reg2681[(4'h9):(1'h0)])};
                    end
                end
              for (forvar2980 = (1'h0); (forvar2980 < (1'h1)); forvar2980 = (forvar2980 + (1'h1)))
                begin
                  for (forvar2981 = (1'h0); (forvar2981 < (1'h0)); forvar2981 = (forvar2981 + (1'h1)))
                    begin
                      reg2982 <= (8'hb7);
                      reg2983 <= reg2812[(4'hc):(3'h4)];
                    end
                end
            end
          else
            begin
              for (forvar2955 = (1'h0); (forvar2955 < (2'h3)); forvar2955 = (forvar2955 + (1'h1)))
                begin
                  for (forvar2956 = (1'h0); (forvar2956 < (1'h0)); forvar2956 = (forvar2956 + (1'h1)))
                    begin
                      reg2957 <= forvar2457[(4'he):(1'h0)];
                      reg2958 <= (~|(reg2912[(3'h4):(1'h0)] >= ((reg2478 & reg2462) >> (8'hb8))));
                      reg2959 <= (~^$signed(reg2450[(4'h8):(2'h3)]));
                      reg2960 <= {(($unsigned(forvar2894) >>> $signed(reg2789)) ?
                              $unsigned((reg2505 ?
                                  forvar2972 : forvar2703)) : (8'hb4))};
                    end
                  for (forvar2961 = (1'h0); (forvar2961 < (2'h3)); forvar2961 = (forvar2961 + (1'h1)))
                    begin
                      reg2962 <= forvar2434;
                    end
                  reg2963 <= $unsigned((^$unsigned($unsigned(forvar2720))));
                end
            end
          for (forvar2984 = (1'h0); (forvar2984 < (1'h1)); forvar2984 = (forvar2984 + (1'h1)))
            begin
              reg2985 <= {(!forvar2967[(3'h4):(2'h2)])};
              for (forvar2986 = (1'h0); (forvar2986 < (1'h1)); forvar2986 = (forvar2986 + (1'h1)))
                begin
                  for (forvar2987 = (1'h0); (forvar2987 < (2'h3)); forvar2987 = (forvar2987 + (1'h1)))
                    begin
                      reg2988 <= (^(8'ha4));
                      reg2989 <= $unsigned((reg2406 ?
                          (&((8'h9d) ? reg2606 : reg2732)) : (8'ha2)));
                      reg2990 <= (8'hb4);
                      reg2991 <= $signed(reg2995);
                    end
                  reg2992 <= reg2497;
                  if (((reg2577 ?
                          (!$signed(reg2899)) : ((reg2848 > reg2740) ?
                              (reg2958 & reg2399) : forvar2450)) ?
                      (~^{reg2594}) : (({(8'had)} ? {reg2652} : reg2389) ?
                          {((8'h9d) ? forvar2642 : (8'ha3))} : (~&reg2428))))
                    begin
                      reg2993 <= $signed((+((reg2407 * wire2373) ?
                          $unsigned(reg2682) : $signed(reg2990))));
                      reg2994 <= (8'ha5);
                      reg2995 <= (!($unsigned({reg2602}) != forvar2810));
                      reg2996 <= reg2506;
                    end
                  else
                    begin
                      reg2993 <= reg2830[(4'h8):(1'h0)];
                    end
                end
              if (reg2707[(1'h0):(1'h0)])
                begin
                  for (forvar2997 = (1'h0); (forvar2997 < (1'h1)); forvar2997 = (forvar2997 + (1'h1)))
                    begin
                      reg2998 <= ($signed($unsigned((reg2947 * reg2843))) ?
                          reg2524 : $unsigned(reg2380[(1'h1):(1'h1)]));
                    end
                  reg2999 <= reg2928[(1'h1):(1'h1)];
                  if ({($unsigned((reg2701 > reg2573)) < $signed((~^(8'hb2))))})
                    begin
                      reg3000 <= wire2825;
                      reg3001 <= forvar2856;
                    end
                  else
                    begin
                      reg3000 <= (-reg2547[(2'h2):(1'h0)]);
                      reg3001 <= (~&{forvar2883});
                    end
                end
              else
                begin
                  for (forvar2997 = (1'h0); (forvar2997 < (2'h3)); forvar2997 = (forvar2997 + (1'h1)))
                    begin
                      reg2998 <= forvar2386;
                      reg2999 <= ((((forvar2714 ?
                                  reg2683 : reg2467) || reg2585) ?
                              reg2421[(1'h1):(1'h0)] : $unsigned(reg2650)) ?
                          (($unsigned(reg2481) ?
                                  reg2660[(2'h3):(2'h2)] : ((8'ha9) << reg2898)) ?
                              $unsigned((wire2543 ?
                                  forvar2641 : reg2743)) : reg2586[(3'h4):(3'h4)]) : (+reg2477[(4'hc):(4'hc)]));
                      reg3000 <= ($unsigned(((reg2454 | reg3001) ?
                          (forvar2939 == reg2471) : $signed(reg2995))) <= forvar2965);
                    end
                  if (($signed((8'hb8)) ?
                      $signed(reg2668[(1'h0):(1'h0)]) : $signed((reg2715 && reg2539))))
                    begin
                      reg3001 <= forvar2904[(3'h5):(2'h3)];
                      reg3002 <= {(-(^(&forvar2681)))};
                      reg3003 <= {(reg2712 ?
                              (~(reg2969 ? reg2999 : reg2893)) : reg2624)};
                      reg3004 <= ((forvar2883 >>> ($unsigned(reg2850) >= $signed(forvar2422))) ?
                          ($signed($signed(reg2971)) ?
                              ((forvar2875 >>> reg3001) != reg2480[(4'he):(3'h6)]) : $unsigned((reg2484 > reg2431))) : (reg2474[(3'h6):(2'h3)] > (~^(8'had))));
                    end
                  else
                    begin
                      reg3001 <= forvar2610[(2'h3):(2'h3)];
                      reg3002 <= $unsigned((!(+((8'ha6) ?
                          reg2589 : forvar2378))));
                    end
                  if ((forvar2965[(1'h0):(1'h0)] ?
                      (reg2786[(2'h3):(2'h2)] << {(8'haa)}) : (8'hb8)))
                    begin
                      reg3005 <= $signed($unsigned($unsigned($unsigned(reg2487))));
                      reg3006 <= (reg2460[(3'h7):(1'h1)] <= {forvar2932});
                    end
                  else
                    begin
                      reg3005 <= reg2432[(3'h4):(2'h2)];
                      reg3006 <= $unsigned(forvar2452);
                      reg3007 <= $signed($signed(reg2785[(4'hc):(4'h8)]));
                      reg3008 <= (forvar2608[(3'h6):(3'h5)] == ({reg2554[(4'h9):(2'h3)]} - $unsigned(reg2435[(3'h6):(2'h3)])));
                    end
                end
            end
          reg3009 <= $unsigned(reg2831);
          if (reg2693[(4'h8):(3'h7)])
            begin
              for (forvar3010 = (1'h0); (forvar3010 < (2'h3)); forvar3010 = (forvar3010 + (1'h1)))
                begin
                  if ($signed((reg3005 & $signed((+reg2434)))))
                    begin
                      reg3011 <= forvar2529[(1'h0):(1'h0)];
                      reg3012 <= ((!forvar2389[(1'h0):(1'h0)]) ?
                          ($unsigned((wire2370 && forvar2856)) ?
                              $unsigned((8'ha6)) : ($unsigned(reg2564) ?
                                  reg2609[(1'h1):(1'h1)] : $unsigned(reg2970))) : ({reg2726[(2'h2):(1'h1)]} >>> $unsigned((forvar2418 ?
                              reg2483 : forvar2649))));
                      reg3013 <= $unsigned({$unsigned({reg2970})});
                    end
                  else
                    begin
                      reg3011 <= (|($signed($signed((8'ha6))) - $signed((forvar2511 > reg2937))));
                      reg3012 <= (+(forvar2909[(4'hd):(4'ha)] ?
                          ({reg2542} & reg2687[(3'h6):(3'h5)]) : ($unsigned(reg2871) - (~wire2372))));
                      reg3013 <= reg2572[(4'ha):(1'h1)];
                    end
                end
            end
          else
            begin
              reg3010 <= (^forvar2797);
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3416  (y, clk, wire3421, wire3420, wire3419, wire3418, wire3417);
  output wire [(32'h31):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire3421;
  input wire signed [(4'ha):(1'h0)] wire3420;
  input wire [(4'hf):(1'h0)] wire3419;
  input wire [(4'ha):(1'h0)] wire3418;
  input wire signed [(2'h3):(1'h0)] wire3417;
  wire [(2'h3):(1'h0)] wire3436;
  reg [(4'h9):(1'h0)] reg3435 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire3434;
  wire signed [(4'hd):(1'h0)] wire3432;
  wire [(4'hf):(1'h0)] wire3422;
  assign y = {wire3436, reg3435, wire3434, wire3432, wire3422, (1'h0)};
  assign wire3422 = wire3421;
  module3423 modinst3433 (wire3432, clk, wire3418, wire3419, wire3421, wire3422);
  assign wire3434 = wire3421;
  always
    @(posedge clk) begin
      reg3435 <= wire3419;
    end
  assign wire3436 = (&$signed({wire3422}));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3423  (y, clk, wire3427, wire3426, wire3425, wire3424);
  output wire [(32'h2e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire3427;
  input wire signed [(3'h6):(1'h0)] wire3426;
  input wire [(5'h10):(1'h0)] wire3425;
  input wire signed [(4'hf):(1'h0)] wire3424;
  wire signed [(3'h5):(1'h0)] wire3431;
  wire [(5'h10):(1'h0)] wire3430;
  wire [(4'ha):(1'h0)] wire3429;
  wire [(4'he):(1'h0)] wire3428;
  assign y = {wire3431, wire3430, wire3429, wire3428, (1'h0)};
  assign wire3428 = ($unsigned(wire3426[(1'h1):(1'h0)]) || (({(8'hb4)} <<< $signed((8'hb3))) << wire3424));
  assign wire3429 = {wire3427};
  assign wire3430 = (~^{wire3429[(1'h0):(1'h0)]});
  assign wire3431 = wire3424[(4'ha):(1'h0)];
endmodule