(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param3107 = (((((8'ha3) == (8'had)) != ((8'ha2) > (8'ha7))) ? ({(8'ha9)} ? (+(8'hba)) : (|(8'ha7))) : (+((8'ha9) ? (8'hac) : (8'hb5)))) ? ((&((8'hb8) << (8'haf))) ~^ (~&(8'haf))) : ((((8'hae) ? (8'hba) : (8'hb1)) | {(8'h9c)}) ~^ {((8'hb9) ? (8'h9e) : (8'hae))})) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h5c3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire3;
  input wire [(4'ha):(1'h0)] wire2;
  input wire [(3'h5):(1'h0)] wire1;
  input wire [(4'he):(1'h0)] wire0;
  wire signed [(3'h5):(1'h0)] wire3105;
  wire signed [(4'ha):(1'h0)] wire144;
  wire [(4'hc):(1'h0)] wire143;
  wire [(3'h6):(1'h0)] wire142;
  wire [(4'hd):(1'h0)] wire141;
  wire signed [(4'he):(1'h0)] wire140;
  wire [(4'he):(1'h0)] wire139;
  reg signed [(4'hd):(1'h0)] reg94 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar84 = (1'h0);
  reg [(4'hf):(1'h0)] forvar76 = (1'h0);
  reg [(3'h6):(1'h0)] forvar70 = (1'h0);
  reg [(2'h2):(1'h0)] reg82 = (1'h0);
  reg [(2'h3):(1'h0)] forvar63 = (1'h0);
  reg [(3'h4):(1'h0)] forvar59 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg57 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg85 = (1'h0);
  reg [(3'h7):(1'h0)] reg138 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg136 = (1'h0);
  reg [(2'h3):(1'h0)] forvar135 = (1'h0);
  reg [(3'h4):(1'h0)] reg134 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg132 = (1'h0);
  reg [(4'ha):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar130 = (1'h0);
  reg [(2'h3):(1'h0)] reg129 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg128 = (1'h0);
  reg [(3'h6):(1'h0)] forvar127 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg125 = (1'h0);
  reg [(4'hc):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg123 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar122 = (1'h0);
  reg [(4'hd):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg119 = (1'h0);
  reg [(3'h5):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar117 = (1'h0);
  reg [(4'hf):(1'h0)] reg116 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg115 = (1'h0);
  reg [(4'hc):(1'h0)] reg114 = (1'h0);
  reg [(4'h8):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar112 = (1'h0);
  reg [(4'h9):(1'h0)] forvar111 = (1'h0);
  reg signed [(4'he):(1'h0)] reg110 = (1'h0);
  reg [(3'h5):(1'h0)] reg109 = (1'h0);
  reg [(4'hb):(1'h0)] reg108 = (1'h0);
  reg signed [(4'he):(1'h0)] reg107 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg106 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg105 = (1'h0);
  reg [(4'hc):(1'h0)] forvar104 = (1'h0);
  reg signed [(4'he):(1'h0)] reg103 = (1'h0);
  reg [(2'h3):(1'h0)] reg102 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar100 = (1'h0);
  reg [(5'h10):(1'h0)] forvar99 = (1'h0);
  reg [(2'h3):(1'h0)] reg98 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg97 = (1'h0);
  reg [(4'hd):(1'h0)] reg96 = (1'h0);
  reg [(4'ha):(1'h0)] reg95 = (1'h0);
  reg [(2'h2):(1'h0)] forvar94 = (1'h0);
  reg [(2'h2):(1'h0)] reg93 = (1'h0);
  reg [(3'h4):(1'h0)] reg92 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg91 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar90 = (1'h0);
  reg signed [(4'he):(1'h0)] reg89 = (1'h0);
  reg [(3'h6):(1'h0)] reg88 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg87 = (1'h0);
  reg [(3'h5):(1'h0)] forvar86 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar85 = (1'h0);
  reg [(5'h10):(1'h0)] reg84 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg83 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar82 = (1'h0);
  reg [(3'h6):(1'h0)] reg81 = (1'h0);
  reg [(2'h3):(1'h0)] reg80 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg79 = (1'h0);
  reg [(4'he):(1'h0)] reg78 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg77 = (1'h0);
  reg signed [(4'he):(1'h0)] reg76 = (1'h0);
  reg [(3'h5):(1'h0)] reg75 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar74 = (1'h0);
  reg [(4'hb):(1'h0)] forvar71 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg68 = (1'h0);
  reg [(2'h3):(1'h0)] forvar67 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar64 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg74 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg71 = (1'h0);
  reg [(2'h2):(1'h0)] reg70 = (1'h0);
  reg [(4'hd):(1'h0)] reg69 = (1'h0);
  reg [(4'h9):(1'h0)] forvar68 = (1'h0);
  reg [(2'h3):(1'h0)] reg67 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg65 = (1'h0);
  reg [(4'h9):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg62 = (1'h0);
  reg [(4'he):(1'h0)] reg61 = (1'h0);
  reg [(4'hd):(1'h0)] reg60 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg59 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar58 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar57 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar54 = (1'h0);
  reg [(2'h3):(1'h0)] reg53 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg52 = (1'h0);
  reg [(3'h6):(1'h0)] reg51 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar50 = (1'h0);
  reg [(4'hf):(1'h0)] reg49 = (1'h0);
  reg [(4'hb):(1'h0)] reg48 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg47 = (1'h0);
  reg [(4'h8):(1'h0)] reg46 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg38 = (1'h0);
  reg [(4'hb):(1'h0)] forvar37 = (1'h0);
  reg [(3'h6):(1'h0)] reg45 = (1'h0);
  reg [(4'h9):(1'h0)] reg44 = (1'h0);
  reg [(2'h3):(1'h0)] reg43 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar42 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg41 = (1'h0);
  reg [(4'hb):(1'h0)] reg40 = (1'h0);
  reg [(4'ha):(1'h0)] reg39 = (1'h0);
  reg [(3'h5):(1'h0)] forvar38 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg37 = (1'h0);
  reg [(4'h8):(1'h0)] reg36 = (1'h0);
  reg [(4'hd):(1'h0)] forvar35 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar34 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg33 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg32 = (1'h0);
  reg [(2'h2):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg30 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar29 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg28 = (1'h0);
  reg [(4'hf):(1'h0)] reg27 = (1'h0);
  reg [(4'hf):(1'h0)] forvar26 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar25 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar11 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar8 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4 = (1'h0);
  reg [(3'h7):(1'h0)] reg24 = (1'h0);
  reg [(3'h5):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar22 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg22 = (1'h0);
  reg [(3'h7):(1'h0)] reg21 = (1'h0);
  reg [(4'hd):(1'h0)] forvar20 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg19 = (1'h0);
  reg [(2'h3):(1'h0)] forvar18 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar15 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar10 = (1'h0);
  reg [(2'h3):(1'h0)] forvar9 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7 = (1'h0);
  reg [(2'h2):(1'h0)] reg6 = (1'h0);
  reg [(4'ha):(1'h0)] reg17 = (1'h0);
  reg [(2'h3):(1'h0)] reg14 = (1'h0);
  reg [(4'hc):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg15 = (1'h0);
  reg [(4'h9):(1'h0)] forvar14 = (1'h0);
  reg [(3'h4):(1'h0)] reg13 = (1'h0);
  reg [(5'h10):(1'h0)] reg12 = (1'h0);
  reg [(5'h10):(1'h0)] reg11 = (1'h0);
  reg [(5'h10):(1'h0)] reg10 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg9 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg8 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6 = (1'h0);
  reg [(5'h10):(1'h0)] reg5 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4 = (1'h0);
  assign y = {wire3105,
                 wire144,
                 wire143,
                 wire142,
                 wire141,
                 wire140,
                 wire139,
                 reg94,
                 reg90,
                 forvar84,
                 forvar76,
                 forvar70,
                 reg82,
                 forvar63,
                 forvar59,
                 reg57,
                 reg85,
                 reg138,
                 reg137,
                 reg136,
                 forvar135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 forvar130,
                 reg129,
                 reg128,
                 forvar127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 forvar122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 forvar117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 forvar112,
                 forvar111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg105,
                 forvar104,
                 reg103,
                 reg102,
                 reg101,
                 forvar100,
                 forvar99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 forvar94,
                 reg93,
                 reg92,
                 reg91,
                 forvar90,
                 reg89,
                 reg88,
                 reg87,
                 forvar86,
                 forvar85,
                 reg84,
                 reg83,
                 forvar82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 forvar74,
                 forvar71,
                 reg68,
                 forvar67,
                 forvar64,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 forvar68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 forvar58,
                 forvar57,
                 reg56,
                 reg55,
                 forvar54,
                 reg53,
                 reg52,
                 reg51,
                 forvar50,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg38,
                 forvar37,
                 reg45,
                 reg44,
                 reg43,
                 forvar42,
                 reg41,
                 reg40,
                 reg39,
                 forvar38,
                 reg37,
                 reg36,
                 forvar35,
                 forvar34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 forvar29,
                 reg28,
                 reg27,
                 forvar26,
                 forvar25,
                 forvar11,
                 forvar8,
                 forvar5,
                 reg4,
                 reg24,
                 reg23,
                 forvar22,
                 reg22,
                 reg21,
                 forvar20,
                 reg19,
                 forvar18,
                 forvar15,
                 forvar10,
                 forvar9,
                 reg7,
                 reg6,
                 reg17,
                 reg14,
                 reg16,
                 reg15,
                 forvar14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar7,
                 forvar6,
                 reg5,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((wire0 <= $unsigned($signed($signed(wire1)))))
        begin
          for (forvar4 = (1'h0); (forvar4 < (1'h0)); forvar4 = (forvar4 + (1'h1)))
            begin
              reg5 <= $unsigned((wire2 ?
                  wire3[(2'h3):(2'h3)] : {(wire3 ? (8'ha7) : (8'ha2))}));
              for (forvar6 = (1'h0); (forvar6 < (1'h0)); forvar6 = (forvar6 + (1'h1)))
                begin
                  for (forvar7 = (1'h0); (forvar7 < (1'h0)); forvar7 = (forvar7 + (1'h1)))
                    begin
                      reg8 <= $unsigned(wire3[(1'h1):(1'h0)]);
                      reg9 <= ($signed(wire0[(4'hd):(4'hb)]) ?
                          ((~|wire2[(2'h3):(1'h0)]) >> wire1[(3'h5):(3'h5)]) : $signed(wire3));
                      reg10 <= (wire1[(2'h3):(1'h1)] << (8'hb2));
                    end
                  if ($unsigned($signed($unsigned((wire0 ? forvar4 : reg5)))))
                    begin
                      reg11 <= $unsigned($signed(wire2));
                      reg12 <= $signed(reg8[(2'h2):(1'h0)]);
                      reg13 <= (~|($signed((wire1 ^ reg10)) ?
                          (~forvar4) : {wire3}));
                    end
                  else
                    begin
                      reg11 <= (^$unsigned({(reg13 <<< (8'hb2))}));
                      reg12 <= reg10;
                      reg13 <= wire3;
                    end
                end
              if ((!({(reg12 ? forvar7 : reg11)} == ((8'ha9) ?
                  (reg9 ? wire2 : reg13) : (wire0 ? reg5 : reg10)))))
                begin
                  for (forvar14 = (1'h0); (forvar14 < (2'h3)); forvar14 = (forvar14 + (1'h1)))
                    begin
                      reg15 <= (&reg9[(4'h8):(2'h2)]);
                      reg16 <= {($signed($unsigned(reg12)) ?
                              $unsigned($signed(forvar7)) : (~&{reg8}))};
                    end
                end
              else
                begin
                  if ((wire2 & $signed(reg12)))
                    begin
                      reg14 <= forvar14;
                    end
                  else
                    begin
                      reg14 <= $unsigned(reg11[(1'h1):(1'h0)]);
                      reg15 <= ((+($signed(reg13) ^~ $unsigned((8'hb3)))) >>> ((~$signed(reg9)) ^ (8'ha1)));
                    end
                end
            end
          reg17 <= ($signed($unsigned($signed(reg14))) ? wire1 : reg5);
        end
      else
        begin
          if ($unsigned(((((8'hb8) || reg8) | (+reg13)) >> reg10[(4'h9):(2'h2)])))
            begin
              if ((^~$unsigned(((reg9 ?
                  (8'ha4) : forvar14) >> ((8'h9c) - reg9)))))
                begin
                  for (forvar4 = (1'h0); (forvar4 < (2'h2)); forvar4 = (forvar4 + (1'h1)))
                    begin
                      reg5 <= $signed((wire2 >= forvar7));
                    end
                end
              else
                begin
                  for (forvar4 = (1'h0); (forvar4 < (1'h1)); forvar4 = (forvar4 + (1'h1)))
                    begin
                      reg5 <= (+reg16[(4'h9):(3'h7)]);
                      reg6 <= (~|($unsigned((+reg17)) >= (reg8[(2'h2):(2'h2)] ?
                          (+reg13) : (wire1 <<< (8'h9d)))));
                      reg7 <= forvar7;
                      reg8 <= $signed((8'hb2));
                    end
                end
              for (forvar9 = (1'h0); (forvar9 < (2'h2)); forvar9 = (forvar9 + (1'h1)))
                begin
                  for (forvar10 = (1'h0); (forvar10 < (1'h1)); forvar10 = (forvar10 + (1'h1)))
                    begin
                      reg11 <= ($signed($unsigned((+reg5))) != {(^reg14)});
                      reg12 <= reg16;
                      reg13 <= $unsigned({({reg16} | (reg9 ?
                              reg9 : forvar10))});
                    end
                  reg14 <= ((+((forvar6 ? (8'h9f) : forvar9) ?
                          $signed(forvar4) : reg6[(1'h0):(1'h0)])) ?
                      $signed({$unsigned(reg17)}) : (($signed(forvar7) ?
                              (-wire1) : (forvar10 < forvar10)) ?
                          reg17 : ({(8'hb5)} ? {forvar14} : (+(8'hb3)))));
                  for (forvar15 = (1'h0); (forvar15 < (1'h0)); forvar15 = (forvar15 + (1'h1)))
                    begin
                      reg16 <= reg11;
                      reg17 <= $unsigned($unsigned(((^~(8'hb7)) || reg14[(2'h3):(2'h2)])));
                    end
                  for (forvar18 = (1'h0); (forvar18 < (1'h1)); forvar18 = (forvar18 + (1'h1)))
                    begin
                      reg19 <= ($signed($signed($unsigned(reg5))) && (reg11[(4'hd):(4'hd)] != {forvar9[(1'h1):(1'h1)]}));
                    end
                end
              for (forvar20 = (1'h0); (forvar20 < (1'h1)); forvar20 = (forvar20 + (1'h1)))
                begin
                  reg21 <= reg17;
                end
              if ({((forvar6 == (~&reg17)) == (^~{wire2}))})
                begin
                  reg22 <= (|$signed(reg15[(4'hb):(3'h4)]));
                end
              else
                begin
                  for (forvar22 = (1'h0); (forvar22 < (1'h1)); forvar22 = (forvar22 + (1'h1)))
                    begin
                      reg23 <= (reg5 ? reg11 : reg19[(1'h1):(1'h0)]);
                      reg24 <= (|reg19);
                    end
                end
            end
          else
            begin
              if (reg24)
                begin
                  reg4 <= ($unsigned($unsigned($unsigned(reg7))) && $unsigned(($unsigned(reg17) - $signed(reg24))));
                  for (forvar5 = (1'h0); (forvar5 < (2'h3)); forvar5 = (forvar5 + (1'h1)))
                    begin
                      reg6 <= (&{reg19});
                      reg7 <= reg19[(2'h3):(2'h2)];
                      reg8 <= (~^$signed(reg14));
                      reg9 <= $signed(forvar4);
                    end
                end
              else
                begin
                  reg4 <= reg8[(1'h1):(1'h1)];
                  reg5 <= forvar7[(4'h9):(2'h2)];
                  for (forvar6 = (1'h0); (forvar6 < (2'h3)); forvar6 = (forvar6 + (1'h1)))
                    begin
                      reg7 <= (^forvar7[(2'h3):(1'h1)]);
                    end
                  for (forvar8 = (1'h0); (forvar8 < (1'h1)); forvar8 = (forvar8 + (1'h1)))
                    begin
                      reg9 <= (~(8'h9f));
                    end
                end
              if ($signed((^~{$signed((8'ha5))})))
                begin
                  for (forvar10 = (1'h0); (forvar10 < (2'h2)); forvar10 = (forvar10 + (1'h1)))
                    begin
                      reg11 <= (8'hb9);
                    end
                end
              else
                begin
                  if (forvar18)
                    begin
                      reg10 <= forvar14;
                    end
                  else
                    begin
                      reg10 <= $signed(forvar18[(2'h2):(1'h0)]);
                    end
                  for (forvar11 = (1'h0); (forvar11 < (1'h1)); forvar11 = (forvar11 + (1'h1)))
                    begin
                      reg12 <= ($unsigned($signed((reg11 ? (8'hb7) : reg17))) ?
                          forvar10[(1'h0):(1'h0)] : forvar10[(2'h3):(2'h3)]);
                      reg13 <= $signed({(^forvar15)});
                      reg14 <= $unsigned($unsigned($signed(reg17[(3'h4):(2'h3)])));
                      reg15 <= $unsigned($signed($unsigned((wire2 ?
                          reg22 : (8'ha4)))));
                    end
                end
            end
          for (forvar25 = (1'h0); (forvar25 < (1'h0)); forvar25 = (forvar25 + (1'h1)))
            begin
              for (forvar26 = (1'h0); (forvar26 < (2'h2)); forvar26 = (forvar26 + (1'h1)))
                begin
                  if (reg5)
                    begin
                      reg27 <= (({$unsigned(reg24)} ?
                          forvar25[(2'h3):(1'h0)] : (reg9[(4'hc):(2'h2)] ?
                              (forvar25 * reg7) : wire3[(3'h6):(2'h2)])) & (&$signed((forvar26 ?
                          (8'hb3) : wire2))));
                      reg28 <= (8'hb1);
                    end
                  else
                    begin
                      reg27 <= reg27[(4'hd):(2'h2)];
                      reg28 <= reg19[(4'hf):(3'h6)];
                    end
                end
              for (forvar29 = (1'h0); (forvar29 < (2'h3)); forvar29 = (forvar29 + (1'h1)))
                begin
                  if ((~forvar25[(4'h9):(3'h6)]))
                    begin
                      reg30 <= $unsigned(reg19);
                      reg31 <= $signed(forvar18);
                      reg32 <= reg11;
                      reg33 <= $signed($unsigned(($unsigned(reg27) && reg21[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg30 <= (^~(+reg17[(4'h9):(3'h4)]));
                    end
                end
            end
          if ((((~|(~&reg22)) ?
                  ({forvar26} ~^ (-reg9)) : ($signed((8'ha1)) ?
                      $signed((8'hb4)) : wire0)) ?
              {$signed((forvar25 || reg17))} : {($signed(reg32) ^~ forvar26)}))
            begin
              for (forvar34 = (1'h0); (forvar34 < (2'h2)); forvar34 = (forvar34 + (1'h1)))
                begin
                  for (forvar35 = (1'h0); (forvar35 < (1'h1)); forvar35 = (forvar35 + (1'h1)))
                    begin
                      reg36 <= forvar22;
                      reg37 <= $unsigned($unsigned(($signed(reg21) < (8'h9c))));
                    end
                  for (forvar38 = (1'h0); (forvar38 < (2'h3)); forvar38 = (forvar38 + (1'h1)))
                    begin
                      reg39 <= reg10[(3'h5):(3'h5)];
                      reg40 <= (&((~^(reg33 > reg7)) ?
                          $signed((-reg30)) : reg30));
                      reg41 <= reg31[(2'h2):(2'h2)];
                    end
                  for (forvar42 = (1'h0); (forvar42 < (2'h2)); forvar42 = (forvar42 + (1'h1)))
                    begin
                      reg43 <= $unsigned(reg37[(3'h5):(2'h2)]);
                      reg44 <= $unsigned((($signed((8'hb6)) > $unsigned(reg41)) ~^ (+(reg27 > (8'h9f)))));
                    end
                  reg45 <= ({(forvar29[(1'h1):(1'h1)] && reg37[(2'h2):(1'h0)])} ?
                      $signed((reg41[(3'h4):(3'h4)] != $unsigned(forvar10))) : $unsigned(((reg13 ?
                              reg31 : reg32) ?
                          $unsigned(forvar26) : (8'hb5))));
                end
            end
          else
            begin
              for (forvar34 = (1'h0); (forvar34 < (1'h1)); forvar34 = (forvar34 + (1'h1)))
                begin
                  for (forvar35 = (1'h0); (forvar35 < (1'h1)); forvar35 = (forvar35 + (1'h1)))
                    begin
                      reg36 <= ($unsigned($unsigned(reg6)) ?
                          (wire2 >> reg12) : $signed(((reg30 ?
                                  (8'hb0) : forvar5) ?
                              $unsigned(forvar29) : {(8'ha9)})));
                    end
                  for (forvar37 = (1'h0); (forvar37 < (1'h1)); forvar37 = (forvar37 + (1'h1)))
                    begin
                      reg38 <= {(forvar34 ^~ ({reg9} ?
                              $signed(reg17) : {reg23}))};
                      reg39 <= $signed($unsigned($unsigned($unsigned(reg41))));
                      reg40 <= ((({reg31} ~^ (reg27 <<< reg4)) || ($signed((8'hb8)) ?
                              (+(8'haa)) : (!reg22))) ?
                          (8'hb7) : ($signed((wire3 - reg9)) + reg21[(3'h6):(3'h6)]));
                      reg41 <= {forvar34};
                    end
                end
              for (forvar42 = (1'h0); (forvar42 < (1'h1)); forvar42 = (forvar42 + (1'h1)))
                begin
                  if ($signed((^reg30[(2'h3):(1'h0)])))
                    begin
                      reg43 <= ($unsigned((+(forvar15 ?
                          (8'ha8) : forvar6))) >>> ((reg45[(3'h6):(1'h1)] * (reg19 ^ (8'haa))) == ((-reg31) ?
                          {reg11} : (^(8'ha7)))));
                    end
                  else
                    begin
                      reg43 <= ((~{(reg39 > reg14)}) ?
                          reg10 : reg13[(1'h1):(1'h1)]);
                      reg44 <= $unsigned(((reg12[(2'h2):(2'h2)] != $unsigned(reg23)) > $unsigned((reg14 & wire2))));
                      reg45 <= $unsigned({(forvar18 ?
                              (forvar10 ?
                                  reg32 : reg27) : reg30[(4'h8):(3'h5)])});
                    end
                  if (forvar8)
                    begin
                      reg46 <= $unsigned($signed((+forvar6[(1'h1):(1'h1)])));
                      reg47 <= {forvar35[(4'hb):(3'h4)]};
                      reg48 <= forvar42;
                    end
                  else
                    begin
                      reg46 <= $signed(wire1);
                      reg47 <= forvar14[(4'h8):(2'h3)];
                      reg48 <= ($signed($unsigned((8'hb7))) ?
                          forvar18[(2'h3):(1'h1)] : reg38[(3'h5):(1'h0)]);
                      reg49 <= ({$unsigned((!forvar34))} ?
                          forvar10[(1'h1):(1'h1)] : $unsigned(((reg38 && forvar20) >>> $signed(reg6))));
                    end
                end
              for (forvar50 = (1'h0); (forvar50 < (2'h3)); forvar50 = (forvar50 + (1'h1)))
                begin
                  if ($unsigned($signed(reg23[(3'h4):(3'h4)])))
                    begin
                      reg51 <= forvar37;
                      reg52 <= $signed(reg39);
                    end
                  else
                    begin
                      reg51 <= reg16;
                      reg52 <= (({reg36} ?
                              ({reg22} ?
                                  reg15[(3'h4):(1'h0)] : $unsigned(reg5)) : reg46[(3'h5):(3'h5)]) ?
                          $signed($unsigned((forvar18 ?
                              forvar18 : reg43))) : $signed(reg32));
                      reg53 <= (|$unsigned((forvar42[(3'h6):(3'h5)] | (reg46 >= reg15))));
                    end
                end
              if (($unsigned($signed(reg16)) < $unsigned({$signed((8'hab))})))
                begin
                  for (forvar54 = (1'h0); (forvar54 < (2'h2)); forvar54 = (forvar54 + (1'h1)))
                    begin
                      reg55 <= $unsigned(($unsigned(reg36) ?
                          (|reg36) : (forvar5 ?
                              $signed(reg21) : forvar18[(2'h3):(2'h3)])));
                      reg56 <= forvar42[(4'h9):(4'h8)];
                    end
                end
              else
                begin
                  for (forvar54 = (1'h0); (forvar54 < (2'h2)); forvar54 = (forvar54 + (1'h1)))
                    begin
                      reg55 <= (forvar42 >= $signed({$signed((8'hb7))}));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ((+$signed(reg46)))
        begin
          if (((~^{$signed(forvar35)}) - {((reg53 ? reg13 : (8'hae)) ?
                  (!wire2) : forvar8)}))
            begin
              for (forvar57 = (1'h0); (forvar57 < (2'h3)); forvar57 = (forvar57 + (1'h1)))
                begin
                  for (forvar58 = (1'h0); (forvar58 < (2'h3)); forvar58 = (forvar58 + (1'h1)))
                    begin
                      reg59 <= reg28;
                      reg60 <= ({reg33} ?
                          $signed((forvar9[(2'h2):(1'h0)] << (reg46 ?
                              reg22 : reg9))) : $signed($signed((reg12 && forvar35))));
                    end
                  if ((8'haf))
                    begin
                      reg61 <= forvar34;
                    end
                  else
                    begin
                      reg61 <= {((~$unsigned(reg36)) ?
                              {(8'had)} : reg28[(1'h0):(1'h0)])};
                      reg62 <= (|reg59);
                    end
                  reg63 <= {{((reg12 ? forvar6 : reg46) ?
                              (8'hb5) : (reg36 ^ reg4))}};
                end
              if (forvar22)
                begin
                  if ($signed(forvar54[(4'hd):(2'h2)]))
                    begin
                      reg64 <= reg37[(2'h3):(1'h0)];
                      reg65 <= (~|(8'ha9));
                    end
                  else
                    begin
                      reg64 <= forvar37;
                      reg65 <= {reg44};
                      reg66 <= ($unsigned($unsigned(reg40)) ^~ (forvar20[(4'hd):(4'hd)] ?
                          (forvar10[(2'h2):(1'h1)] ?
                              $signed(reg12) : (reg16 || reg55)) : ((reg27 ?
                                  reg7 : forvar4) ?
                              reg63[(1'h0):(1'h0)] : $signed(forvar18))));
                      reg67 <= (^(^$signed((reg32 ~^ forvar22))));
                    end
                  for (forvar68 = (1'h0); (forvar68 < (2'h3)); forvar68 = (forvar68 + (1'h1)))
                    begin
                      reg69 <= reg16[(3'h7):(2'h3)];
                      reg70 <= (~|reg21[(1'h0):(1'h0)]);
                      reg71 <= $unsigned($unsigned($signed(forvar42[(2'h2):(1'h1)])));
                      reg72 <= forvar34;
                    end
                  if ($unsigned((!forvar8[(1'h0):(1'h0)])))
                    begin
                      reg73 <= $signed(reg28);
                      reg74 <= reg24[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg73 <= reg67[(2'h2):(1'h0)];
                    end
                end
              else
                begin
                  if ((~^forvar34[(3'h6):(3'h5)]))
                    begin
                      reg64 <= (^($unsigned(reg62[(3'h6):(3'h5)]) >>> (forvar35 << $unsigned((8'h9f)))));
                      reg65 <= $unsigned(reg66[(3'h4):(1'h0)]);
                      reg66 <= forvar20[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg64 <= forvar34[(3'h6):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar57 = (1'h0); (forvar57 < (1'h0)); forvar57 = (forvar57 + (1'h1)))
                begin
                  for (forvar58 = (1'h0); (forvar58 < (2'h3)); forvar58 = (forvar58 + (1'h1)))
                    begin
                      reg59 <= $unsigned($signed($unsigned(((8'ha9) ?
                          (8'hb0) : reg62))));
                      reg60 <= (forvar6[(1'h0):(1'h0)] ?
                          (^(-$signed(forvar14))) : forvar25[(3'h7):(2'h2)]);
                      reg61 <= (8'h9e);
                      reg62 <= reg36;
                    end
                  reg63 <= ((&forvar8) ? (-(^~wire3)) : reg11);
                end
              if (reg38[(2'h3):(1'h0)])
                begin
                  for (forvar64 = (1'h0); (forvar64 < (2'h3)); forvar64 = (forvar64 + (1'h1)))
                    begin
                      reg65 <= {((forvar10[(1'h0):(1'h0)] ?
                                  $unsigned(reg37) : (&forvar20)) ?
                              (((8'h9c) ^ (8'h9f)) ?
                                  (reg12 ?
                                      reg19 : reg15) : (8'h9d)) : forvar9)};
                      reg66 <= ($unsigned(reg73) ?
                          $unsigned(((reg41 & reg48) >= {reg36})) : {$signed({(8'haa)})});
                    end
                  for (forvar67 = (1'h0); (forvar67 < (1'h1)); forvar67 = (forvar67 + (1'h1)))
                    begin
                      reg68 <= $signed(reg66[(2'h2):(1'h1)]);
                      reg69 <= (8'ha2);
                      reg70 <= $unsigned(($signed(forvar5[(1'h0):(1'h0)]) * ((reg9 ~^ (8'haf)) ^~ ((8'hb1) ?
                          reg71 : reg14))));
                    end
                end
              else
                begin
                  for (forvar64 = (1'h0); (forvar64 < (2'h3)); forvar64 = (forvar64 + (1'h1)))
                    begin
                      reg65 <= reg47[(3'h6):(1'h1)];
                      reg66 <= (8'ha2);
                    end
                end
              if (forvar50[(3'h4):(2'h2)])
                begin
                  for (forvar71 = (1'h0); (forvar71 < (2'h3)); forvar71 = (forvar71 + (1'h1)))
                    begin
                      reg72 <= ($unsigned(reg46[(1'h1):(1'h1)]) ^~ $signed((reg10 <= (8'hb3))));
                      reg73 <= (+$unsigned(($signed(reg10) ~^ (forvar15 <= forvar71))));
                    end
                  for (forvar74 = (1'h0); (forvar74 < (2'h2)); forvar74 = (forvar74 + (1'h1)))
                    begin
                      reg75 <= ($signed(((~|reg30) + $signed(forvar67))) < reg22[(1'h0):(1'h0)]);
                      reg76 <= $unsigned(($signed((reg48 ? (8'hb7) : reg31)) ?
                          forvar42[(4'h8):(2'h3)] : {$unsigned(forvar7)}));
                      reg77 <= ((reg19 ?
                              ((reg6 ? reg62 : forvar11) ?
                                  (reg46 <<< forvar11) : (8'hb0)) : (8'hab)) ?
                          $signed((!(reg65 ? forvar9 : reg14))) : (~reg69));
                      reg78 <= $unsigned((forvar64 & {$unsigned(reg62)}));
                    end
                  if (({reg75} + (reg30[(3'h4):(3'h4)] < $unsigned(reg70[(2'h2):(2'h2)]))))
                    begin
                      reg79 <= forvar35[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg79 <= (($signed((forvar5 && forvar26)) && $unsigned($unsigned(reg33))) ?
                          reg73 : (^((forvar18 && wire0) || reg77)));
                      reg80 <= $unsigned((|((&(8'h9d)) < $signed(forvar38))));
                      reg81 <= $unsigned((((reg11 * (8'haa)) + (reg28 ?
                              reg30 : forvar22)) ?
                          forvar18[(1'h1):(1'h1)] : forvar34[(4'h8):(1'h0)]));
                    end
                end
              else
                begin
                  if ((($signed($signed(forvar74)) ?
                      $unsigned((!(8'hae))) : $signed($signed(reg9))) >= (!{$signed(reg44)})))
                    begin
                      reg71 <= (-(^~((|forvar4) ?
                          {forvar50} : (forvar26 >>> reg36))));
                    end
                  else
                    begin
                      reg71 <= forvar10;
                      reg72 <= ({(-$signed(forvar8))} ?
                          ((~|$signed(forvar8)) <= $unsigned(reg44)) : $signed(($signed(reg48) ?
                              (~(8'ha8)) : reg48)));
                    end
                  reg73 <= ((forvar15[(4'hd):(1'h1)] ?
                          ((forvar18 > reg79) ?
                              (wire3 ?
                                  reg9 : (8'hb8)) : $unsigned(reg24)) : $unsigned((reg16 <<< (8'hb7)))) ?
                      $signed(reg17) : $unsigned(reg43[(1'h0):(1'h0)]));
                end
              for (forvar82 = (1'h0); (forvar82 < (2'h2)); forvar82 = (forvar82 + (1'h1)))
                begin
                  reg83 <= (reg6[(1'h1):(1'h1)] ?
                      (!{(reg45 ? (8'ha0) : reg47)}) : $signed((&(^reg63))));
                  reg84 <= ($signed($unsigned((+reg15))) >>> ((reg7[(2'h3):(2'h2)] ?
                      $unsigned((8'hb7)) : reg63) == $unsigned($unsigned(reg8))));
                end
            end
          if ({reg70})
            begin
              for (forvar85 = (1'h0); (forvar85 < (1'h1)); forvar85 = (forvar85 + (1'h1)))
                begin
                  for (forvar86 = (1'h0); (forvar86 < (2'h3)); forvar86 = (forvar86 + (1'h1)))
                    begin
                      reg87 <= forvar15;
                      reg88 <= $unsigned($unsigned($signed((~^reg87))));
                      reg89 <= reg48;
                    end
                  for (forvar90 = (1'h0); (forvar90 < (2'h3)); forvar90 = (forvar90 + (1'h1)))
                    begin
                      reg91 <= ((&forvar37) ~^ $unsigned(wire2[(1'h1):(1'h1)]));
                      reg92 <= reg88[(3'h4):(1'h0)];
                      reg93 <= (~^$signed((8'h9e)));
                    end
                  for (forvar94 = (1'h0); (forvar94 < (2'h3)); forvar94 = (forvar94 + (1'h1)))
                    begin
                      reg95 <= (|{(reg84[(4'h9):(4'h8)] ?
                              (reg10 ? reg55 : reg59) : (reg15 == reg93))});
                      reg96 <= forvar22[(4'ha):(3'h4)];
                    end
                  if (((reg53 >= reg27[(4'hf):(3'h7)]) ?
                      reg89 : forvar37[(3'h7):(2'h3)]))
                    begin
                      reg97 <= forvar26;
                    end
                  else
                    begin
                      reg97 <= {$signed(($signed(reg67) ?
                              ((8'hb6) != reg38) : (wire3 * forvar14)))};
                      reg98 <= ((forvar10 ?
                          $signed((~&forvar64)) : forvar94) >>> (&($unsigned(wire0) ?
                          {forvar18} : $signed(reg15))));
                    end
                end
              for (forvar99 = (1'h0); (forvar99 < (2'h2)); forvar99 = (forvar99 + (1'h1)))
                begin
                  for (forvar100 = (1'h0); (forvar100 < (2'h3)); forvar100 = (forvar100 + (1'h1)))
                    begin
                      reg101 <= {(~$signed($signed(reg77)))};
                      reg102 <= reg24;
                      reg103 <= (8'haa);
                    end
                  for (forvar104 = (1'h0); (forvar104 < (2'h3)); forvar104 = (forvar104 + (1'h1)))
                    begin
                      reg105 <= $unsigned(forvar8[(3'h4):(2'h3)]);
                      reg106 <= {{(reg59[(1'h1):(1'h0)] ?
                                  (wire3 ^~ reg76) : (reg10 << forvar100))}};
                      reg107 <= forvar90[(1'h1):(1'h1)];
                      reg108 <= ((~((reg88 ? forvar64 : reg96) ?
                              (forvar8 ? reg68 : reg76) : forvar15)) ?
                          ({(~&(8'hb9))} != forvar4[(1'h1):(1'h1)]) : (($signed(forvar29) > reg27[(4'h9):(1'h0)]) >> $signed((~reg61))));
                    end
                  if ({reg36[(3'h6):(1'h1)]})
                    begin
                      reg109 <= $signed({(reg45[(2'h2):(1'h0)] ?
                              $unsigned(forvar8) : (forvar11 ?
                                  reg103 : reg55))});
                    end
                  else
                    begin
                      reg109 <= (~$signed(reg8[(2'h3):(2'h2)]));
                      reg110 <= forvar58[(3'h4):(3'h4)];
                    end
                end
              for (forvar111 = (1'h0); (forvar111 < (2'h3)); forvar111 = (forvar111 + (1'h1)))
                begin
                  for (forvar112 = (1'h0); (forvar112 < (1'h0)); forvar112 = (forvar112 + (1'h1)))
                    begin
                      reg113 <= {reg67};
                      reg114 <= ((~|reg65) ?
                          (reg19 ?
                              ($signed((8'h9f)) * $signed(forvar29)) : forvar8) : $signed(forvar22[(1'h0):(1'h0)]));
                      reg115 <= (reg83 ?
                          forvar94[(2'h2):(1'h1)] : reg55[(1'h1):(1'h1)]);
                      reg116 <= ((~^reg43) == $signed($signed(reg63[(2'h2):(1'h1)])));
                    end
                  for (forvar117 = (1'h0); (forvar117 < (1'h0)); forvar117 = (forvar117 + (1'h1)))
                    begin
                      reg118 <= (({(reg109 ? reg63 : reg110)} ?
                          reg31[(2'h2):(1'h1)] : (reg41 | reg89)) ~^ reg38[(2'h3):(1'h1)]);
                      reg119 <= $unsigned($unsigned(reg15[(4'hc):(3'h7)]));
                      reg120 <= ($unsigned(reg13) ?
                          {reg13} : reg93[(1'h1):(1'h1)]);
                      reg121 <= forvar71;
                    end
                end
              for (forvar122 = (1'h0); (forvar122 < (1'h1)); forvar122 = (forvar122 + (1'h1)))
                begin
                  if (forvar54[(4'h9):(4'h8)])
                    begin
                      reg123 <= reg4;
                      reg124 <= (+{(forvar58[(4'h9):(4'h8)] | ((8'hb4) ~^ reg38))});
                      reg125 <= $unsigned({reg23[(2'h2):(1'h0)]});
                      reg126 <= {$signed(reg32)};
                    end
                  else
                    begin
                      reg123 <= reg27;
                      reg124 <= {{reg19}};
                      reg125 <= reg12;
                    end
                  for (forvar127 = (1'h0); (forvar127 < (1'h1)); forvar127 = (forvar127 + (1'h1)))
                    begin
                      reg128 <= reg11;
                      reg129 <= $signed((reg5[(4'h9):(3'h4)] > $signed($unsigned(reg45))));
                    end
                  for (forvar130 = (1'h0); (forvar130 < (2'h2)); forvar130 = (forvar130 + (1'h1)))
                    begin
                      reg131 <= ((^~$signed((|reg75))) == $signed((8'ha3)));
                      reg132 <= reg91[(1'h0):(1'h0)];
                      reg133 <= ($unsigned((((8'h9c) ?
                          reg30 : reg6) | (8'hb0))) * (($unsigned(reg89) ^ (forvar14 ?
                          reg76 : forvar90)) <= forvar99[(4'hc):(4'h9)]));
                      reg134 <= reg30;
                    end
                  for (forvar135 = (1'h0); (forvar135 < (2'h3)); forvar135 = (forvar135 + (1'h1)))
                    begin
                      reg136 <= (!wire3);
                      reg137 <= (8'hac);
                      reg138 <= $unsigned({$unsigned((|reg52))});
                    end
                end
            end
          else
            begin
              reg85 <= ({forvar29[(3'h4):(2'h3)]} != (reg15[(4'hd):(4'hb)] ?
                  reg81[(1'h0):(1'h0)] : reg47));
            end
        end
      else
        begin
          reg57 <= {({(8'h9e)} ^ $signed((8'ha7)))};
          for (forvar58 = (1'h0); (forvar58 < (1'h1)); forvar58 = (forvar58 + (1'h1)))
            begin
              for (forvar59 = (1'h0); (forvar59 < (2'h3)); forvar59 = (forvar59 + (1'h1)))
                begin
                  reg60 <= ((~&((wire0 ? reg57 : (8'hb1)) ?
                      reg13 : reg15[(4'h9):(3'h4)])) | reg22);
                  if (forvar42[(3'h4):(1'h1)])
                    begin
                      reg61 <= (8'h9e);
                    end
                  else
                    begin
                      reg61 <= $unsigned(reg59);
                      reg62 <= {$unsigned($signed((^reg66)))};
                    end
                  for (forvar63 = (1'h0); (forvar63 < (1'h1)); forvar63 = (forvar63 + (1'h1)))
                    begin
                      reg64 <= (8'h9c);
                      reg65 <= $signed($unsigned($signed((reg41 ?
                          reg79 : reg88))));
                      reg66 <= ($unsigned($signed(reg63)) ?
                          $unsigned($unsigned($signed(reg71))) : forvar37);
                    end
                  for (forvar67 = (1'h0); (forvar67 < (2'h2)); forvar67 = (forvar67 + (1'h1)))
                    begin
                      reg68 <= (&$unsigned(reg15[(2'h3):(1'h1)]));
                      reg69 <= $signed($signed((~^(wire2 ? reg4 : reg67))));
                    end
                end
              if ($signed((reg53[(2'h3):(2'h2)] ?
                  reg116[(3'h7):(2'h2)] : {reg16[(3'h7):(3'h6)]})))
                begin
                  if (($signed(wire0) << ($unsigned(reg5) >= ($unsigned(reg27) << reg137))))
                    begin
                      reg70 <= reg98[(1'h1):(1'h0)];
                      reg71 <= $unsigned(wire1);
                    end
                  else
                    begin
                      reg70 <= reg106;
                      reg71 <= reg70[(1'h1):(1'h1)];
                      reg72 <= reg63[(3'h5):(1'h1)];
                      reg73 <= forvar127;
                    end
                  for (forvar74 = (1'h0); (forvar74 < (2'h2)); forvar74 = (forvar74 + (1'h1)))
                    begin
                      reg75 <= {reg57};
                      reg76 <= forvar7;
                    end
                  if ((&$unsigned(((~(8'hb0)) ~^ $unsigned(reg78)))))
                    begin
                      reg77 <= reg118[(3'h4):(3'h4)];
                      reg78 <= reg132[(3'h5):(2'h3)];
                      reg79 <= (($signed(reg46) ?
                          $signed((~^(8'h9e))) : reg27) || ($unsigned((reg75 ?
                              reg4 : reg48)) ?
                          wire3[(1'h0):(1'h0)] : (~reg118[(2'h3):(1'h1)])));
                    end
                  else
                    begin
                      reg77 <= forvar54;
                      reg78 <= reg126;
                      reg79 <= ((reg14 ?
                          $unsigned($unsigned(reg44)) : $unsigned((8'h9c))) != $unsigned($unsigned((reg11 ?
                          reg114 : reg85))));
                      reg80 <= $signed((~^$unsigned(reg118[(3'h4):(2'h3)])));
                    end
                  if (reg69)
                    begin
                      reg81 <= (reg103[(3'h6):(3'h4)] - reg97);
                    end
                  else
                    begin
                      reg81 <= $unsigned((reg16[(2'h2):(1'h0)] ?
                          $signed(((8'h9d) * reg115)) : (!$unsigned(forvar34))));
                      reg82 <= forvar58[(4'ha):(3'h6)];
                      reg83 <= ($unsigned((8'haa)) & (((forvar99 ?
                              forvar35 : forvar59) ?
                          $signed((8'hb7)) : $unsigned((8'hb5))) ^~ {$signed(forvar10)}));
                    end
                end
              else
                begin
                  for (forvar70 = (1'h0); (forvar70 < (1'h0)); forvar70 = (forvar70 + (1'h1)))
                    begin
                      reg71 <= (reg114[(3'h5):(3'h4)] & (({reg138} ?
                              reg66 : (reg98 ? reg59 : (8'hb4))) ?
                          ($unsigned(reg23) ?
                              (+reg72) : $unsigned(reg88)) : reg71));
                    end
                  if (reg93[(1'h0):(1'h0)])
                    begin
                      reg72 <= (8'ha9);
                      reg73 <= ((~|((+reg75) ? (8'hb2) : (!reg128))) ?
                          $unsigned(((-reg136) ?
                              (!reg66) : {reg93})) : $signed($unsigned((reg95 >= reg56))));
                      reg74 <= forvar10[(2'h3):(2'h2)];
                      reg75 <= $signed((+$signed($signed(forvar85))));
                    end
                  else
                    begin
                      reg72 <= (8'hb4);
                      reg73 <= reg133;
                      reg74 <= $unsigned($unsigned(reg30[(1'h1):(1'h0)]));
                    end
                  for (forvar76 = (1'h0); (forvar76 < (1'h0)); forvar76 = (forvar76 + (1'h1)))
                    begin
                      reg77 <= forvar50;
                      reg78 <= (+reg64);
                      reg79 <= forvar4;
                      reg80 <= ((reg125 ?
                              (reg39[(4'h9):(2'h3)] ?
                                  (reg39 - forvar9) : (reg75 == forvar10)) : forvar59[(3'h4):(1'h1)]) ?
                          ((~^$signed((8'hb8))) ?
                              $signed($unsigned((8'ha3))) : ($unsigned(reg65) <<< (reg6 ^ reg38))) : ((((8'ha3) ?
                                      forvar20 : forvar58) ?
                                  ((8'hb6) << forvar135) : $signed(reg30)) ?
                              (reg129 >> $unsigned(forvar99)) : reg109[(2'h2):(1'h0)]));
                    end
                end
              for (forvar84 = (1'h0); (forvar84 < (1'h0)); forvar84 = (forvar84 + (1'h1)))
                begin
                  reg85 <= ($unsigned(reg52) == reg40);
                  for (forvar86 = (1'h0); (forvar86 < (2'h3)); forvar86 = (forvar86 + (1'h1)))
                    begin
                      reg87 <= (-$signed(($unsigned((8'ha6)) ?
                          (reg84 ? reg70 : (8'hb3)) : forvar8[(2'h3):(1'h0)])));
                      reg88 <= {(forvar9[(1'h1):(1'h0)] ?
                              $unsigned((reg92 >= forvar67)) : reg7[(1'h0):(1'h0)])};
                      reg89 <= (8'hb2);
                      reg90 <= ({$signed($signed(reg53))} ?
                          $unsigned(reg52) : (&reg125));
                    end
                  if ((forvar50 & reg102[(2'h2):(1'h1)]))
                    begin
                      reg91 <= $unsigned($unsigned($unsigned({reg47})));
                      reg92 <= (forvar127[(3'h5):(2'h3)] ?
                          reg103 : $signed(reg9));
                    end
                  else
                    begin
                      reg91 <= (reg4[(2'h3):(1'h1)] - $signed(reg134[(1'h1):(1'h1)]));
                      reg92 <= ($unsigned($unsigned((reg21 >> forvar82))) ?
                          $unsigned(forvar22) : forvar82);
                      reg93 <= (~&$unsigned(reg49));
                      reg94 <= reg15[(4'hc):(3'h6)];
                    end
                end
            end
        end
    end
  assign wire139 = (reg90 ?
                       (~&$signed((reg16 ?
                           reg79 : reg88))) : $unsigned($signed((reg103 ?
                           (8'ha3) : forvar54))));
  assign wire140 = $unsigned($unsigned($signed((+wire1))));
  assign wire141 = {reg131[(4'h8):(3'h5)]};
  assign wire142 = (forvar104[(2'h2):(1'h0)] ?
                       $signed($unsigned((reg118 ?
                           reg113 : reg70))) : ($signed((8'hb9)) ?
                           reg4[(1'h0):(1'h0)] : $signed({reg113})));
  assign wire143 = {(($unsigned(reg56) ?
                               reg93[(1'h0):(1'h0)] : $signed(reg67)) ?
                           forvar82[(2'h2):(1'h0)] : ((reg22 ?
                                   reg33 : forvar57) ?
                               reg69 : (reg12 ? (8'hb0) : reg108)))};
  assign wire144 = $signed($unsigned(reg24[(3'h6):(2'h3)]));
  module145 modinst3106 (.y(wire3105), .wire149(reg107), .wire148(forvar54), .wire147(reg120), .wire146(reg125), .clk(clk));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module145
#(parameter param3104 = (~((^(~|(8'hb3))) ? (^~(8'hba)) : (8'hba))))
(y, clk, wire149, wire148, wire147, wire146);
  output wire [(32'h143a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire149;
  input wire signed [(4'ha):(1'h0)] wire148;
  input wire signed [(3'h4):(1'h0)] wire147;
  input wire [(3'h7):(1'h0)] wire146;
  wire [(3'h5):(1'h0)] wire3103;
  wire [(4'hd):(1'h0)] wire3102;
  reg signed [(5'h10):(1'h0)] reg3101 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3100 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3099 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3098 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3097 = (1'h0);
  reg [(4'ha):(1'h0)] reg3096 = (1'h0);
  reg [(2'h3):(1'h0)] reg3095 = (1'h0);
  reg [(4'he):(1'h0)] forvar3094 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3093 = (1'h0);
  reg [(4'h9):(1'h0)] reg3092 = (1'h0);
  reg [(3'h5):(1'h0)] reg3091 = (1'h0);
  reg [(4'hf):(1'h0)] reg3090 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3089 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3088 = (1'h0);
  reg [(4'ha):(1'h0)] reg3087 = (1'h0);
  reg [(3'h7):(1'h0)] reg3086 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3085 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3084 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3083 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3082 = (1'h0);
  reg [(4'he):(1'h0)] reg3081 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3080 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3079 = (1'h0);
  reg [(4'hb):(1'h0)] reg3078 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3077 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3076 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3073 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3076 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3075 = (1'h0);
  reg [(4'hc):(1'h0)] reg3074 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3073 = (1'h0);
  reg [(5'h10):(1'h0)] reg3072 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3071 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3070 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3069 = (1'h0);
  reg [(4'hc):(1'h0)] reg3068 = (1'h0);
  reg [(4'ha):(1'h0)] reg3067 = (1'h0);
  reg [(4'he):(1'h0)] reg3066 = (1'h0);
  reg [(3'h4):(1'h0)] reg3065 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3064 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3063 = (1'h0);
  reg [(4'h8):(1'h0)] reg3062 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3061 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3060 = (1'h0);
  reg [(3'h7):(1'h0)] reg3059 = (1'h0);
  reg [(4'hd):(1'h0)] reg3058 = (1'h0);
  reg [(3'h5):(1'h0)] reg3057 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3056 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3053 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3048 = (1'h0);
  reg [(3'h7):(1'h0)] reg3056 = (1'h0);
  reg [(4'ha):(1'h0)] reg3055 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3054 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3053 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3052 = (1'h0);
  reg [(4'ha):(1'h0)] reg3051 = (1'h0);
  reg [(2'h3):(1'h0)] reg3050 = (1'h0);
  reg [(3'h4):(1'h0)] reg3049 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3048 = (1'h0);
  reg [(4'he):(1'h0)] forvar3047 = (1'h0);
  reg [(2'h3):(1'h0)] reg3046 = (1'h0);
  reg [(4'hb):(1'h0)] reg3045 = (1'h0);
  reg [(3'h4):(1'h0)] reg3044 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3043 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3042 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3037 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3041 = (1'h0);
  reg [(3'h5):(1'h0)] reg3040 = (1'h0);
  reg [(2'h2):(1'h0)] reg3039 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3038 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3037 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3036 = (1'h0);
  reg [(4'hd):(1'h0)] reg3035 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3034 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3029 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3033 = (1'h0);
  reg [(4'h9):(1'h0)] reg3032 = (1'h0);
  reg [(4'hb):(1'h0)] reg3031 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3030 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3029 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3028 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3027 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3026 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3024 = (1'h0);
  reg [(4'hf):(1'h0)] reg3023 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3019 = (1'h0);
  reg [(4'hb):(1'h0)] reg3018 = (1'h0);
  reg [(3'h6):(1'h0)] reg3013 = (1'h0);
  reg [(4'ha):(1'h0)] reg3025 = (1'h0);
  reg [(4'hc):(1'h0)] reg3024 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3023 = (1'h0);
  reg [(3'h5):(1'h0)] reg3022 = (1'h0);
  reg [(3'h4):(1'h0)] reg3021 = (1'h0);
  reg [(3'h4):(1'h0)] reg3020 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3019 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3018 = (1'h0);
  reg [(2'h3):(1'h0)] reg3017 = (1'h0);
  reg [(2'h3):(1'h0)] reg3016 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3015 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3014 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3013 = (1'h0);
  reg [(4'ha):(1'h0)] reg3012 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3011 = (1'h0);
  reg [(3'h5):(1'h0)] reg3010 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3009 = (1'h0);
  reg [(4'hb):(1'h0)] reg3008 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3007 = (1'h0);
  reg [(4'ha):(1'h0)] reg3006 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3005 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3004 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3003 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3002 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3001 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3000 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2999 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2996 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2998 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2997 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2996 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2995 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2994 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2993 = (1'h0);
  reg [(3'h7):(1'h0)] reg2992 = (1'h0);
  reg [(3'h6):(1'h0)] reg2991 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2990 = (1'h0);
  reg [(3'h5):(1'h0)] reg2989 = (1'h0);
  reg [(4'ha):(1'h0)] reg2988 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2987 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2986 = (1'h0);
  reg [(4'hd):(1'h0)] reg2985 = (1'h0);
  reg [(4'hd):(1'h0)] reg2984 = (1'h0);
  reg [(4'h8):(1'h0)] reg2983 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2982 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2981 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2980 = (1'h0);
  reg [(5'h10):(1'h0)] reg2979 = (1'h0);
  reg [(4'he):(1'h0)] forvar2978 = (1'h0);
  reg [(4'hb):(1'h0)] reg2977 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2976 = (1'h0);
  reg [(4'h9):(1'h0)] reg2975 = (1'h0);
  reg [(4'hd):(1'h0)] reg2974 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2973 = (1'h0);
  reg [(4'h9):(1'h0)] reg2972 = (1'h0);
  reg [(4'h8):(1'h0)] reg2964 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2971 = (1'h0);
  reg [(2'h2):(1'h0)] reg2970 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2969 = (1'h0);
  reg [(4'hc):(1'h0)] reg2968 = (1'h0);
  reg [(3'h5):(1'h0)] reg2967 = (1'h0);
  reg [(4'ha):(1'h0)] reg2966 = (1'h0);
  reg [(3'h5):(1'h0)] reg2965 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2964 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2963 = (1'h0);
  reg [(3'h7):(1'h0)] reg2962 = (1'h0);
  reg [(4'hf):(1'h0)] reg2961 = (1'h0);
  reg [(2'h2):(1'h0)] reg2960 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2959 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2958 = (1'h0);
  reg [(3'h7):(1'h0)] reg2952 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2951 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2957 = (1'h0);
  reg [(4'hf):(1'h0)] reg2956 = (1'h0);
  reg [(4'h8):(1'h0)] reg2955 = (1'h0);
  reg [(4'h8):(1'h0)] reg2954 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2953 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2952 = (1'h0);
  reg [(4'hc):(1'h0)] reg2951 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2950 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2949 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2948 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2947 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2946 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2945 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2944 = (1'h0);
  reg [(3'h4):(1'h0)] reg2943 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2942 = (1'h0);
  reg [(3'h4):(1'h0)] reg2941 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2940 = (1'h0);
  reg [(4'he):(1'h0)] reg2939 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2938 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2937 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2936 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2935 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2934 = (1'h0);
  reg [(4'he):(1'h0)] reg2933 = (1'h0);
  reg [(2'h2):(1'h0)] reg2932 = (1'h0);
  reg [(2'h2):(1'h0)] reg2931 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2930 = (1'h0);
  reg [(4'he):(1'h0)] reg2929 = (1'h0);
  reg [(4'hd):(1'h0)] reg2928 = (1'h0);
  reg [(3'h5):(1'h0)] reg2927 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2926 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2925 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2924 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2923 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2922 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2921 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2919 = (1'h0);
  reg [(4'hb):(1'h0)] reg2921 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2918 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2912 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2914 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2910 = (1'h0);
  reg [(4'hd):(1'h0)] reg2906 = (1'h0);
  reg [(4'hd):(1'h0)] reg2905 = (1'h0);
  reg [(4'he):(1'h0)] forvar2917 = (1'h0);
  reg [(4'ha):(1'h0)] reg2916 = (1'h0);
  reg [(4'hb):(1'h0)] reg2920 = (1'h0);
  reg [(4'ha):(1'h0)] reg2919 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2918 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2917 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2916 = (1'h0);
  reg [(2'h3):(1'h0)] reg2915 = (1'h0);
  reg [(2'h3):(1'h0)] reg2914 = (1'h0);
  reg [(4'h8):(1'h0)] reg2913 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2912 = (1'h0);
  reg [(4'ha):(1'h0)] reg2911 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2910 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2909 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2908 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2907 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2906 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2905 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2904 = (1'h0);
  reg [(4'he):(1'h0)] reg2903 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2902 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2901 = (1'h0);
  reg [(2'h2):(1'h0)] reg2900 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2899 = (1'h0);
  reg [(2'h2):(1'h0)] reg2898 = (1'h0);
  reg [(2'h3):(1'h0)] reg2897 = (1'h0);
  reg [(3'h5):(1'h0)] reg2896 = (1'h0);
  reg [(4'he):(1'h0)] reg2895 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2894 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2893 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2892 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2891 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2890 = (1'h0);
  reg [(3'h7):(1'h0)] reg2889 = (1'h0);
  reg [(4'h9):(1'h0)] reg2888 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2887 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2886 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2885 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2884 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2883 = (1'h0);
  reg [(3'h6):(1'h0)] reg2882 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2881 = (1'h0);
  reg [(2'h3):(1'h0)] reg2880 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2879 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2878 = (1'h0);
  reg [(4'hd):(1'h0)] reg2877 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2876 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2875 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2874 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2873 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2872 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2871 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2870 = (1'h0);
  reg [(4'he):(1'h0)] forvar2869 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2868 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2867 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2866 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2865 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2864 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2863 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2862 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2861 = (1'h0);
  reg [(4'hd):(1'h0)] reg2860 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2859 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2854 = (1'h0);
  reg [(4'ha):(1'h0)] reg2851 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2850 = (1'h0);
  reg [(2'h3):(1'h0)] reg2859 = (1'h0);
  reg [(5'h10):(1'h0)] reg2858 = (1'h0);
  reg [(4'h9):(1'h0)] reg2857 = (1'h0);
  reg [(4'ha):(1'h0)] reg2856 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2855 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2854 = (1'h0);
  reg [(2'h2):(1'h0)] reg2853 = (1'h0);
  reg [(2'h3):(1'h0)] reg2852 = (1'h0);
  reg [(4'he):(1'h0)] forvar2851 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2849 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2850 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2849 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2848 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2847 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2846 = (1'h0);
  reg [(4'h8):(1'h0)] reg2845 = (1'h0);
  reg [(2'h2):(1'h0)] reg2844 = (1'h0);
  reg [(4'h9):(1'h0)] reg2843 = (1'h0);
  reg [(4'hf):(1'h0)] reg2842 = (1'h0);
  reg [(2'h2):(1'h0)] reg2841 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2840 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2839 = (1'h0);
  reg [(4'hb):(1'h0)] reg2838 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2837 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2836 = (1'h0);
  reg [(4'ha):(1'h0)] reg2833 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2835 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2834 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2833 = (1'h0);
  reg [(4'hf):(1'h0)] reg2832 = (1'h0);
  reg [(4'hf):(1'h0)] reg2831 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2830 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2829 = (1'h0);
  reg [(4'hb):(1'h0)] reg2828 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2827 = (1'h0);
  reg [(5'h10):(1'h0)] reg2826 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2825 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2794 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2813 = (1'h0);
  reg [(3'h7):(1'h0)] reg2812 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2811 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2824 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2823 = (1'h0);
  reg [(3'h5):(1'h0)] reg2822 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2821 = (1'h0);
  reg [(4'hb):(1'h0)] reg2820 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2819 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2818 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2817 = (1'h0);
  reg [(3'h4):(1'h0)] reg2816 = (1'h0);
  reg [(3'h5):(1'h0)] reg2815 = (1'h0);
  reg [(4'he):(1'h0)] reg2814 = (1'h0);
  reg [(2'h2):(1'h0)] reg2813 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2812 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2811 = (1'h0);
  reg [(2'h3):(1'h0)] reg2810 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2809 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2808 = (1'h0);
  reg [(2'h3):(1'h0)] reg2807 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2806 = (1'h0);
  reg [(4'ha):(1'h0)] reg2805 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2804 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2802 = (1'h0);
  reg [(3'h6):(1'h0)] reg2803 = (1'h0);
  reg [(4'ha):(1'h0)] reg2802 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2801 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2800 = (1'h0);
  reg [(3'h6):(1'h0)] reg2799 = (1'h0);
  reg [(3'h6):(1'h0)] reg2798 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2797 = (1'h0);
  reg [(4'hd):(1'h0)] reg2796 = (1'h0);
  reg [(4'ha):(1'h0)] reg2795 = (1'h0);
  reg [(4'he):(1'h0)] forvar2794 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2793 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2792 = (1'h0);
  reg [(4'h9):(1'h0)] reg2791 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2790 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2789 = (1'h0);
  reg [(4'hb):(1'h0)] reg2788 = (1'h0);
  reg [(4'h9):(1'h0)] reg2787 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2786 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2785 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2784 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2783 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2782 = (1'h0);
  reg [(4'he):(1'h0)] forvar2781 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2780 = (1'h0);
  reg [(3'h7):(1'h0)] reg2779 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2778 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2777 = (1'h0);
  reg [(4'ha):(1'h0)] reg2776 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2775 = (1'h0);
  reg [(4'he):(1'h0)] forvar2774 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2773 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2772 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2771 = (1'h0);
  reg [(3'h5):(1'h0)] reg2770 = (1'h0);
  reg [(5'h10):(1'h0)] reg2769 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2768 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2767 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2766 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2765 = (1'h0);
  reg [(4'hf):(1'h0)] reg2764 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2763 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2762 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2761 = (1'h0);
  reg [(5'h10):(1'h0)] reg2760 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2759 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2758 = (1'h0);
  reg [(4'hd):(1'h0)] reg2757 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2756 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2755 = (1'h0);
  reg [(4'he):(1'h0)] forvar2754 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2753 = (1'h0);
  reg [(4'hf):(1'h0)] reg2752 = (1'h0);
  reg [(4'hf):(1'h0)] reg2751 = (1'h0);
  reg [(2'h3):(1'h0)] reg2750 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2749 = (1'h0);
  reg [(4'h8):(1'h0)] reg2748 = (1'h0);
  reg [(4'hf):(1'h0)] reg2747 = (1'h0);
  reg [(3'h7):(1'h0)] reg2746 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2745 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2744 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2743 = (1'h0);
  reg [(3'h5):(1'h0)] reg2742 = (1'h0);
  reg [(4'ha):(1'h0)] reg2741 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2740 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2739 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2738 = (1'h0);
  reg [(4'he):(1'h0)] reg2737 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2736 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2735 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2734 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2733 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2732 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2726 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2723 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2718 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2715 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2710 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2731 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2730 = (1'h0);
  reg [(4'hb):(1'h0)] reg2729 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2728 = (1'h0);
  reg [(3'h6):(1'h0)] reg2727 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2726 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2719 = (1'h0);
  reg [(3'h7):(1'h0)] reg2725 = (1'h0);
  reg [(4'ha):(1'h0)] reg2724 = (1'h0);
  reg [(5'h10):(1'h0)] reg2723 = (1'h0);
  reg [(4'hf):(1'h0)] reg2722 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2721 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2720 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2719 = (1'h0);
  reg [(3'h7):(1'h0)] reg2718 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2717 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2716 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2715 = (1'h0);
  reg [(4'hb):(1'h0)] reg2714 = (1'h0);
  reg [(3'h5):(1'h0)] reg2713 = (1'h0);
  reg [(4'hd):(1'h0)] reg2712 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2711 = (1'h0);
  reg [(4'hc):(1'h0)] reg2710 = (1'h0);
  reg [(3'h7):(1'h0)] reg2709 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2708 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2686 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2676 = (1'h0);
  reg [(3'h4):(1'h0)] reg2707 = (1'h0);
  reg [(4'hb):(1'h0)] reg2706 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2705 = (1'h0);
  reg [(3'h7):(1'h0)] reg2704 = (1'h0);
  reg [(3'h6):(1'h0)] reg2703 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2702 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2687 = (1'h0);
  reg [(3'h7):(1'h0)] reg2688 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2683 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2682 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2681 = (1'h0);
  reg [(3'h4):(1'h0)] reg2678 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2701 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2700 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2699 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2698 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2697 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2695 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2692 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2689 = (1'h0);
  reg [(4'ha):(1'h0)] reg2696 = (1'h0);
  reg [(2'h3):(1'h0)] reg2695 = (1'h0);
  reg [(4'hc):(1'h0)] reg2694 = (1'h0);
  reg [(4'hf):(1'h0)] reg2693 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2692 = (1'h0);
  reg [(3'h7):(1'h0)] reg2691 = (1'h0);
  reg [(2'h3):(1'h0)] reg2690 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2689 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2688 = (1'h0);
  reg [(2'h3):(1'h0)] reg2687 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2686 = (1'h0);
  reg [(4'he):(1'h0)] reg2685 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2684 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2683 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2682 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2681 = (1'h0);
  reg [(5'h10):(1'h0)] reg2680 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2679 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2678 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2677 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2676 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire2675;
  wire signed [(4'hc):(1'h0)] wire581;
  wire signed [(5'h10):(1'h0)] wire285;
  wire [(4'hc):(1'h0)] wire226;
  wire signed [(4'hb):(1'h0)] wire225;
  wire [(4'ha):(1'h0)] wire224;
  reg signed [(4'ha):(1'h0)] reg223 = (1'h0);
  reg [(3'h5):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg221 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg219 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar218 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar217 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar216 = (1'h0);
  reg [(5'h10):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg214 = (1'h0);
  reg [(4'hd):(1'h0)] reg213 = (1'h0);
  reg [(4'he):(1'h0)] reg212 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg211 = (1'h0);
  reg [(4'he):(1'h0)] reg210 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg209 = (1'h0);
  reg [(4'h8):(1'h0)] forvar208 = (1'h0);
  reg [(4'ha):(1'h0)] reg207 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar206 = (1'h0);
  reg [(4'hf):(1'h0)] forvar205 = (1'h0);
  reg signed [(4'he):(1'h0)] reg204 = (1'h0);
  reg [(4'hf):(1'h0)] reg203 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg202 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(3'h7):(1'h0)] reg200 = (1'h0);
  reg [(2'h2):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar198 = (1'h0);
  reg [(4'h9):(1'h0)] forvar197 = (1'h0);
  reg [(3'h6):(1'h0)] forvar196 = (1'h0);
  reg [(4'ha):(1'h0)] forvar172 = (1'h0);
  reg [(4'hb):(1'h0)] forvar169 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar164 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar161 = (1'h0);
  reg [(3'h5):(1'h0)] forvar157 = (1'h0);
  reg [(4'h9):(1'h0)] forvar156 = (1'h0);
  reg [(4'h9):(1'h0)] forvar153 = (1'h0);
  reg [(4'hb):(1'h0)] reg195 = (1'h0);
  reg [(4'hc):(1'h0)] reg194 = (1'h0);
  reg signed [(4'he):(1'h0)] reg193 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg192 = (1'h0);
  reg [(4'hb):(1'h0)] forvar191 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg190 = (1'h0);
  reg [(5'h10):(1'h0)] reg189 = (1'h0);
  reg [(4'hf):(1'h0)] reg188 = (1'h0);
  reg [(4'hf):(1'h0)] reg187 = (1'h0);
  reg signed [(4'he):(1'h0)] reg186 = (1'h0);
  reg [(4'hf):(1'h0)] reg185 = (1'h0);
  reg [(5'h10):(1'h0)] forvar184 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg183 = (1'h0);
  reg [(3'h4):(1'h0)] reg182 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg180 = (1'h0);
  reg [(4'h8):(1'h0)] forvar179 = (1'h0);
  reg [(3'h5):(1'h0)] reg178 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar176 = (1'h0);
  reg [(2'h3):(1'h0)] reg175 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg174 = (1'h0);
  reg [(3'h7):(1'h0)] reg173 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg172 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg171 = (1'h0);
  reg [(4'hb):(1'h0)] forvar170 = (1'h0);
  reg [(5'h10):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar168 = (1'h0);
  reg [(4'hf):(1'h0)] reg167 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg166 = (1'h0);
  reg [(4'h8):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg164 = (1'h0);
  reg [(4'ha):(1'h0)] reg163 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg162 = (1'h0);
  reg [(5'h10):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg160 = (1'h0);
  reg [(3'h6):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg158 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg157 = (1'h0);
  reg [(3'h6):(1'h0)] reg156 = (1'h0);
  reg [(4'ha):(1'h0)] reg155 = (1'h0);
  reg [(4'h9):(1'h0)] reg154 = (1'h0);
  reg [(3'h5):(1'h0)] reg153 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar152 = (1'h0);
  reg [(5'h10):(1'h0)] forvar151 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire150;
  wire [(2'h3):(1'h0)] wire583;
  wire signed [(4'hd):(1'h0)] wire2673;
  assign y = {wire3103,
                 wire3102,
                 reg3101,
                 reg3100,
                 reg3099,
                 forvar3098,
                 reg3097,
                 reg3096,
                 reg3095,
                 forvar3094,
                 reg3093,
                 reg3092,
                 reg3091,
                 reg3090,
                 forvar3089,
                 reg3088,
                 reg3087,
                 reg3086,
                 reg3085,
                 forvar3084,
                 forvar3083,
                 reg3082,
                 reg3081,
                 reg3080,
                 reg3079,
                 reg3078,
                 reg3077,
                 forvar3076,
                 reg3073,
                 reg3076,
                 reg3075,
                 reg3074,
                 forvar3073,
                 reg3072,
                 forvar3071,
                 reg3070,
                 reg3069,
                 reg3068,
                 reg3067,
                 reg3066,
                 reg3065,
                 reg3064,
                 reg3063,
                 reg3062,
                 forvar3061,
                 forvar3060,
                 reg3059,
                 reg3058,
                 reg3057,
                 forvar3056,
                 forvar3053,
                 forvar3048,
                 reg3056,
                 reg3055,
                 reg3054,
                 reg3053,
                 reg3052,
                 reg3051,
                 reg3050,
                 reg3049,
                 reg3048,
                 forvar3047,
                 reg3046,
                 reg3045,
                 reg3044,
                 reg3043,
                 reg3042,
                 reg3037,
                 reg3041,
                 reg3040,
                 reg3039,
                 reg3038,
                 forvar3037,
                 reg3036,
                 reg3035,
                 reg3034,
                 reg3029,
                 reg3033,
                 reg3032,
                 reg3031,
                 reg3030,
                 forvar3029,
                 reg3028,
                 forvar3027,
                 forvar3026,
                 forvar3024,
                 reg3023,
                 forvar3019,
                 reg3018,
                 reg3013,
                 reg3025,
                 reg3024,
                 forvar3023,
                 reg3022,
                 reg3021,
                 reg3020,
                 reg3019,
                 forvar3018,
                 reg3017,
                 reg3016,
                 reg3015,
                 reg3014,
                 forvar3013,
                 reg3012,
                 reg3011,
                 reg3010,
                 reg3009,
                 reg3008,
                 forvar3007,
                 reg3006,
                 forvar3005,
                 reg3004,
                 reg3003,
                 forvar3002,
                 forvar3001,
                 reg3000,
                 forvar2999,
                 forvar2996,
                 reg2998,
                 reg2997,
                 reg2996,
                 reg2995,
                 reg2994,
                 reg2993,
                 reg2992,
                 reg2991,
                 reg2990,
                 reg2989,
                 reg2988,
                 reg2987,
                 reg2986,
                 reg2985,
                 reg2984,
                 reg2983,
                 reg2982,
                 forvar2981,
                 forvar2980,
                 reg2979,
                 forvar2978,
                 reg2977,
                 reg2976,
                 reg2975,
                 reg2974,
                 reg2973,
                 reg2972,
                 reg2964,
                 reg2971,
                 reg2970,
                 reg2969,
                 reg2968,
                 reg2967,
                 reg2966,
                 reg2965,
                 forvar2964,
                 reg2963,
                 reg2962,
                 reg2961,
                 reg2960,
                 forvar2959,
                 forvar2958,
                 reg2952,
                 forvar2951,
                 reg2957,
                 reg2956,
                 reg2955,
                 reg2954,
                 reg2953,
                 forvar2952,
                 reg2951,
                 forvar2950,
                 reg2949,
                 reg2948,
                 reg2947,
                 reg2946,
                 forvar2945,
                 reg2944,
                 reg2943,
                 reg2942,
                 reg2941,
                 forvar2940,
                 reg2939,
                 reg2938,
                 reg2937,
                 reg2936,
                 forvar2935,
                 forvar2934,
                 reg2933,
                 reg2932,
                 reg2931,
                 forvar2930,
                 reg2929,
                 reg2928,
                 reg2927,
                 reg2926,
                 forvar2925,
                 reg2924,
                 reg2923,
                 reg2922,
                 forvar2921,
                 forvar2919,
                 reg2921,
                 forvar2918,
                 reg2912,
                 forvar2914,
                 reg2910,
                 reg2906,
                 reg2905,
                 forvar2917,
                 reg2916,
                 reg2920,
                 reg2919,
                 reg2918,
                 reg2917,
                 forvar2916,
                 reg2915,
                 reg2914,
                 reg2913,
                 forvar2912,
                 reg2911,
                 forvar2910,
                 reg2909,
                 reg2908,
                 reg2907,
                 forvar2906,
                 forvar2905,
                 forvar2904,
                 reg2903,
                 reg2902,
                 reg2901,
                 reg2900,
                 reg2899,
                 reg2898,
                 reg2897,
                 reg2896,
                 reg2895,
                 reg2894,
                 reg2893,
                 reg2892,
                 forvar2891,
                 reg2890,
                 reg2889,
                 reg2888,
                 reg2887,
                 reg2886,
                 forvar2885,
                 forvar2884,
                 reg2883,
                 reg2882,
                 reg2881,
                 reg2880,
                 reg2879,
                 forvar2878,
                 reg2877,
                 reg2876,
                 reg2875,
                 reg2874,
                 forvar2873,
                 reg2872,
                 forvar2871,
                 forvar2870,
                 forvar2869,
                 forvar2868,
                 reg2867,
                 reg2866,
                 forvar2865,
                 forvar2864,
                 reg2863,
                 reg2862,
                 reg2861,
                 reg2860,
                 forvar2859,
                 forvar2854,
                 reg2851,
                 forvar2850,
                 reg2859,
                 reg2858,
                 reg2857,
                 reg2856,
                 forvar2855,
                 reg2854,
                 reg2853,
                 reg2852,
                 forvar2851,
                 forvar2849,
                 reg2850,
                 reg2849,
                 reg2848,
                 reg2847,
                 reg2846,
                 reg2845,
                 reg2844,
                 reg2843,
                 reg2842,
                 reg2841,
                 forvar2840,
                 forvar2839,
                 reg2838,
                 forvar2837,
                 forvar2836,
                 reg2833,
                 reg2835,
                 reg2834,
                 forvar2833,
                 reg2832,
                 reg2831,
                 forvar2830,
                 forvar2829,
                 reg2828,
                 reg2827,
                 reg2826,
                 forvar2825,
                 reg2794,
                 forvar2813,
                 reg2812,
                 forvar2811,
                 reg2824,
                 reg2823,
                 reg2822,
                 forvar2821,
                 reg2820,
                 reg2819,
                 reg2818,
                 forvar2817,
                 reg2816,
                 reg2815,
                 reg2814,
                 reg2813,
                 forvar2812,
                 reg2811,
                 reg2810,
                 reg2809,
                 reg2808,
                 reg2807,
                 reg2806,
                 reg2805,
                 forvar2804,
                 forvar2802,
                 reg2803,
                 reg2802,
                 reg2801,
                 reg2800,
                 reg2799,
                 reg2798,
                 reg2797,
                 reg2796,
                 reg2795,
                 forvar2794,
                 forvar2793,
                 reg2792,
                 reg2791,
                 reg2790,
                 forvar2789,
                 reg2788,
                 reg2787,
                 forvar2786,
                 forvar2785,
                 forvar2784,
                 reg2783,
                 reg2782,
                 forvar2781,
                 forvar2780,
                 reg2779,
                 reg2778,
                 reg2777,
                 reg2776,
                 forvar2775,
                 forvar2774,
                 forvar2773,
                 reg2772,
                 reg2771,
                 reg2770,
                 reg2769,
                 reg2768,
                 reg2767,
                 reg2766,
                 forvar2765,
                 reg2764,
                 reg2763,
                 forvar2762,
                 forvar2761,
                 reg2760,
                 reg2759,
                 reg2758,
                 reg2757,
                 reg2756,
                 forvar2755,
                 forvar2754,
                 reg2753,
                 reg2752,
                 reg2751,
                 reg2750,
                 forvar2749,
                 reg2748,
                 reg2747,
                 reg2746,
                 reg2745,
                 reg2744,
                 reg2743,
                 reg2742,
                 reg2741,
                 forvar2740,
                 forvar2739,
                 forvar2738,
                 reg2737,
                 forvar2736,
                 reg2735,
                 forvar2734,
                 forvar2733,
                 reg2732,
                 reg2726,
                 forvar2723,
                 forvar2718,
                 forvar2715,
                 forvar2710,
                 reg2731,
                 reg2730,
                 reg2729,
                 reg2728,
                 reg2727,
                 forvar2726,
                 forvar2719,
                 reg2725,
                 reg2724,
                 reg2723,
                 reg2722,
                 reg2721,
                 reg2720,
                 reg2719,
                 reg2718,
                 reg2717,
                 reg2716,
                 reg2715,
                 reg2714,
                 reg2713,
                 reg2712,
                 reg2711,
                 reg2710,
                 reg2709,
                 forvar2708,
                 forvar2686,
                 reg2676,
                 reg2707,
                 reg2706,
                 reg2705,
                 reg2704,
                 reg2703,
                 forvar2702,
                 forvar2687,
                 reg2688,
                 reg2683,
                 forvar2682,
                 reg2681,
                 reg2678,
                 reg2701,
                 reg2700,
                 reg2699,
                 reg2698,
                 reg2697,
                 forvar2695,
                 reg2692,
                 forvar2689,
                 reg2696,
                 reg2695,
                 reg2694,
                 reg2693,
                 forvar2692,
                 reg2691,
                 reg2690,
                 reg2689,
                 forvar2688,
                 reg2687,
                 reg2686,
                 reg2685,
                 reg2684,
                 forvar2683,
                 reg2682,
                 forvar2681,
                 reg2680,
                 reg2679,
                 forvar2678,
                 forvar2677,
                 forvar2676,
                 wire2675,
                 wire581,
                 wire285,
                 wire226,
                 wire225,
                 wire224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 forvar218,
                 forvar217,
                 forvar216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 forvar208,
                 reg207,
                 forvar206,
                 forvar205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 forvar198,
                 forvar197,
                 forvar196,
                 forvar172,
                 forvar169,
                 reg168,
                 forvar164,
                 forvar161,
                 forvar157,
                 forvar156,
                 forvar153,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 forvar191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 forvar184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 forvar179,
                 reg178,
                 reg177,
                 forvar176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 forvar170,
                 reg169,
                 forvar168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 forvar152,
                 forvar151,
                 wire150,
                 wire583,
                 wire2673,
                 (1'h0)};
  assign wire150 = (wire149 ?
                       {$unsigned($unsigned(wire148))} : $signed({$signed(wire149)}));
  always
    @(posedge clk) begin
      for (forvar151 = (1'h0); (forvar151 < (2'h3)); forvar151 = (forvar151 + (1'h1)))
        begin
          if (((wire150[(3'h5):(3'h5)] != (wire149[(4'ha):(2'h3)] - wire147)) ?
              $signed((!$signed(wire146))) : forvar151[(1'h1):(1'h1)]))
            begin
              for (forvar152 = (1'h0); (forvar152 < (2'h2)); forvar152 = (forvar152 + (1'h1)))
                begin
                  if ($unsigned((((|forvar152) != (forvar151 < (8'hb7))) ?
                      (wire146 >> forvar151[(3'h5):(3'h5)]) : $unsigned($unsigned((8'hb0))))))
                    begin
                      reg153 <= $unsigned(((+wire147[(2'h3):(1'h1)]) >>> $unsigned($unsigned(wire148))));
                      reg154 <= $unsigned((wire146[(2'h3):(2'h2)] ?
                          (-{wire147}) : wire147));
                      reg155 <= forvar152[(1'h1):(1'h1)];
                      reg156 <= reg153[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg153 <= $signed((($unsigned(wire149) ?
                          reg153[(1'h0):(1'h0)] : (^~forvar151)) - reg155));
                      reg154 <= $unsigned((((wire148 ? reg156 : wire149) ?
                              (!reg153) : (reg155 ? wire147 : reg153)) ?
                          $unsigned((^reg155)) : wire146[(2'h3):(1'h1)]));
                    end
                  if ((wire150 ? {wire146[(2'h3):(1'h1)]} : wire147))
                    begin
                      reg157 <= (!{$unsigned((|reg156))});
                      reg158 <= wire146;
                      reg159 <= wire148[(2'h3):(2'h2)];
                      reg160 <= $signed(($signed((wire146 >>> wire147)) ?
                          reg153[(3'h5):(3'h5)] : (8'h9f)));
                    end
                  else
                    begin
                      reg157 <= reg157;
                      reg158 <= $unsigned(reg153);
                    end
                  if (((^wire148) ?
                      (~wire146[(2'h2):(2'h2)]) : (&$signed($unsigned(wire148)))))
                    begin
                      reg161 <= {$unsigned(reg157[(3'h7):(1'h0)])};
                    end
                  else
                    begin
                      reg161 <= $unsigned(($unsigned($unsigned(reg155)) ?
                          {reg157} : (~(reg154 ? reg159 : reg154))));
                      reg162 <= ((($signed((8'haf)) ?
                                  $unsigned(wire146) : ((8'hb2) ?
                                      (8'hb7) : reg159)) ?
                              reg161 : $signed($unsigned(reg154))) ?
                          {wire148} : wire146);
                      reg163 <= ($unsigned(reg162) ?
                          reg154[(3'h7):(3'h5)] : reg155);
                    end
                  if ((((~(wire150 <<< (8'ha3))) - {$signed(reg156)}) ?
                      $unsigned(forvar152[(2'h3):(2'h2)]) : reg154[(3'h4):(3'h4)]))
                    begin
                      reg164 <= $unsigned((wire150 & (~^$signed(reg163))));
                      reg165 <= ({(~&{wire146})} <= (8'haf));
                      reg166 <= (((reg157 ~^ (reg159 < reg161)) ?
                              ((reg158 || forvar151) >> wire146[(3'h4):(1'h0)]) : reg161[(4'he):(3'h4)]) ?
                          reg154 : (+($unsigned(reg161) & forvar152)));
                    end
                  else
                    begin
                      reg164 <= $signed($unsigned($unsigned({reg160})));
                      reg165 <= $signed($unsigned(((+reg162) >= (reg166 ?
                          (8'ha0) : (8'h9e)))));
                      reg166 <= $signed($unsigned(reg162[(3'h6):(1'h1)]));
                      reg167 <= reg159[(3'h6):(3'h5)];
                    end
                end
              for (forvar168 = (1'h0); (forvar168 < (1'h0)); forvar168 = (forvar168 + (1'h1)))
                begin
                  if ((&(^(|(~&reg160)))))
                    begin
                      reg169 <= $unsigned($signed(reg158[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg169 <= $signed($signed(wire149));
                    end
                end
              for (forvar170 = (1'h0); (forvar170 < (1'h0)); forvar170 = (forvar170 + (1'h1)))
                begin
                  if ($signed(reg155[(3'h6):(3'h6)]))
                    begin
                      reg171 <= forvar168;
                      reg172 <= reg165;
                      reg173 <= $signed($unsigned(reg163[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg171 <= $signed($unsigned($unsigned($unsigned(wire148))));
                      reg172 <= ((8'ha9) ?
                          $signed((reg167 || reg169)) : ($unsigned(reg157) << reg160[(1'h0):(1'h0)]));
                      reg173 <= (^~reg166[(1'h1):(1'h1)]);
                      reg174 <= $signed((~|reg156));
                    end
                  if ((reg165 ?
                      $signed(((reg171 ? wire149 : wire146) ?
                          reg173[(2'h2):(1'h1)] : $unsigned(wire150))) : (+reg159)))
                    begin
                      reg175 <= (forvar151[(4'hf):(2'h2)] ?
                          reg165[(2'h2):(1'h1)] : $unsigned(wire150[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg175 <= (-(({reg175} && forvar168[(1'h1):(1'h1)]) || {{reg157}}));
                    end
                  for (forvar176 = (1'h0); (forvar176 < (2'h3)); forvar176 = (forvar176 + (1'h1)))
                    begin
                      reg177 <= (reg160 << reg167[(4'hd):(1'h0)]);
                      reg178 <= reg172;
                    end
                  for (forvar179 = (1'h0); (forvar179 < (1'h1)); forvar179 = (forvar179 + (1'h1)))
                    begin
                      reg180 <= reg163;
                    end
                end
              if ((((reg174 - (~&wire150)) ?
                  reg177[(2'h2):(1'h1)] : reg175[(1'h1):(1'h0)]) * ((~(~&reg173)) || (reg172[(1'h1):(1'h0)] ?
                  (reg166 ? (8'haf) : reg157) : $unsigned(reg174)))))
                begin
                  if (reg160)
                    begin
                      reg181 <= (8'ha0);
                      reg182 <= $unsigned((^(~^(!reg169))));
                      reg183 <= ((reg171 >>> wire148) ?
                          (|(^~reg169)) : $signed($signed({wire147})));
                    end
                  else
                    begin
                      reg181 <= $signed(($signed($unsigned(reg162)) ?
                          reg156 : reg169));
                      reg182 <= $unsigned(wire148[(3'h6):(1'h0)]);
                    end
                  for (forvar184 = (1'h0); (forvar184 < (1'h1)); forvar184 = (forvar184 + (1'h1)))
                    begin
                      reg185 <= $unsigned($unsigned((+wire150[(2'h3):(2'h3)])));
                      reg186 <= $signed(reg153[(2'h3):(2'h3)]);
                    end
                  if ((~|reg172))
                    begin
                      reg187 <= ((-$unsigned($unsigned(reg177))) ?
                          $unsigned($signed(forvar151)) : $unsigned(reg186[(3'h4):(1'h0)]));
                      reg188 <= (reg153 ?
                          {$unsigned((reg162 < reg159))} : $unsigned(($signed(reg181) + (reg156 ?
                              (8'ha9) : reg161))));
                      reg189 <= reg165[(2'h2):(2'h2)];
                      reg190 <= (-($unsigned(reg160[(3'h4):(1'h1)]) ?
                          reg160 : wire146));
                    end
                  else
                    begin
                      reg187 <= $unsigned(({(reg169 ? wire150 : reg187)} ?
                          {forvar176[(2'h2):(1'h0)]} : ($unsigned(reg155) > (|reg165))));
                    end
                  for (forvar191 = (1'h0); (forvar191 < (2'h3)); forvar191 = (forvar191 + (1'h1)))
                    begin
                      reg192 <= {{((reg173 >> reg178) ?
                                  reg155[(3'h6):(1'h0)] : {reg166})}};
                      reg193 <= $unsigned(($signed((!reg158)) & ((reg172 || forvar151) ?
                          ((8'ha8) ? (8'ha3) : reg192) : ((8'hba) ?
                              forvar184 : reg188))));
                      reg194 <= (-((((8'ha1) | reg171) >> (wire147 > reg174)) ?
                          reg187 : $signed($unsigned(reg190))));
                      reg195 <= (^(((|forvar176) == $signed((8'hac))) ?
                          reg181[(2'h2):(1'h1)] : {$signed(reg171)}));
                    end
                end
              else
                begin
                  if (($signed((^~(8'ha5))) ~^ (&$signed($unsigned(reg195)))))
                    begin
                      reg181 <= forvar179;
                    end
                  else
                    begin
                      reg181 <= reg185[(1'h0):(1'h0)];
                      reg182 <= $signed((~^(^reg171[(1'h0):(1'h0)])));
                    end
                end
            end
          else
            begin
              for (forvar152 = (1'h0); (forvar152 < (2'h2)); forvar152 = (forvar152 + (1'h1)))
                begin
                  for (forvar153 = (1'h0); (forvar153 < (2'h3)); forvar153 = (forvar153 + (1'h1)))
                    begin
                      reg154 <= reg174;
                    end
                end
              reg155 <= {((~^(wire150 ? (8'ha3) : wire148)) <<< (^~(forvar170 ?
                      reg192 : (8'haa))))};
              for (forvar156 = (1'h0); (forvar156 < (2'h2)); forvar156 = (forvar156 + (1'h1)))
                begin
                  for (forvar157 = (1'h0); (forvar157 < (1'h1)); forvar157 = (forvar157 + (1'h1)))
                    begin
                      reg158 <= $signed(reg167[(1'h1):(1'h1)]);
                      reg159 <= (8'hab);
                      reg160 <= $signed($unsigned($signed(forvar152[(2'h3):(1'h1)])));
                    end
                  for (forvar161 = (1'h0); (forvar161 < (2'h3)); forvar161 = (forvar161 + (1'h1)))
                    begin
                      reg162 <= (&(((forvar176 ?
                          forvar179 : forvar179) >> reg154[(3'h5):(3'h5)]) ^ (forvar151[(3'h5):(2'h2)] ?
                          wire150 : wire146)));
                    end
                  reg163 <= (+{reg166});
                  for (forvar164 = (1'h0); (forvar164 < (2'h3)); forvar164 = (forvar164 + (1'h1)))
                    begin
                      reg165 <= forvar157[(2'h3):(1'h1)];
                      reg166 <= $unsigned($unsigned(((wire150 | reg164) < (forvar170 ?
                          reg182 : (8'hb1)))));
                      reg167 <= {(reg178[(3'h5):(2'h3)] >> (~|(|forvar157)))};
                      reg168 <= {(((~^reg187) ?
                                  wire148[(3'h5):(2'h2)] : (forvar151 ?
                                      reg187 : forvar161)) ?
                              ($signed(reg187) ?
                                  (reg154 >> reg180) : (reg183 && reg154)) : (reg166 ?
                                  ((8'hb0) ?
                                      reg157 : reg169) : $unsigned((8'hb0))))};
                    end
                end
              for (forvar169 = (1'h0); (forvar169 < (2'h3)); forvar169 = (forvar169 + (1'h1)))
                begin
                  for (forvar170 = (1'h0); (forvar170 < (1'h0)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= reg163[(3'h5):(3'h5)];
                    end
                  for (forvar172 = (1'h0); (forvar172 < (1'h1)); forvar172 = (forvar172 + (1'h1)))
                    begin
                      reg173 <= $unsigned($signed(({reg188} + $signed(forvar170))));
                    end
                end
            end
          for (forvar196 = (1'h0); (forvar196 < (2'h3)); forvar196 = (forvar196 + (1'h1)))
            begin
              for (forvar197 = (1'h0); (forvar197 < (2'h2)); forvar197 = (forvar197 + (1'h1)))
                begin
                  for (forvar198 = (1'h0); (forvar198 < (2'h2)); forvar198 = (forvar198 + (1'h1)))
                    begin
                      reg199 <= (forvar151 ?
                          $signed(((~&reg164) ?
                              (forvar172 > reg193) : ((8'h9c) ^ forvar191))) : (~^{$unsigned(forvar169)}));
                      reg200 <= $unsigned((^{reg171}));
                      reg201 <= (((((8'hb2) ?
                          (8'ha5) : reg193) || (~&(8'hb5))) == $unsigned(reg168[(1'h0):(1'h0)])) ^ $signed((&forvar198[(3'h5):(1'h0)])));
                      reg202 <= ({($signed(forvar172) ? {reg177} : reg167)} ?
                          (8'h9e) : $signed(reg201));
                    end
                  reg203 <= forvar152;
                  reg204 <= reg202;
                end
              for (forvar205 = (1'h0); (forvar205 < (1'h1)); forvar205 = (forvar205 + (1'h1)))
                begin
                  for (forvar206 = (1'h0); (forvar206 < (2'h2)); forvar206 = (forvar206 + (1'h1)))
                    begin
                      reg207 <= $unsigned(($unsigned($signed(reg174)) ?
                          (8'haa) : $signed(wire147[(2'h3):(1'h1)])));
                    end
                end
              for (forvar208 = (1'h0); (forvar208 < (1'h0)); forvar208 = (forvar208 + (1'h1)))
                begin
                  if ((((reg172 * (reg187 ?
                      reg194 : (8'ha1))) || forvar161) + wire146))
                    begin
                      reg209 <= ($unsigned(forvar161) ? (8'hb0) : reg195);
                      reg210 <= ((forvar176 ^ reg201[(2'h2):(1'h1)]) ?
                          reg190 : reg160);
                    end
                  else
                    begin
                      reg209 <= ((($unsigned((8'hb5)) ~^ (~forvar196)) ?
                          $signed((|forvar205)) : $unsigned(((8'had) ?
                              wire147 : reg175))) ~^ reg207);
                      reg210 <= {(forvar197[(4'h8):(1'h0)] ?
                              (!(+reg160)) : forvar169)};
                    end
                  if (reg168[(1'h1):(1'h0)])
                    begin
                      reg211 <= ((reg204[(4'hd):(3'h5)] - {forvar208[(3'h6):(3'h6)]}) ?
                          (-forvar170[(1'h1):(1'h0)]) : (reg190[(2'h3):(2'h2)] >>> $unsigned({forvar161})));
                      reg212 <= (forvar161 | ({$signed(forvar198)} ?
                          wire147 : reg209));
                    end
                  else
                    begin
                      reg211 <= ({(~|(8'hb4))} ?
                          (~^({reg189} <<< ((8'hb9) ?
                              reg209 : forvar151))) : ((reg207 ?
                                  $signed(reg165) : (&reg167)) ?
                              {(^~forvar198)} : $signed((reg183 ?
                                  (8'hb1) : forvar164))));
                      reg212 <= ((8'had) ?
                          ($unsigned((reg209 ?
                              wire150 : forvar169)) >> wire147) : reg171[(4'hb):(2'h2)]);
                      reg213 <= $unsigned({reg168[(2'h2):(1'h0)]});
                    end
                  reg214 <= (^~$signed(reg168));
                end
            end
        end
      reg215 <= reg173;
      for (forvar216 = (1'h0); (forvar216 < (1'h1)); forvar216 = (forvar216 + (1'h1)))
        begin
          for (forvar217 = (1'h0); (forvar217 < (1'h1)); forvar217 = (forvar217 + (1'h1)))
            begin
              for (forvar218 = (1'h0); (forvar218 < (2'h2)); forvar218 = (forvar218 + (1'h1)))
                begin
                  if (($signed((~&reg153[(2'h3):(1'h0)])) ?
                      reg159 : {(|(~^forvar152))}))
                    begin
                      reg219 <= $unsigned(({(8'ha0)} ?
                          {(^wire148)} : $unsigned($signed((8'hb5)))));
                      reg220 <= forvar172[(1'h0):(1'h0)];
                      reg221 <= $unsigned((reg165 ?
                          (-forvar168[(3'h4):(3'h4)]) : (~^(|wire149))));
                      reg222 <= reg173[(3'h7):(2'h3)];
                    end
                  else
                    begin
                      reg219 <= (~($unsigned(reg210) ?
                          ($signed(forvar218) && (reg195 ?
                              reg165 : forvar217)) : ((reg209 ^~ forvar172) ?
                              wire149[(2'h3):(2'h3)] : (-forvar153))));
                    end
                end
            end
          reg223 <= ((forvar170[(1'h0):(1'h0)] ?
                  $signed(reg182) : $unsigned((reg190 ? reg162 : forvar176))) ?
              (+$unsigned($unsigned(forvar164))) : {((+forvar205) ?
                      (+forvar161) : reg186[(1'h1):(1'h0)])});
        end
    end
  assign wire224 = (&reg188[(4'hf):(3'h5)]);
  assign wire225 = (($unsigned((8'h9e)) ?
                           ($unsigned(reg178) + {reg164}) : ($unsigned(reg213) << forvar196[(2'h3):(2'h2)])) ?
                       $signed($signed({reg204})) : (({reg193} ?
                               reg171 : $unsigned(reg189)) ?
                           reg222 : ($signed(reg186) ^ (|reg195))));
  assign wire226 = $signed((-(~&$unsigned(forvar216))));
  module227 modinst286 (.wire230(reg193), .wire228(reg195), .y(wire285), .clk(clk), .wire231(reg189), .wire229(wire146));
  module287 modinst582 (wire581, clk, wire150, reg192, reg189, forvar172, reg220);
  assign wire583 = (((8'hb9) + {$signed(forvar196)}) ~^ reg164[(3'h4):(1'h0)]);
  module584 modinst2674 (.wire589(wire581), .wire586(forvar170), .wire587(reg193), .wire585(reg185), .wire588(reg190), .y(wire2673), .clk(clk));
  assign wire2675 = forvar151[(4'hd):(4'hb)];
  always
    @(posedge clk) begin
      if (reg160[(3'h4):(1'h0)])
        begin
          for (forvar2676 = (1'h0); (forvar2676 < (1'h0)); forvar2676 = (forvar2676 + (1'h1)))
            begin
              for (forvar2677 = (1'h0); (forvar2677 < (2'h2)); forvar2677 = (forvar2677 + (1'h1)))
                begin
                  for (forvar2678 = (1'h0); (forvar2678 < (2'h3)); forvar2678 = (forvar2678 + (1'h1)))
                    begin
                      reg2679 <= reg204;
                      reg2680 <= (((8'ha4) + {reg160[(4'hb):(3'h5)]}) <= (|$unsigned(reg174[(3'h4):(3'h4)])));
                    end
                  for (forvar2681 = (1'h0); (forvar2681 < (2'h3)); forvar2681 = (forvar2681 + (1'h1)))
                    begin
                      reg2682 <= (^~{(~&{reg154})});
                    end
                  for (forvar2683 = (1'h0); (forvar2683 < (2'h2)); forvar2683 = (forvar2683 + (1'h1)))
                    begin
                      reg2684 <= $unsigned($unsigned((reg177[(2'h2):(1'h0)] - (forvar164 ?
                          reg181 : (8'hb3)))));
                      reg2685 <= reg193;
                      reg2686 <= {(!(&forvar217[(1'h1):(1'h1)]))};
                      reg2687 <= $unsigned(reg2682[(2'h2):(1'h1)]);
                    end
                end
            end
          if ($unsigned({$unsigned((8'ha1))}))
            begin
              for (forvar2688 = (1'h0); (forvar2688 < (2'h2)); forvar2688 = (forvar2688 + (1'h1)))
                begin
                  if (reg220)
                    begin
                      reg2689 <= forvar218[(3'h6):(2'h2)];
                      reg2690 <= reg203[(4'ha):(4'ha)];
                      reg2691 <= {reg174};
                    end
                  else
                    begin
                      reg2689 <= $signed((8'hb9));
                      reg2690 <= (((&{forvar156}) >>> (^(reg187 ?
                              reg202 : forvar217))) ?
                          reg183[(4'hb):(3'h7)] : (((-forvar196) ?
                              forvar196 : forvar2676[(1'h1):(1'h1)]) && $unsigned((forvar2681 * reg207))));
                    end
                  for (forvar2692 = (1'h0); (forvar2692 < (2'h2)); forvar2692 = (forvar2692 + (1'h1)))
                    begin
                      reg2693 <= $unsigned($unsigned($signed((wire148 ^~ reg183))));
                    end
                  if (($signed($signed($signed(forvar196))) ?
                      $signed((~|forvar172)) : {reg2680}))
                    begin
                      reg2694 <= {forvar218[(1'h0):(1'h0)]};
                      reg2695 <= wire583[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2694 <= reg166;
                      reg2695 <= forvar205;
                      reg2696 <= ((forvar191 * wire146[(2'h2):(2'h2)]) ^~ {(!forvar184)});
                    end
                end
            end
          else
            begin
              for (forvar2688 = (1'h0); (forvar2688 < (2'h3)); forvar2688 = (forvar2688 + (1'h1)))
                begin
                  for (forvar2689 = (1'h0); (forvar2689 < (2'h2)); forvar2689 = (forvar2689 + (1'h1)))
                    begin
                      reg2690 <= $unsigned($signed(({reg2684} + reg194)));
                      reg2691 <= (+reg211[(4'ha):(2'h3)]);
                      reg2692 <= ({reg169[(4'hd):(2'h2)]} ^ (+(forvar2676 ?
                          (!(8'h9e)) : $signed(reg189))));
                      reg2693 <= (|$signed(reg174[(3'h5):(1'h1)]));
                    end
                  reg2694 <= (forvar2678[(3'h5):(1'h0)] & forvar198[(3'h4):(2'h2)]);
                  for (forvar2695 = (1'h0); (forvar2695 < (1'h0)); forvar2695 = (forvar2695 + (1'h1)))
                    begin
                      reg2696 <= (wire2675 ^ forvar2676[(3'h4):(2'h3)]);
                      reg2697 <= (reg210[(4'he):(3'h7)] >= $signed((~^(~|reg203))));
                    end
                  if ($unsigned(($signed((reg2696 >>> (8'hb2))) > $signed($unsigned(wire146)))))
                    begin
                      reg2698 <= ({reg160} ?
                          reg212 : {(+forvar205[(1'h0):(1'h0)])});
                      reg2699 <= $signed(reg212);
                    end
                  else
                    begin
                      reg2698 <= ((~^forvar161) + (~^forvar164));
                      reg2699 <= ((forvar196[(2'h2):(1'h0)] ?
                              reg163 : ((+reg183) ^~ $signed(forvar170))) ?
                          $unsigned({forvar206}) : $unsigned(reg172));
                      reg2700 <= (~^reg161);
                      reg2701 <= $signed(($signed(((8'hab) ?
                              wire147 : reg192)) ?
                          $unsigned((&reg2695)) : $unsigned((reg155 & wire225))));
                    end
                end
            end
        end
      else
        begin
          if (((^~$unsigned($unsigned(forvar2689))) ?
              ((|wire226) ?
                  ((reg207 >= wire149) ? {reg212} : (&reg212)) : (((8'hb5) ?
                          reg183 : reg209) ?
                      $unsigned(reg165) : reg192[(4'ha):(1'h0)])) : $signed(forvar2681[(4'he):(3'h5)])))
            begin
              for (forvar2676 = (1'h0); (forvar2676 < (1'h1)); forvar2676 = (forvar2676 + (1'h1)))
                begin
                  for (forvar2677 = (1'h0); (forvar2677 < (1'h1)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= (reg2696[(1'h0):(1'h0)] ?
                          $unsigned((~reg2700)) : forvar196[(3'h4):(2'h3)]);
                      reg2679 <= reg210;
                      reg2680 <= $signed(($unsigned({(8'hb8)}) ?
                          ((&(8'ha1)) ?
                              forvar205[(2'h3):(2'h3)] : $signed(reg207)) : $unsigned({(8'h9c)})));
                      reg2681 <= (reg2685 | $signed((&(reg194 ?
                          forvar170 : forvar2695))));
                    end
                  for (forvar2682 = (1'h0); (forvar2682 < (1'h0)); forvar2682 = (forvar2682 + (1'h1)))
                    begin
                      reg2683 <= {((reg204 ?
                                  reg2693[(4'hb):(1'h1)] : (wire146 ?
                                      reg182 : (8'h9e))) ?
                              $unsigned($unsigned(reg175)) : forvar156)};
                      reg2684 <= ($signed((+{(8'hb2)})) ^~ ($signed(reg214) ?
                          {(reg213 - forvar2689)} : (~|$unsigned((8'had)))));
                      reg2685 <= (~reg2694);
                    end
                  reg2686 <= ((+{$signed(reg202)}) ?
                      ($unsigned((&(8'hb7))) >= $unsigned(forvar152[(4'h8):(3'h5)])) : forvar184[(4'hd):(3'h4)]);
                end
              if (($unsigned({forvar2678}) ?
                  (^~wire581[(4'hc):(4'hc)]) : (wire285 ?
                      forvar179 : $unsigned(reg172[(3'h4):(3'h4)]))))
                begin
                  if (forvar198)
                    begin
                      reg2687 <= reg161[(2'h3):(1'h1)];
                      reg2688 <= (((+reg190) && $unsigned($signed(reg166))) <= reg162[(4'hd):(4'hc)]);
                      reg2689 <= ($signed({((8'hb6) ? reg171 : reg200)}) ?
                          ($unsigned((&reg215)) ?
                              reg2679[(1'h1):(1'h1)] : $signed($unsigned(reg214))) : $unsigned(($signed(reg173) || reg222[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg2687 <= $unsigned({(^~$unsigned(reg154))});
                      reg2688 <= (~reg220);
                    end
                  if ((($signed((reg220 & wire146)) >>> {(8'hae)}) ?
                      (~(~(~^forvar2677))) : (reg2681 ?
                          $unsigned((reg193 << forvar206)) : (~&reg2690))))
                    begin
                      reg2690 <= (~|(^~reg2691));
                      reg2691 <= ((forvar169 | reg2700) | (($signed(reg2688) ?
                          forvar161[(2'h3):(2'h2)] : (~&forvar2678)) == ((~|reg169) && reg203[(4'hb):(3'h6)])));
                      reg2692 <= $signed($unsigned(reg177));
                      reg2693 <= forvar216;
                    end
                  else
                    begin
                      reg2690 <= $unsigned(forvar2689);
                    end
                  reg2694 <= $unsigned($unsigned(((reg2680 ? reg167 : reg173) ?
                      reg167 : (^reg164))));
                end
              else
                begin
                  for (forvar2687 = (1'h0); (forvar2687 < (2'h2)); forvar2687 = (forvar2687 + (1'h1)))
                    begin
                      reg2688 <= ($signed((reg2690[(1'h0):(1'h0)] ?
                          (reg173 == reg154) : (reg175 ?
                              (8'had) : (8'had)))) ^~ $signed((reg2684[(3'h5):(2'h2)] ~^ forvar152)));
                      reg2689 <= ($unsigned({reg199[(1'h1):(1'h0)]}) * reg220[(2'h2):(1'h1)]);
                      reg2690 <= reg203;
                    end
                end
              for (forvar2695 = (1'h0); (forvar2695 < (2'h3)); forvar2695 = (forvar2695 + (1'h1)))
                begin
                  if ((~&reg194))
                    begin
                      reg2696 <= ($signed((reg188[(4'ha):(1'h0)] ?
                          (forvar217 ?
                              (8'hac) : (8'hb7)) : $signed((8'hb7)))) - (8'had));
                      reg2697 <= (((|(^reg180)) >>> $signed((~|reg161))) ?
                          reg210 : (((~^(8'hae)) < (reg212 ?
                                  reg181 : forvar2695)) ?
                              (8'ha3) : $signed($unsigned(wire226))));
                    end
                  else
                    begin
                      reg2696 <= reg2682;
                    end
                  if ($signed((^$signed((forvar208 < reg207)))))
                    begin
                      reg2698 <= $signed(reg201);
                    end
                  else
                    begin
                      reg2698 <= forvar2678;
                      reg2699 <= $unsigned((+reg2683[(2'h2):(1'h0)]));
                      reg2700 <= reg173;
                      reg2701 <= ((~&(reg161[(2'h3):(1'h0)] <<< (reg2689 ?
                          reg164 : reg220))) ~^ $unsigned((~{reg214})));
                    end
                  for (forvar2702 = (1'h0); (forvar2702 < (1'h0)); forvar2702 = (forvar2702 + (1'h1)))
                    begin
                      reg2703 <= (|$unsigned($signed($signed((8'had)))));
                      reg2704 <= {($unsigned($signed(reg164)) < $signed($unsigned(reg207)))};
                      reg2705 <= $unsigned(reg207[(2'h3):(1'h1)]);
                      reg2706 <= (reg215 ?
                          ($signed($signed(reg158)) ?
                              (~|(&(8'h9f))) : (8'h9d)) : forvar2682);
                    end
                end
              reg2707 <= (forvar216 >= (($unsigned(forvar179) | {reg210}) ?
                  reg158 : (reg2695 ?
                      $signed(reg202) : (reg166 ? reg187 : reg188))));
            end
          else
            begin
              if ((~|(~|((forvar152 <= reg2692) ^~ reg202[(3'h7):(3'h6)]))))
                begin
                  reg2676 <= {($signed($signed(reg2689)) == (^(reg183 ?
                          reg210 : reg185)))};
                  for (forvar2677 = (1'h0); (forvar2677 < (1'h0)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= $signed($signed($unsigned({(8'hb9)})));
                    end
                  if (reg2700)
                    begin
                      reg2679 <= (((~&(reg200 > reg165)) ?
                              $unsigned(reg2676[(1'h0):(1'h0)]) : {(reg203 ?
                                      reg166 : (8'hb8))}) ?
                          $signed($signed((forvar206 + reg2686))) : {$signed(((8'ha1) ?
                                  reg223 : forvar2682))});
                      reg2680 <= (forvar151 <<< reg178[(3'h5):(2'h2)]);
                      reg2681 <= $unsigned((reg180 ^~ (reg200 ?
                          $signed(reg159) : reg209)));
                    end
                  else
                    begin
                      reg2679 <= (~(&reg212));
                      reg2680 <= {(((|(8'ha2)) ?
                              (-reg2689) : (-reg187)) != ((reg183 || forvar2695) >> (reg166 | wire146)))};
                      reg2681 <= $unsigned(reg159);
                    end
                end
              else
                begin
                  reg2676 <= (&wire149[(4'he):(1'h1)]);
                  for (forvar2677 = (1'h0); (forvar2677 < (2'h2)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= forvar2682;
                      reg2679 <= reg220;
                      reg2680 <= reg2705;
                      reg2681 <= reg171;
                    end
                  if (((({(8'haa)} ? reg2688[(1'h0):(1'h0)] : forvar2681) ?
                      reg167 : $unsigned($unsigned(reg209))) != ((|forvar2688[(1'h0):(1'h0)]) ?
                      reg175[(2'h3):(2'h3)] : ((forvar2688 ^ forvar170) ?
                          wire285 : $signed((8'hb7))))))
                    begin
                      reg2682 <= reg213;
                    end
                  else
                    begin
                      reg2682 <= $unsigned($unsigned(forvar2676[(1'h1):(1'h0)]));
                      reg2683 <= wire583[(2'h3):(1'h1)];
                      reg2684 <= (wire146[(2'h3):(2'h2)] ?
                          $unsigned((~{forvar206})) : ((~&$signed(reg154)) ?
                              {(~|reg203)} : reg210));
                      reg2685 <= reg200[(1'h1):(1'h0)];
                    end
                end
              for (forvar2686 = (1'h0); (forvar2686 < (2'h3)); forvar2686 = (forvar2686 + (1'h1)))
                begin
                  for (forvar2687 = (1'h0); (forvar2687 < (2'h3)); forvar2687 = (forvar2687 + (1'h1)))
                    begin
                      reg2688 <= (~|(|reg209));
                    end
                  for (forvar2689 = (1'h0); (forvar2689 < (2'h3)); forvar2689 = (forvar2689 + (1'h1)))
                    begin
                      reg2690 <= $signed(($signed($unsigned((8'ha9))) <= $unsigned(reg201[(1'h1):(1'h1)])));
                    end
                  reg2691 <= (reg163[(2'h2):(1'h1)] * (reg192 & ($unsigned(forvar217) && ((8'hb5) <<< reg214))));
                  for (forvar2692 = (1'h0); (forvar2692 < (1'h1)); forvar2692 = (forvar2692 + (1'h1)))
                    begin
                      reg2693 <= $unsigned((|(^~(reg167 ?
                          reg178 : forvar197))));
                      reg2694 <= reg2696[(4'h9):(3'h6)];
                      reg2695 <= forvar2688;
                    end
                end
              reg2696 <= reg222[(2'h3):(2'h3)];
            end
          if ($signed(forvar197[(4'h8):(3'h5)]))
            begin
              for (forvar2708 = (1'h0); (forvar2708 < (2'h3)); forvar2708 = (forvar2708 + (1'h1)))
                begin
                  if ($unsigned(forvar179[(2'h2):(1'h0)]))
                    begin
                      reg2709 <= (8'ha3);
                      reg2710 <= reg2681;
                      reg2711 <= reg213;
                      reg2712 <= reg200[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg2709 <= reg2711;
                      reg2710 <= ((((~&reg220) ?
                              (~^reg156) : wire150) | $unsigned((reg180 ^~ wire2673))) ?
                          {reg153} : (forvar2688[(2'h3):(2'h3)] ?
                              $unsigned((8'hab)) : (forvar2708[(4'h9):(4'h9)] ?
                                  reg2695 : $unsigned(reg2710))));
                      reg2711 <= (reg2681[(3'h5):(2'h3)] ?
                          (reg163[(4'ha):(4'h8)] >= ((|reg212) ?
                              (!forvar196) : {reg199})) : $unsigned($signed($signed((8'hb7)))));
                    end
                  if ((reg2709 ?
                      $unsigned((&(reg2679 * reg2710))) : reg204[(3'h4):(1'h0)]))
                    begin
                      reg2713 <= {$signed(((~^reg159) <<< $unsigned(forvar170)))};
                      reg2714 <= wire225;
                      reg2715 <= ($signed({reg186[(4'h9):(3'h4)]}) * ((!$unsigned(reg2698)) && reg2687));
                      reg2716 <= (!($signed((forvar205 ?
                          reg213 : (8'h9f))) >= ((reg2686 ?
                          (8'hb1) : forvar206) >= (~(8'hb0)))));
                    end
                  else
                    begin
                      reg2713 <= ((($signed(forvar218) ?
                                  $unsigned(reg189) : (^~reg2710)) ?
                              ($signed(reg160) != (reg182 ?
                                  wire583 : reg174)) : reg2690) ?
                          forvar206[(2'h3):(1'h1)] : forvar2681);
                      reg2714 <= ((8'h9d) << (~reg2690[(2'h3):(2'h3)]));
                    end
                end
              reg2717 <= (~|$signed((+{forvar2687})));
              if (((reg211 ? {(reg2713 & reg2692)} : forvar2683) ?
                  reg192[(2'h2):(1'h1)] : (reg2681 ?
                      $signed($signed(reg2712)) : ($unsigned(reg193) ?
                          {wire2675} : (reg159 ? (8'haf) : reg2716)))))
                begin
                  if (($unsigned(({(8'hac)} ?
                      (reg2693 ?
                          forvar2688 : reg219) : (reg220 && (8'hb4)))) ~^ $signed((+reg199))))
                    begin
                      reg2718 <= {reg2685};
                      reg2719 <= reg2697;
                      reg2720 <= (($signed(wire581) <<< (!(forvar2681 ^~ reg2712))) >>> ((-(reg2709 ^ reg158)) - $unsigned((~reg161))));
                      reg2721 <= ((((reg154 ? reg175 : reg168) ?
                          $unsigned(forvar2683) : forvar197) | $signed($unsigned(wire225))) <<< $signed(forvar2683[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg2718 <= reg2700[(3'h4):(1'h0)];
                      reg2719 <= forvar153[(4'h9):(1'h1)];
                    end
                  if (((~&{$signed((8'h9e))}) ?
                      ((wire224 ? (^(8'hb9)) : (~&reg2703)) ?
                          ((reg174 ? forvar2702 : reg212) ?
                              $signed(reg2701) : $signed(forvar216)) : (reg2690[(2'h2):(2'h2)] ?
                              $signed(reg181) : (wire285 >> reg166))) : forvar2683[(1'h1):(1'h1)]))
                    begin
                      reg2722 <= (&((8'hba) ?
                          reg166 : $unsigned($signed((8'hb0)))));
                      reg2723 <= $signed(reg192[(4'hb):(3'h4)]);
                    end
                  else
                    begin
                      reg2722 <= ($unsigned((8'ha4)) ?
                          $unsigned(wire224) : {reg2676[(2'h3):(1'h0)]});
                      reg2723 <= (-(($unsigned(reg171) ~^ forvar2688[(4'h8):(2'h3)]) <= reg2689[(2'h2):(1'h0)]));
                      reg2724 <= (~^$unsigned($signed(reg2692)));
                    end
                  reg2725 <= (~reg158);
                end
              else
                begin
                  reg2718 <= ((forvar196[(2'h2):(1'h0)] ?
                      reg168 : forvar153) >> $signed($signed((reg2699 ^ reg2698))));
                  for (forvar2719 = (1'h0); (forvar2719 < (2'h3)); forvar2719 = (forvar2719 + (1'h1)))
                    begin
                      reg2720 <= {$unsigned(forvar157[(2'h2):(2'h2)])};
                      reg2721 <= $unsigned($unsigned(reg2692[(1'h1):(1'h0)]));
                      reg2722 <= $unsigned({(8'ha3)});
                      reg2723 <= forvar218[(2'h2):(1'h1)];
                    end
                  reg2724 <= {{$unsigned((8'ha5))}};
                  reg2725 <= ((((reg221 ? reg214 : reg156) ?
                          $signed((8'hb0)) : reg213) ?
                      (^~(!reg202)) : ((reg203 ? reg154 : wire149) ?
                          forvar218 : $unsigned(reg163))) >= forvar184);
                end
              for (forvar2726 = (1'h0); (forvar2726 < (2'h3)); forvar2726 = (forvar2726 + (1'h1)))
                begin
                  if (reg159)
                    begin
                      reg2727 <= (forvar2688 >> reg162[(4'hd):(1'h1)]);
                      reg2728 <= (~{forvar156[(4'h9):(4'h8)]});
                    end
                  else
                    begin
                      reg2727 <= {forvar196[(3'h4):(1'h1)]};
                      reg2728 <= ($signed(($signed((8'hb8)) ?
                          $signed(forvar184) : reg169[(4'h8):(3'h6)])) == {$unsigned($signed(reg207))});
                      reg2729 <= {(^~{$unsigned((8'ha9))})};
                    end
                  reg2730 <= reg214[(1'h1):(1'h1)];
                  reg2731 <= ((8'hb5) & {forvar157[(1'h0):(1'h0)]});
                end
            end
          else
            begin
              for (forvar2708 = (1'h0); (forvar2708 < (2'h2)); forvar2708 = (forvar2708 + (1'h1)))
                begin
                  if ((8'hab))
                    begin
                      reg2709 <= (~reg2717[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg2709 <= (^~reg2676[(2'h2):(1'h0)]);
                    end
                end
              for (forvar2710 = (1'h0); (forvar2710 < (1'h1)); forvar2710 = (forvar2710 + (1'h1)))
                begin
                  if (reg156)
                    begin
                      reg2711 <= $unsigned((~^(-$signed((8'haf)))));
                      reg2712 <= $unsigned($unsigned(reg168[(1'h1):(1'h0)]));
                      reg2713 <= (8'hb9);
                      reg2714 <= (((!(-forvar161)) - (reg168 ?
                          (|forvar152) : $unsigned(reg166))) > $signed(reg2701[(4'hb):(1'h1)]));
                    end
                  else
                    begin
                      reg2711 <= $signed(((^~reg163[(4'h8):(1'h0)]) ?
                          ((8'hb5) ?
                              (8'haf) : $unsigned(reg214)) : $unsigned($signed(reg177))));
                      reg2712 <= (({(reg2705 != reg195)} ?
                          {$signed(reg221)} : forvar168[(3'h4):(1'h0)]) || reg2689);
                    end
                  for (forvar2715 = (1'h0); (forvar2715 < (2'h3)); forvar2715 = (forvar2715 + (1'h1)))
                    begin
                      reg2716 <= (8'had);
                      reg2717 <= reg172[(2'h3):(2'h3)];
                    end
                end
              for (forvar2718 = (1'h0); (forvar2718 < (2'h2)); forvar2718 = (forvar2718 + (1'h1)))
                begin
                  for (forvar2719 = (1'h0); (forvar2719 < (2'h2)); forvar2719 = (forvar2719 + (1'h1)))
                    begin
                      reg2720 <= forvar152;
                      reg2721 <= ($signed($signed({reg220})) <= (^forvar179));
                    end
                  reg2722 <= (~^forvar161[(2'h2):(1'h1)]);
                end
              for (forvar2723 = (1'h0); (forvar2723 < (2'h3)); forvar2723 = (forvar2723 + (1'h1)))
                begin
                  reg2724 <= (+$signed(((forvar161 ~^ reg195) - $unsigned(reg160))));
                  if ((^~$unsigned((8'haf))))
                    begin
                      reg2725 <= {reg162};
                      reg2726 <= forvar2686;
                      reg2727 <= (!$unsigned((~$signed(wire583))));
                      reg2728 <= {$signed((wire148 != forvar2683[(2'h2):(1'h1)]))};
                    end
                  else
                    begin
                      reg2725 <= ($signed(reg2729[(3'h4):(3'h4)]) || reg2704[(2'h3):(1'h1)]);
                      reg2726 <= ({$unsigned({(8'h9f)})} & $signed(reg2715[(2'h3):(1'h1)]));
                      reg2727 <= $unsigned((reg2714[(1'h0):(1'h0)] ?
                          reg174 : (reg2729[(2'h3):(1'h0)] >> reg2707[(2'h2):(1'h1)])));
                      reg2728 <= {reg2687};
                    end
                  reg2729 <= wire225[(4'ha):(4'h8)];
                end
            end
          if (((reg2714 ?
                  $unsigned($signed(reg177)) : $signed(reg185[(3'h7):(2'h2)])) ?
              reg2698[(2'h2):(1'h1)] : {(forvar2710 ?
                      (reg190 ? reg181 : reg2723) : (^~reg203))}))
            begin
              reg2732 <= reg2711[(4'ha):(4'ha)];
              for (forvar2733 = (1'h0); (forvar2733 < (1'h0)); forvar2733 = (forvar2733 + (1'h1)))
                begin
                  for (forvar2734 = (1'h0); (forvar2734 < (2'h2)); forvar2734 = (forvar2734 + (1'h1)))
                    begin
                      reg2735 <= reg157[(3'h7):(1'h1)];
                    end
                end
              for (forvar2736 = (1'h0); (forvar2736 < (1'h1)); forvar2736 = (forvar2736 + (1'h1)))
                begin
                  reg2737 <= (reg2725 ?
                      ((|(reg2682 ?
                          reg194 : forvar157)) <<< $signed($unsigned((8'hb9)))) : ($signed($signed(reg213)) ?
                          (reg2728[(3'h6):(3'h5)] | (forvar2726 >= reg194)) : reg2676[(1'h0):(1'h0)]));
                end
            end
          else
            begin
              reg2732 <= reg171;
            end
        end
      for (forvar2738 = (1'h0); (forvar2738 < (1'h1)); forvar2738 = (forvar2738 + (1'h1)))
        begin
          for (forvar2739 = (1'h0); (forvar2739 < (1'h0)); forvar2739 = (forvar2739 + (1'h1)))
            begin
              for (forvar2740 = (1'h0); (forvar2740 < (1'h1)); forvar2740 = (forvar2740 + (1'h1)))
                begin
                  if ((~&$unsigned((forvar205 ?
                      wire224[(3'h7):(3'h6)] : (reg160 ? reg2709 : reg158)))))
                    begin
                      reg2741 <= (!(reg168 ?
                          $signed($unsigned((8'hb9))) : ($signed(forvar2687) & (forvar2677 ?
                              reg2703 : (8'hb3)))));
                      reg2742 <= ($signed($signed($signed((8'ha3)))) + $signed(($signed((8'h9e)) | (wire226 ?
                          reg167 : forvar156))));
                      reg2743 <= $signed((^~(((8'hae) != reg165) ?
                          $unsigned(reg173) : $signed(forvar2734))));
                      reg2744 <= $signed((($signed(reg2680) == (^~forvar151)) ?
                          ($unsigned(reg2718) ?
                              (reg2687 && forvar2687) : $unsigned(reg2728)) : $unsigned((reg2700 ?
                              reg2714 : reg164))));
                    end
                  else
                    begin
                      reg2741 <= forvar2719;
                      reg2742 <= forvar2702[(3'h4):(3'h4)];
                      reg2743 <= $unsigned((((reg2718 ?
                                  forvar2708 : forvar2738) ?
                              reg153[(1'h1):(1'h1)] : (reg2712 ?
                                  (8'ha3) : forvar2734)) ?
                          $unsigned($signed(forvar2736)) : $signed($unsigned(reg2704))));
                    end
                  if (reg201)
                    begin
                      reg2745 <= ((!$signed((reg174 ?
                          reg188 : reg2698))) * (^wire148[(3'h4):(3'h4)]));
                      reg2746 <= (forvar2678[(3'h5):(3'h5)] < $signed($unsigned(reg2691)));
                      reg2747 <= $unsigned($unsigned(forvar2734));
                      reg2748 <= $signed(($unsigned(((8'haf) ?
                              reg207 : reg220)) ?
                          reg2728 : reg181));
                    end
                  else
                    begin
                      reg2745 <= reg2720;
                      reg2746 <= (&(8'hac));
                    end
                  for (forvar2749 = (1'h0); (forvar2749 < (1'h1)); forvar2749 = (forvar2749 + (1'h1)))
                    begin
                      reg2750 <= (~&forvar2739);
                      reg2751 <= ((reg2731[(4'hc):(3'h4)] ?
                          {(reg2685 + (8'hb0))} : ($unsigned(forvar2715) != forvar217[(1'h1):(1'h0)])) + forvar2681);
                      reg2752 <= $unsigned((^((reg2684 ?
                          forvar2708 : forvar2708) >= $unsigned(reg172))));
                    end
                  reg2753 <= (^~reg2703);
                end
              for (forvar2754 = (1'h0); (forvar2754 < (2'h3)); forvar2754 = (forvar2754 + (1'h1)))
                begin
                  for (forvar2755 = (1'h0); (forvar2755 < (1'h0)); forvar2755 = (forvar2755 + (1'h1)))
                    begin
                      reg2756 <= (-({(+reg2679)} & (!(forvar157 < (8'h9e)))));
                    end
                  if ($unsigned($unsigned(forvar184[(2'h3):(2'h3)])))
                    begin
                      reg2757 <= {((8'ha8) || reg200)};
                      reg2758 <= wire149[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg2757 <= ((-(|(reg158 >>> (8'hb7)))) == $unsigned(reg165));
                      reg2758 <= ({((8'ha8) * (forvar2677 >>> reg177))} ?
                          reg2687 : (($unsigned(reg2715) ? reg169 : forvar196) ?
                              ((reg189 ? (8'had) : reg209) ?
                                  (reg200 - (8'ha4)) : reg159) : {reg159[(2'h3):(2'h2)]}));
                      reg2759 <= (~(^reg169[(4'h9):(3'h5)]));
                    end
                  reg2760 <= $unsigned((($signed((8'hb6)) | (reg2732 - reg157)) ?
                      forvar2719[(2'h3):(1'h1)] : $unsigned(reg2726)));
                end
              for (forvar2761 = (1'h0); (forvar2761 < (2'h2)); forvar2761 = (forvar2761 + (1'h1)))
                begin
                  for (forvar2762 = (1'h0); (forvar2762 < (2'h2)); forvar2762 = (forvar2762 + (1'h1)))
                    begin
                      reg2763 <= {$unsigned($signed({wire2673}))};
                    end
                  reg2764 <= $signed((+($unsigned((8'hb4)) >>> (~|reg215))));
                end
              for (forvar2765 = (1'h0); (forvar2765 < (2'h2)); forvar2765 = (forvar2765 + (1'h1)))
                begin
                  if ($signed({$unsigned((~^forvar179))}))
                    begin
                      reg2766 <= $unsigned(reg2757);
                      reg2767 <= ({forvar191[(4'hb):(3'h5)]} == ((&reg195) ?
                          reg185 : (^$signed(forvar198))));
                      reg2768 <= $unsigned($unsigned(reg222));
                      reg2769 <= (($unsigned((~&reg203)) ?
                          reg2737[(2'h2):(1'h0)] : (reg160 ?
                              $unsigned((8'ha4)) : (~^reg2719))) <= $unsigned(reg2690));
                    end
                  else
                    begin
                      reg2766 <= ((8'hb5) ?
                          {reg214[(3'h5):(2'h3)]} : $unsigned(forvar217));
                      reg2767 <= forvar176[(1'h1):(1'h1)];
                      reg2768 <= (reg156[(3'h5):(1'h1)] + $unsigned(reg219));
                    end
                  if ((!$signed(((reg166 ? reg2727 : reg212) ?
                      reg182[(1'h0):(1'h0)] : (reg2735 >>> forvar2733)))))
                    begin
                      reg2770 <= reg2748[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2770 <= forvar164[(4'hb):(4'ha)];
                      reg2771 <= (8'ha5);
                      reg2772 <= (8'hb0);
                    end
                end
            end
          for (forvar2773 = (1'h0); (forvar2773 < (2'h2)); forvar2773 = (forvar2773 + (1'h1)))
            begin
              for (forvar2774 = (1'h0); (forvar2774 < (1'h1)); forvar2774 = (forvar2774 + (1'h1)))
                begin
                  for (forvar2775 = (1'h0); (forvar2775 < (2'h2)); forvar2775 = (forvar2775 + (1'h1)))
                    begin
                      reg2776 <= (!$signed($signed($unsigned((8'ha9)))));
                      reg2777 <= ((+reg174) != reg185);
                      reg2778 <= (forvar2738 ?
                          $unsigned(reg2772[(3'h4):(1'h1)]) : ({(-reg220)} <<< (~^forvar198[(1'h1):(1'h1)])));
                    end
                end
              reg2779 <= ((8'ha6) + (~|({reg2763} != $signed(reg212))));
              for (forvar2780 = (1'h0); (forvar2780 < (2'h2)); forvar2780 = (forvar2780 + (1'h1)))
                begin
                  for (forvar2781 = (1'h0); (forvar2781 < (1'h0)); forvar2781 = (forvar2781 + (1'h1)))
                    begin
                      reg2782 <= $unsigned((reg2720[(2'h3):(2'h2)] + (reg2753 && (reg203 && reg220))));
                      reg2783 <= (&(8'hb7));
                    end
                end
            end
          for (forvar2784 = (1'h0); (forvar2784 < (1'h0)); forvar2784 = (forvar2784 + (1'h1)))
            begin
              for (forvar2785 = (1'h0); (forvar2785 < (2'h2)); forvar2785 = (forvar2785 + (1'h1)))
                begin
                  for (forvar2786 = (1'h0); (forvar2786 < (2'h3)); forvar2786 = (forvar2786 + (1'h1)))
                    begin
                      reg2787 <= forvar169;
                      reg2788 <= $unsigned((($signed(forvar2734) ^~ (&forvar169)) * ({reg2684} ?
                          reg2758[(4'ha):(4'h9)] : (reg2763 ?
                              reg203 : reg207))));
                    end
                  for (forvar2789 = (1'h0); (forvar2789 < (1'h0)); forvar2789 = (forvar2789 + (1'h1)))
                    begin
                      reg2790 <= $signed($signed(((~(8'h9c)) + $unsigned(forvar156))));
                      reg2791 <= reg2769;
                      reg2792 <= (^~reg207[(3'h5):(1'h1)]);
                    end
                end
            end
          if (reg2745[(3'h5):(3'h4)])
            begin
              for (forvar2793 = (1'h0); (forvar2793 < (2'h2)); forvar2793 = (forvar2793 + (1'h1)))
                begin
                  for (forvar2794 = (1'h0); (forvar2794 < (2'h2)); forvar2794 = (forvar2794 + (1'h1)))
                    begin
                      reg2795 <= ({$unsigned(forvar2686[(4'ha):(3'h4)])} ?
                          (+wire150[(1'h1):(1'h1)]) : reg202);
                      reg2796 <= $signed($unsigned(wire226[(1'h0):(1'h0)]));
                      reg2797 <= reg2720[(3'h7):(3'h4)];
                    end
                  if ($unsigned(((((8'ha4) ^ reg2725) ?
                          ((8'ha7) ?
                              reg2790 : (8'ha2)) : forvar151[(4'he):(3'h7)]) ?
                      (~|$unsigned(reg2704)) : (+$signed((8'ha5))))))
                    begin
                      reg2798 <= wire226[(3'h7):(1'h0)];
                      reg2799 <= (8'hab);
                      reg2800 <= $signed((~|reg2747));
                    end
                  else
                    begin
                      reg2798 <= ((((^~reg2776) >>> $signed((8'ha6))) ?
                              $signed((!forvar2683)) : {forvar2755}) ?
                          (reg2691 ?
                              ($unsigned(reg166) ?
                                  $signed(reg180) : (reg199 + wire150)) : $unsigned((~^reg178))) : (((reg155 && reg2701) << (reg2783 << (8'ha7))) - $signed($unsigned(reg2681))));
                      reg2799 <= forvar2784;
                    end
                end
              reg2801 <= {(reg2711 ?
                      ((-(8'ha7)) + (wire224 ?
                          (8'ha2) : wire147)) : $signed($signed(reg2716)))};
              if ($unsigned($signed(wire149[(3'h4):(1'h0)])))
                begin
                  if (forvar216)
                    begin
                      reg2802 <= $unsigned(forvar2765);
                      reg2803 <= forvar205;
                    end
                  else
                    begin
                      reg2802 <= ($signed($signed($unsigned(reg2778))) ?
                          {((-reg2758) ?
                                  {reg203} : $signed(reg166))} : $signed((forvar179 * $unsigned(wire226))));
                      reg2803 <= ($unsigned($unsigned($unsigned(reg2719))) ?
                          (^({reg2714} >> $unsigned((8'ha4)))) : ((~|$signed(reg2741)) ?
                              reg213[(3'h6):(1'h0)] : ((~reg2680) ?
                                  reg2730 : (8'ha0))));
                    end
                end
              else
                begin
                  for (forvar2802 = (1'h0); (forvar2802 < (1'h0)); forvar2802 = (forvar2802 + (1'h1)))
                    begin
                      reg2803 <= ((&$signed(reg2722[(2'h3):(1'h1)])) ?
                          $unsigned($signed(reg2797[(3'h4):(1'h1)])) : forvar2755);
                    end
                  for (forvar2804 = (1'h0); (forvar2804 < (2'h2)); forvar2804 = (forvar2804 + (1'h1)))
                    begin
                      reg2805 <= {{(reg2787 ? (~|reg2710) : (^forvar2761))}};
                      reg2806 <= wire226[(4'h8):(2'h3)];
                      reg2807 <= ((8'ha8) ? {reg2751} : reg2692[(3'h5):(1'h0)]);
                    end
                  if ({(((reg160 >> wire285) ?
                          reg2678 : (~|(8'hb3))) >> $signed({(8'hb3)}))})
                    begin
                      reg2808 <= $unsigned($signed(((forvar2784 >>> reg2796) ?
                          $unsigned(reg2678) : (~forvar2695))));
                      reg2809 <= reg2682[(1'h0):(1'h0)];
                      reg2810 <= forvar2762;
                    end
                  else
                    begin
                      reg2808 <= ((($unsigned(reg2801) || ((8'ha0) ?
                                  reg2690 : reg2741)) ?
                              reg2730[(4'hb):(4'hb)] : (|$unsigned(reg2799))) ?
                          (-((reg223 != reg2709) ?
                              reg211[(1'h0):(1'h0)] : (reg178 <= (8'hb8)))) : (({forvar2785} ?
                                  (+forvar2738) : ((8'ha0) ?
                                      forvar2762 : (8'hac))) ?
                              reg2756[(3'h7):(1'h0)] : ((reg2687 - reg2747) ~^ wire150)));
                      reg2809 <= forvar191;
                      reg2810 <= ((reg187 ^~ $unsigned($unsigned(reg2753))) ?
                          (forvar2681[(1'h0):(1'h0)] ?
                              (~^reg2692[(1'h0):(1'h0)]) : $signed($signed(reg2771))) : reg2687);
                    end
                end
              if ((|(~&reg153)))
                begin
                  reg2811 <= ((|(reg2757[(1'h1):(1'h0)] ^ forvar208[(3'h7):(3'h5)])) >>> forvar176[(1'h1):(1'h0)]);
                  for (forvar2812 = (1'h0); (forvar2812 < (1'h1)); forvar2812 = (forvar2812 + (1'h1)))
                    begin
                      reg2813 <= (^~(reg212 ?
                          {$unsigned(reg213)} : ((reg2725 & reg209) ?
                              (reg188 == reg2731) : (-reg160))));
                      reg2814 <= reg2730;
                      reg2815 <= $signed(reg2730[(2'h3):(2'h2)]);
                      reg2816 <= ($signed(forvar2695[(1'h0):(1'h0)]) ?
                          reg2760 : {forvar153});
                    end
                  for (forvar2817 = (1'h0); (forvar2817 < (2'h2)); forvar2817 = (forvar2817 + (1'h1)))
                    begin
                      reg2818 <= ({(|(&forvar2695))} ?
                          {{$unsigned((8'ha0))}} : ((!reg173[(2'h2):(2'h2)]) | ($signed(reg213) ?
                              (reg193 >= reg2753) : $signed(reg2681))));
                      reg2819 <= ({(~&(|(8'hb8)))} ?
                          $unsigned(reg223) : reg2686);
                      reg2820 <= (+(~&$unsigned((forvar2695 - reg2813))));
                    end
                  for (forvar2821 = (1'h0); (forvar2821 < (2'h3)); forvar2821 = (forvar2821 + (1'h1)))
                    begin
                      reg2822 <= (8'ha0);
                      reg2823 <= ($signed((((8'hae) << reg174) >>> (^~forvar184))) - $signed(reg160));
                      reg2824 <= reg2763;
                    end
                end
              else
                begin
                  for (forvar2811 = (1'h0); (forvar2811 < (2'h3)); forvar2811 = (forvar2811 + (1'h1)))
                    begin
                      reg2812 <= (~($signed(reg2701) ?
                          reg2735 : forvar2793[(2'h2):(2'h2)]));
                    end
                  for (forvar2813 = (1'h0); (forvar2813 < (1'h0)); forvar2813 = (forvar2813 + (1'h1)))
                    begin
                      reg2814 <= (forvar2739[(3'h5):(1'h0)] ?
                          (+$unsigned({(8'hab)})) : reg2744[(4'hd):(3'h6)]);
                      reg2815 <= $unsigned($unsigned($unsigned($signed(reg173))));
                      reg2816 <= {((-$unsigned(reg222)) ?
                              forvar2686 : ((reg2694 >> reg2758) >= reg204))};
                    end
                  for (forvar2817 = (1'h0); (forvar2817 < (2'h3)); forvar2817 = (forvar2817 + (1'h1)))
                    begin
                      reg2818 <= reg165;
                      reg2819 <= reg2768;
                    end
                  reg2820 <= $unsigned({(reg200 ?
                          $unsigned((8'haa)) : (forvar2702 && (8'hb1)))});
                end
            end
          else
            begin
              for (forvar2793 = (1'h0); (forvar2793 < (2'h3)); forvar2793 = (forvar2793 + (1'h1)))
                begin
                  if ({{reg2823}})
                    begin
                      reg2794 <= (8'ha9);
                      reg2795 <= reg2751[(4'hc):(2'h3)];
                      reg2796 <= $signed((8'ha7));
                    end
                  else
                    begin
                      reg2794 <= forvar205[(3'h6):(1'h1)];
                      reg2795 <= reg2707[(3'h4):(2'h2)];
                      reg2796 <= (!forvar2710[(4'h8):(3'h4)]);
                    end
                end
            end
        end
      for (forvar2825 = (1'h0); (forvar2825 < (2'h3)); forvar2825 = (forvar2825 + (1'h1)))
        begin
          reg2826 <= (reg2693[(4'hd):(1'h1)] ? reg178 : reg200);
          reg2827 <= (|(8'hb7));
          reg2828 <= (~|$unsigned(($signed((8'hb3)) ?
              $unsigned((8'hb1)) : (reg2798 - reg2716))));
          for (forvar2829 = (1'h0); (forvar2829 < (1'h1)); forvar2829 = (forvar2829 + (1'h1)))
            begin
              if ((|((reg2689 ? ((8'ha7) | (8'h9c)) : $unsigned(reg2752)) ?
                  reg2722 : reg2689[(1'h1):(1'h0)])))
                begin
                  for (forvar2830 = (1'h0); (forvar2830 < (2'h2)); forvar2830 = (forvar2830 + (1'h1)))
                    begin
                      reg2831 <= $signed(((-(wire2675 ^~ forvar2775)) ?
                          (^~(^~reg2715)) : $signed((!reg2687))));
                      reg2832 <= $unsigned({($unsigned(reg2769) > (reg2689 - forvar2736))});
                    end
                  for (forvar2833 = (1'h0); (forvar2833 < (1'h0)); forvar2833 = (forvar2833 + (1'h1)))
                    begin
                      reg2834 <= $unsigned(reg203[(1'h1):(1'h0)]);
                      reg2835 <= reg2714[(4'h9):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar2830 = (1'h0); (forvar2830 < (2'h2)); forvar2830 = (forvar2830 + (1'h1)))
                    begin
                      reg2831 <= (~&reg2826);
                    end
                  if ($unsigned(($signed((~reg201)) ?
                      reg2757 : ($unsigned(reg2759) ?
                          $signed(reg2819) : (8'ha8)))))
                    begin
                      reg2832 <= ($signed($signed((reg2729 <= (8'ha0)))) >> $signed($unsigned((forvar156 ?
                          forvar2733 : forvar2718))));
                      reg2833 <= reg2744;
                      reg2834 <= (~($signed((&reg2684)) ^~ $signed(reg2728[(3'h6):(2'h3)])));
                      reg2835 <= ((($signed(forvar184) | (reg2741 && wire2673)) | (8'ha0)) || (~^{((8'h9e) ?
                              reg2772 : forvar2794)}));
                    end
                  else
                    begin
                      reg2832 <= $signed((~&reg2704[(3'h5):(3'h4)]));
                      reg2833 <= reg2687[(2'h2):(2'h2)];
                      reg2834 <= reg2760;
                    end
                end
            end
        end
      for (forvar2836 = (1'h0); (forvar2836 < (1'h0)); forvar2836 = (forvar2836 + (1'h1)))
        begin
          for (forvar2837 = (1'h0); (forvar2837 < (2'h2)); forvar2837 = (forvar2837 + (1'h1)))
            begin
              reg2838 <= (8'hb1);
              for (forvar2839 = (1'h0); (forvar2839 < (2'h2)); forvar2839 = (forvar2839 + (1'h1)))
                begin
                  for (forvar2840 = (1'h0); (forvar2840 < (1'h0)); forvar2840 = (forvar2840 + (1'h1)))
                    begin
                      reg2841 <= $signed((~|((+forvar161) >>> (forvar196 ?
                          forvar2687 : (8'hb2)))));
                      reg2842 <= reg2811[(1'h1):(1'h1)];
                      reg2843 <= reg2831[(4'hf):(3'h7)];
                    end
                  if ($signed(((+reg169) ? {reg2788[(4'ha):(4'h9)]} : reg162)))
                    begin
                      reg2844 <= reg2720[(3'h7):(3'h5)];
                      reg2845 <= ((8'hb9) ?
                          (reg182[(3'h4):(3'h4)] ?
                              $signed((reg2778 <<< forvar2682)) : ((reg2802 ?
                                  wire148 : (8'hb9)) != ((8'h9f) ?
                                  reg2711 : forvar2688))) : (8'ha2));
                    end
                  else
                    begin
                      reg2844 <= $signed($signed($unsigned((reg2788 >= forvar2836))));
                      reg2845 <= forvar218[(4'hf):(4'hd)];
                      reg2846 <= $unsigned((reg2808[(3'h4):(2'h2)] * {(~|(8'ha9))}));
                      reg2847 <= (^{(-(~^forvar2755))});
                    end
                  reg2848 <= $unsigned(forvar184[(4'hc):(1'h0)]);
                end
            end
          if (($unsigned(((~^(8'ha9)) ?
              ((8'ha7) == reg2848) : $unsigned(reg174))) ^~ (~|(|(~reg165)))))
            begin
              if (wire150)
                begin
                  reg2849 <= forvar2738[(4'hb):(3'h4)];
                  reg2850 <= $unsigned(($signed($signed(wire225)) ?
                      $unsigned(forvar2812[(1'h1):(1'h1)]) : $signed($unsigned(forvar2836))));
                end
              else
                begin
                  for (forvar2849 = (1'h0); (forvar2849 < (1'h0)); forvar2849 = (forvar2849 + (1'h1)))
                    begin
                      reg2850 <= (reg2757 ?
                          $signed((!$signed(reg2794))) : (8'had));
                    end
                  for (forvar2851 = (1'h0); (forvar2851 < (2'h2)); forvar2851 = (forvar2851 + (1'h1)))
                    begin
                      reg2852 <= (reg2828 * (8'had));
                      reg2853 <= {(((reg2752 || reg2849) + $unsigned(wire148)) >= $signed((reg222 != reg2816)))};
                      reg2854 <= (($signed($signed(reg2843)) ?
                          ((8'hae) | (forvar216 ?
                              (8'ha3) : reg2727)) : $unsigned(reg2752)) * reg2690[(2'h3):(2'h3)]);
                    end
                  for (forvar2855 = (1'h0); (forvar2855 < (1'h1)); forvar2855 = (forvar2855 + (1'h1)))
                    begin
                      reg2856 <= forvar2780;
                      reg2857 <= (((reg2790[(4'hb):(3'h5)] ?
                                  (reg2751 - forvar2849) : {(8'h9f)}) ?
                              $unsigned($unsigned(forvar176)) : forvar2687) ?
                          reg2681 : $signed($signed((reg2764 - (8'hac)))));
                      reg2858 <= {{$unsigned($signed(reg2724))}};
                      reg2859 <= (^~(forvar208[(3'h5):(3'h4)] ?
                          ((reg2697 << reg195) - {reg2799}) : $signed($signed((8'hb4)))));
                    end
                end
            end
          else
            begin
              for (forvar2849 = (1'h0); (forvar2849 < (1'h1)); forvar2849 = (forvar2849 + (1'h1)))
                begin
                  for (forvar2850 = (1'h0); (forvar2850 < (2'h3)); forvar2850 = (forvar2850 + (1'h1)))
                    begin
                      reg2851 <= reg2763;
                      reg2852 <= reg2753;
                      reg2853 <= ((reg153[(3'h5):(3'h5)] ?
                          $unsigned((reg2841 ?
                              forvar2839 : forvar2784)) : ($unsigned(reg2809) && forvar2781)) || (+($unsigned(reg155) ?
                          reg2776 : $signed(reg2844))));
                    end
                end
              for (forvar2854 = (1'h0); (forvar2854 < (2'h3)); forvar2854 = (forvar2854 + (1'h1)))
                begin
                  for (forvar2855 = (1'h0); (forvar2855 < (1'h0)); forvar2855 = (forvar2855 + (1'h1)))
                    begin
                      reg2856 <= (^reg2791);
                      reg2857 <= $unsigned(forvar168[(2'h2):(1'h0)]);
                      reg2858 <= (reg2795 + $unsigned((!$unsigned(reg2808))));
                    end
                  for (forvar2859 = (1'h0); (forvar2859 < (1'h1)); forvar2859 = (forvar2859 + (1'h1)))
                    begin
                      reg2860 <= $unsigned((((~^forvar152) & reg2730[(4'ha):(1'h0)]) & ((reg2844 + (8'hb3)) ?
                          (|reg2689) : forvar2855)));
                      reg2861 <= reg2853[(1'h1):(1'h0)];
                      reg2862 <= $signed(forvar152);
                    end
                  reg2863 <= {$unsigned(($unsigned(reg2766) ?
                          (~reg2688) : (reg172 ? forvar2689 : reg2846)))};
                end
              for (forvar2864 = (1'h0); (forvar2864 < (1'h1)); forvar2864 = (forvar2864 + (1'h1)))
                begin
                  for (forvar2865 = (1'h0); (forvar2865 < (1'h1)); forvar2865 = (forvar2865 + (1'h1)))
                    begin
                      reg2866 <= reg2730[(4'h8):(2'h3)];
                      reg2867 <= $unsigned((forvar191 ?
                          reg2741 : ((^reg2767) ?
                              forvar2726[(3'h5):(1'h1)] : (~&(8'h9d)))));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2868 = (1'h0); (forvar2868 < (1'h1)); forvar2868 = (forvar2868 + (1'h1)))
        begin
          for (forvar2869 = (1'h0); (forvar2869 < (1'h1)); forvar2869 = (forvar2869 + (1'h1)))
            begin
              for (forvar2870 = (1'h0); (forvar2870 < (2'h2)); forvar2870 = (forvar2870 + (1'h1)))
                begin
                  for (forvar2871 = (1'h0); (forvar2871 < (1'h1)); forvar2871 = (forvar2871 + (1'h1)))
                    begin
                      reg2872 <= forvar2804[(3'h5):(3'h4)];
                    end
                  for (forvar2873 = (1'h0); (forvar2873 < (2'h2)); forvar2873 = (forvar2873 + (1'h1)))
                    begin
                      reg2874 <= (!forvar2740[(1'h0):(1'h0)]);
                    end
                  if ((|reg2766))
                    begin
                      reg2875 <= {reg2863[(3'h6):(1'h1)]};
                      reg2876 <= $unsigned(reg2845);
                      reg2877 <= ($signed(({(8'hac)} ?
                              (reg2835 * reg2807) : (&reg204))) ?
                          reg157 : forvar2733);
                    end
                  else
                    begin
                      reg2875 <= $unsigned(forvar2692);
                    end
                  for (forvar2878 = (1'h0); (forvar2878 < (1'h1)); forvar2878 = (forvar2878 + (1'h1)))
                    begin
                      reg2879 <= (forvar2682 ?
                          reg2741 : $signed($unsigned(forvar2710[(2'h2):(1'h1)])));
                      reg2880 <= ($unsigned(((reg2751 < forvar2761) * {wire226})) <<< (~reg2787[(3'h4):(2'h2)]));
                      reg2881 <= $signed({{forvar2829[(4'h8):(3'h6)]}});
                      reg2882 <= ((~|$signed(reg2768[(3'h6):(3'h5)])) ?
                          reg2695 : (-$signed((reg2812 ?
                              reg2715 : forvar2811))));
                    end
                end
              reg2883 <= (^~($unsigned((reg2735 ? (8'ha2) : reg2841)) ?
                  $signed({reg2803}) : (reg203 & (reg2703 <= forvar2817))));
            end
          for (forvar2884 = (1'h0); (forvar2884 < (1'h1)); forvar2884 = (forvar2884 + (1'h1)))
            begin
              for (forvar2885 = (1'h0); (forvar2885 < (1'h0)); forvar2885 = (forvar2885 + (1'h1)))
                begin
                  reg2886 <= $unsigned($signed(($signed(reg2705) ?
                      (reg2806 != forvar2784) : (reg2842 ?
                          forvar2871 : reg2861))));
                  if ((8'hab))
                    begin
                      reg2887 <= {$signed(($signed((8'hb1)) ?
                              (~|(8'ha9)) : reg2768[(3'h6):(3'h5)]))};
                      reg2888 <= ((+reg2856) + $signed(((forvar2840 > reg2772) ?
                          reg2875 : (^reg2763))));
                    end
                  else
                    begin
                      reg2887 <= reg2824;
                      reg2888 <= reg2722;
                      reg2889 <= forvar172[(4'h8):(1'h1)];
                      reg2890 <= $signed((((^~(8'hb5)) ?
                          $signed((8'hb5)) : $unsigned(forvar179)) ^~ (|(forvar156 ?
                          reg2857 : reg2741))));
                    end
                  for (forvar2891 = (1'h0); (forvar2891 < (2'h3)); forvar2891 = (forvar2891 + (1'h1)))
                    begin
                      reg2892 <= $signed({$signed((~&(8'hba)))});
                      reg2893 <= $unsigned({(8'hac)});
                      reg2894 <= (~|(!$signed(reg2724)));
                      reg2895 <= (reg2685 ?
                          $unsigned(($unsigned(reg2816) < (reg2820 ?
                              reg153 : reg2693))) : $signed({(forvar197 >= reg165)}));
                    end
                end
              if (reg2694)
                begin
                  if (reg2862)
                    begin
                      reg2896 <= reg200;
                      reg2897 <= reg223;
                    end
                  else
                    begin
                      reg2896 <= ((~&$signed((forvar191 ? reg2792 : reg157))) ?
                          (((forvar2891 ?
                              forvar2891 : reg2822) != $unsigned(forvar156)) > (^(forvar2884 ?
                              reg2748 : forvar2687))) : (&{$unsigned((8'h9c))}));
                      reg2897 <= (8'ha6);
                      reg2898 <= (($unsigned((reg2889 != reg2693)) * (-(reg2811 < reg2824))) != forvar2687);
                    end
                  if ({{reg215}})
                    begin
                      reg2899 <= reg2856;
                    end
                  else
                    begin
                      reg2899 <= ((~^reg2728) != ($signed(forvar161) ?
                          {(reg185 * reg201)} : ((reg2827 ?
                                  forvar2686 : reg2712) ?
                              {(8'ha4)} : (reg2682 << reg2826))));
                    end
                  if (($unsigned(reg2751) ?
                      $unsigned(($signed(reg220) >>> (|forvar2775))) : reg2706))
                    begin
                      reg2900 <= reg2806;
                      reg2901 <= (8'hb0);
                      reg2902 <= ($unsigned($unsigned(((8'hab) ?
                          (8'ha3) : reg2729))) << forvar2784[(3'h4):(3'h4)]);
                      reg2903 <= $signed(reg2732[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg2900 <= $unsigned((~&(~wire2673)));
                      reg2901 <= reg2744;
                    end
                end
              else
                begin
                  if ($unsigned((forvar169 ?
                      ($signed(reg2893) ^ reg2826[(1'h0):(1'h0)]) : $unsigned($signed(reg2724)))))
                    begin
                      reg2896 <= {reg2684[(3'h4):(1'h1)]};
                      reg2897 <= (($signed($signed((8'ha9))) ?
                          forvar2682[(1'h1):(1'h0)] : ((^~forvar2708) ?
                              $unsigned(reg2726) : $unsigned((8'ha7)))) && wire150[(4'h8):(2'h2)]);
                      reg2898 <= (((forvar2830 ?
                              {(8'hb4)} : ((8'ha4) ^~ reg2819)) ?
                          {((8'hb3) || reg2844)} : {(!reg2787)}) <= {(~|$unsigned(forvar2715))});
                    end
                  else
                    begin
                      reg2896 <= {(&(8'haa))};
                    end
                  reg2899 <= ($signed(reg2759) ?
                      $signed(((!reg2705) ~^ reg2899[(1'h1):(1'h1)])) : $signed(wire285[(3'h7):(2'h2)]));
                end
            end
        end
      if ((!((~&(reg2809 ? reg2848 : forvar2811)) ?
          $unsigned(reg2802) : forvar170)))
        begin
          for (forvar2904 = (1'h0); (forvar2904 < (2'h2)); forvar2904 = (forvar2904 + (1'h1)))
            begin
              for (forvar2905 = (1'h0); (forvar2905 < (1'h1)); forvar2905 = (forvar2905 + (1'h1)))
                begin
                  for (forvar2906 = (1'h0); (forvar2906 < (2'h2)); forvar2906 = (forvar2906 + (1'h1)))
                    begin
                      reg2907 <= reg223[(2'h3):(1'h0)];
                      reg2908 <= reg2834;
                    end
                  reg2909 <= ({(!reg2688)} >= $unsigned($unsigned(((8'hac) && reg201))));
                  for (forvar2910 = (1'h0); (forvar2910 < (1'h1)); forvar2910 = (forvar2910 + (1'h1)))
                    begin
                      reg2911 <= (8'had);
                    end
                  for (forvar2912 = (1'h0); (forvar2912 < (2'h3)); forvar2912 = (forvar2912 + (1'h1)))
                    begin
                      reg2913 <= (reg2813 ?
                          $unsigned((~&$signed(forvar2738))) : $signed((((8'ha3) <= reg2746) ?
                              reg2725 : (forvar2692 > reg2901))));
                      reg2914 <= reg214;
                      reg2915 <= (((~$signed(forvar2830)) || (-(~&(8'hae)))) - (reg2854 ?
                          $signed((~^(8'ha9))) : (!forvar2829[(1'h1):(1'h1)])));
                    end
                end
              if (forvar2749)
                begin
                  for (forvar2916 = (1'h0); (forvar2916 < (2'h3)); forvar2916 = (forvar2916 + (1'h1)))
                    begin
                      reg2917 <= reg2698;
                      reg2918 <= (reg2861 ?
                          $unsigned((8'hb5)) : (~$signed(forvar176[(1'h1):(1'h0)])));
                      reg2919 <= ((((^(8'h9f)) != (reg2845 + reg2742)) > $signed($signed(wire226))) ?
                          $unsigned({{reg2767}}) : (~reg2787));
                      reg2920 <= ((!(~&reg2812)) && (+$unsigned(forvar196[(3'h6):(2'h2)])));
                    end
                end
              else
                begin
                  reg2916 <= (reg2896 <<< {(^reg2712[(4'h9):(2'h3)])});
                  for (forvar2917 = (1'h0); (forvar2917 < (1'h1)); forvar2917 = (forvar2917 + (1'h1)))
                    begin
                      reg2918 <= {(^(^~(reg2907 - forvar2710)))};
                      reg2919 <= $unsigned($signed(reg2679));
                      reg2920 <= $signed(reg2816[(2'h3):(2'h3)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar2904 = (1'h0); (forvar2904 < (1'h0)); forvar2904 = (forvar2904 + (1'h1)))
            begin
              if ({(-$signed((reg2834 ? reg2701 : reg2816)))})
                begin
                  if (forvar2904[(4'h9):(3'h4)])
                    begin
                      reg2905 <= {{((^~reg174) ?
                                  (~|forvar2802) : (+forvar168))}};
                      reg2906 <= (^(({reg214} ?
                          reg2824[(3'h4):(3'h4)] : {reg2850}) | ($unsigned((8'ha6)) != (forvar2837 & reg2920))));
                      reg2907 <= reg2898[(2'h2):(2'h2)];
                      reg2908 <= reg2818;
                    end
                  else
                    begin
                      reg2905 <= ($signed((forvar2762 ?
                              forvar198[(3'h6):(3'h4)] : (|reg193))) ?
                          reg2823 : (reg2801 ?
                              (~|$unsigned(reg2842)) : forvar172[(1'h0):(1'h0)]));
                    end
                  if ({$unsigned(reg2893)})
                    begin
                      reg2909 <= {((~|wire581) - $signed((8'ha0)))};
                      reg2910 <= reg2803;
                      reg2911 <= reg2743;
                    end
                  else
                    begin
                      reg2909 <= ({$signed(reg180[(1'h1):(1'h0)])} ?
                          $signed($unsigned((reg2777 ^ reg2875))) : ((8'haa) ?
                              (!(wire226 ?
                                  reg213 : reg2777)) : reg2692[(1'h0):(1'h0)]));
                      reg2910 <= {{reg2721}};
                    end
                  for (forvar2912 = (1'h0); (forvar2912 < (2'h3)); forvar2912 = (forvar2912 + (1'h1)))
                    begin
                      reg2913 <= reg2787;
                    end
                  for (forvar2914 = (1'h0); (forvar2914 < (1'h0)); forvar2914 = (forvar2914 + (1'h1)))
                    begin
                      reg2915 <= forvar2821;
                      reg2916 <= {(reg2769[(4'hf):(1'h0)] > ($unsigned(reg2881) <<< (&forvar2761)))};
                      reg2917 <= (^forvar152[(3'h7):(3'h7)]);
                    end
                end
              else
                begin
                  if (($signed($signed($unsigned(forvar2833))) ?
                      {reg213} : (forvar151 ?
                          ($unsigned(reg2783) > $signed(reg2858)) : reg2767[(1'h0):(1'h0)])))
                    begin
                      reg2905 <= (^forvar2715[(2'h2):(2'h2)]);
                      reg2906 <= $signed(forvar2865);
                    end
                  else
                    begin
                      reg2905 <= (-$unsigned($signed($signed(reg2683))));
                      reg2906 <= (!(~$signed($signed((8'hab)))));
                      reg2907 <= (~^(reg2730 ?
                          {(reg2681 ? forvar2829 : reg2906)} : (((8'hb9) ?
                              reg202 : (8'ha3)) > $unsigned((8'ha8)))));
                      reg2908 <= (8'ha4);
                    end
                  reg2909 <= reg2831[(4'he):(1'h1)];
                  if ((8'haf))
                    begin
                      reg2910 <= (^~(~|(8'hb6)));
                      reg2911 <= ($signed($signed((reg2908 ^~ reg186))) ?
                          $signed($unsigned({reg153})) : (~^$unsigned($unsigned(reg2812))));
                      reg2912 <= (!{(~^(^(8'hb0)))});
                      reg2913 <= reg2722;
                    end
                  else
                    begin
                      reg2910 <= $signed(($signed(((8'hab) != reg2791)) ?
                          {{reg2690}} : $unsigned(forvar2775[(3'h6):(1'h0)])));
                      reg2911 <= reg2820;
                      reg2912 <= reg2794;
                    end
                  for (forvar2914 = (1'h0); (forvar2914 < (2'h2)); forvar2914 = (forvar2914 + (1'h1)))
                    begin
                      reg2915 <= (!$signed(($unsigned(reg2684) ?
                          reg2681 : {(8'ha4)})));
                      reg2916 <= $signed((reg2828 ?
                          (~&$unsigned(wire226)) : (&(forvar2813 ^ reg2847))));
                    end
                end
            end
          for (forvar2918 = (1'h0); (forvar2918 < (1'h1)); forvar2918 = (forvar2918 + (1'h1)))
            begin
              if ($unsigned((reg2772 == (reg2771[(2'h3):(1'h0)] | $signed(forvar2855)))))
                begin
                  if ((~((reg158 ?
                      $signed(forvar2849) : (~^(8'ha0))) && ((!reg2826) ?
                      {(8'hb5)} : $signed((8'hb9))))))
                    begin
                      reg2919 <= ((forvar2738[(1'h0):(1'h0)] ?
                              {$unsigned(forvar152)} : (~&forvar2749)) ?
                          reg2725[(1'h1):(1'h1)] : $signed((8'hb1)));
                      reg2920 <= $unsigned(forvar2723);
                      reg2921 <= (~reg2824);
                    end
                  else
                    begin
                      reg2919 <= reg2872;
                      reg2920 <= ((((reg2771 - (8'hb6)) ^~ forvar2678) ~^ (~^(forvar2761 == forvar2802))) ?
                          $unsigned(($signed(reg154) ?
                              (reg2908 ?
                                  reg2743 : reg171) : {reg2798})) : $unsigned(forvar2865[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar2919 = (1'h0); (forvar2919 < (2'h2)); forvar2919 = (forvar2919 + (1'h1)))
                    begin
                      reg2920 <= ((~&$signed($signed((8'hac)))) ?
                          forvar2794[(3'h7):(3'h5)] : $signed($signed(reg2694[(3'h5):(3'h4)])));
                    end
                  for (forvar2921 = (1'h0); (forvar2921 < (2'h2)); forvar2921 = (forvar2921 + (1'h1)))
                    begin
                      reg2922 <= (&reg2848[(1'h1):(1'h1)]);
                      reg2923 <= (~^reg2799);
                      reg2924 <= ((^($signed((8'haf)) ?
                              (-reg2842) : $signed(forvar2761))) ?
                          (|(!reg182)) : (((^~forvar2689) ?
                                  $unsigned((8'hb1)) : $signed(reg2751)) ?
                              ($unsigned(forvar2910) - reg2704) : ($signed(reg2705) ?
                                  (reg222 ?
                                      forvar2829 : reg159) : $unsigned(reg221))));
                    end
                  for (forvar2925 = (1'h0); (forvar2925 < (1'h0)); forvar2925 = (forvar2925 + (1'h1)))
                    begin
                      reg2926 <= (reg2850[(2'h3):(1'h0)] & forvar216[(3'h6):(3'h6)]);
                      reg2927 <= $signed($signed($unsigned((|reg2883))));
                    end
                  if (reg2806[(4'h8):(1'h1)])
                    begin
                      reg2928 <= (($unsigned(reg2745[(3'h5):(2'h3)]) < ($unsigned((8'hae)) * {reg165})) ?
                          (&$unsigned((reg2877 >>> forvar2688))) : (&(forvar2868[(1'h0):(1'h0)] ?
                              reg2715[(1'h1):(1'h0)] : $signed(forvar216))));
                      reg2929 <= (forvar2708 ?
                          {reg2803} : $unsigned($signed(((8'hb5) ?
                              reg2772 : reg2848))));
                    end
                  else
                    begin
                      reg2928 <= ((wire285[(4'ha):(4'h9)] ?
                              forvar156[(3'h5):(3'h5)] : $signed(reg2706[(3'h5):(3'h4)])) ?
                          $signed({reg2679}) : $unsigned((forvar169[(4'ha):(3'h6)] || (reg2813 ?
                              forvar2910 : (8'had)))));
                    end
                end
              for (forvar2930 = (1'h0); (forvar2930 < (2'h3)); forvar2930 = (forvar2930 + (1'h1)))
                begin
                  if ($unsigned(($signed(forvar2836) ?
                      (reg2787 ? {(8'hac)} : reg2815) : (reg209 ?
                          (-reg2918) : reg222[(3'h4):(2'h3)]))))
                    begin
                      reg2931 <= (8'h9c);
                      reg2932 <= $unsigned((8'ha9));
                      reg2933 <= ((forvar196[(1'h1):(1'h1)] < (forvar2761 == (^~reg2816))) ?
                          (reg223[(2'h3):(2'h3)] << ({reg2706} ?
                              reg2766 : $signed(reg2826))) : $signed(reg200[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg2931 <= $unsigned($unsigned(({forvar2749} > $signed(forvar2762))));
                      reg2932 <= (~|{$unsigned($unsigned(reg2843))});
                    end
                end
              for (forvar2934 = (1'h0); (forvar2934 < (2'h3)); forvar2934 = (forvar2934 + (1'h1)))
                begin
                  for (forvar2935 = (1'h0); (forvar2935 < (1'h1)); forvar2935 = (forvar2935 + (1'h1)))
                    begin
                      reg2936 <= (reg2929[(2'h2):(2'h2)] ^~ (!(8'had)));
                      reg2937 <= $signed((forvar205 > reg207));
                    end
                  if ({(-$unsigned(forvar157))})
                    begin
                      reg2938 <= $unsigned((8'hb0));
                    end
                  else
                    begin
                      reg2938 <= forvar2836[(2'h3):(1'h0)];
                    end
                  reg2939 <= ((+reg2938[(1'h1):(1'h1)]) >> ((+((8'hb4) ^ forvar2921)) ?
                      reg2910 : reg2921[(4'h9):(3'h4)]));
                end
            end
          for (forvar2940 = (1'h0); (forvar2940 < (2'h2)); forvar2940 = (forvar2940 + (1'h1)))
            begin
              reg2941 <= $unsigned(reg221[(3'h4):(1'h1)]);
              if ($unsigned($unsigned($unsigned({reg2748}))))
                begin
                  if (reg155)
                    begin
                      reg2942 <= (8'h9e);
                      reg2943 <= $signed(forvar2916[(2'h3):(2'h3)]);
                      reg2944 <= $unsigned((reg2720[(3'h7):(3'h6)] ?
                          (^~(reg2895 + forvar2925)) : ({(8'hb5)} & (reg2753 ?
                              reg2721 : reg2911))));
                    end
                  else
                    begin
                      reg2942 <= reg2767;
                      reg2943 <= reg2807;
                      reg2944 <= (forvar2710 ?
                          (&$signed(reg178[(2'h3):(1'h1)])) : {$unsigned(reg188[(3'h7):(1'h1)])});
                    end
                end
              else
                begin
                  if (wire226[(4'hb):(1'h1)])
                    begin
                      reg2942 <= (^((^$signed(reg2776)) ?
                          reg2808 : (+(forvar2906 ? reg2796 : forvar2871))));
                    end
                  else
                    begin
                      reg2942 <= $signed($unsigned(forvar2849[(1'h0):(1'h0)]));
                      reg2943 <= reg2912[(1'h0):(1'h0)];
                      reg2944 <= forvar2836;
                    end
                  for (forvar2945 = (1'h0); (forvar2945 < (2'h2)); forvar2945 = (forvar2945 + (1'h1)))
                    begin
                      reg2946 <= $signed((~&$unsigned($unsigned(reg2744))));
                      reg2947 <= {(forvar197 | (-((8'haa) ?
                              reg2783 : reg156)))};
                      reg2948 <= $unsigned((+($unsigned(forvar2773) >= (forvar2755 <= reg2938))));
                      reg2949 <= ($unsigned({forvar2733[(2'h3):(1'h0)]}) >= $signed((forvar2775 - forvar216[(1'h0):(1'h0)])));
                    end
                end
            end
          for (forvar2950 = (1'h0); (forvar2950 < (1'h1)); forvar2950 = (forvar2950 + (1'h1)))
            begin
              if (($unsigned(reg2801[(3'h6):(2'h3)]) ?
                  reg161 : (forvar2681[(2'h3):(2'h3)] ?
                      $unsigned((^reg2693)) : (~&reg172[(3'h5):(2'h3)]))))
                begin
                  reg2951 <= ((((forvar2870 >= reg2746) - (8'hb5)) ~^ (+{reg2937})) != {(!forvar2710)});
                  for (forvar2952 = (1'h0); (forvar2952 < (1'h0)); forvar2952 = (forvar2952 + (1'h1)))
                    begin
                      reg2953 <= (forvar2804 ?
                          reg2894 : (&(^~forvar2813[(2'h2):(1'h0)])));
                      reg2954 <= ($unsigned(((reg2746 ~^ forvar2950) ?
                              $signed(forvar2736) : (^(8'ha2)))) ?
                          reg2801 : ({reg2810[(2'h2):(2'h2)]} ?
                              (8'h9e) : (forvar2950 - (~&(8'hab)))));
                      reg2955 <= $unsigned({(-$signed(reg154))});
                      reg2956 <= (&reg2842);
                    end
                  reg2957 <= reg2916[(3'h4):(1'h0)];
                end
              else
                begin
                  for (forvar2951 = (1'h0); (forvar2951 < (1'h0)); forvar2951 = (forvar2951 + (1'h1)))
                    begin
                      reg2952 <= reg2916;
                      reg2953 <= $signed($unsigned($unsigned($unsigned(reg2753))));
                      reg2954 <= $unsigned(wire225);
                    end
                  if ($unsigned($signed(reg2703[(3'h6):(3'h6)])))
                    begin
                      reg2955 <= (^$unsigned($unsigned((reg2911 && reg2689))));
                    end
                  else
                    begin
                      reg2955 <= forvar2891;
                    end
                end
              for (forvar2958 = (1'h0); (forvar2958 < (2'h3)); forvar2958 = (forvar2958 + (1'h1)))
                begin
                  for (forvar2959 = (1'h0); (forvar2959 < (2'h2)); forvar2959 = (forvar2959 + (1'h1)))
                    begin
                      reg2960 <= (~|(-(forvar2916[(2'h3):(1'h0)] ?
                          (reg2851 <<< (8'hb8)) : (reg2843 * forvar206))));
                      reg2961 <= $unsigned(reg2715[(2'h2):(1'h0)]);
                      reg2962 <= forvar2914[(2'h3):(2'h2)];
                      reg2963 <= reg2688;
                    end
                end
              if (((-((~&reg2880) ?
                  (forvar2784 << reg2806) : {reg2768})) >> wire2673[(4'h8):(3'h5)]))
                begin
                  for (forvar2964 = (1'h0); (forvar2964 < (1'h1)); forvar2964 = (forvar2964 + (1'h1)))
                    begin
                      reg2965 <= (&{((forvar2925 ?
                              reg2687 : (8'hae)) && (reg200 ^~ reg2693))});
                      reg2966 <= reg2688;
                      reg2967 <= ((!$signed({forvar2719})) ?
                          forvar2786[(4'h9):(3'h6)] : {forvar2951});
                    end
                  reg2968 <= $unsigned(reg2779[(3'h6):(3'h4)]);
                  if ({(~&reg2782[(1'h0):(1'h0)])})
                    begin
                      reg2969 <= $signed(reg2689[(3'h5):(3'h5)]);
                      reg2970 <= (reg2849 & wire583[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2969 <= ({$signed($unsigned(forvar2940))} ?
                          (+forvar2906) : ((&{forvar2917}) ?
                              reg2872[(2'h2):(1'h0)] : (|$unsigned(reg2922))));
                      reg2970 <= (forvar151[(1'h0):(1'h0)] ?
                          (forvar2719[(2'h3):(1'h0)] ?
                              ($unsigned(forvar2910) ^~ $signed(reg2805)) : ($unsigned(reg2764) - reg2902)) : reg2743[(2'h3):(2'h3)]);
                      reg2971 <= forvar2687;
                    end
                end
              else
                begin
                  if (($signed((-reg2805)) >>> (8'hac)))
                    begin
                      reg2964 <= (&$unsigned(((forvar2726 != forvar2904) << reg2928[(1'h1):(1'h1)])));
                      reg2965 <= ((~&forvar2733[(2'h3):(2'h2)]) ~^ forvar2749[(1'h1):(1'h0)]);
                      reg2966 <= $signed(reg2694[(4'h9):(4'h8)]);
                    end
                  else
                    begin
                      reg2964 <= reg175;
                      reg2965 <= forvar2773[(3'h5):(3'h4)];
                      reg2966 <= {$signed((~|$signed(reg2937)))};
                      reg2967 <= (($unsigned({reg2771}) - ((reg2699 ?
                              reg2783 : reg2834) ?
                          $unsigned(reg2915) : (reg2896 ?
                              forvar2715 : reg2797))) ^~ (reg2895[(4'hc):(3'h7)] ?
                          (~|$unsigned(wire225)) : (!wire146[(3'h7):(2'h2)])));
                    end
                  if ($unsigned({$signed($unsigned(reg2861))}))
                    begin
                      reg2968 <= (((~&$unsigned(forvar196)) + forvar191[(2'h3):(1'h0)]) || (^~((reg2906 ?
                              reg189 : reg2906) ?
                          $signed(reg2802) : reg2872[(2'h2):(2'h2)])));
                      reg2969 <= ($unsigned($signed((forvar2682 + (8'hb6)))) ^ $signed((reg182[(2'h3):(2'h2)] && {(8'hab)})));
                      reg2970 <= $unsigned(reg2851);
                    end
                  else
                    begin
                      reg2968 <= {$unsigned($signed((reg2906 ?
                              reg2970 : reg2729)))};
                      reg2969 <= $unsigned({(~|(~forvar2868))});
                    end
                  if (reg2689)
                    begin
                      reg2971 <= reg2705;
                    end
                  else
                    begin
                      reg2971 <= (!reg2797[(1'h0):(1'h0)]);
                      reg2972 <= $unsigned(($signed($unsigned(forvar2945)) >> (~reg2877)));
                      reg2973 <= $signed((^~{reg2750}));
                    end
                  if ($signed((reg2912 ? (+(-reg2726)) : forvar2878)))
                    begin
                      reg2974 <= (((reg2716 >= (reg2795 + forvar2687)) ~^ ((reg2688 ?
                                  reg2818 : forvar2871) ?
                              ((8'hb4) >>> reg2943) : reg2735)) ?
                          ($unsigned((reg193 <<< (8'hb9))) ?
                              {{reg166}} : reg164[(3'h5):(3'h4)]) : $signed((reg177[(1'h1):(1'h0)] ?
                              reg2892 : $unsigned(reg2943))));
                      reg2975 <= $signed(reg2849[(3'h7):(1'h1)]);
                      reg2976 <= (8'had);
                      reg2977 <= (|($signed({reg2699}) ?
                          {(|reg2838)} : $unsigned((forvar161 ?
                              forvar2917 : (8'haa)))));
                    end
                  else
                    begin
                      reg2974 <= (-$signed({reg2806}));
                      reg2975 <= $signed(reg2744[(4'he):(1'h1)]);
                      reg2976 <= (reg183 ?
                          ({forvar2761[(1'h0):(1'h0)]} ?
                              $signed(reg2948[(4'h9):(3'h6)]) : (^(^(8'h9c)))) : (^~((!reg2741) != (~^forvar2891))));
                    end
                end
            end
        end
      for (forvar2978 = (1'h0); (forvar2978 < (2'h2)); forvar2978 = (forvar2978 + (1'h1)))
        begin
          reg2979 <= $signed($unsigned(($signed((8'hb5)) | reg2838[(2'h3):(2'h3)])));
          for (forvar2980 = (1'h0); (forvar2980 < (2'h3)); forvar2980 = (forvar2980 + (1'h1)))
            begin
              for (forvar2981 = (1'h0); (forvar2981 < (1'h1)); forvar2981 = (forvar2981 + (1'h1)))
                begin
                  if ($signed((8'ha1)))
                    begin
                      reg2982 <= ((({reg173} ~^ $unsigned(forvar2775)) ?
                          ((~^reg2883) << reg2872) : (((8'ha6) >= reg2963) < (+forvar2851))) + $unsigned(forvar2715));
                      reg2983 <= $unsigned(({(reg2710 ? reg2973 : reg2843)} ?
                          (|(forvar2871 >= forvar2676)) : reg200[(3'h6):(3'h6)]));
                      reg2984 <= $unsigned($signed({reg2822}));
                    end
                  else
                    begin
                      reg2982 <= ((forvar198[(2'h2):(2'h2)] <<< {(reg2692 ?
                              reg2922 : (8'ha8))}) || forvar2945);
                      reg2983 <= reg2815;
                      reg2984 <= (~^(((reg2877 ? reg201 : (8'h9c)) ?
                          reg2796[(4'hc):(2'h3)] : (8'hb5)) >= (^$unsigned(reg2972))));
                    end
                  if (((forvar2804[(3'h6):(3'h4)] >> reg2683[(1'h1):(1'h1)]) - ($signed(reg2720[(2'h3):(2'h3)]) ?
                      reg2812 : (reg2879[(3'h7):(3'h6)] ?
                          reg2876 : $signed((8'haf))))))
                    begin
                      reg2985 <= ($unsigned(wire226[(4'hc):(1'h1)]) * $signed(((~|reg2699) >= (-reg2915))));
                      reg2986 <= {(^~(((8'hb6) ?
                              reg2937 : reg2971) + {reg2918}))};
                    end
                  else
                    begin
                      reg2985 <= forvar2702;
                      reg2986 <= (|(+$unsigned((^~reg2802))));
                    end
                  if ($signed(((8'had) ?
                      ((~reg2901) ? reg2692 : {(8'hb5)}) : ($signed((8'ha9)) ?
                          $signed(forvar2734) : (~reg2949)))))
                    begin
                      reg2987 <= (!(!(((8'hac) ? reg2688 : reg210) || (reg2911 ?
                          reg157 : forvar216))));
                      reg2988 <= $unsigned(reg2946);
                      reg2989 <= (({(reg2932 ? reg2942 : reg2711)} ?
                          forvar205[(1'h1):(1'h0)] : reg2841) || (reg2947[(3'h4):(2'h2)] >= ((reg220 < forvar157) ?
                          (8'ha3) : (^~(8'hb4)))));
                      reg2990 <= ($signed((forvar2865 ?
                          (^reg153) : {(8'h9f)})) <<< forvar2676[(3'h5):(2'h3)]);
                    end
                  else
                    begin
                      reg2987 <= $signed((reg2843 ?
                          ($signed((8'h9c)) >>> (reg2745 || reg2979)) : {(^reg2764)}));
                      reg2988 <= ((-$unsigned($signed((8'h9c)))) ?
                          reg2806 : ($unsigned(reg2886[(3'h4):(1'h0)]) | $signed((reg2831 ^ forvar184))));
                    end
                  if (({reg203} + (|forvar2683)))
                    begin
                      reg2991 <= ({(|(reg2772 ? reg209 : reg2909))} ?
                          reg2896[(2'h2):(1'h0)] : $unsigned((reg2711[(2'h2):(1'h0)] > (^reg2697))));
                      reg2992 <= {{forvar2802[(3'h7):(3'h6)]}};
                      reg2993 <= $signed(($signed({forvar2789}) <<< (wire2675[(2'h3):(2'h3)] ?
                          (^reg211) : (reg2790 << reg2905))));
                      reg2994 <= reg2874[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2991 <= (~reg154[(3'h7):(3'h6)]);
                      reg2992 <= reg2882;
                    end
                end
              if ($unsigned((~reg210[(2'h2):(2'h2)])))
                begin
                  if ((|$unsigned((reg2820 ?
                      (reg2722 ? reg2812 : reg213) : (forvar2749 ?
                          reg2795 : (8'h9c))))))
                    begin
                      reg2995 <= $unsigned((reg2790[(2'h2):(1'h0)] ?
                          ($unsigned((8'h9f)) ?
                              reg2682 : ((8'hb5) ?
                                  reg2745 : (8'haa))) : ((forvar2917 <= forvar2916) ?
                              $unsigned(reg2875) : $signed(forvar2978))));
                      reg2996 <= forvar2980[(1'h1):(1'h0)];
                      reg2997 <= $signed(($signed($signed(forvar2855)) ?
                          (forvar2692[(2'h3):(2'h2)] ?
                              (+forvar2749) : (reg2972 && reg2802)) : (~(reg2703 ?
                              reg2691 : forvar179))));
                      reg2998 <= (~{$signed((-reg2901))});
                    end
                  else
                    begin
                      reg2995 <= $signed((((8'hb4) ?
                          (!forvar2719) : {wire2675}) ^ $unsigned((+reg2842))));
                    end
                end
              else
                begin
                  reg2995 <= reg2863[(3'h5):(2'h2)];
                  for (forvar2996 = (1'h0); (forvar2996 < (1'h1)); forvar2996 = (forvar2996 + (1'h1)))
                    begin
                      reg2997 <= $unsigned((reg2756 ?
                          $unsigned((~&reg2900)) : {$signed(forvar2859)}));
                      reg2998 <= reg213[(3'h6):(3'h4)];
                    end
                  for (forvar2999 = (1'h0); (forvar2999 < (2'h3)); forvar2999 = (forvar2999 + (1'h1)))
                    begin
                      reg3000 <= reg2859;
                    end
                end
              for (forvar3001 = (1'h0); (forvar3001 < (2'h2)); forvar3001 = (forvar3001 + (1'h1)))
                begin
                  for (forvar3002 = (1'h0); (forvar3002 < (1'h1)); forvar3002 = (forvar3002 + (1'h1)))
                    begin
                      reg3003 <= ({($signed(reg2828) ?
                              $signed(forvar196) : (reg2889 ^~ reg2994))} && forvar2917);
                      reg3004 <= $unsigned(forvar2865);
                    end
                  for (forvar3005 = (1'h0); (forvar3005 < (1'h1)); forvar3005 = (forvar3005 + (1'h1)))
                    begin
                      reg3006 <= reg2895[(4'he):(3'h5)];
                    end
                  for (forvar3007 = (1'h0); (forvar3007 < (1'h0)); forvar3007 = (forvar3007 + (1'h1)))
                    begin
                      reg3008 <= $signed((|$signed($signed(reg2970))));
                      reg3009 <= $signed(reg2743);
                      reg3010 <= reg2974[(2'h3):(2'h2)];
                      reg3011 <= {{($signed(reg2860) != (reg2743 ?
                                  reg2976 : reg2831))}};
                    end
                  reg3012 <= $unsigned(reg2919[(4'h9):(3'h4)]);
                end
              if (($signed((reg2866[(4'ha):(3'h5)] ?
                  (~&reg2684) : $signed(reg2716))) < (forvar217 <<< (reg2920[(2'h3):(1'h0)] ?
                  reg2849 : $signed(forvar2884)))))
                begin
                  for (forvar3013 = (1'h0); (forvar3013 < (1'h1)); forvar3013 = (forvar3013 + (1'h1)))
                    begin
                      reg3014 <= (~&$unsigned($unsigned(reg2859[(2'h2):(1'h0)])));
                      reg3015 <= $unsigned($signed(({(8'haa)} ?
                          (reg183 * reg2924) : $signed(forvar2780))));
                      reg3016 <= $signed(reg2866);
                      reg3017 <= $signed((~^(&reg2691)));
                    end
                  for (forvar3018 = (1'h0); (forvar3018 < (2'h3)); forvar3018 = (forvar3018 + (1'h1)))
                    begin
                      reg3019 <= reg2695[(2'h2):(1'h1)];
                      reg3020 <= ($unsigned($unsigned((-reg2805))) ?
                          (8'h9d) : reg190);
                      reg3021 <= forvar179[(3'h7):(3'h6)];
                    end
                  reg3022 <= ({forvar2959} ?
                      $signed(((reg2906 > (8'h9e)) ?
                          $signed(forvar2695) : reg2720[(1'h0):(1'h0)])) : forvar172[(3'h6):(2'h2)]);
                  for (forvar3023 = (1'h0); (forvar3023 < (2'h2)); forvar3023 = (forvar3023 + (1'h1)))
                    begin
                      reg3024 <= (forvar2738 && $unsigned($unsigned((&reg195))));
                      reg3025 <= {forvar2733};
                    end
                end
              else
                begin
                  if ($signed(($signed((wire146 ? forvar2687 : forvar197)) ?
                      $signed({reg3004}) : $signed($signed(reg2698)))))
                    begin
                      reg3013 <= {forvar2951};
                    end
                  else
                    begin
                      reg3013 <= (^reg2833[(1'h0):(1'h0)]);
                      reg3014 <= $unsigned((((forvar2855 ?
                          forvar2878 : reg3024) << (-forvar2755)) + ((&(8'hb2)) ?
                          {forvar2884} : $signed(reg3014))));
                      reg3015 <= reg3021;
                    end
                  if ({{(~$unsigned((8'h9f)))}})
                    begin
                      reg3016 <= (+reg2943[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg3016 <= ($unsigned(reg204[(1'h1):(1'h1)]) ?
                          forvar2676[(2'h3):(1'h0)] : ((8'had) != $unsigned(forvar2830)));
                      reg3017 <= reg2747;
                      reg3018 <= $unsigned(reg2948);
                    end
                  for (forvar3019 = (1'h0); (forvar3019 < (2'h3)); forvar3019 = (forvar3019 + (1'h1)))
                    begin
                      reg3020 <= $signed($signed(($signed((8'hb7)) & forvar2864[(2'h2):(1'h0)])));
                      reg3021 <= $unsigned($signed($unsigned((forvar2793 ?
                          reg2694 : reg171))));
                      reg3022 <= forvar2677;
                      reg3023 <= reg2929[(1'h0):(1'h0)];
                    end
                  for (forvar3024 = (1'h0); (forvar3024 < (1'h0)); forvar3024 = (forvar3024 + (1'h1)))
                    begin
                      reg3025 <= (reg2875[(3'h6):(3'h5)] ~^ reg165);
                    end
                end
            end
        end
      for (forvar3026 = (1'h0); (forvar3026 < (2'h2)); forvar3026 = (forvar3026 + (1'h1)))
        begin
          for (forvar3027 = (1'h0); (forvar3027 < (2'h2)); forvar3027 = (forvar3027 + (1'h1)))
            begin
              reg3028 <= forvar2959;
              if (forvar2773[(1'h0):(1'h0)])
                begin
                  for (forvar3029 = (1'h0); (forvar3029 < (1'h1)); forvar3029 = (forvar3029 + (1'h1)))
                    begin
                      reg3030 <= (&reg2993[(2'h2):(1'h1)]);
                      reg3031 <= reg2876[(3'h7):(1'h1)];
                      reg3032 <= (forvar2999[(5'h10):(4'h8)] + $unsigned(reg2790[(4'h8):(3'h4)]));
                      reg3033 <= $signed(reg2907);
                    end
                end
              else
                begin
                  if ($unsigned((($unsigned(reg2975) ?
                      (!(8'h9f)) : $unsigned((8'ha4))) <= $signed(reg2943[(1'h1):(1'h0)]))))
                    begin
                      reg3029 <= $signed(reg2926);
                      reg3030 <= {reg2835[(3'h7):(3'h7)]};
                      reg3031 <= reg3011[(4'h8):(1'h0)];
                      reg3032 <= reg2678;
                    end
                  else
                    begin
                      reg3029 <= $unsigned(((forvar2916[(1'h1):(1'h0)] || $signed((8'hab))) ?
                          $unsigned((reg2823 ?
                              reg2843 : reg3018)) : reg2961[(4'ha):(3'h7)]));
                      reg3030 <= ($signed(reg2892) ? reg2750 : forvar2854);
                    end
                  if ((reg2714[(3'h5):(1'h1)] && reg2969))
                    begin
                      reg3033 <= (reg2700 != (((reg209 ?
                          wire226 : forvar169) && (reg2709 ?
                          reg2792 : reg2691)) & (-reg2852[(1'h0):(1'h0)])));
                      reg3034 <= $unsigned(reg2862);
                      reg3035 <= (^{{{reg173}}});
                    end
                  else
                    begin
                      reg3033 <= $signed({(((8'ha7) <<< (8'ha1)) ?
                              ((8'ha4) - reg2735) : (wire2673 ?
                                  reg2939 : reg2750))});
                      reg3034 <= (!((8'hb4) * forvar218));
                      reg3035 <= reg183[(4'hf):(1'h0)];
                      reg3036 <= $unsigned(($signed({reg2718}) ^ reg2923));
                    end
                end
              if ($signed((((reg2729 ?
                      reg2843 : (8'hb4)) <<< forvar3002[(3'h4):(3'h4)]) ?
                  forvar2739[(4'hc):(3'h7)] : (8'haa))))
                begin
                  for (forvar3037 = (1'h0); (forvar3037 < (1'h0)); forvar3037 = (forvar3037 + (1'h1)))
                    begin
                      reg3038 <= (+reg158);
                      reg3039 <= ((&reg2826) ^ $signed(forvar2686[(4'h8):(3'h4)]));
                      reg3040 <= (^~(^{(reg2957 << forvar2952)}));
                    end
                  reg3041 <= (~&(!(((8'ha8) ? reg2886 : reg2847) ?
                      (^~reg2994) : $unsigned(reg2853))));
                end
              else
                begin
                  if (reg2866[(2'h3):(1'h1)])
                    begin
                      reg3037 <= {reg2835};
                    end
                  else
                    begin
                      reg3037 <= reg2974[(2'h2):(2'h2)];
                      reg3038 <= (-reg2806);
                    end
                  if ((forvar2708 | $unsigned($signed($signed(reg2982)))))
                    begin
                      reg3039 <= forvar151[(4'he):(4'h9)];
                      reg3040 <= ((reg2844[(1'h0):(1'h0)] ?
                          forvar2884 : $signed($signed(forvar2695))) >= (8'haf));
                      reg3041 <= ((~((forvar2825 * reg203) ^~ {reg2707})) >>> reg2701);
                    end
                  else
                    begin
                      reg3039 <= ($signed($unsigned(reg2741[(3'h5):(3'h4)])) ?
                          $signed($unsigned($signed(forvar2765))) : ((((8'hb9) ?
                                      reg3029 : reg2905) ?
                                  $unsigned(reg2927) : (reg2676 ?
                                      reg2912 : reg167)) ?
                              ($unsigned(reg3020) ?
                                  forvar191[(2'h3):(1'h0)] : (~reg2790)) : (forvar2689[(2'h3):(2'h2)] ?
                                  reg2679[(3'h6):(2'h3)] : ((8'hab) ^ (8'ha2)))));
                      reg3040 <= {(|(!$signed(reg2956)))};
                      reg3041 <= $unsigned(({(reg2684 ? (8'ha8) : reg2895)} ?
                          $unsigned((~^forvar2940)) : $signed(reg2834)));
                    end
                  if ((forvar2804[(2'h3):(1'h1)] || (+reg2729)))
                    begin
                      reg3042 <= reg2847;
                      reg3043 <= (^(~|$unsigned((reg157 ? reg3037 : reg2938))));
                      reg3044 <= $unsigned((reg2975 ?
                          reg2856[(4'h8):(2'h2)] : ({(8'hab)} ?
                              (reg3032 ?
                                  forvar2829 : reg2893) : $unsigned(reg2737))));
                      reg3045 <= (forvar2773 ?
                          reg2924 : ({$signed(forvar2774)} ?
                              $unsigned((reg212 ?
                                  forvar2708 : reg162)) : forvar2726[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg3042 <= ($unsigned(((forvar2736 ?
                              reg2991 : reg2744) < (reg2800 ?
                              (8'ha6) : forvar2959))) ?
                          $unsigned((&reg2696[(4'ha):(3'h5)])) : (reg178 >>> $unsigned({forvar2849})));
                      reg3043 <= $signed((wire285 >>> (8'hb4)));
                    end
                end
            end
          reg3046 <= (8'haf);
          if (reg180[(2'h2):(1'h0)])
            begin
              if ((!(+(^~(^~reg2968)))))
                begin
                  for (forvar3047 = (1'h0); (forvar3047 < (2'h2)); forvar3047 = (forvar3047 + (1'h1)))
                    begin
                      reg3048 <= $unsigned(reg2994);
                      reg3049 <= $signed(reg2895);
                      reg3050 <= (8'ha5);
                      reg3051 <= (forvar2837 ?
                          $unsigned((~^wire583)) : reg2725);
                    end
                  if (($signed(reg2987) != (|reg2897[(1'h0):(1'h0)])))
                    begin
                      reg3052 <= reg2849;
                      reg3053 <= (($signed((^forvar3001)) ?
                          (!$unsigned(forvar2802)) : (reg2915[(2'h2):(2'h2)] == (reg2806 >= (8'hb5)))) ^ $unsigned($unsigned((forvar3027 ?
                          (8'hb0) : forvar206))));
                      reg3054 <= $signed(forvar216[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg3052 <= ((|(wire226 ?
                              (~|reg2798) : reg2715[(2'h2):(1'h1)])) ?
                          $signed(((-(8'h9d)) ?
                              (reg2937 ^~ reg2686) : (&reg2759))) : reg2721);
                    end
                  reg3055 <= (~&reg162[(4'hb):(3'h5)]);
                end
              else
                begin
                  for (forvar3047 = (1'h0); (forvar3047 < (2'h2)); forvar3047 = (forvar3047 + (1'h1)))
                    begin
                      reg3048 <= ({$signed($unsigned(reg2926))} ~^ ($unsigned(forvar2817[(2'h3):(1'h1)]) ?
                          reg190 : ($unsigned(forvar191) ? reg180 : reg200)));
                      reg3049 <= (~^$signed((reg2976 == (-reg2769))));
                    end
                  if (($unsigned((~&reg2857[(3'h6):(1'h1)])) && reg2832))
                    begin
                      reg3050 <= reg2691;
                    end
                  else
                    begin
                      reg3050 <= (-({(reg180 && forvar151)} ?
                          (+(forvar2925 >= reg161)) : ($unsigned(forvar172) ^ (^reg2704))));
                    end
                  reg3051 <= ((~|wire225[(2'h3):(2'h2)]) ?
                      ($signed((reg2833 == reg2861)) >>> $signed((8'hb1))) : (reg2812 ?
                          $unsigned($unsigned(reg2915)) : (!((8'h9e) || reg200))));
                end
              reg3056 <= $signed(reg2879[(2'h2):(2'h2)]);
            end
          else
            begin
              for (forvar3047 = (1'h0); (forvar3047 < (2'h3)); forvar3047 = (forvar3047 + (1'h1)))
                begin
                  for (forvar3048 = (1'h0); (forvar3048 < (1'h1)); forvar3048 = (forvar3048 + (1'h1)))
                    begin
                      reg3049 <= reg3043[(3'h7):(2'h3)];
                      reg3050 <= $unsigned(((~|forvar2904[(1'h0):(1'h0)]) ~^ ($signed(reg2682) << (~|reg2767))));
                      reg3051 <= (|{$unsigned((reg2957 ^ reg2796))});
                      reg3052 <= (~&($unsigned($unsigned(reg2782)) < forvar2904[(1'h1):(1'h1)]));
                    end
                  for (forvar3053 = (1'h0); (forvar3053 < (2'h2)); forvar3053 = (forvar3053 + (1'h1)))
                    begin
                      reg3054 <= $signed(reg2747);
                      reg3055 <= (reg2875[(3'h6):(2'h3)] >> ((~^(reg3016 || reg2797)) ?
                          ((reg2917 ? forvar2830 : reg2971) ?
                              (8'hb8) : forvar2951[(1'h1):(1'h0)]) : $signed((reg2911 < reg160))));
                    end
                end
              if (reg2876[(2'h3):(2'h3)])
                begin
                  for (forvar3056 = (1'h0); (forvar3056 < (2'h3)); forvar3056 = (forvar3056 + (1'h1)))
                    begin
                      reg3057 <= forvar2780;
                    end
                end
              else
                begin
                  for (forvar3056 = (1'h0); (forvar3056 < (1'h1)); forvar3056 = (forvar3056 + (1'h1)))
                    begin
                      reg3057 <= $unsigned(($signed($unsigned(reg2833)) & reg3010[(1'h0):(1'h0)]));
                      reg3058 <= reg2798[(3'h6):(1'h1)];
                      reg3059 <= forvar2681[(4'hd):(4'h9)];
                    end
                end
              for (forvar3060 = (1'h0); (forvar3060 < (2'h2)); forvar3060 = (forvar3060 + (1'h1)))
                begin
                  for (forvar3061 = (1'h0); (forvar3061 < (2'h2)); forvar3061 = (forvar3061 + (1'h1)))
                    begin
                      reg3062 <= (wire150 >> forvar2793[(2'h2):(1'h0)]);
                      reg3063 <= ($unsigned(((-reg2777) | ((8'ha1) ?
                              reg2682 : reg159))) ?
                          forvar3047[(4'hb):(3'h7)] : ($signed($unsigned(reg2862)) >>> (8'ha5)));
                      reg3064 <= ((^{$signed(reg2866)}) - (((8'hb9) || (reg2699 | reg2732)) >= $signed((~reg2744))));
                    end
                  if (($signed($unsigned($unsigned(forvar2925))) ?
                      ((((8'hb3) ? reg3063 : forvar206) ?
                              {(8'hb2)} : (reg2872 ? reg2962 : reg169)) ?
                          reg2687[(1'h1):(1'h0)] : ((reg3034 ~^ forvar164) ?
                              {(8'ha6)} : (~&(8'ha6)))) : {(~&reg2763)}))
                    begin
                      reg3065 <= (({reg2815[(2'h3):(2'h2)]} ?
                          {$signed((8'h9d))} : {{reg2735}}) == forvar2740);
                    end
                  else
                    begin
                      reg3065 <= {((|$unsigned(reg2911)) << $signed((forvar3027 ?
                              (8'ha1) : reg161)))};
                      reg3066 <= ($signed($unsigned(reg2901[(3'h5):(3'h5)])) << (8'hae));
                      reg3067 <= ((~^$unsigned(reg2883[(3'h4):(2'h2)])) != $unsigned($unsigned($signed(reg3028))));
                    end
                  if ((-{wire224}))
                    begin
                      reg3068 <= reg2937[(2'h2):(1'h0)];
                      reg3069 <= $signed((~|($unsigned(reg220) ?
                          reg2936 : (forvar198 ? reg2756 : (8'h9d)))));
                      reg3070 <= (!reg2875);
                    end
                  else
                    begin
                      reg3068 <= reg194[(2'h3):(2'h3)];
                      reg3069 <= forvar2878[(2'h3):(1'h0)];
                      reg3070 <= reg193;
                    end
                end
              if (($unsigned(reg2848[(2'h3):(1'h1)]) < reg3033[(4'ha):(3'h7)]))
                begin
                  for (forvar3071 = (1'h0); (forvar3071 < (2'h3)); forvar3071 = (forvar3071 + (1'h1)))
                    begin
                      reg3072 <= $unsigned(reg204[(4'h9):(2'h2)]);
                    end
                  for (forvar3073 = (1'h0); (forvar3073 < (2'h2)); forvar3073 = (forvar3073 + (1'h1)))
                    begin
                      reg3074 <= (~reg3033[(4'hb):(1'h1)]);
                      reg3075 <= $unsigned(((|{reg2931}) && ({forvar2773} ?
                          $signed((8'ha1)) : (reg3028 ? reg2763 : reg2769))));
                      reg3076 <= reg2687;
                    end
                end
              else
                begin
                  for (forvar3071 = (1'h0); (forvar3071 < (2'h3)); forvar3071 = (forvar3071 + (1'h1)))
                    begin
                      reg3072 <= reg219;
                      reg3073 <= reg2877;
                      reg3074 <= (8'hb9);
                      reg3075 <= $signed($unsigned((|$signed(forvar2891))));
                    end
                  for (forvar3076 = (1'h0); (forvar3076 < (1'h0)); forvar3076 = (forvar3076 + (1'h1)))
                    begin
                      reg3077 <= (|(+reg2782));
                      reg3078 <= (reg3014[(1'h0):(1'h0)] ?
                          (reg2685 & forvar2794[(3'h5):(2'h2)]) : (8'ha8));
                    end
                  if (reg3053)
                    begin
                      reg3079 <= ((^{(-forvar2676)}) ?
                          ($signed($unsigned(reg2896)) ?
                              (~$signed(reg2962)) : reg2893) : ((~&reg2853) ?
                              $signed($signed(reg201)) : reg2947[(2'h3):(1'h0)]));
                      reg3080 <= (forvar3019[(1'h1):(1'h0)] ?
                          reg3015 : $signed(forvar2708));
                    end
                  else
                    begin
                      reg3079 <= reg3049[(2'h2):(2'h2)];
                      reg3080 <= (~forvar3056[(4'h8):(3'h4)]);
                      reg3081 <= $signed((&$unsigned($signed(reg3056))));
                      reg3082 <= reg192[(4'hb):(3'h4)];
                    end
                end
            end
          for (forvar3083 = (1'h0); (forvar3083 < (1'h1)); forvar3083 = (forvar3083 + (1'h1)))
            begin
              if ({(~|$unsigned((^forvar2840)))})
                begin
                  for (forvar3084 = (1'h0); (forvar3084 < (1'h0)); forvar3084 = (forvar3084 + (1'h1)))
                    begin
                      reg3085 <= forvar2682[(1'h1):(1'h1)];
                      reg3086 <= ($signed(forvar2945) ?
                          (8'hb8) : ($unsigned(forvar191[(1'h0):(1'h0)]) ?
                              $unsigned((!reg2719)) : reg3070[(3'h5):(2'h2)]));
                      reg3087 <= ($unsigned({$unsigned((8'hb1))}) ~^ $signed(((+reg2745) ?
                          $unsigned(reg2876) : (~|reg2707))));
                    end
                end
              else
                begin
                  for (forvar3084 = (1'h0); (forvar3084 < (2'h2)); forvar3084 = (forvar3084 + (1'h1)))
                    begin
                      reg3085 <= wire147[(1'h0):(1'h0)];
                      reg3086 <= (8'hb8);
                      reg3087 <= {(^reg2955)};
                      reg3088 <= ((~|(forvar2780 >= $unsigned(reg2903))) && forvar2839);
                    end
                end
              for (forvar3089 = (1'h0); (forvar3089 < (1'h0)); forvar3089 = (forvar3089 + (1'h1)))
                begin
                  if ($unsigned(((|(reg2705 >> forvar3061)) << (&reg167[(1'h0):(1'h0)]))))
                    begin
                      reg3090 <= $unsigned(reg211[(3'h7):(1'h1)]);
                      reg3091 <= ((!(~{(8'ha1)})) <= {$signed((forvar2829 ?
                              (8'hb4) : reg3040))});
                      reg3092 <= $unsigned($signed(($signed(reg164) ?
                          $signed((8'hab)) : $unsigned(reg2751))));
                      reg3093 <= ($signed($unsigned((wire2675 || forvar2785))) > reg2952[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg3090 <= ((reg2889[(3'h5):(3'h4)] * reg2851) * (&((8'ha5) && (reg3079 ?
                          reg3012 : (8'hab)))));
                    end
                  for (forvar3094 = (1'h0); (forvar3094 < (1'h1)); forvar3094 = (forvar3094 + (1'h1)))
                    begin
                      reg3095 <= (~reg2924[(4'hc):(4'h9)]);
                      reg3096 <= $signed(reg2938[(4'ha):(3'h5)]);
                      reg3097 <= reg2972;
                    end
                  for (forvar3098 = (1'h0); (forvar3098 < (2'h2)); forvar3098 = (forvar3098 + (1'h1)))
                    begin
                      reg3099 <= (8'hb7);
                      reg3100 <= (wire224[(4'ha):(3'h7)] ?
                          (~^reg2850[(3'h5):(1'h0)]) : (((-reg2824) ?
                              (reg2947 && reg3024) : $signed(reg2828)) != forvar2774[(1'h1):(1'h0)]));
                      reg3101 <= {reg2778};
                    end
                end
            end
        end
    end
  assign wire3102 = forvar2780[(2'h3):(2'h3)];
  assign wire3103 = (-reg207[(4'h9):(4'h9)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module584
#( parameter param2672 = (^~{(((8'hac) ? (8'had) : (8'hb0)) ? {(8'ha6)} : (!(8'ha7)))}) )
(y, clk, wire589, wire588, wire587, wire586, wire585);
  output wire [(32'h181e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire589;
  input wire [(5'h10):(1'h0)] wire588;
  input wire signed [(4'he):(1'h0)] wire587;
  input wire [(4'hb):(1'h0)] wire586;
  input wire signed [(4'h9):(1'h0)] wire585;
  wire [(4'h9):(1'h0)] wire2671;
  wire signed [(4'hf):(1'h0)] wire2670;
  wire signed [(4'h9):(1'h0)] wire2669;
  wire [(3'h5):(1'h0)] wire1145;
  wire signed [(3'h7):(1'h0)] wire590;
  wire [(4'he):(1'h0)] wire1147;
  reg signed [(3'h7):(1'h0)] reg1148 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1149 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1150 = (1'h0);
  reg [(3'h6):(1'h0)] reg1151 = (1'h0);
  reg [(3'h4):(1'h0)] reg1152 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1153 = (1'h0);
  reg [(3'h4):(1'h0)] reg1154 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1155 = (1'h0);
  reg [(3'h5):(1'h0)] reg1156 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1157 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1158 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1159 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1160 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1161 = (1'h0);
  reg [(3'h6):(1'h0)] reg1149 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1150 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1156 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1158 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1162 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1163 = (1'h0);
  reg [(3'h4):(1'h0)] reg1164 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1165 = (1'h0);
  reg [(3'h6):(1'h0)] reg1166 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1167 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1169 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1170 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1151 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1153 = (1'h0);
  reg [(4'hc):(1'h0)] reg1163 = (1'h0);
  reg [(4'hf):(1'h0)] reg1165 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1166 = (1'h0);
  reg [(4'hc):(1'h0)] reg1167 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1171 = (1'h0);
  reg [(4'h8):(1'h0)] reg1172 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1173 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1174 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1175 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1177 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1178 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1179 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1180 = (1'h0);
  reg [(3'h6):(1'h0)] reg1181 = (1'h0);
  reg [(5'h10):(1'h0)] reg1182 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1183 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1184 = (1'h0);
  reg [(2'h3):(1'h0)] reg1185 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1186 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1187 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1178 = (1'h0);
  reg [(3'h7):(1'h0)] reg1179 = (1'h0);
  reg [(3'h5):(1'h0)] reg1180 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1183 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1186 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1188 = (1'h0);
  reg [(4'ha):(1'h0)] reg1189 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1190 = (1'h0);
  reg [(3'h6):(1'h0)] reg1191 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1192 = (1'h0);
  reg [(4'he):(1'h0)] reg1193 = (1'h0);
  reg [(2'h2):(1'h0)] reg1194 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1195 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1152 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1154 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1157 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1159 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1162 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1161 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1168 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1169 = (1'h0);
  reg [(4'ha):(1'h0)] reg1171 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1177 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1148 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1196 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1197 = (1'h0);
  reg [(5'h10):(1'h0)] reg1198 = (1'h0);
  reg [(5'h10):(1'h0)] reg1199 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1200 = (1'h0);
  reg [(3'h6):(1'h0)] reg1201 = (1'h0);
  reg [(5'h10):(1'h0)] reg1202 = (1'h0);
  reg [(4'he):(1'h0)] reg1203 = (1'h0);
  reg [(4'hc):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1205 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1206 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1207 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1208 = (1'h0);
  reg [(3'h4):(1'h0)] reg1209 = (1'h0);
  reg [(2'h3):(1'h0)] reg1210 = (1'h0);
  reg [(3'h7):(1'h0)] reg1211 = (1'h0);
  reg [(4'ha):(1'h0)] reg1212 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1213 = (1'h0);
  reg [(4'hf):(1'h0)] reg1214 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1215 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1205 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1207 = (1'h0);
  reg [(4'h9):(1'h0)] reg1216 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1217 = (1'h0);
  reg [(4'hb):(1'h0)] reg1218 = (1'h0);
  reg [(5'h10):(1'h0)] reg1219 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1220 = (1'h0);
  reg [(4'hc):(1'h0)] reg1221 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1216 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1218 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1222 = (1'h0);
  reg [(4'hc):(1'h0)] reg1197 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1202 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1209 = (1'h0);
  reg [(4'he):(1'h0)] reg1213 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1214 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1219 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1221 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1201 = (1'h0);
  reg [(4'hd):(1'h0)] reg1196 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1210 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1212 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1223 = (1'h0);
  reg [(3'h4):(1'h0)] reg1224 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1225 = (1'h0);
  reg [(4'hb):(1'h0)] reg1226 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1227 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1228 = (1'h0);
  reg [(2'h2):(1'h0)] reg1229 = (1'h0);
  reg [(3'h6):(1'h0)] reg1230 = (1'h0);
  reg [(4'hd):(1'h0)] reg1231 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1232 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1233 = (1'h0);
  reg [(4'hf):(1'h0)] reg1234 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1235 = (1'h0);
  reg [(3'h6):(1'h0)] reg1236 = (1'h0);
  reg [(2'h3):(1'h0)] reg1237 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1238 = (1'h0);
  reg [(4'hc):(1'h0)] reg1239 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1240 = (1'h0);
  reg [(3'h4):(1'h0)] reg1241 = (1'h0);
  reg [(4'he):(1'h0)] reg1242 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1243 = (1'h0);
  reg [(5'h10):(1'h0)] reg1244 = (1'h0);
  reg [(3'h6):(1'h0)] reg1245 = (1'h0);
  reg [(4'ha):(1'h0)] reg1246 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1247 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1248 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1249 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1250 = (1'h0);
  reg [(4'ha):(1'h0)] reg1251 = (1'h0);
  reg [(3'h5):(1'h0)] reg1252 = (1'h0);
  reg [(4'ha):(1'h0)] reg1238 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1243 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1246 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1251 = (1'h0);
  reg [(4'h8):(1'h0)] reg1253 = (1'h0);
  reg [(4'hd):(1'h0)] reg1254 = (1'h0);
  reg [(4'hc):(1'h0)] reg1255 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1256 = (1'h0);
  reg [(5'h10):(1'h0)] reg1257 = (1'h0);
  reg [(5'h10):(1'h0)] reg1258 = (1'h0);
  reg [(4'hf):(1'h0)] reg1259 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1260 = (1'h0);
  reg [(4'hb):(1'h0)] reg1261 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1262 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1263 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1264 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1265 = (1'h0);
  reg [(4'hd):(1'h0)] reg1266 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1267 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1268 = (1'h0);
  reg [(3'h7):(1'h0)] reg1269 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1270 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1271 = (1'h0);
  reg [(4'he):(1'h0)] forvar1265 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1229 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1232 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1272 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1273 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1274 = (1'h0);
  reg [(2'h2):(1'h0)] reg1275 = (1'h0);
  reg [(2'h2):(1'h0)] reg1276 = (1'h0);
  reg [(4'he):(1'h0)] reg1277 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1278 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1279 = (1'h0);
  reg [(5'h10):(1'h0)] reg1280 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1281 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1282 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1283 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1284 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1286 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1287 = (1'h0);
  reg [(4'hd):(1'h0)] reg1288 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1289 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1290 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1291 = (1'h0);
  reg [(2'h3):(1'h0)] reg1292 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1293 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1294 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1295 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1296 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1297 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1290 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1291 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1298 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1299 = (1'h0);
  reg [(3'h7):(1'h0)] reg1300 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1301 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1302 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1303 = (1'h0);
  reg [(4'hb):(1'h0)] reg1304 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1305 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1306 = (1'h0);
  reg [(4'hd):(1'h0)] reg1307 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1308 = (1'h0);
  reg [(3'h6):(1'h0)] reg1309 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1310 = (1'h0);
  reg [(4'hb):(1'h0)] reg1311 = (1'h0);
  reg [(2'h3):(1'h0)] reg1312 = (1'h0);
  reg [(3'h6):(1'h0)] reg1313 = (1'h0);
  reg [(3'h7):(1'h0)] reg1305 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1306 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1310 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1314 = (1'h0);
  reg [(3'h5):(1'h0)] reg1315 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1316 = (1'h0);
  reg [(4'he):(1'h0)] reg1314 = (1'h0);
  reg [(5'h10):(1'h0)] reg1317 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1318 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1319 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1320 = (1'h0);
  reg [(3'h5):(1'h0)] reg1321 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1322 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1323 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1324 = (1'h0);
  reg [(4'ha):(1'h0)] reg1325 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1326 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1323 = (1'h0);
  reg [(4'hd):(1'h0)] reg1327 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1304 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1309 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1328 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1329 = (1'h0);
  reg [(4'h8):(1'h0)] reg1330 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1331 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1332 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1333 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1335 = (1'h0);
  reg [(3'h7):(1'h0)] reg1336 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1337 = (1'h0);
  reg [(2'h2):(1'h0)] reg1338 = (1'h0);
  reg [(4'hf):(1'h0)] reg1339 = (1'h0);
  reg [(2'h2):(1'h0)] reg1340 = (1'h0);
  reg [(5'h10):(1'h0)] reg1341 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1342 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1343 = (1'h0);
  reg [(3'h7):(1'h0)] reg1344 = (1'h0);
  reg [(3'h4):(1'h0)] reg1345 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1341 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1346 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1347 = (1'h0);
  reg [(3'h6):(1'h0)] reg1348 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1349 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1350 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1351 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1352 = (1'h0);
  reg [(2'h2):(1'h0)] reg1353 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1354 = (1'h0);
  reg [(4'hb):(1'h0)] reg1355 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1356 = (1'h0);
  reg [(4'he):(1'h0)] reg1357 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1358 = (1'h0);
  reg [(4'he):(1'h0)] forvar1348 = (1'h0);
  reg [(4'ha):(1'h0)] reg1350 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1351 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1354 = (1'h0);
  reg [(4'ha):(1'h0)] reg1359 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1360 = (1'h0);
  reg [(2'h2):(1'h0)] reg1361 = (1'h0);
  reg [(2'h2):(1'h0)] reg1362 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1363 = (1'h0);
  reg [(2'h2):(1'h0)] reg1364 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1365 = (1'h0);
  reg [(4'h9):(1'h0)] reg1366 = (1'h0);
  reg [(3'h5):(1'h0)] reg1367 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1328 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1330 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1332 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1334 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1337 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1224 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1228 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1231 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1233 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1223 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1226 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1239 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1241 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1247 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1248 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1250 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1252 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1256 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1258 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1259 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1261 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1262 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1260 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1264 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1269 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1271 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1272 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1273 = (1'h0);
  reg [(2'h3):(1'h0)] reg1274 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1368 = (1'h0);
  reg [(3'h6):(1'h0)] reg1369 = (1'h0);
  reg [(4'h8):(1'h0)] reg1370 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1371 = (1'h0);
  reg [(2'h2):(1'h0)] reg1372 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1373 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1374 = (1'h0);
  reg [(4'hd):(1'h0)] reg1375 = (1'h0);
  reg [(4'h8):(1'h0)] reg1376 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1377 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1378 = (1'h0);
  reg [(4'he):(1'h0)] reg1379 = (1'h0);
  reg [(3'h5):(1'h0)] reg1380 = (1'h0);
  reg [(3'h7):(1'h0)] reg1381 = (1'h0);
  reg [(4'hd):(1'h0)] reg1382 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1383 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1373 = (1'h0);
  reg [(4'hf):(1'h0)] reg1378 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1370 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1371 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1384 = (1'h0);
  reg [(4'he):(1'h0)] reg1385 = (1'h0);
  reg [(4'h9):(1'h0)] reg1386 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1387 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1388 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1389 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1390 = (1'h0);
  reg [(2'h3):(1'h0)] reg1384 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1391 = (1'h0);
  reg [(4'h8):(1'h0)] reg1392 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1393 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1394 = (1'h0);
  reg [(4'ha):(1'h0)] reg1395 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1396 = (1'h0);
  reg [(4'hf):(1'h0)] reg1397 = (1'h0);
  reg [(4'ha):(1'h0)] reg1398 = (1'h0);
  reg [(4'ha):(1'h0)] reg1394 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1395 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1399 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1400 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1401 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1402 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1403 = (1'h0);
  reg [(4'h8):(1'h0)] reg1404 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1405 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1406 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1407 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1408 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1409 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1410 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1411 = (1'h0);
  reg [(3'h7):(1'h0)] reg1412 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1413 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1414 = (1'h0);
  reg [(2'h2):(1'h0)] reg1415 = (1'h0);
  reg [(4'hd):(1'h0)] reg1416 = (1'h0);
  reg [(5'h10):(1'h0)] reg1417 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1418 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1419 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1420 = (1'h0);
  reg [(5'h10):(1'h0)] reg1421 = (1'h0);
  reg [(2'h2):(1'h0)] reg1422 = (1'h0);
  reg [(4'h9):(1'h0)] reg1423 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1424 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1425 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1426 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1427 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1428 = (1'h0);
  reg [(5'h10):(1'h0)] reg1429 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1430 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1431 = (1'h0);
  reg [(4'he):(1'h0)] reg1432 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1433 = (1'h0);
  reg [(5'h10):(1'h0)] reg1434 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1435 = (1'h0);
  reg [(4'hb):(1'h0)] reg1436 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1437 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1438 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1439 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1440 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1438 = (1'h0);
  reg [(4'ha):(1'h0)] reg1441 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1442 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1443 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1444 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1445 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1446 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1447 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1448 = (1'h0);
  reg [(4'hc):(1'h0)] reg1449 = (1'h0);
  reg [(4'hf):(1'h0)] reg1450 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1446 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1448 = (1'h0);
  reg [(3'h6):(1'h0)] reg1451 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1450 = (1'h0);
  reg [(4'hd):(1'h0)] reg1452 = (1'h0);
  reg [(4'hb):(1'h0)] reg1453 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1454 = (1'h0);
  reg [(2'h3):(1'h0)] reg1455 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1456 = (1'h0);
  reg [(2'h3):(1'h0)] reg1457 = (1'h0);
  reg [(3'h5):(1'h0)] reg1458 = (1'h0);
  reg [(4'hd):(1'h0)] reg1459 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1460 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1461 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1462 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1463 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1464 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1465 = (1'h0);
  reg [(5'h10):(1'h0)] reg1466 = (1'h0);
  reg [(3'h4):(1'h0)] reg1467 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1468 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1469 = (1'h0);
  reg [(4'hc):(1'h0)] reg1470 = (1'h0);
  reg [(2'h2):(1'h0)] reg1471 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1472 = (1'h0);
  reg [(4'hb):(1'h0)] reg1473 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1474 = (1'h0);
  reg [(4'h8):(1'h0)] reg1475 = (1'h0);
  reg [(4'h9):(1'h0)] reg1476 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1477 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1478 = (1'h0);
  reg [(4'hc):(1'h0)] reg1479 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1480 = (1'h0);
  reg [(4'hc):(1'h0)] reg1481 = (1'h0);
  reg [(2'h2):(1'h0)] reg1482 = (1'h0);
  reg [(4'hc):(1'h0)] reg1469 = (1'h0);
  reg [(3'h5):(1'h0)] reg1472 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1479 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1480 = (1'h0);
  reg [(2'h2):(1'h0)] reg1483 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1484 = (1'h0);
  reg [(3'h7):(1'h0)] reg1485 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1486 = (1'h0);
  reg [(3'h4):(1'h0)] reg1487 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1488 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1489 = (1'h0);
  reg [(4'hc):(1'h0)] reg1490 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1484 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1491 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1492 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1493 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1494 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1495 = (1'h0);
  reg [(4'hf):(1'h0)] reg1496 = (1'h0);
  reg [(4'ha):(1'h0)] reg1497 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1498 = (1'h0);
  reg [(4'hc):(1'h0)] reg1499 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1500 = (1'h0);
  reg [(4'h8):(1'h0)] reg1501 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1502 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1495 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1496 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1503 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1504 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1505 = (1'h0);
  reg [(3'h6):(1'h0)] reg1506 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1507 = (1'h0);
  reg [(3'h6):(1'h0)] reg1508 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1504 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire1735;
  reg signed [(3'h4):(1'h0)] forvar1737 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1738 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1739 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1740 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1741 = (1'h0);
  reg [(3'h7):(1'h0)] reg1742 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1743 = (1'h0);
  reg [(2'h2):(1'h0)] reg1744 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1745 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1746 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1747 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1748 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1749 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1750 = (1'h0);
  reg [(4'hc):(1'h0)] reg1751 = (1'h0);
  reg [(3'h6):(1'h0)] reg1752 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1753 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1754 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1755 = (1'h0);
  reg [(4'hd):(1'h0)] reg1756 = (1'h0);
  reg [(2'h3):(1'h0)] reg1757 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1758 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1759 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1760 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1761 = (1'h0);
  reg [(4'h8):(1'h0)] reg1762 = (1'h0);
  reg [(5'h10):(1'h0)] reg1763 = (1'h0);
  reg [(4'hd):(1'h0)] reg1764 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1765 = (1'h0);
  reg [(3'h4):(1'h0)] reg1766 = (1'h0);
  reg [(4'hc):(1'h0)] reg1767 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1768 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1769 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1770 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1771 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1772 = (1'h0);
  reg [(4'hf):(1'h0)] reg1773 = (1'h0);
  reg [(3'h7):(1'h0)] reg1774 = (1'h0);
  reg [(3'h6):(1'h0)] reg1775 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1776 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1777 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1778 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1779 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1780 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1781 = (1'h0);
  reg [(4'hd):(1'h0)] reg1782 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1783 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1784 = (1'h0);
  reg [(4'ha):(1'h0)] reg1785 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1786 = (1'h0);
  reg [(3'h4):(1'h0)] reg1787 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1788 = (1'h0);
  reg [(4'hb):(1'h0)] reg1789 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1790 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1791 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1792 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1793 = (1'h0);
  reg [(4'he):(1'h0)] reg1794 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1795 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1796 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1797 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1798 = (1'h0);
  reg [(2'h3):(1'h0)] reg1799 = (1'h0);
  reg [(4'he):(1'h0)] reg1800 = (1'h0);
  reg [(4'hd):(1'h0)] reg1801 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1802 = (1'h0);
  reg [(4'h8):(1'h0)] reg1803 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1804 = (1'h0);
  reg [(4'hd):(1'h0)] reg1805 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1806 = (1'h0);
  reg [(2'h3):(1'h0)] reg1807 = (1'h0);
  reg [(2'h2):(1'h0)] reg1808 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1809 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1810 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1811 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1812 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1813 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1814 = (1'h0);
  reg [(3'h7):(1'h0)] reg1815 = (1'h0);
  reg [(5'h10):(1'h0)] reg1816 = (1'h0);
  reg [(3'h4):(1'h0)] reg1817 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1813 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1816 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1818 = (1'h0);
  reg [(3'h7):(1'h0)] reg1819 = (1'h0);
  reg [(4'hb):(1'h0)] reg1820 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1803 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1807 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1808 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1809 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1821 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1822 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1823 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1824 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1825 = (1'h0);
  reg [(4'hd):(1'h0)] reg1826 = (1'h0);
  reg [(2'h3):(1'h0)] reg1827 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1828 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1829 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1830 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1831 = (1'h0);
  reg [(5'h10):(1'h0)] reg1832 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1833 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1834 = (1'h0);
  reg [(2'h2):(1'h0)] reg1831 = (1'h0);
  reg [(4'h8):(1'h0)] reg1835 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1836 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1837 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1838 = (1'h0);
  reg [(4'ha):(1'h0)] reg1839 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1828 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1830 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1835 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1836 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1837 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1839 = (1'h0);
  reg [(4'he):(1'h0)] reg1840 = (1'h0);
  reg [(4'hd):(1'h0)] reg1841 = (1'h0);
  reg [(3'h6):(1'h0)] reg1842 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1840 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1843 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1844 = (1'h0);
  reg [(4'hd):(1'h0)] reg1845 = (1'h0);
  reg [(2'h2):(1'h0)] reg1846 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1844 = (1'h0);
  reg [(3'h5):(1'h0)] reg1847 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1848 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1849 = (1'h0);
  reg [(4'h8):(1'h0)] reg1850 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1833 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1851 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1852 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1853 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1854 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1855 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1856 = (1'h0);
  reg [(4'hb):(1'h0)] reg1857 = (1'h0);
  reg [(4'he):(1'h0)] reg1858 = (1'h0);
  reg [(4'hb):(1'h0)] reg1859 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1860 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1861 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1862 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1863 = (1'h0);
  reg [(4'hb):(1'h0)] reg1864 = (1'h0);
  reg [(5'h10):(1'h0)] reg1865 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1866 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1867 = (1'h0);
  reg [(4'h9):(1'h0)] reg1868 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1863 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1869 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1870 = (1'h0);
  reg [(2'h2):(1'h0)] reg1871 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1872 = (1'h0);
  reg [(3'h7):(1'h0)] reg1873 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1874 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1875 = (1'h0);
  reg [(3'h5):(1'h0)] reg1876 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1877 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1878 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1879 = (1'h0);
  reg [(4'hb):(1'h0)] reg1880 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1881 = (1'h0);
  reg [(3'h6):(1'h0)] reg1882 = (1'h0);
  reg [(2'h3):(1'h0)] reg1883 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1884 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1885 = (1'h0);
  reg [(2'h3):(1'h0)] reg1886 = (1'h0);
  reg [(5'h10):(1'h0)] reg1887 = (1'h0);
  reg [(2'h3):(1'h0)] reg1888 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1889 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1890 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1891 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1892 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1893 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1894 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1895 = (1'h0);
  reg [(4'he):(1'h0)] reg1896 = (1'h0);
  reg [(3'h7):(1'h0)] reg1897 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1898 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1899 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1900 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1901 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1902 = (1'h0);
  reg [(4'h9):(1'h0)] reg1903 = (1'h0);
  reg [(4'he):(1'h0)] reg1904 = (1'h0);
  reg [(4'h8):(1'h0)] reg1905 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1906 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1907 = (1'h0);
  reg [(4'h9):(1'h0)] reg1908 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1909 = (1'h0);
  reg [(4'hb):(1'h0)] reg1910 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1911 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1912 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1913 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1914 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1915 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1916 = (1'h0);
  reg [(4'ha):(1'h0)] reg1917 = (1'h0);
  reg [(3'h4):(1'h0)] reg1918 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1919 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1920 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1921 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire1922;
  wire [(2'h2):(1'h0)] wire2667;
  assign y = {wire2671,
                 wire2670,
                 wire2669,
                 wire1145,
                 wire590,
                 wire1147,
                 reg1148,
                 forvar1149,
                 reg1150,
                 reg1151,
                 reg1152,
                 reg1153,
                 reg1154,
                 reg1155,
                 reg1156,
                 reg1157,
                 forvar1158,
                 reg1159,
                 reg1160,
                 reg1161,
                 reg1149,
                 forvar1150,
                 forvar1156,
                 reg1158,
                 forvar1162,
                 forvar1163,
                 reg1164,
                 forvar1165,
                 reg1166,
                 forvar1167,
                 reg1168,
                 reg1169,
                 reg1170,
                 forvar1151,
                 forvar1153,
                 reg1163,
                 reg1165,
                 forvar1166,
                 reg1167,
                 forvar1171,
                 reg1172,
                 reg1173,
                 reg1174,
                 reg1175,
                 reg1176,
                 forvar1177,
                 reg1178,
                 forvar1179,
                 forvar1180,
                 reg1181,
                 reg1182,
                 reg1183,
                 reg1184,
                 reg1185,
                 reg1186,
                 reg1187,
                 forvar1178,
                 reg1179,
                 reg1180,
                 forvar1183,
                 forvar1186,
                 forvar1188,
                 reg1189,
                 reg1190,
                 reg1191,
                 forvar1192,
                 reg1193,
                 reg1194,
                 reg1195,
                 forvar1152,
                 forvar1154,
                 forvar1157,
                 forvar1159,
                 reg1162,
                 forvar1161,
                 forvar1168,
                 forvar1169,
                 reg1171,
                 reg1177,
                 forvar1148,
                 forvar1196,
                 forvar1197,
                 reg1198,
                 reg1199,
                 reg1200,
                 reg1201,
                 reg1202,
                 reg1203,
                 reg1204,
                 forvar1205,
                 reg1206,
                 reg1207,
                 reg1208,
                 reg1209,
                 reg1210,
                 reg1211,
                 reg1212,
                 forvar1213,
                 reg1214,
                 reg1215,
                 reg1205,
                 forvar1207,
                 reg1216,
                 reg1217,
                 reg1218,
                 reg1219,
                 reg1220,
                 reg1221,
                 forvar1216,
                 forvar1218,
                 reg1222,
                 reg1197,
                 forvar1202,
                 forvar1209,
                 reg1213,
                 forvar1214,
                 forvar1219,
                 forvar1221,
                 forvar1201,
                 reg1196,
                 forvar1210,
                 forvar1212,
                 forvar1223,
                 reg1224,
                 reg1225,
                 reg1226,
                 reg1227,
                 reg1228,
                 reg1229,
                 reg1230,
                 reg1231,
                 forvar1232,
                 reg1233,
                 reg1234,
                 reg1235,
                 reg1236,
                 reg1237,
                 forvar1238,
                 reg1239,
                 reg1240,
                 reg1241,
                 reg1242,
                 forvar1243,
                 reg1244,
                 reg1245,
                 reg1246,
                 reg1247,
                 reg1248,
                 reg1249,
                 reg1250,
                 reg1251,
                 reg1252,
                 reg1238,
                 reg1243,
                 forvar1246,
                 forvar1251,
                 reg1253,
                 reg1254,
                 reg1255,
                 forvar1256,
                 reg1257,
                 reg1258,
                 reg1259,
                 reg1260,
                 reg1261,
                 forvar1262,
                 reg1263,
                 reg1264,
                 reg1265,
                 reg1266,
                 reg1267,
                 reg1268,
                 reg1269,
                 reg1270,
                 reg1271,
                 forvar1265,
                 forvar1229,
                 reg1232,
                 forvar1272,
                 forvar1273,
                 forvar1274,
                 reg1275,
                 reg1276,
                 reg1277,
                 reg1278,
                 reg1279,
                 reg1280,
                 forvar1281,
                 forvar1282,
                 reg1283,
                 reg1284,
                 forvar1285,
                 reg1286,
                 reg1287,
                 reg1288,
                 reg1289,
                 reg1290,
                 forvar1291,
                 reg1292,
                 reg1293,
                 reg1294,
                 forvar1295,
                 reg1296,
                 reg1297,
                 forvar1290,
                 reg1291,
                 forvar1298,
                 forvar1299,
                 reg1300,
                 reg1301,
                 reg1302,
                 reg1303,
                 reg1304,
                 forvar1305,
                 reg1306,
                 reg1307,
                 reg1308,
                 reg1309,
                 forvar1310,
                 reg1311,
                 reg1312,
                 reg1313,
                 reg1305,
                 forvar1306,
                 reg1310,
                 forvar1314,
                 reg1315,
                 reg1316,
                 reg1314,
                 reg1317,
                 reg1318,
                 reg1319,
                 reg1320,
                 reg1321,
                 reg1322,
                 forvar1323,
                 reg1324,
                 reg1325,
                 reg1326,
                 reg1323,
                 reg1327,
                 forvar1304,
                 forvar1309,
                 reg1328,
                 reg1329,
                 reg1330,
                 reg1331,
                 forvar1332,
                 reg1333,
                 forvar1334,
                 reg1335,
                 reg1336,
                 reg1337,
                 reg1338,
                 reg1339,
                 reg1340,
                 reg1341,
                 reg1342,
                 reg1343,
                 reg1344,
                 reg1345,
                 forvar1341,
                 reg1346,
                 reg1347,
                 reg1348,
                 reg1349,
                 forvar1350,
                 reg1351,
                 reg1352,
                 reg1353,
                 reg1354,
                 reg1355,
                 reg1356,
                 reg1357,
                 reg1358,
                 forvar1348,
                 reg1350,
                 forvar1351,
                 forvar1354,
                 reg1359,
                 reg1360,
                 reg1361,
                 reg1362,
                 forvar1363,
                 reg1364,
                 forvar1365,
                 reg1366,
                 reg1367,
                 forvar1328,
                 forvar1330,
                 reg1332,
                 reg1334,
                 forvar1337,
                 forvar1224,
                 forvar1228,
                 forvar1231,
                 forvar1233,
                 reg1223,
                 forvar1226,
                 forvar1239,
                 forvar1241,
                 forvar1247,
                 forvar1248,
                 forvar1250,
                 forvar1252,
                 reg1256,
                 forvar1258,
                 forvar1259,
                 forvar1261,
                 reg1262,
                 forvar1260,
                 forvar1264,
                 forvar1269,
                 forvar1271,
                 reg1272,
                 reg1273,
                 reg1274,
                 forvar1368,
                 reg1369,
                 reg1370,
                 reg1371,
                 reg1372,
                 reg1373,
                 reg1374,
                 reg1375,
                 reg1376,
                 reg1377,
                 forvar1378,
                 reg1379,
                 reg1380,
                 reg1381,
                 reg1382,
                 reg1383,
                 forvar1373,
                 reg1378,
                 forvar1370,
                 forvar1371,
                 forvar1384,
                 reg1385,
                 reg1386,
                 reg1387,
                 reg1388,
                 reg1389,
                 reg1390,
                 reg1384,
                 forvar1391,
                 reg1392,
                 forvar1393,
                 forvar1394,
                 reg1395,
                 reg1396,
                 reg1397,
                 reg1398,
                 reg1394,
                 forvar1395,
                 reg1399,
                 reg1400,
                 reg1401,
                 reg1402,
                 forvar1403,
                 reg1404,
                 reg1405,
                 reg1406,
                 reg1407,
                 forvar1408,
                 forvar1409,
                 reg1410,
                 reg1411,
                 reg1412,
                 forvar1413,
                 forvar1414,
                 reg1415,
                 reg1416,
                 reg1417,
                 reg1418,
                 forvar1419,
                 reg1420,
                 reg1421,
                 reg1422,
                 reg1423,
                 forvar1424,
                 reg1425,
                 forvar1426,
                 reg1427,
                 forvar1428,
                 reg1429,
                 forvar1430,
                 reg1431,
                 reg1432,
                 forvar1433,
                 reg1434,
                 reg1435,
                 reg1436,
                 reg1437,
                 reg1438,
                 reg1439,
                 reg1440,
                 forvar1438,
                 reg1441,
                 reg1442,
                 forvar1443,
                 reg1444,
                 reg1445,
                 forvar1446,
                 reg1447,
                 forvar1448,
                 reg1449,
                 reg1450,
                 reg1446,
                 reg1448,
                 reg1451,
                 forvar1450,
                 reg1452,
                 reg1453,
                 forvar1454,
                 reg1455,
                 forvar1456,
                 reg1457,
                 reg1458,
                 reg1459,
                 reg1460,
                 reg1461,
                 forvar1462,
                 forvar1463,
                 reg1464,
                 reg1465,
                 reg1466,
                 reg1467,
                 reg1468,
                 forvar1469,
                 reg1470,
                 reg1471,
                 forvar1472,
                 reg1473,
                 reg1474,
                 reg1475,
                 reg1476,
                 reg1477,
                 reg1478,
                 reg1479,
                 forvar1480,
                 reg1481,
                 reg1482,
                 reg1469,
                 reg1472,
                 forvar1479,
                 reg1480,
                 reg1483,
                 forvar1484,
                 reg1485,
                 reg1486,
                 reg1487,
                 forvar1488,
                 reg1489,
                 reg1490,
                 reg1484,
                 reg1491,
                 reg1492,
                 reg1493,
                 reg1494,
                 forvar1495,
                 reg1496,
                 reg1497,
                 reg1498,
                 reg1499,
                 forvar1500,
                 reg1501,
                 reg1502,
                 reg1495,
                 forvar1496,
                 reg1503,
                 forvar1504,
                 reg1505,
                 reg1506,
                 reg1507,
                 reg1508,
                 reg1504,
                 wire1735,
                 forvar1737,
                 reg1738,
                 forvar1739,
                 forvar1740,
                 forvar1741,
                 reg1742,
                 reg1743,
                 reg1744,
                 reg1745,
                 forvar1746,
                 reg1747,
                 reg1748,
                 reg1749,
                 reg1750,
                 reg1751,
                 reg1752,
                 reg1753,
                 forvar1754,
                 forvar1755,
                 reg1756,
                 reg1757,
                 reg1758,
                 reg1759,
                 forvar1760,
                 reg1761,
                 reg1762,
                 reg1763,
                 reg1764,
                 forvar1765,
                 reg1766,
                 reg1767,
                 forvar1768,
                 reg1769,
                 reg1770,
                 reg1771,
                 forvar1772,
                 reg1773,
                 reg1774,
                 reg1775,
                 forvar1776,
                 reg1777,
                 reg1778,
                 reg1779,
                 reg1780,
                 forvar1781,
                 reg1782,
                 reg1783,
                 reg1784,
                 reg1785,
                 forvar1786,
                 reg1787,
                 reg1788,
                 reg1789,
                 forvar1790,
                 reg1791,
                 forvar1792,
                 reg1793,
                 reg1794,
                 reg1795,
                 reg1796,
                 reg1797,
                 reg1798,
                 reg1799,
                 reg1800,
                 reg1801,
                 forvar1802,
                 reg1803,
                 reg1804,
                 reg1805,
                 reg1806,
                 reg1807,
                 reg1808,
                 forvar1809,
                 reg1810,
                 reg1811,
                 reg1812,
                 forvar1813,
                 reg1814,
                 reg1815,
                 reg1816,
                 reg1817,
                 reg1813,
                 forvar1816,
                 reg1818,
                 reg1819,
                 reg1820,
                 forvar1803,
                 forvar1807,
                 forvar1808,
                 reg1809,
                 forvar1821,
                 forvar1822,
                 reg1823,
                 reg1824,
                 reg1825,
                 reg1826,
                 reg1827,
                 reg1828,
                 reg1829,
                 reg1830,
                 forvar1831,
                 reg1832,
                 reg1833,
                 reg1834,
                 reg1831,
                 reg1835,
                 forvar1836,
                 forvar1837,
                 reg1838,
                 reg1839,
                 forvar1828,
                 forvar1830,
                 forvar1835,
                 reg1836,
                 reg1837,
                 forvar1839,
                 reg1840,
                 reg1841,
                 reg1842,
                 forvar1840,
                 reg1843,
                 forvar1844,
                 reg1845,
                 reg1846,
                 reg1844,
                 reg1847,
                 reg1848,
                 reg1849,
                 reg1850,
                 forvar1833,
                 forvar1851,
                 reg1852,
                 forvar1853,
                 reg1854,
                 reg1855,
                 reg1856,
                 reg1857,
                 reg1858,
                 reg1859,
                 reg1860,
                 reg1861,
                 reg1862,
                 reg1863,
                 reg1864,
                 reg1865,
                 reg1866,
                 reg1867,
                 reg1868,
                 forvar1863,
                 forvar1869,
                 forvar1870,
                 reg1871,
                 forvar1872,
                 reg1873,
                 forvar1874,
                 reg1875,
                 reg1876,
                 forvar1877,
                 forvar1878,
                 forvar1879,
                 reg1880,
                 reg1881,
                 reg1882,
                 reg1883,
                 forvar1884,
                 reg1885,
                 reg1886,
                 reg1887,
                 reg1888,
                 forvar1889,
                 reg1890,
                 forvar1891,
                 reg1892,
                 reg1893,
                 reg1894,
                 reg1895,
                 reg1896,
                 reg1897,
                 forvar1898,
                 reg1899,
                 reg1900,
                 reg1901,
                 reg1902,
                 reg1903,
                 reg1904,
                 reg1905,
                 reg1906,
                 reg1907,
                 reg1908,
                 reg1909,
                 reg1910,
                 forvar1911,
                 reg1912,
                 reg1913,
                 forvar1914,
                 forvar1915,
                 forvar1916,
                 reg1917,
                 reg1918,
                 reg1919,
                 reg1920,
                 reg1921,
                 wire1922,
                 wire2667,
                 (1'h0)};
  assign wire590 = (^~(8'hba));
  module591 modinst1146 (wire1145, clk, wire585, wire589, wire586, wire590, wire588);
  assign wire1147 = wire589[(4'h8):(1'h1)];
  always
    @(posedge clk) begin
      if (($signed($signed($signed(wire588))) ?
          (|wire586[(4'ha):(4'h9)]) : {(!{(8'ha1)})}))
        begin
          if (wire590[(3'h5):(3'h5)])
            begin
              reg1148 <= wire590[(1'h0):(1'h0)];
              if ($signed((^~(~&(~|wire588)))))
                begin
                  for (forvar1149 = (1'h0); (forvar1149 < (2'h3)); forvar1149 = (forvar1149 + (1'h1)))
                    begin
                      reg1150 <= ((8'hb2) <<< ((wire586[(3'h5):(1'h0)] && (wire1145 < wire586)) >>> ({wire585} ?
                          (8'ha2) : (~wire1147))));
                      reg1151 <= (wire1147 >>> (|$unsigned((wire586 ?
                          wire585 : wire588))));
                      reg1152 <= ((8'hb6) ?
                          ((&$unsigned(forvar1149)) >> (~|{wire1145})) : wire588);
                      reg1153 <= $signed($unsigned(wire1145));
                    end
                  if ($unsigned($unsigned((wire1145[(3'h4):(3'h4)] + wire589[(2'h3):(1'h1)]))))
                    begin
                      reg1154 <= {(&((reg1151 ?
                              reg1151 : reg1148) <= (wire586 >= reg1152)))};
                      reg1155 <= $signed($signed(((reg1153 ^~ wire588) > (~&reg1151))));
                      reg1156 <= (wire1147 & (reg1153 + $signed((reg1152 << forvar1149))));
                      reg1157 <= {((-(reg1155 ? (8'ha2) : wire590)) ?
                              $signed($unsigned(wire590)) : ($signed(reg1150) << $signed(forvar1149)))};
                    end
                  else
                    begin
                      reg1154 <= (($signed((~^reg1148)) ?
                          reg1152[(1'h0):(1'h0)] : (reg1156 >>> (-wire589))) < $signed(wire1145));
                      reg1155 <= forvar1149;
                      reg1156 <= ((+{$unsigned(wire587)}) ?
                          ($unsigned(wire589[(2'h3):(1'h1)]) ?
                              reg1157[(3'h4):(1'h1)] : $signed($signed(reg1150))) : reg1152[(3'h4):(2'h2)]);
                    end
                  for (forvar1158 = (1'h0); (forvar1158 < (2'h2)); forvar1158 = (forvar1158 + (1'h1)))
                    begin
                      reg1159 <= ((wire590[(2'h2):(1'h1)] ?
                              $signed({reg1151}) : (reg1155 != $unsigned(wire1147))) ?
                          wire587[(2'h3):(1'h1)] : (~^(^~wire1147[(4'hc):(4'h9)])));
                      reg1160 <= (+(forvar1158 ?
                          {(reg1152 ? reg1159 : (8'ha9))} : $signed(wire1145)));
                    end
                  if ($signed($unsigned($signed((reg1157 ?
                      wire589 : wire586)))))
                    begin
                      reg1161 <= wire1145[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg1161 <= $signed(reg1156[(2'h3):(2'h3)]);
                    end
                end
              else
                begin
                  if ((wire1147 >>> (&$unsigned((wire588 ?
                      reg1154 : wire590)))))
                    begin
                      reg1149 <= $signed($signed($unsigned((reg1150 > reg1157))));
                    end
                  else
                    begin
                      reg1149 <= $unsigned(reg1151[(3'h6):(3'h4)]);
                    end
                  for (forvar1150 = (1'h0); (forvar1150 < (2'h3)); forvar1150 = (forvar1150 + (1'h1)))
                    begin
                      reg1151 <= reg1151[(3'h4):(2'h3)];
                      reg1152 <= $signed(reg1156);
                      reg1153 <= (wire589[(4'hc):(3'h7)] ?
                          $unsigned($unsigned($signed(wire585))) : reg1155);
                      reg1154 <= ({{$unsigned((8'hb8))}} ?
                          forvar1150[(1'h1):(1'h0)] : {wire586});
                    end
                  reg1155 <= $signed(($signed((8'hb4)) - ($signed(reg1159) ?
                      $signed(wire587) : (wire588 * (8'h9e)))));
                  for (forvar1156 = (1'h0); (forvar1156 < (2'h3)); forvar1156 = (forvar1156 + (1'h1)))
                    begin
                      reg1157 <= ((~^{reg1148[(2'h3):(2'h3)]}) != (~reg1161[(3'h5):(2'h2)]));
                      reg1158 <= wire1147;
                      reg1159 <= reg1161[(3'h4):(1'h1)];
                      reg1160 <= reg1157[(1'h0):(1'h0)];
                    end
                end
              for (forvar1162 = (1'h0); (forvar1162 < (2'h3)); forvar1162 = (forvar1162 + (1'h1)))
                begin
                  for (forvar1163 = (1'h0); (forvar1163 < (2'h3)); forvar1163 = (forvar1163 + (1'h1)))
                    begin
                      reg1164 <= reg1149;
                    end
                  for (forvar1165 = (1'h0); (forvar1165 < (2'h3)); forvar1165 = (forvar1165 + (1'h1)))
                    begin
                      reg1166 <= ((^forvar1158) >= $unsigned(wire587[(4'ha):(4'ha)]));
                    end
                  for (forvar1167 = (1'h0); (forvar1167 < (1'h1)); forvar1167 = (forvar1167 + (1'h1)))
                    begin
                      reg1168 <= forvar1158;
                    end
                  if ((((+forvar1149) ?
                          (|(wire588 ? reg1164 : reg1164)) : (((8'had) ?
                              forvar1163 : (8'hb4)) + $signed(wire587))) ?
                      wire589 : $unsigned({(~^reg1161)})))
                    begin
                      reg1169 <= $unsigned(($signed(forvar1149) ?
                          $signed(wire590) : $unsigned(wire590[(3'h5):(2'h2)])));
                      reg1170 <= forvar1163[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg1169 <= $unsigned(($unsigned((forvar1158 ?
                          wire589 : reg1151)) >>> (+forvar1165)));
                      reg1170 <= {$unsigned((-$signed(wire1145)))};
                    end
                end
            end
          else
            begin
              reg1148 <= wire588;
              for (forvar1149 = (1'h0); (forvar1149 < (1'h0)); forvar1149 = (forvar1149 + (1'h1)))
                begin
                  reg1150 <= {reg1157};
                  for (forvar1151 = (1'h0); (forvar1151 < (1'h0)); forvar1151 = (forvar1151 + (1'h1)))
                    begin
                      reg1152 <= $signed(($unsigned(reg1164) ?
                          forvar1165 : {$signed(reg1169)}));
                    end
                  for (forvar1153 = (1'h0); (forvar1153 < (1'h0)); forvar1153 = (forvar1153 + (1'h1)))
                    begin
                      reg1154 <= (&(^{$unsigned(forvar1167)}));
                      reg1155 <= ($signed(((reg1150 ? reg1156 : (8'h9f)) ?
                          reg1154[(3'h4):(1'h1)] : $unsigned((8'hb0)))) <<< reg1155[(3'h6):(2'h3)]);
                      reg1156 <= (~&((~^(reg1161 ?
                          forvar1162 : reg1157)) ~^ {(forvar1156 >> reg1161)}));
                      reg1157 <= ($unsigned($signed(reg1164[(2'h2):(1'h1)])) || ((reg1161[(3'h5):(3'h5)] << forvar1156[(4'hb):(1'h1)]) == ({reg1160} ?
                          wire589 : wire588)));
                    end
                  if ({reg1154[(3'h4):(1'h0)]})
                    begin
                      reg1158 <= (^$signed((forvar1163 ?
                          (~|reg1151) : (reg1148 + wire589))));
                      reg1159 <= ((&{$signed(forvar1158)}) <<< {reg1150[(4'hb):(1'h0)]});
                      reg1160 <= $unsigned(wire1147[(2'h3):(2'h3)]);
                      reg1161 <= reg1164[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg1158 <= $unsigned($unsigned($unsigned($signed(reg1164))));
                      reg1159 <= {$signed((~^(-reg1159)))};
                    end
                end
              if (($signed(((~&reg1150) && reg1153)) <= reg1164[(3'h4):(2'h3)]))
                begin
                  for (forvar1162 = (1'h0); (forvar1162 < (1'h1)); forvar1162 = (forvar1162 + (1'h1)))
                    begin
                      reg1163 <= (($signed(reg1166[(2'h2):(1'h1)]) >>> $signed(forvar1158[(3'h5):(3'h4)])) ?
                          (|reg1153) : reg1154);
                    end
                  if (((((forvar1162 ? (8'ha9) : reg1169) & $signed(reg1153)) ?
                          wire588 : $unsigned((^~(8'h9d)))) ?
                      (~^(forvar1151[(4'h8):(3'h5)] ?
                          forvar1153 : $unsigned(reg1148))) : ($signed({reg1169}) ~^ reg1150)))
                    begin
                      reg1164 <= (|{(^~{reg1149})});
                    end
                  else
                    begin
                      reg1164 <= (reg1166 ?
                          $unsigned((8'hb5)) : $unsigned(wire590[(2'h2):(2'h2)]));
                      reg1165 <= wire590;
                    end
                  for (forvar1166 = (1'h0); (forvar1166 < (2'h2)); forvar1166 = (forvar1166 + (1'h1)))
                    begin
                      reg1167 <= {wire585[(3'h6):(3'h5)]};
                    end
                end
              else
                begin
                  for (forvar1162 = (1'h0); (forvar1162 < (2'h2)); forvar1162 = (forvar1162 + (1'h1)))
                    begin
                      reg1163 <= (wire586 ?
                          reg1161[(2'h3):(1'h1)] : (-$signed($unsigned(forvar1166))));
                      reg1164 <= $unsigned($unsigned((wire587 >= $unsigned(reg1148))));
                    end
                  for (forvar1165 = (1'h0); (forvar1165 < (2'h2)); forvar1165 = (forvar1165 + (1'h1)))
                    begin
                      reg1166 <= ({reg1168[(2'h3):(1'h1)]} >> $signed($unsigned($unsigned(wire1147))));
                      reg1167 <= (~|((|(reg1159 < wire585)) ?
                          (wire1147 >> (reg1154 * forvar1167)) : $unsigned((wire587 >> reg1156))));
                      reg1168 <= $signed({($signed((8'ha4)) ?
                              $unsigned(reg1150) : ((8'hb3) + reg1157))});
                    end
                  reg1169 <= ({wire1145[(2'h2):(1'h1)]} > reg1148[(1'h1):(1'h1)]);
                end
            end
          for (forvar1171 = (1'h0); (forvar1171 < (1'h1)); forvar1171 = (forvar1171 + (1'h1)))
            begin
              if (($unsigned({$unsigned(reg1158)}) ?
                  (((&forvar1149) ?
                      $unsigned(wire1145) : (~wire588)) >= ((forvar1153 ?
                          reg1156 : wire590) ?
                      (reg1167 - (8'ha4)) : $signed(wire585))) : {wire589}))
                begin
                  reg1172 <= $unsigned($signed($signed((reg1159 ?
                      wire587 : wire585))));
                end
              else
                begin
                  reg1172 <= $signed((^~{(reg1152 - forvar1167)}));
                  if ($unsigned(forvar1151))
                    begin
                      reg1173 <= (wire586 ? (8'hab) : (~|wire589));
                      reg1174 <= reg1168;
                      reg1175 <= {forvar1162};
                      reg1176 <= forvar1171[(4'hc):(2'h3)];
                    end
                  else
                    begin
                      reg1173 <= $signed(((+(reg1150 >>> wire1147)) ?
                          ((^(8'ha3)) ?
                              (reg1175 >>> reg1154) : ((8'hb3) << reg1173)) : $unsigned((forvar1153 ?
                              reg1158 : forvar1163))));
                    end
                end
            end
          if ((&$unsigned(wire590[(3'h5):(2'h2)])))
            begin
              for (forvar1177 = (1'h0); (forvar1177 < (1'h1)); forvar1177 = (forvar1177 + (1'h1)))
                begin
                  reg1178 <= (reg1158 >> $unsigned(reg1158));
                end
              for (forvar1179 = (1'h0); (forvar1179 < (2'h3)); forvar1179 = (forvar1179 + (1'h1)))
                begin
                  for (forvar1180 = (1'h0); (forvar1180 < (1'h1)); forvar1180 = (forvar1180 + (1'h1)))
                    begin
                      reg1181 <= ({reg1153[(4'hb):(3'h5)]} == reg1161[(3'h4):(2'h3)]);
                      reg1182 <= $unsigned(reg1160[(3'h7):(1'h0)]);
                      reg1183 <= $unsigned($unsigned(forvar1156[(4'ha):(4'h8)]));
                    end
                  if ($signed(wire1147[(4'h8):(2'h3)]))
                    begin
                      reg1184 <= reg1163[(2'h2):(2'h2)];
                      reg1185 <= {{$signed((~|reg1181))}};
                      reg1186 <= (|{$signed(reg1157[(4'h8):(4'h8)])});
                    end
                  else
                    begin
                      reg1184 <= (reg1178 ?
                          reg1182[(1'h0):(1'h0)] : (({forvar1163} ^ $unsigned(reg1155)) >= (reg1176 ^~ {(8'ha5)})));
                      reg1185 <= (((~{forvar1180}) ?
                              ($unsigned((8'ha1)) >= (8'ha9)) : $signed(((8'hb0) ?
                                  reg1153 : reg1173))) ?
                          $signed((^~$unsigned(reg1168))) : (((|reg1185) << $signed((8'hab))) ?
                              $signed(reg1181) : $unsigned(reg1148)));
                      reg1186 <= {forvar1167[(1'h0):(1'h0)]};
                      reg1187 <= $unsigned((~forvar1158));
                    end
                end
            end
          else
            begin
              for (forvar1177 = (1'h0); (forvar1177 < (2'h2)); forvar1177 = (forvar1177 + (1'h1)))
                begin
                  for (forvar1178 = (1'h0); (forvar1178 < (1'h1)); forvar1178 = (forvar1178 + (1'h1)))
                    begin
                      reg1179 <= ($signed(reg1164) ^ $unsigned((&(forvar1166 | forvar1180))));
                      reg1180 <= reg1175[(3'h6):(3'h4)];
                      reg1181 <= reg1154[(2'h2):(1'h1)];
                      reg1182 <= $signed((forvar1158 ?
                          reg1166 : $signed($unsigned(reg1160))));
                    end
                  for (forvar1183 = (1'h0); (forvar1183 < (2'h2)); forvar1183 = (forvar1183 + (1'h1)))
                    begin
                      reg1184 <= (wire1145[(2'h3):(2'h2)] ?
                          reg1174[(2'h2):(1'h1)] : (($unsigned(forvar1156) + ((8'ha7) ?
                              wire1147 : reg1160)) < reg1183[(2'h3):(1'h0)]));
                      reg1185 <= $signed($unsigned(reg1179[(3'h4):(1'h1)]));
                    end
                end
              for (forvar1186 = (1'h0); (forvar1186 < (1'h0)); forvar1186 = (forvar1186 + (1'h1)))
                begin
                  reg1187 <= forvar1171[(4'hc):(2'h3)];
                  for (forvar1188 = (1'h0); (forvar1188 < (2'h3)); forvar1188 = (forvar1188 + (1'h1)))
                    begin
                      reg1189 <= wire586[(2'h2):(2'h2)];
                      reg1190 <= {$signed({$unsigned(reg1185)})};
                      reg1191 <= ($unsigned(reg1158) ?
                          (|((forvar1151 ? (8'haf) : reg1180) ?
                              $unsigned(wire586) : (reg1175 ?
                                  reg1181 : wire1145))) : forvar1165[(1'h1):(1'h0)]);
                    end
                end
              for (forvar1192 = (1'h0); (forvar1192 < (2'h3)); forvar1192 = (forvar1192 + (1'h1)))
                begin
                  if (reg1186[(3'h4):(2'h3)])
                    begin
                      reg1193 <= (reg1168 ^~ reg1156);
                      reg1194 <= forvar1158;
                    end
                  else
                    begin
                      reg1193 <= (reg1185[(1'h1):(1'h0)] >= $unsigned(({forvar1150} + reg1187[(1'h0):(1'h0)])));
                    end
                end
              reg1195 <= forvar1150;
            end
        end
      else
        begin
          if (reg1153[(4'hd):(1'h0)])
            begin
              if ($signed(reg1165))
                begin
                  if (($signed($signed($signed(reg1152))) ?
                      $signed($unsigned((8'hb4))) : reg1183))
                    begin
                      reg1148 <= reg1155[(1'h1):(1'h1)];
                      reg1149 <= ((($unsigned((8'hb4)) ?
                                  $signed(reg1180) : {reg1178}) ?
                              forvar1178 : (~&forvar1177[(3'h6):(3'h6)])) ?
                          ({$unsigned(forvar1178)} ?
                              (^(+reg1157)) : (^~(reg1161 ?
                                  reg1161 : reg1179))) : ((reg1184[(2'h3):(1'h1)] ?
                                  (8'ha7) : (forvar1179 && forvar1165)) ?
                              $signed(reg1170[(3'h6):(1'h1)]) : (+(reg1182 ?
                                  reg1150 : (8'haa)))));
                    end
                  else
                    begin
                      reg1148 <= reg1169[(3'h6):(2'h3)];
                    end
                end
              else
                begin
                  reg1148 <= reg1180[(3'h4):(2'h2)];
                end
              for (forvar1150 = (1'h0); (forvar1150 < (2'h2)); forvar1150 = (forvar1150 + (1'h1)))
                begin
                  reg1151 <= {reg1170};
                  for (forvar1152 = (1'h0); (forvar1152 < (2'h3)); forvar1152 = (forvar1152 + (1'h1)))
                    begin
                      reg1153 <= (($unsigned(forvar1156[(4'h8):(2'h3)]) ?
                              reg1155[(1'h0):(1'h0)] : reg1170) ?
                          forvar1165 : $signed({$signed(wire588)}));
                    end
                  for (forvar1154 = (1'h0); (forvar1154 < (2'h3)); forvar1154 = (forvar1154 + (1'h1)))
                    begin
                      reg1155 <= reg1195[(4'hb):(4'hb)];
                      reg1156 <= forvar1156;
                    end
                end
              if ($signed(forvar1192[(2'h2):(1'h0)]))
                begin
                  for (forvar1157 = (1'h0); (forvar1157 < (1'h0)); forvar1157 = (forvar1157 + (1'h1)))
                    begin
                      reg1158 <= reg1170[(3'h5):(1'h1)];
                    end
                  for (forvar1159 = (1'h0); (forvar1159 < (2'h2)); forvar1159 = (forvar1159 + (1'h1)))
                    begin
                      reg1160 <= reg1160[(3'h5):(1'h1)];
                      reg1161 <= ((forvar1171[(4'hd):(4'h9)] ?
                          (&$signed(reg1183)) : $unsigned(wire588)) >> reg1156);
                      reg1162 <= reg1178;
                      reg1163 <= ((~&$signed($unsigned(reg1170))) ?
                          ($unsigned($unsigned(wire1147)) ?
                              reg1156 : {$signed(reg1186)}) : (~^((forvar1157 ?
                              reg1153 : reg1172) << ((8'had) ?
                              forvar1179 : reg1157))));
                    end
                  if ((($signed((-reg1178)) ^~ (|$signed(wire588))) <<< $signed($signed((reg1149 ?
                      reg1172 : reg1169)))))
                    begin
                      reg1164 <= ((({forvar1153} <= ((8'h9d) + forvar1153)) != ((~|reg1161) >= reg1168[(3'h4):(1'h1)])) ?
                          ($unsigned($unsigned(wire1145)) ~^ forvar1153) : reg1157);
                      reg1165 <= reg1155[(4'hb):(3'h7)];
                      reg1166 <= reg1169[(3'h7):(3'h7)];
                    end
                  else
                    begin
                      reg1164 <= $unsigned($signed(((~^reg1194) ?
                          wire588 : reg1179[(2'h2):(2'h2)])));
                      reg1165 <= $unsigned($unsigned(reg1184));
                      reg1166 <= ((((reg1191 <<< reg1174) > reg1156[(1'h0):(1'h0)]) - forvar1163) + $signed(({reg1182} ?
                          $signed(reg1184) : forvar1150[(1'h1):(1'h1)])));
                      reg1167 <= wire588;
                    end
                end
              else
                begin
                  if ((~({(reg1153 ?
                          forvar1153 : (8'ha2))} == $unsigned(reg1158[(3'h7):(2'h2)]))))
                    begin
                      reg1157 <= $unsigned(reg1179);
                      reg1158 <= ($signed(((forvar1149 ? (8'ha5) : forvar1162) ?
                              (wire1147 ?
                                  (8'hb7) : forvar1167) : reg1184[(2'h3):(1'h0)])) ?
                          (|((reg1189 + reg1180) ?
                              reg1185 : (reg1189 <<< reg1190))) : (((forvar1163 | reg1172) ?
                                  (~^forvar1153) : $unsigned(reg1151)) ?
                              $unsigned(forvar1159) : $unsigned($signed(reg1185))));
                      reg1159 <= $signed($signed(((reg1157 ?
                              (8'hb6) : reg1169) ?
                          (reg1179 + wire590) : (-reg1169))));
                      reg1160 <= $unsigned({(&{(8'ha4)})});
                    end
                  else
                    begin
                      reg1157 <= $unsigned((~&forvar1178[(3'h4):(1'h0)]));
                      reg1158 <= $signed((^~((^~reg1189) + {forvar1192})));
                      reg1159 <= $signed(reg1166[(3'h6):(2'h2)]);
                      reg1160 <= ($unsigned({(+reg1168)}) ?
                          (reg1186[(3'h5):(3'h4)] ?
                              ($unsigned(reg1158) * $unsigned(reg1175)) : (8'hae)) : reg1164);
                    end
                  for (forvar1161 = (1'h0); (forvar1161 < (1'h1)); forvar1161 = (forvar1161 + (1'h1)))
                    begin
                      reg1162 <= reg1190;
                      reg1163 <= $unsigned($unsigned(forvar1156[(1'h0):(1'h0)]));
                      reg1164 <= $unsigned($signed(($signed(forvar1178) >> (reg1185 >> reg1170))));
                      reg1165 <= forvar1178;
                    end
                end
              for (forvar1168 = (1'h0); (forvar1168 < (2'h3)); forvar1168 = (forvar1168 + (1'h1)))
                begin
                  for (forvar1169 = (1'h0); (forvar1169 < (2'h2)); forvar1169 = (forvar1169 + (1'h1)))
                    begin
                      reg1170 <= forvar1163;
                      reg1171 <= (&reg1175[(2'h2):(1'h1)]);
                      reg1172 <= reg1191[(3'h6):(2'h3)];
                      reg1173 <= $unsigned(reg1172);
                    end
                  reg1174 <= ($signed(forvar1159) != forvar1165[(3'h7):(2'h2)]);
                  reg1175 <= wire590;
                  if (((reg1184[(3'h4):(2'h3)] ?
                      (8'hb0) : ((|reg1189) ?
                          $unsigned(reg1183) : wire588[(3'h6):(3'h6)])) < ($signed(reg1180) != ((8'hb3) ?
                      (reg1153 ? reg1166 : reg1152) : $unsigned(reg1191)))))
                    begin
                      reg1176 <= (|(^((~^(8'hb2)) <= (reg1155 >>> forvar1167))));
                      reg1177 <= $signed((reg1155[(1'h0):(1'h0)] ?
                          $signed({(8'hb6)}) : ($signed(forvar1165) < forvar1180[(4'hb):(4'h8)])));
                      reg1178 <= ($unsigned($unsigned(wire587)) + reg1189[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1176 <= reg1160;
                    end
                end
            end
          else
            begin
              for (forvar1148 = (1'h0); (forvar1148 < (1'h0)); forvar1148 = (forvar1148 + (1'h1)))
                begin
                  for (forvar1149 = (1'h0); (forvar1149 < (1'h1)); forvar1149 = (forvar1149 + (1'h1)))
                    begin
                      reg1150 <= ((reg1161[(1'h0):(1'h0)] ?
                              ({wire586} ?
                                  ((8'hb3) ?
                                      forvar1148 : reg1163) : $unsigned((8'had))) : reg1191) ?
                          (~|(8'haf)) : {{(reg1155 ?
                                      forvar1165 : forvar1156)}});
                      reg1151 <= ((8'hae) >>> reg1178[(3'h7):(3'h4)]);
                    end
                  reg1152 <= $unsigned({$signed($signed(forvar1171))});
                  for (forvar1153 = (1'h0); (forvar1153 < (1'h1)); forvar1153 = (forvar1153 + (1'h1)))
                    begin
                      reg1154 <= ($unsigned($signed($signed(reg1175))) ?
                          {($signed(reg1151) ?
                                  (forvar1163 ~^ (8'hb3)) : forvar1150[(1'h1):(1'h1)])} : $unsigned(forvar1157));
                      reg1155 <= forvar1152[(2'h2):(1'h0)];
                      reg1156 <= reg1162;
                      reg1157 <= reg1174[(3'h7):(2'h3)];
                    end
                end
            end
          reg1179 <= $unsigned($signed(((reg1181 - forvar1149) ?
              {forvar1179} : $unsigned(reg1177))));
        end
      if ((!forvar1161))
        begin
          for (forvar1196 = (1'h0); (forvar1196 < (1'h0)); forvar1196 = (forvar1196 + (1'h1)))
            begin
              for (forvar1197 = (1'h0); (forvar1197 < (2'h2)); forvar1197 = (forvar1197 + (1'h1)))
                begin
                  if ((8'ha7))
                    begin
                      reg1198 <= ((&($signed((8'ha8)) ^~ reg1176)) & reg1176[(2'h3):(2'h3)]);
                      reg1199 <= (($signed(reg1151[(2'h3):(2'h3)]) ?
                          $signed($signed(forvar1161)) : (~&$unsigned(reg1164))) && $signed((^~reg1191)));
                      reg1200 <= $signed((~|(~|(reg1165 ? reg1195 : (8'hb1)))));
                    end
                  else
                    begin
                      reg1198 <= (&reg1150);
                    end
                  reg1201 <= ($unsigned(((+forvar1166) ?
                          $unsigned(reg1174) : (-reg1177))) ?
                      {wire1147[(2'h2):(2'h2)]} : forvar1159);
                  if ({reg1162[(3'h7):(2'h2)]})
                    begin
                      reg1202 <= $signed((|$signed((~reg1151))));
                    end
                  else
                    begin
                      reg1202 <= (|reg1157);
                      reg1203 <= forvar1153[(4'hd):(4'hc)];
                      reg1204 <= {(~&$unsigned((forvar1166 ?
                              wire587 : forvar1178)))};
                    end
                end
              if ($signed((&reg1202)))
                begin
                  for (forvar1205 = (1'h0); (forvar1205 < (1'h1)); forvar1205 = (forvar1205 + (1'h1)))
                    begin
                      reg1206 <= (((-reg1187[(1'h1):(1'h1)]) ?
                          ((forvar1158 ?
                              reg1157 : forvar1159) != (~&wire586)) : forvar1205[(3'h6):(2'h3)]) != forvar1188[(3'h5):(1'h1)]);
                      reg1207 <= reg1150[(1'h0):(1'h0)];
                      reg1208 <= {($unsigned(wire587[(2'h3):(1'h1)]) < $unsigned(((8'hae) <= reg1159)))};
                      reg1209 <= wire1147;
                    end
                  if (reg1185[(2'h3):(1'h0)])
                    begin
                      reg1210 <= forvar1165;
                      reg1211 <= (!{{(reg1177 ^ forvar1165)}});
                    end
                  else
                    begin
                      reg1210 <= (~^forvar1157[(3'h5):(1'h0)]);
                    end
                  reg1212 <= ({(~|forvar1178[(1'h1):(1'h1)])} ?
                      (reg1149 == $signed(reg1154)) : $unsigned((!$unsigned(forvar1179))));
                  for (forvar1213 = (1'h0); (forvar1213 < (1'h0)); forvar1213 = (forvar1213 + (1'h1)))
                    begin
                      reg1214 <= wire590[(2'h2):(2'h2)];
                      reg1215 <= $signed((+$unsigned((reg1212 ?
                          reg1158 : forvar1166))));
                    end
                end
              else
                begin
                  reg1205 <= (forvar1163[(2'h2):(1'h1)] ^~ {((wire1147 >>> wire1145) ?
                          wire588 : (!reg1149))});
                  reg1206 <= (&wire590);
                  for (forvar1207 = (1'h0); (forvar1207 < (1'h0)); forvar1207 = (forvar1207 + (1'h1)))
                    begin
                      reg1208 <= $signed(reg1161[(3'h5):(1'h0)]);
                      reg1209 <= ((((reg1151 ? forvar1213 : (8'hba)) ?
                              reg1211 : reg1212[(1'h0):(1'h0)]) <= ($signed(reg1189) <= (+reg1183))) ?
                          forvar1213[(3'h7):(2'h3)] : $signed(wire587[(2'h3):(2'h3)]));
                      reg1210 <= $unsigned((^forvar1197));
                      reg1211 <= $signed($unsigned(forvar1154));
                    end
                  reg1212 <= $unsigned((|((forvar1197 ?
                      reg1162 : (8'hb0)) >> (reg1210 ? reg1210 : reg1176))));
                end
              if (reg1179[(1'h0):(1'h0)])
                begin
                  if (forvar1154[(1'h1):(1'h1)])
                    begin
                      reg1216 <= wire1145;
                      reg1217 <= $unsigned(reg1169[(4'h8):(3'h7)]);
                      reg1218 <= (|$signed(({reg1182} ?
                          {forvar1159} : (~|reg1165))));
                      reg1219 <= (+$signed(((!reg1153) - (~^(8'ha9)))));
                    end
                  else
                    begin
                      reg1216 <= (~|$signed($unsigned($unsigned(reg1208))));
                      reg1217 <= ((|(&(reg1160 >> (8'ha5)))) == ((forvar1180 ?
                              {(8'ha8)} : reg1184) ?
                          forvar1177[(3'h7):(1'h1)] : $signed((reg1161 <= forvar1188))));
                      reg1218 <= (forvar1177[(1'h1):(1'h0)] ?
                          $signed(forvar1177) : (reg1163 >>> {$unsigned(reg1166)}));
                      reg1219 <= (+((forvar1166 ?
                              reg1184[(2'h3):(1'h1)] : (|reg1181)) ?
                          wire1145 : forvar1188[(2'h2):(2'h2)]));
                    end
                  reg1220 <= forvar1171[(1'h1):(1'h0)];
                  reg1221 <= forvar1205[(1'h0):(1'h0)];
                end
              else
                begin
                  for (forvar1216 = (1'h0); (forvar1216 < (2'h2)); forvar1216 = (forvar1216 + (1'h1)))
                    begin
                      reg1217 <= $signed(forvar1148[(3'h6):(3'h6)]);
                    end
                  for (forvar1218 = (1'h0); (forvar1218 < (2'h3)); forvar1218 = (forvar1218 + (1'h1)))
                    begin
                      reg1219 <= (8'hb4);
                      reg1220 <= ($unsigned(forvar1188) ?
                          reg1219[(3'h5):(1'h0)] : (({reg1182} ~^ $unsigned(wire590)) ?
                              $unsigned(reg1177[(3'h4):(2'h3)]) : $signed((reg1151 ?
                                  (8'ha2) : (8'ha2)))));
                    end
                end
              reg1222 <= forvar1177;
            end
        end
      else
        begin
          if ((^~($unsigned((forvar1169 ? (8'ha0) : reg1171)) && ((-reg1203) ?
              (~(8'hae)) : (-(8'had))))))
            begin
              if (($signed(((reg1214 == reg1187) ?
                      reg1198[(4'he):(3'h5)] : reg1218)) ?
                  $unsigned(($unsigned(forvar1165) & $signed(reg1212))) : $signed({(8'hb2)})))
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (2'h3)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= (^~$signed({forvar1151}));
                    end
                  if ({$signed($unsigned((reg1183 ^~ reg1203)))})
                    begin
                      reg1198 <= $unsigned(reg1180[(3'h4):(2'h2)]);
                      reg1199 <= reg1198[(4'hc):(4'hc)];
                      reg1200 <= $unsigned((reg1181[(3'h6):(1'h0)] ?
                          (^reg1155) : forvar1165));
                      reg1201 <= $signed(($unsigned((forvar1197 ?
                              forvar1213 : reg1160)) ?
                          $unsigned(reg1214[(3'h6):(2'h3)]) : (reg1169 ?
                              forvar1168 : $unsigned(forvar1159))));
                    end
                  else
                    begin
                      reg1198 <= reg1150;
                    end
                  for (forvar1202 = (1'h0); (forvar1202 < (1'h0)); forvar1202 = (forvar1202 + (1'h1)))
                    begin
                      reg1203 <= ((8'haa) || forvar1157[(2'h3):(1'h0)]);
                      reg1204 <= wire588;
                    end
                  if ((~^($signed((~reg1168)) ?
                      (reg1148[(1'h0):(1'h0)] ?
                          ((8'ha0) ?
                              reg1200 : reg1185) : $signed(reg1222)) : $signed((forvar1205 ?
                          reg1163 : forvar1180)))))
                    begin
                      reg1205 <= {(($signed(wire589) ?
                              forvar1161[(3'h4):(1'h0)] : forvar1178[(1'h1):(1'h1)]) < reg1153[(3'h6):(2'h3)])};
                      reg1206 <= (^~(~|reg1204));
                      reg1207 <= (^~reg1197);
                    end
                  else
                    begin
                      reg1205 <= (~|{({wire585} * {(8'hab)})});
                      reg1206 <= reg1215[(3'h6):(1'h0)];
                      reg1207 <= {$unsigned($unsigned({reg1181}))};
                      reg1208 <= reg1162[(3'h4):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (2'h2)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= $signed($unsigned(forvar1161));
                    end
                  reg1198 <= $unsigned($signed(($unsigned(reg1173) == $signed((8'hb2)))));
                end
              if ($unsigned(reg1214[(2'h3):(1'h1)]))
                begin
                  for (forvar1209 = (1'h0); (forvar1209 < (2'h2)); forvar1209 = (forvar1209 + (1'h1)))
                    begin
                      reg1210 <= (~reg1212);
                    end
                end
              else
                begin
                  for (forvar1209 = (1'h0); (forvar1209 < (1'h1)); forvar1209 = (forvar1209 + (1'h1)))
                    begin
                      reg1210 <= (($unsigned((|forvar1171)) ?
                          reg1190 : (~&reg1157)) * $unsigned(reg1185[(1'h0):(1'h0)]));
                      reg1211 <= (+reg1157);
                      reg1212 <= (-((forvar1161[(4'h9):(4'h9)] ?
                              (-reg1205) : {reg1161}) ?
                          (~^$unsigned(reg1216)) : (reg1195 || forvar1205[(3'h4):(2'h2)])));
                      reg1213 <= ($signed({reg1198}) >>> (-reg1205));
                    end
                  for (forvar1214 = (1'h0); (forvar1214 < (1'h0)); forvar1214 = (forvar1214 + (1'h1)))
                    begin
                      reg1215 <= ((~|$signed(forvar1158)) * {((^reg1191) ?
                              (-forvar1186) : (reg1220 ?
                                  forvar1183 : forvar1148))});
                      reg1216 <= $signed($signed(forvar1154));
                      reg1217 <= forvar1186;
                      reg1218 <= {(&reg1215)};
                    end
                  for (forvar1219 = (1'h0); (forvar1219 < (1'h0)); forvar1219 = (forvar1219 + (1'h1)))
                    begin
                      reg1220 <= (((8'ha8) ^~ {{forvar1179}}) ?
                          {$signed($unsigned(reg1189))} : reg1149[(1'h0):(1'h0)]);
                    end
                  for (forvar1221 = (1'h0); (forvar1221 < (1'h0)); forvar1221 = (forvar1221 + (1'h1)))
                    begin
                      reg1222 <= (($signed(reg1153[(1'h0):(1'h0)]) & reg1204) <<< $unsigned($unsigned((reg1193 && (8'ha1)))));
                    end
                end
            end
          else
            begin
              if (reg1178)
                begin
                  for (forvar1196 = (1'h0); (forvar1196 < (2'h3)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= (forvar1168 + $unsigned($unsigned(((8'ha5) ~^ (8'h9f)))));
                      reg1198 <= reg1216[(3'h5):(1'h1)];
                    end
                  reg1199 <= reg1208[(3'h7):(3'h4)];
                  reg1200 <= forvar1188[(2'h3):(1'h0)];
                  for (forvar1201 = (1'h0); (forvar1201 < (1'h0)); forvar1201 = (forvar1201 + (1'h1)))
                    begin
                      reg1202 <= reg1160;
                      reg1203 <= wire590[(3'h6):(2'h3)];
                    end
                end
              else
                begin
                  reg1196 <= $signed($signed(forvar1183));
                  for (forvar1197 = (1'h0); (forvar1197 < (1'h0)); forvar1197 = (forvar1197 + (1'h1)))
                    begin
                      reg1198 <= reg1174[(3'h6):(3'h4)];
                      reg1199 <= ((((&(8'ha3)) ^~ reg1175) << $unsigned((8'hb4))) ?
                          {($unsigned(reg1213) ?
                                  reg1172[(4'h8):(3'h4)] : (reg1162 < forvar1148))} : ((|(forvar1216 ?
                              reg1210 : forvar1167)) > ((wire590 << forvar1159) >>> forvar1165)));
                    end
                end
              reg1204 <= $unsigned({reg1154});
              if ((forvar1221 * ($unsigned((reg1208 ? forvar1216 : reg1180)) ?
                  $unsigned($signed(forvar1162)) : $unsigned(reg1207))))
                begin
                  if ($unsigned((reg1185 ?
                      reg1219 : ({reg1201} && reg1196[(1'h0):(1'h0)]))))
                    begin
                      reg1205 <= forvar1178;
                      reg1206 <= ((~&((^~forvar1218) != $signed(forvar1166))) <<< (reg1189[(4'h9):(3'h6)] >> reg1200));
                      reg1207 <= ($unsigned(reg1159) ?
                          (~|reg1209[(3'h4):(3'h4)]) : ((~^(reg1212 < forvar1192)) ?
                              reg1219[(4'hc):(1'h1)] : $unsigned($signed(reg1184))));
                    end
                  else
                    begin
                      reg1205 <= (reg1221 ?
                          forvar1219[(4'ha):(3'h7)] : reg1193[(3'h5):(3'h4)]);
                    end
                end
              else
                begin
                  for (forvar1205 = (1'h0); (forvar1205 < (2'h3)); forvar1205 = (forvar1205 + (1'h1)))
                    begin
                      reg1206 <= ($unsigned(reg1216) >>> (^$signed(forvar1192)));
                    end
                  for (forvar1207 = (1'h0); (forvar1207 < (1'h0)); forvar1207 = (forvar1207 + (1'h1)))
                    begin
                      reg1208 <= wire588;
                      reg1209 <= wire588[(2'h3):(2'h2)];
                    end
                  for (forvar1210 = (1'h0); (forvar1210 < (1'h0)); forvar1210 = (forvar1210 + (1'h1)))
                    begin
                      reg1211 <= (&((-forvar1188) ?
                          (reg1219[(4'h8):(2'h3)] ?
                              (forvar1183 + wire588) : (&reg1202)) : $unsigned((reg1207 >= reg1210))));
                    end
                  for (forvar1212 = (1'h0); (forvar1212 < (1'h1)); forvar1212 = (forvar1212 + (1'h1)))
                    begin
                      reg1213 <= $signed($signed($signed($unsigned(reg1158))));
                    end
                end
              reg1214 <= ((forvar1167 <= reg1217) * (^~(~^(reg1150 == forvar1196))));
            end
        end
      if ((&(^~forvar1178[(2'h2):(1'h1)])))
        begin
          if ($signed((reg1187 << reg1205)))
            begin
              for (forvar1223 = (1'h0); (forvar1223 < (2'h2)); forvar1223 = (forvar1223 + (1'h1)))
                begin
                  if ((8'hb0))
                    begin
                      reg1224 <= ((reg1172[(1'h1):(1'h0)] ?
                              $signed($signed(forvar1169)) : $unsigned(reg1215[(3'h5):(1'h1)])) ?
                          $signed(forvar1186) : ((forvar1162 ?
                                  reg1149 : (forvar1221 < reg1157)) ?
                              {(^reg1162)} : $signed($signed(wire586))));
                    end
                  else
                    begin
                      reg1224 <= $unsigned($signed((forvar1188[(3'h5):(3'h5)] ?
                          $unsigned(reg1189) : {forvar1168})));
                      reg1225 <= forvar1161;
                      reg1226 <= ((wire1145[(1'h0):(1'h0)] >>> (^(reg1171 ?
                              (8'haa) : (8'hae)))) ?
                          reg1157 : $unsigned(forvar1166));
                      reg1227 <= reg1194;
                    end
                  if (forvar1177)
                    begin
                      reg1228 <= ((reg1222 ?
                              forvar1150 : ((reg1214 ?
                                  forvar1162 : reg1166) >>> {forvar1221})) ?
                          ((&(8'had)) ?
                              $signed((reg1180 ?
                                  reg1211 : forvar1201)) : {(reg1208 ^ reg1211)}) : {{{(8'ha6)}}});
                      reg1229 <= $signed($signed($unsigned(reg1195)));
                      reg1230 <= {$unsigned($unsigned($signed((8'ha5))))};
                    end
                  else
                    begin
                      reg1228 <= {((reg1184[(2'h2):(1'h1)] ?
                              forvar1196 : $signed(forvar1152)) * (+(~forvar1205)))};
                      reg1229 <= $signed(((+(reg1205 ? (8'ha9) : reg1201)) ?
                          forvar1213[(4'ha):(2'h3)] : ((reg1167 >= forvar1202) >= forvar1158)));
                      reg1230 <= $signed($signed(reg1160));
                      reg1231 <= (&{((reg1206 <<< forvar1214) ?
                              (reg1208 < reg1157) : (|reg1160))});
                    end
                  for (forvar1232 = (1'h0); (forvar1232 < (1'h0)); forvar1232 = (forvar1232 + (1'h1)))
                    begin
                      reg1233 <= reg1164[(1'h1):(1'h1)];
                      reg1234 <= $unsigned(reg1210);
                    end
                  if ((((8'hb6) ?
                          ($unsigned(reg1184) ?
                              reg1180 : $signed(reg1204)) : $unsigned((reg1233 * reg1198))) ?
                      $unsigned($unsigned(reg1178[(4'hd):(3'h4)])) : ($signed(forvar1188[(3'h4):(1'h1)]) >>> (~(reg1217 ?
                          (8'hae) : forvar1209)))))
                    begin
                      reg1235 <= $unsigned($signed($unsigned((reg1217 && reg1196))));
                    end
                  else
                    begin
                      reg1235 <= $signed({reg1207});
                      reg1236 <= $unsigned(reg1196);
                      reg1237 <= $signed(($unsigned($signed(reg1211)) ?
                          ((reg1152 * forvar1152) ?
                              {reg1218} : reg1228[(2'h3):(2'h3)]) : (8'ha2)));
                    end
                end
              if (({((forvar1188 + (8'had)) << ((8'ha4) >> reg1197))} & wire1147))
                begin
                  for (forvar1238 = (1'h0); (forvar1238 < (1'h0)); forvar1238 = (forvar1238 + (1'h1)))
                    begin
                      reg1239 <= $signed((|({forvar1202} <<< forvar1167)));
                      reg1240 <= $unsigned((((reg1194 ? (8'hb0) : reg1152) ?
                              reg1171[(1'h0):(1'h0)] : (reg1163 ?
                                  reg1209 : (8'ha4))) ?
                          (reg1158[(3'h7):(1'h0)] ?
                              reg1167 : (+reg1199)) : (|$signed((8'haf)))));
                      reg1241 <= (^reg1193[(3'h6):(2'h2)]);
                      reg1242 <= reg1209;
                    end
                  for (forvar1243 = (1'h0); (forvar1243 < (2'h2)); forvar1243 = (forvar1243 + (1'h1)))
                    begin
                      reg1244 <= reg1183[(2'h2):(1'h1)];
                    end
                  if ((-(8'ha2)))
                    begin
                      reg1245 <= $signed($signed(forvar1218[(2'h3):(1'h0)]));
                      reg1246 <= forvar1186;
                      reg1247 <= $unsigned(forvar1205);
                    end
                  else
                    begin
                      reg1245 <= $unsigned((~reg1194[(2'h2):(2'h2)]));
                      reg1246 <= {forvar1207};
                      reg1247 <= (^(|$signed(reg1159[(3'h6):(1'h1)])));
                      reg1248 <= (reg1246 ?
                          $unsigned(($unsigned(reg1171) ?
                              reg1213 : (|(8'ha8)))) : reg1187[(1'h0):(1'h0)]);
                    end
                  if ($unsigned(($unsigned($signed(forvar1168)) & $signed((reg1199 ?
                      reg1203 : reg1182)))))
                    begin
                      reg1249 <= {(reg1227[(4'h9):(2'h2)] ?
                              $unsigned((forvar1205 >>> reg1241)) : $signed($unsigned((8'h9d))))};
                      reg1250 <= reg1200;
                      reg1251 <= ((wire586 ?
                          $unsigned((~&reg1212)) : reg1248[(2'h3):(2'h2)]) > (!reg1187));
                      reg1252 <= (forvar1183 <<< reg1216[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg1249 <= (reg1148 >> (|{reg1176[(2'h2):(1'h1)]}));
                      reg1250 <= $unsigned(({forvar1219} | ((reg1226 << forvar1186) ?
                          (&reg1241) : (reg1207 < reg1180))));
                    end
                end
              else
                begin
                  if (({(|(|(8'h9c)))} ?
                      ($unsigned((!(8'h9c))) ?
                          reg1149 : (((8'ha2) ? reg1174 : forvar1207) ?
                              $unsigned(forvar1161) : (forvar1192 != reg1231))) : $signed(forvar1154[(1'h0):(1'h0)])))
                    begin
                      reg1238 <= ($signed((|(~|reg1214))) <<< (($unsigned(reg1251) ?
                              reg1201 : forvar1166) ?
                          reg1155 : wire1145));
                      reg1239 <= (reg1156[(1'h0):(1'h0)] <<< reg1186);
                    end
                  else
                    begin
                      reg1238 <= reg1205;
                      reg1239 <= reg1210[(1'h0):(1'h0)];
                      reg1240 <= $signed($signed($unsigned($signed(reg1208))));
                      reg1241 <= (($unsigned($unsigned(reg1154)) * $unsigned(reg1189)) ~^ (|$signed($signed(reg1225))));
                    end
                  if (((-forvar1196) ?
                      ($signed((^~(8'ha4))) && (forvar1202 ?
                          $unsigned(reg1186) : $signed(forvar1216))) : {$unsigned((reg1216 ?
                              (8'hb2) : reg1174))}))
                    begin
                      reg1242 <= (reg1208 ? {reg1152} : reg1190[(1'h1):(1'h0)]);
                      reg1243 <= reg1247[(3'h6):(3'h6)];
                      reg1244 <= (-{{{forvar1186}}});
                      reg1245 <= $signed({($unsigned((8'hab)) * forvar1202[(1'h1):(1'h0)])});
                    end
                  else
                    begin
                      reg1242 <= (^~reg1243);
                    end
                  for (forvar1246 = (1'h0); (forvar1246 < (1'h0)); forvar1246 = (forvar1246 + (1'h1)))
                    begin
                      reg1247 <= forvar1188[(3'h4):(3'h4)];
                      reg1248 <= reg1197[(4'hc):(2'h2)];
                      reg1249 <= forvar1186;
                      reg1250 <= $signed((8'h9c));
                    end
                  for (forvar1251 = (1'h0); (forvar1251 < (1'h0)); forvar1251 = (forvar1251 + (1'h1)))
                    begin
                      reg1252 <= $unsigned((-$signed((&reg1229))));
                      reg1253 <= ((^reg1184) ?
                          {$signed((&forvar1153))} : reg1247[(1'h1):(1'h1)]);
                      reg1254 <= (reg1163[(1'h1):(1'h1)] ?
                          $unsigned({$signed(reg1162)}) : $unsigned(forvar1162[(3'h5):(1'h0)]));
                      reg1255 <= $unsigned($signed($unsigned((reg1193 ?
                          forvar1168 : (8'ha7)))));
                    end
                end
              for (forvar1256 = (1'h0); (forvar1256 < (1'h0)); forvar1256 = (forvar1256 + (1'h1)))
                begin
                  if ((~({$signed((8'hab))} ?
                      {(reg1159 | (8'ha5))} : (^~(^~reg1175)))))
                    begin
                      reg1257 <= reg1246;
                      reg1258 <= (($unsigned((reg1208 ?
                              reg1186 : reg1207)) != $unsigned($unsigned((8'ha1)))) ?
                          $signed((~|(^~reg1187))) : (|wire590[(2'h2):(1'h1)]));
                      reg1259 <= ($signed(reg1176) != (~|((reg1193 && reg1253) ^~ (reg1243 >= reg1238))));
                    end
                  else
                    begin
                      reg1257 <= (reg1156[(1'h1):(1'h0)] ?
                          $unsigned(reg1151[(2'h2):(2'h2)]) : ((~|wire586[(4'hb):(3'h4)]) ?
                              ($signed((8'hb0)) ?
                                  reg1174 : (&(8'ha2))) : $unsigned(reg1154)));
                    end
                  if ((+(8'hb0)))
                    begin
                      reg1260 <= $unsigned($unsigned({$unsigned(reg1196)}));
                    end
                  else
                    begin
                      reg1260 <= ((^$signed((reg1156 ?
                          forvar1201 : reg1158))) != {forvar1156[(4'hb):(3'h6)]});
                      reg1261 <= $signed($signed($signed((reg1166 ?
                          forvar1232 : forvar1196))));
                    end
                  for (forvar1262 = (1'h0); (forvar1262 < (2'h3)); forvar1262 = (forvar1262 + (1'h1)))
                    begin
                      reg1263 <= reg1168;
                      reg1264 <= $unsigned((^~(~|(forvar1183 + reg1174))));
                    end
                end
              if ((8'ha8))
                begin
                  if ($signed((~$signed(forvar1165))))
                    begin
                      reg1265 <= (($signed((reg1180 <<< reg1181)) << $signed((&(8'ha5)))) ?
                          $signed($signed($signed(reg1198))) : $unsigned(forvar1148[(3'h7):(1'h1)]));
                      reg1266 <= ((($unsigned(forvar1159) > reg1151) * $signed((!reg1190))) <= reg1225[(2'h2):(2'h2)]);
                      reg1267 <= reg1151[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg1265 <= ($signed($signed(reg1216)) ?
                          ((reg1184[(1'h0):(1'h0)] >= reg1228[(3'h6):(1'h1)]) ?
                              reg1187[(1'h0):(1'h0)] : ((reg1246 ?
                                  reg1177 : forvar1243) && (^forvar1159))) : ((reg1240[(3'h7):(1'h0)] || $signed(reg1226)) || (8'ha9)));
                      reg1266 <= ($signed($unsigned({reg1166})) ?
                          reg1187 : {$signed((8'hb5))});
                      reg1267 <= reg1182[(4'hf):(2'h3)];
                      reg1268 <= reg1226;
                    end
                  if (reg1242[(3'h7):(3'h6)])
                    begin
                      reg1269 <= reg1196[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg1269 <= ({reg1177[(4'hd):(4'hb)]} > ({forvar1202[(3'h6):(3'h5)]} ?
                          forvar1216 : {$unsigned(forvar1177)}));
                      reg1270 <= reg1264[(2'h2):(1'h0)];
                      reg1271 <= (($signed($unsigned(reg1156)) ?
                              reg1196 : (!(8'hae))) ?
                          $signed(wire588[(4'hb):(3'h5)]) : $signed(reg1211[(2'h3):(2'h2)]));
                    end
                end
              else
                begin
                  for (forvar1265 = (1'h0); (forvar1265 < (2'h2)); forvar1265 = (forvar1265 + (1'h1)))
                    begin
                      reg1266 <= (&(reg1255 || {(wire588 ?
                              reg1251 : (8'hb6))}));
                      reg1267 <= forvar1180;
                      reg1268 <= $unsigned((reg1252[(2'h3):(2'h2)] == $signed(reg1171[(2'h2):(2'h2)])));
                    end
                end
            end
          else
            begin
              for (forvar1223 = (1'h0); (forvar1223 < (1'h0)); forvar1223 = (forvar1223 + (1'h1)))
                begin
                  reg1224 <= (8'hb2);
                  if ({(8'hb2)})
                    begin
                      reg1225 <= reg1190;
                      reg1226 <= reg1215;
                      reg1227 <= $unsigned((^~$unsigned($unsigned((8'hb0)))));
                    end
                  else
                    begin
                      reg1225 <= (~forvar1154[(2'h2):(2'h2)]);
                      reg1226 <= (({wire590} > forvar1246) || (((reg1251 ?
                                  reg1175 : reg1264) ?
                              (reg1237 <= (8'hb4)) : (reg1239 ?
                                  forvar1148 : forvar1192)) ?
                          ($unsigned(wire586) ?
                              (forvar1202 ?
                                  reg1201 : (8'h9f)) : $unsigned(reg1267)) : reg1175));
                      reg1227 <= (reg1189[(1'h0):(1'h0)] ^~ {$unsigned({reg1166})});
                      reg1228 <= reg1209;
                    end
                end
              for (forvar1229 = (1'h0); (forvar1229 < (1'h1)); forvar1229 = (forvar1229 + (1'h1)))
                begin
                  if ((^~$unsigned($unsigned(reg1202))))
                    begin
                      reg1230 <= $signed(reg1199[(4'hd):(3'h5)]);
                      reg1231 <= reg1250[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg1230 <= reg1183[(1'h1):(1'h1)];
                      reg1231 <= ((wire589[(1'h0):(1'h0)] ?
                          ($unsigned(reg1240) < (^forvar1158)) : $signed((forvar1178 >>> reg1170))) >> $unsigned(reg1237[(2'h2):(1'h1)]));
                      reg1232 <= {({$signed(reg1176)} ?
                              (~|reg1212[(4'ha):(3'h5)]) : ((~|reg1194) > {reg1157}))};
                    end
                end
            end
          for (forvar1272 = (1'h0); (forvar1272 < (2'h3)); forvar1272 = (forvar1272 + (1'h1)))
            begin
              for (forvar1273 = (1'h0); (forvar1273 < (2'h2)); forvar1273 = (forvar1273 + (1'h1)))
                begin
                  for (forvar1274 = (1'h0); (forvar1274 < (2'h2)); forvar1274 = (forvar1274 + (1'h1)))
                    begin
                      reg1275 <= {(^~((~|(8'ha7)) ? reg1234 : (^~reg1243)))};
                      reg1276 <= $signed((-$unsigned($signed(reg1245))));
                      reg1277 <= ((+$unsigned((~&reg1184))) <<< reg1178);
                    end
                  if ((^$signed($signed((forvar1210 - reg1218)))))
                    begin
                      reg1278 <= reg1239[(4'h8):(3'h7)];
                    end
                  else
                    begin
                      reg1278 <= {reg1221};
                      reg1279 <= $unsigned(forvar1178);
                      reg1280 <= (~^$unsigned($signed($signed((8'hb1)))));
                    end
                end
              for (forvar1281 = (1'h0); (forvar1281 < (1'h1)); forvar1281 = (forvar1281 + (1'h1)))
                begin
                  for (forvar1282 = (1'h0); (forvar1282 < (2'h2)); forvar1282 = (forvar1282 + (1'h1)))
                    begin
                      reg1283 <= reg1151[(3'h4):(1'h0)];
                      reg1284 <= (8'hb9);
                    end
                  for (forvar1285 = (1'h0); (forvar1285 < (1'h0)); forvar1285 = (forvar1285 + (1'h1)))
                    begin
                      reg1286 <= reg1251;
                      reg1287 <= (forvar1154[(1'h0):(1'h0)] || $unsigned(reg1283[(1'h1):(1'h0)]));
                    end
                  reg1288 <= (!reg1200);
                end
              if ((reg1250[(2'h2):(1'h1)] ?
                  (~^{{reg1179}}) : {reg1258[(4'h8):(3'h4)]}))
                begin
                  reg1289 <= (reg1230 ?
                      forvar1272 : $unsigned(({forvar1210} >= $signed((8'ha1)))));
                  reg1290 <= {reg1181};
                  for (forvar1291 = (1'h0); (forvar1291 < (1'h1)); forvar1291 = (forvar1291 + (1'h1)))
                    begin
                      reg1292 <= $signed(((~&forvar1214) != reg1225));
                      reg1293 <= (-forvar1246);
                      reg1294 <= (forvar1216 ^~ forvar1281);
                    end
                  for (forvar1295 = (1'h0); (forvar1295 < (1'h0)); forvar1295 = (forvar1295 + (1'h1)))
                    begin
                      reg1296 <= $unsigned(reg1183);
                      reg1297 <= $signed((reg1215[(2'h2):(2'h2)] ~^ reg1228));
                    end
                end
              else
                begin
                  reg1289 <= ((8'ha0) << {{(8'hb2)}});
                  for (forvar1290 = (1'h0); (forvar1290 < (2'h3)); forvar1290 = (forvar1290 + (1'h1)))
                    begin
                      reg1291 <= ((reg1162[(4'hc):(3'h5)] ?
                          ((forvar1163 + forvar1177) <= $unsigned(reg1156)) : reg1276) != reg1250[(3'h7):(3'h4)]);
                      reg1292 <= ($signed($unsigned((|reg1230))) ?
                          forvar1156 : $signed(reg1250[(1'h1):(1'h0)]));
                      reg1293 <= forvar1265[(3'h5):(1'h0)];
                    end
                end
              for (forvar1298 = (1'h0); (forvar1298 < (2'h2)); forvar1298 = (forvar1298 + (1'h1)))
                begin
                  for (forvar1299 = (1'h0); (forvar1299 < (1'h1)); forvar1299 = (forvar1299 + (1'h1)))
                    begin
                      reg1300 <= {(((reg1264 ?
                                  forvar1150 : (8'haf)) >>> ((8'hb7) - wire588)) ?
                              (!$unsigned(reg1244)) : reg1181)};
                      reg1301 <= (|(^~forvar1183[(1'h0):(1'h0)]));
                      reg1302 <= (~|forvar1221);
                      reg1303 <= (~|$signed(reg1284[(4'h8):(4'h8)]));
                    end
                end
            end
          if (($signed({(reg1280 ?
                  reg1194 : (8'hb4))}) >= (($unsigned(reg1156) ?
                  ((8'hb9) ^~ reg1261) : (forvar1162 ?
                      forvar1295 : forvar1272)) ?
              (reg1283[(3'h4):(2'h2)] ?
                  forvar1212[(3'h6):(2'h2)] : (~^(8'haa))) : (reg1173[(1'h0):(1'h0)] ?
                  {reg1201} : reg1181))))
            begin
              if (reg1207)
                begin
                  reg1304 <= (|$signed((~|(~reg1170))));
                  for (forvar1305 = (1'h0); (forvar1305 < (1'h0)); forvar1305 = (forvar1305 + (1'h1)))
                    begin
                      reg1306 <= {(&reg1211[(2'h2):(1'h0)])};
                      reg1307 <= reg1216;
                      reg1308 <= {reg1263[(3'h5):(2'h2)]};
                      reg1309 <= $unsigned($signed({(forvar1151 ?
                              reg1284 : forvar1232)}));
                    end
                  for (forvar1310 = (1'h0); (forvar1310 < (2'h2)); forvar1310 = (forvar1310 + (1'h1)))
                    begin
                      reg1311 <= (+reg1304[(3'h5):(1'h1)]);
                      reg1312 <= {(reg1296 ?
                              $unsigned((+reg1196)) : ($unsigned((8'h9e)) && (~^forvar1229)))};
                      reg1313 <= reg1228;
                    end
                end
              else
                begin
                  reg1304 <= (forvar1246 ?
                      $signed($unsigned((!wire590))) : ($unsigned(reg1176) + (reg1248 <= $signed(reg1289))));
                  reg1305 <= ((((reg1254 ?
                      reg1215 : reg1261) > forvar1161) | ($unsigned(reg1275) + (!reg1240))) ^ (((reg1175 ?
                          (8'ha6) : (8'hb8)) ~^ $signed((8'ha9))) ?
                      ((~&reg1247) << forvar1196) : (~$signed(reg1306))));
                  for (forvar1306 = (1'h0); (forvar1306 < (1'h0)); forvar1306 = (forvar1306 + (1'h1)))
                    begin
                      reg1307 <= $signed(reg1242[(2'h2):(1'h1)]);
                      reg1308 <= forvar1216[(3'h7):(3'h5)];
                      reg1309 <= reg1189;
                    end
                  if ($unsigned($unsigned($unsigned($unsigned((8'h9f))))))
                    begin
                      reg1310 <= $signed(((forvar1310 + $unsigned(reg1199)) ?
                          (forvar1282 >> reg1165[(4'ha):(1'h1)]) : reg1211[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg1310 <= reg1249[(2'h3):(1'h1)];
                      reg1311 <= reg1165[(4'hf):(2'h3)];
                    end
                end
              if (reg1202)
                begin
                  for (forvar1314 = (1'h0); (forvar1314 < (1'h1)); forvar1314 = (forvar1314 + (1'h1)))
                    begin
                      reg1315 <= (reg1194[(1'h1):(1'h0)] ?
                          forvar1213[(1'h1):(1'h1)] : reg1239);
                    end
                  reg1316 <= (((~&$signed(reg1309)) <= forvar1161) ?
                      (wire587 && reg1271[(3'h4):(1'h1)]) : ($signed(reg1193) < reg1248));
                end
              else
                begin
                  if (reg1237)
                    begin
                      reg1314 <= wire1145;
                      reg1315 <= (|wire586[(3'h4):(2'h3)]);
                      reg1316 <= $unsigned((($unsigned(reg1210) <<< forvar1148[(2'h2):(1'h1)]) ?
                          (((8'h9f) ? reg1148 : forvar1197) ?
                              (^~reg1224) : (forvar1213 <<< reg1209)) : $signed(reg1308)));
                    end
                  else
                    begin
                      reg1314 <= (forvar1156 >> reg1221[(2'h2):(1'h0)]);
                    end
                  if (reg1271[(2'h2):(1'h0)])
                    begin
                      reg1317 <= (~&reg1199);
                      reg1318 <= reg1180[(2'h2):(1'h0)];
                      reg1319 <= ($signed((~|((8'ha2) ?
                              (8'h9f) : forvar1251))) ?
                          forvar1153[(3'h7):(2'h2)] : $signed(((8'hb2) ?
                              $signed(wire1145) : $signed(reg1206))));
                    end
                  else
                    begin
                      reg1317 <= $signed({forvar1197[(3'h7):(3'h6)]});
                      reg1318 <= {(($signed(forvar1305) ?
                              $unsigned(reg1222) : ((8'h9f) ?
                                  reg1172 : reg1217)) <= $unsigned((8'hb5)))};
                      reg1319 <= (+{$signed(reg1230[(2'h2):(1'h0)])});
                    end
                  if ((-$unsigned(({reg1303} + $unsigned(reg1306)))))
                    begin
                      reg1320 <= $signed($unsigned(($signed(reg1254) - reg1279[(3'h4):(2'h3)])));
                      reg1321 <= (reg1187[(1'h0):(1'h0)] ?
                          $signed(((&reg1268) | reg1204[(1'h0):(1'h0)])) : {reg1208});
                    end
                  else
                    begin
                      reg1320 <= {wire588[(4'h8):(1'h0)]};
                      reg1321 <= (^~$signed($signed(reg1277)));
                    end
                  reg1322 <= $unsigned({forvar1148[(3'h4):(2'h3)]});
                end
              if ((~|$signed($signed(reg1316[(3'h4):(1'h0)]))))
                begin
                  for (forvar1323 = (1'h0); (forvar1323 < (1'h1)); forvar1323 = (forvar1323 + (1'h1)))
                    begin
                      reg1324 <= (|(|$signed(forvar1151)));
                      reg1325 <= $signed(reg1265[(3'h7):(3'h7)]);
                      reg1326 <= {forvar1188};
                    end
                end
              else
                begin
                  reg1323 <= $unsigned($signed((-$unsigned(reg1229))));
                  if ($signed(forvar1179[(4'ha):(3'h4)]))
                    begin
                      reg1324 <= $signed((reg1148 ?
                          (((8'haa) >= (8'ha5)) >= (reg1232 + forvar1153)) : $signed({(8'hb2)})));
                      reg1325 <= reg1195;
                      reg1326 <= {reg1289[(2'h2):(2'h2)]};
                      reg1327 <= ({reg1320[(4'h8):(1'h1)]} ?
                          $unsigned($signed({wire590})) : $signed(reg1155[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1324 <= (forvar1214 ?
                          $unsigned($signed((+reg1235))) : $signed({(reg1167 ?
                                  reg1229 : reg1261)}));
                      reg1325 <= (~&reg1199[(4'h8):(2'h2)]);
                      reg1326 <= forvar1151[(4'hb):(3'h6)];
                    end
                end
            end
          else
            begin
              if ($signed($unsigned(reg1284[(4'ha):(3'h4)])))
                begin
                  for (forvar1304 = (1'h0); (forvar1304 < (2'h3)); forvar1304 = (forvar1304 + (1'h1)))
                    begin
                      reg1305 <= (~|reg1196);
                      reg1306 <= $signed(reg1236[(2'h3):(1'h1)]);
                      reg1307 <= (forvar1251 ?
                          $unsigned(($signed(reg1221) ~^ reg1201[(2'h3):(1'h0)])) : $unsigned((!(-reg1222))));
                      reg1308 <= $unsigned((wire1145 && {(reg1194 <= reg1254)}));
                    end
                  for (forvar1309 = (1'h0); (forvar1309 < (1'h0)); forvar1309 = (forvar1309 + (1'h1)))
                    begin
                      reg1310 <= {{($unsigned(forvar1158) | $signed((8'hba)))}};
                      reg1311 <= reg1296[(2'h2):(2'h2)];
                    end
                  if (reg1221[(3'h7):(3'h4)])
                    begin
                      reg1312 <= ((&(8'hb3)) ~^ reg1196);
                      reg1313 <= ($signed($signed((forvar1207 ?
                          reg1214 : reg1162))) ~^ {$signed((forvar1186 ?
                              reg1275 : reg1208))});
                      reg1314 <= $signed($unsigned((^$unsigned((8'hba)))));
                      reg1315 <= (forvar1214[(1'h0):(1'h0)] ?
                          reg1254 : reg1154[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg1312 <= (reg1248[(1'h1):(1'h1)] ?
                          (^forvar1243) : (+(reg1237[(1'h0):(1'h0)] ?
                              reg1149[(1'h0):(1'h0)] : ((8'had) ^ (8'ha1)))));
                    end
                  if (forvar1205[(2'h2):(1'h1)])
                    begin
                      reg1316 <= $unsigned($unsigned($signed(forvar1168)));
                      reg1317 <= reg1288[(2'h3):(1'h1)];
                      reg1318 <= $signed((~$unsigned((|forvar1150))));
                    end
                  else
                    begin
                      reg1316 <= reg1206;
                      reg1317 <= (^(reg1290 ?
                          $signed($signed(forvar1153)) : (!(reg1317 ?
                              reg1209 : reg1220))));
                      reg1318 <= (|(8'h9e));
                    end
                end
              else
                begin
                  for (forvar1304 = (1'h0); (forvar1304 < (1'h0)); forvar1304 = (forvar1304 + (1'h1)))
                    begin
                      reg1305 <= ($unsigned((~&(forvar1153 ?
                              reg1165 : (8'hba)))) ?
                          reg1184[(1'h0):(1'h0)] : {$signed(reg1315[(3'h5):(3'h5)])});
                    end
                  for (forvar1306 = (1'h0); (forvar1306 < (1'h0)); forvar1306 = (forvar1306 + (1'h1)))
                    begin
                      reg1307 <= forvar1285;
                      reg1308 <= (($signed((forvar1179 + forvar1298)) ?
                          reg1149 : reg1155[(3'h7):(3'h7)]) && forvar1177[(4'hc):(4'h8)]);
                    end
                  reg1309 <= ({$unsigned((reg1174 ? reg1211 : forvar1209))} ?
                      (+$signed({reg1267})) : reg1243[(2'h3):(2'h2)]);
                  if ((+(~$signed(reg1254[(4'h9):(2'h2)]))))
                    begin
                      reg1310 <= $unsigned((reg1149 * $unsigned((reg1304 ?
                          forvar1192 : reg1278))));
                      reg1311 <= ($unsigned(((&(8'hb7)) >>> $unsigned(reg1280))) ?
                          ((+forvar1157[(2'h2):(2'h2)]) | reg1226) : $signed({$signed(forvar1157)}));
                      reg1312 <= (^$unsigned((~|{reg1296})));
                      reg1313 <= ($signed(forvar1323[(2'h3):(1'h1)]) && (reg1216[(2'h2):(1'h1)] ~^ ({reg1237} >= $signed(reg1300))));
                    end
                  else
                    begin
                      reg1310 <= $unsigned(reg1216);
                      reg1311 <= (8'haf);
                      reg1312 <= (~(reg1233 >>> $unsigned((+reg1226))));
                      reg1313 <= reg1242;
                    end
                end
              reg1319 <= (|(~|reg1316[(3'h4):(1'h0)]));
            end
          if ($signed({reg1148}))
            begin
              if ((~(($unsigned(reg1220) ?
                  forvar1310 : (reg1182 ?
                      (8'ha8) : forvar1148)) || {$signed((8'hb1))})))
                begin
                  reg1328 <= {(~^$unsigned({forvar1219}))};
                  reg1329 <= (forvar1151[(3'h5):(3'h5)] ?
                      $signed(((reg1149 <<< (8'hab)) * reg1237[(1'h0):(1'h0)])) : reg1300[(3'h5):(1'h0)]);
                end
              else
                begin
                  if (((((8'ha6) << $signed((8'h9c))) * {$signed(reg1240)}) < (8'hb3)))
                    begin
                      reg1328 <= $signed(reg1266[(1'h1):(1'h1)]);
                      reg1329 <= ((($signed(forvar1167) ?
                              forvar1158[(3'h4):(2'h2)] : (~|forvar1180)) > $signed(reg1176)) ?
                          ((forvar1178[(1'h1):(1'h0)] ?
                                  forvar1154 : $signed(reg1250)) ?
                              ((reg1186 << reg1265) ?
                                  (reg1181 ^ reg1232) : (reg1199 ?
                                      forvar1323 : forvar1310)) : (forvar1168 & (reg1201 ?
                                  reg1306 : reg1229))) : (!$unsigned((reg1315 > reg1150))));
                      reg1330 <= ((!$signed((reg1202 ? forvar1219 : reg1300))) ?
                          $signed($unsigned((forvar1201 ?
                              reg1149 : reg1164))) : {(reg1230[(1'h0):(1'h0)] ?
                                  forvar1216[(1'h0):(1'h0)] : reg1185[(2'h3):(1'h0)])});
                      reg1331 <= $signed((^~reg1149[(3'h5):(3'h5)]));
                    end
                  else
                    begin
                      reg1328 <= ($unsigned(reg1225) + (forvar1159[(4'h8):(2'h2)] ?
                          $unsigned(forvar1209[(1'h1):(1'h0)]) : (^(reg1268 ?
                              reg1315 : reg1284))));
                      reg1329 <= (forvar1149[(1'h1):(1'h0)] == (|reg1303));
                      reg1330 <= (((reg1239 > forvar1304) ?
                              $unsigned($signed(reg1261)) : (8'hac)) ?
                          (($unsigned(forvar1188) && (8'hb4)) ^ $signed((!reg1268))) : reg1160[(2'h2):(1'h1)]);
                    end
                  for (forvar1332 = (1'h0); (forvar1332 < (2'h2)); forvar1332 = (forvar1332 + (1'h1)))
                    begin
                      reg1333 <= ({reg1178} ?
                          (reg1199[(5'h10):(3'h6)] ?
                              $unsigned(reg1198[(1'h0):(1'h0)]) : $signed((reg1179 ?
                                  reg1241 : (8'haf)))) : (^wire1147[(4'hb):(4'h8)]));
                    end
                  for (forvar1334 = (1'h0); (forvar1334 < (2'h2)); forvar1334 = (forvar1334 + (1'h1)))
                    begin
                      reg1335 <= forvar1161[(3'h7):(2'h2)];
                      reg1336 <= ($signed(reg1217) ?
                          forvar1251[(2'h3):(2'h2)] : $unsigned((~|(reg1263 ?
                              reg1177 : (8'ha7)))));
                      reg1337 <= (!$signed(($signed(reg1291) ?
                          reg1237 : $unsigned(reg1243))));
                    end
                  if (reg1163)
                    begin
                      reg1338 <= (-reg1153);
                      reg1339 <= {wire587};
                    end
                  else
                    begin
                      reg1338 <= ((~|($signed((8'ha0)) | forvar1274)) <= (8'hb6));
                      reg1339 <= $signed(($unsigned($unsigned((8'hb7))) && reg1316[(1'h1):(1'h1)]));
                      reg1340 <= reg1214[(4'ha):(3'h4)];
                    end
                end
              if ((!(reg1237 ?
                  reg1244[(4'h8):(3'h6)] : forvar1282[(4'h9):(3'h6)])))
                begin
                  if ((forvar1168[(1'h1):(1'h1)] && reg1215[(2'h2):(2'h2)]))
                    begin
                      reg1341 <= forvar1221[(3'h5):(3'h5)];
                      reg1342 <= ($unsigned($unsigned($signed(reg1196))) << (&{(forvar1157 ?
                              forvar1216 : (8'ha6))}));
                      reg1343 <= ({(reg1287 ?
                                  (wire588 + reg1229) : $unsigned(wire587))} ?
                          reg1287 : $signed((8'had)));
                      reg1344 <= ({($signed(reg1315) ?
                              (~&reg1320) : reg1162)} | reg1293[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg1341 <= reg1166;
                      reg1342 <= reg1327;
                      reg1343 <= $unsigned($signed(reg1291));
                    end
                  reg1345 <= $unsigned(($unsigned((forvar1167 ^ (8'hae))) - reg1261[(4'h8):(2'h2)]));
                end
              else
                begin
                  for (forvar1341 = (1'h0); (forvar1341 < (2'h3)); forvar1341 = (forvar1341 + (1'h1)))
                    begin
                      reg1342 <= $signed((reg1196 | {reg1244}));
                      reg1343 <= $signed($signed((((8'ha1) || reg1210) ?
                          reg1210[(1'h1):(1'h0)] : reg1283[(3'h4):(2'h2)])));
                      reg1344 <= $signed(($unsigned((^~reg1237)) ^ reg1297));
                      reg1345 <= $unsigned(($unsigned($unsigned(reg1179)) >> reg1229[(1'h0):(1'h0)]));
                    end
                  if ($unsigned(reg1340[(2'h2):(1'h1)]))
                    begin
                      reg1346 <= forvar1299;
                      reg1347 <= {(-(forvar1310 ?
                              {reg1311} : ((8'had) ? forvar1156 : reg1226)))};
                    end
                  else
                    begin
                      reg1346 <= {wire590[(3'h6):(2'h3)]};
                      reg1347 <= ($signed(forvar1167[(2'h3):(2'h2)]) > ($signed((forvar1161 && reg1162)) ^~ reg1165[(2'h3):(1'h1)]));
                    end
                end
              if ((-$signed(((reg1333 ? reg1199 : reg1171) ?
                  (reg1289 ? reg1160 : (8'ha6)) : {forvar1177}))))
                begin
                  if ($signed((((reg1172 ? reg1171 : reg1161) ?
                          forvar1162[(3'h4):(1'h1)] : $unsigned(reg1200)) ?
                      (!(reg1340 ? (8'ha0) : reg1168)) : {{forvar1183}})))
                    begin
                      reg1348 <= ($signed($unsigned($signed(forvar1157))) || $signed(forvar1157[(3'h4):(3'h4)]));
                    end
                  else
                    begin
                      reg1348 <= (~$signed({(&reg1267)}));
                      reg1349 <= (((&(&reg1255)) + ($unsigned(reg1209) ?
                              $unsigned(wire587) : reg1238[(4'h8):(2'h3)])) ?
                          $unsigned(reg1271[(1'h0):(1'h0)]) : reg1239);
                    end
                  for (forvar1350 = (1'h0); (forvar1350 < (2'h3)); forvar1350 = (forvar1350 + (1'h1)))
                    begin
                      reg1351 <= (|($signed(reg1346) ?
                          (~^(forvar1216 ?
                              reg1243 : reg1269)) : $signed($unsigned(reg1175))));
                      reg1352 <= $signed(reg1345);
                      reg1353 <= reg1236[(3'h6):(3'h5)];
                    end
                  if (reg1293)
                    begin
                      reg1354 <= ((+(^(|reg1269))) >> $signed((~|(forvar1305 ?
                          reg1207 : reg1198))));
                      reg1355 <= ($signed(reg1338) ~^ $signed($unsigned((^~reg1261))));
                    end
                  else
                    begin
                      reg1354 <= wire589;
                      reg1355 <= ($unsigned(($unsigned(reg1351) ?
                          $signed(reg1240) : (^reg1244))) + reg1170);
                      reg1356 <= {$signed(reg1221)};
                      reg1357 <= $signed($signed($unsigned((reg1294 ?
                          reg1318 : reg1257))));
                    end
                  reg1358 <= forvar1149;
                end
              else
                begin
                  for (forvar1348 = (1'h0); (forvar1348 < (2'h2)); forvar1348 = (forvar1348 + (1'h1)))
                    begin
                      reg1349 <= ((^~forvar1350[(1'h0):(1'h0)]) || (&((^~reg1189) & $unsigned(forvar1207))));
                      reg1350 <= (&($unsigned(reg1172[(3'h7):(3'h4)]) ?
                          {$unsigned(reg1171)} : $signed(forvar1221)));
                    end
                  for (forvar1351 = (1'h0); (forvar1351 < (1'h1)); forvar1351 = (forvar1351 + (1'h1)))
                    begin
                      reg1352 <= reg1276[(2'h2):(1'h0)];
                      reg1353 <= $signed((&reg1310));
                    end
                  for (forvar1354 = (1'h0); (forvar1354 < (1'h0)); forvar1354 = (forvar1354 + (1'h1)))
                    begin
                      reg1355 <= reg1198;
                      reg1356 <= forvar1332[(2'h3):(1'h1)];
                      reg1357 <= ($signed($signed((reg1225 ?
                              forvar1161 : (8'haf)))) ?
                          {(reg1166[(1'h1):(1'h0)] ?
                                  (forvar1214 ?
                                      reg1358 : reg1169) : {(8'ha1)})} : $unsigned($signed((^~reg1314))));
                      reg1358 <= wire586;
                    end
                  if (reg1344)
                    begin
                      reg1359 <= $signed(reg1349);
                      reg1360 <= $signed((8'hb8));
                    end
                  else
                    begin
                      reg1359 <= ((&reg1277) ?
                          $unsigned($signed((reg1212 <= reg1294))) : $unsigned(((reg1196 ?
                                  (8'hb3) : reg1291) ?
                              reg1357[(4'h9):(4'h8)] : $unsigned((8'hb8)))));
                      reg1360 <= {(^~({reg1220} ?
                              (forvar1148 | forvar1310) : forvar1163))};
                      reg1361 <= ($unsigned(($unsigned(forvar1161) ?
                              reg1335[(3'h7):(2'h2)] : $unsigned(forvar1153))) ?
                          forvar1295 : (((reg1234 ? reg1313 : (8'haf)) ?
                              (reg1287 ^~ (8'ha7)) : (forvar1221 ?
                                  (8'ha3) : reg1347)) + (~{reg1185})));
                      reg1362 <= {$unsigned({$unsigned((8'ha8))})};
                    end
                end
              for (forvar1363 = (1'h0); (forvar1363 < (1'h1)); forvar1363 = (forvar1363 + (1'h1)))
                begin
                  reg1364 <= reg1198[(3'h5):(3'h4)];
                  for (forvar1365 = (1'h0); (forvar1365 < (2'h2)); forvar1365 = (forvar1365 + (1'h1)))
                    begin
                      reg1366 <= reg1220;
                      reg1367 <= (($unsigned((&forvar1178)) * $unsigned({reg1197})) ?
                          $signed((((8'h9e) * reg1224) && $signed((8'haa)))) : (^wire585));
                    end
                end
            end
          else
            begin
              for (forvar1328 = (1'h0); (forvar1328 < (1'h0)); forvar1328 = (forvar1328 + (1'h1)))
                begin
                  reg1329 <= reg1336[(1'h1):(1'h1)];
                end
              for (forvar1330 = (1'h0); (forvar1330 < (2'h2)); forvar1330 = (forvar1330 + (1'h1)))
                begin
                  if (((reg1306 ?
                          ((!reg1315) ?
                              ((8'hb2) | (8'h9d)) : $unsigned(reg1242)) : $signed(reg1303[(1'h1):(1'h1)])) ?
                      $signed($signed((!reg1172))) : $unsigned(((reg1361 << reg1170) ?
                          forvar1149[(2'h2):(1'h1)] : ((8'ha5) == (8'ha4))))))
                    begin
                      reg1331 <= reg1300[(1'h0):(1'h0)];
                      reg1332 <= reg1353[(1'h0):(1'h0)];
                      reg1333 <= $unsigned($signed((reg1228[(1'h0):(1'h0)] ?
                          reg1176[(2'h3):(1'h0)] : (reg1264 && (8'hb4)))));
                    end
                  else
                    begin
                      reg1331 <= $unsigned($unsigned((8'h9c)));
                    end
                  if (($unsigned(((^~(8'ha6)) & (reg1313 ?
                      (8'h9d) : reg1271))) * forvar1213))
                    begin
                      reg1334 <= ({forvar1232} - $signed(reg1230));
                    end
                  else
                    begin
                      reg1334 <= (forvar1238 ?
                          reg1336[(2'h2):(2'h2)] : (^~({forvar1265} <<< ((8'ha6) ?
                              forvar1162 : forvar1171))));
                      reg1335 <= {(reg1317 ?
                              (~^((8'h9c) && forvar1183)) : (8'hba))};
                      reg1336 <= reg1164;
                    end
                  for (forvar1337 = (1'h0); (forvar1337 < (1'h0)); forvar1337 = (forvar1337 + (1'h1)))
                    begin
                      reg1338 <= $unsigned(reg1339[(4'he):(3'h5)]);
                    end
                end
            end
        end
      else
        begin
          if (($unsigned($signed($unsigned(forvar1291))) ?
              ((&(8'h9e)) <<< forvar1167[(1'h1):(1'h1)]) : $unsigned(((reg1268 ?
                      reg1277 : reg1352) ?
                  {reg1321} : (+reg1260)))))
            begin
              for (forvar1223 = (1'h0); (forvar1223 < (2'h2)); forvar1223 = (forvar1223 + (1'h1)))
                begin
                  for (forvar1224 = (1'h0); (forvar1224 < (2'h3)); forvar1224 = (forvar1224 + (1'h1)))
                    begin
                      reg1225 <= $unsigned((~&($unsigned(reg1224) ?
                          {(8'hb4)} : {forvar1213})));
                      reg1226 <= reg1176;
                      reg1227 <= (~{reg1251[(3'h7):(2'h3)]});
                    end
                  for (forvar1228 = (1'h0); (forvar1228 < (1'h1)); forvar1228 = (forvar1228 + (1'h1)))
                    begin
                      reg1229 <= $unsigned($unsigned(forvar1205));
                    end
                  reg1230 <= $signed($signed(reg1345[(1'h0):(1'h0)]));
                  for (forvar1231 = (1'h0); (forvar1231 < (2'h3)); forvar1231 = (forvar1231 + (1'h1)))
                    begin
                      reg1232 <= ($signed($unsigned($unsigned(reg1167))) ?
                          (forvar1365[(1'h0):(1'h0)] ^ $signed($unsigned(forvar1341))) : ($signed($signed(forvar1196)) == forvar1224));
                    end
                end
              for (forvar1233 = (1'h0); (forvar1233 < (2'h3)); forvar1233 = (forvar1233 + (1'h1)))
                begin
                  if ($signed(reg1327[(3'h7):(1'h0)]))
                    begin
                      reg1234 <= $unsigned($unsigned($unsigned(reg1337)));
                      reg1235 <= reg1158;
                    end
                  else
                    begin
                      reg1234 <= ({(-((8'h9f) ?
                              forvar1152 : forvar1365))} ~^ (|(reg1338 || (~wire587))));
                      reg1235 <= ($unsigned({$signed(reg1241)}) >> ($unsigned(reg1297) < reg1364));
                    end
                  reg1236 <= forvar1299;
                end
            end
          else
            begin
              if ((!(((reg1252 ? reg1279 : (8'ha2)) << reg1283) - reg1217)))
                begin
                  reg1223 <= (~&reg1184);
                  for (forvar1224 = (1'h0); (forvar1224 < (1'h1)); forvar1224 = (forvar1224 + (1'h1)))
                    begin
                      reg1225 <= $unsigned(reg1230);
                      reg1226 <= reg1348;
                      reg1227 <= $unsigned((forvar1256 ?
                          ((~reg1326) + $unsigned(wire588)) : (^~(reg1202 | forvar1179))));
                      reg1228 <= ($unsigned({reg1297}) >> forvar1151);
                    end
                  reg1229 <= $unsigned((~^(!{forvar1246})));
                end
              else
                begin
                  if (reg1199[(2'h3):(1'h1)])
                    begin
                      reg1223 <= ($unsigned((~|reg1367)) ?
                          (reg1259 + reg1357[(4'h9):(1'h0)]) : (reg1238 < reg1258));
                      reg1224 <= ({(~&(reg1178 ? forvar1162 : (8'ha1)))} ?
                          reg1193[(4'hd):(1'h1)] : reg1347);
                      reg1225 <= (reg1223 ~^ reg1180);
                    end
                  else
                    begin
                      reg1223 <= forvar1232[(2'h2):(1'h1)];
                      reg1224 <= (~^$unsigned((forvar1178 >> $signed(reg1175))));
                      reg1225 <= forvar1304;
                    end
                  for (forvar1226 = (1'h0); (forvar1226 < (2'h3)); forvar1226 = (forvar1226 + (1'h1)))
                    begin
                      reg1227 <= reg1283[(2'h2):(2'h2)];
                      reg1228 <= (-$unsigned($unsigned($signed(forvar1179))));
                    end
                  for (forvar1229 = (1'h0); (forvar1229 < (2'h3)); forvar1229 = (forvar1229 + (1'h1)))
                    begin
                      reg1230 <= reg1152[(1'h1):(1'h0)];
                      reg1231 <= $unsigned((|(!forvar1224)));
                      reg1232 <= reg1156[(1'h1):(1'h0)];
                    end
                  for (forvar1233 = (1'h0); (forvar1233 < (1'h1)); forvar1233 = (forvar1233 + (1'h1)))
                    begin
                      reg1234 <= ((forvar1169 * {$unsigned((8'ha4))}) == (^~(~|reg1164[(1'h0):(1'h0)])));
                    end
                end
              if (($signed(($unsigned(reg1359) + (reg1210 << (8'hba)))) | reg1238))
                begin
                  if ((-(($unsigned(reg1352) ?
                          reg1257[(4'ha):(4'h8)] : (reg1149 ?
                              reg1194 : reg1196)) ?
                      (reg1306 ? forvar1218 : (8'had)) : ((reg1321 ?
                          reg1252 : reg1167) * reg1238))))
                    begin
                      reg1235 <= (~|$unsigned($signed({forvar1304})));
                      reg1236 <= (+reg1248[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg1235 <= (-forvar1282);
                      reg1236 <= {(reg1221[(1'h0):(1'h0)] ?
                              {(forvar1202 >>> reg1200)} : reg1224[(2'h3):(2'h3)])};
                      reg1237 <= ({reg1349} ?
                          $unsigned(reg1307[(3'h6):(2'h2)]) : $signed(((8'haa) << (|(8'hb3)))));
                      reg1238 <= reg1290;
                    end
                  for (forvar1239 = (1'h0); (forvar1239 < (2'h3)); forvar1239 = (forvar1239 + (1'h1)))
                    begin
                      reg1240 <= (&($signed((+forvar1354)) ?
                          reg1330 : reg1159[(2'h2):(1'h1)]));
                    end
                  for (forvar1241 = (1'h0); (forvar1241 < (1'h0)); forvar1241 = (forvar1241 + (1'h1)))
                    begin
                      reg1242 <= {(((reg1218 ? reg1250 : reg1317) ?
                              $signed(forvar1150) : (^forvar1196)) <<< $signed($signed(reg1300)))};
                    end
                  for (forvar1243 = (1'h0); (forvar1243 < (2'h2)); forvar1243 = (forvar1243 + (1'h1)))
                    begin
                      reg1244 <= $signed((forvar1216[(1'h1):(1'h0)] ~^ (8'h9e)));
                      reg1245 <= $signed((((~&reg1259) ?
                          reg1166[(3'h6):(1'h1)] : (~&forvar1334)) >> forvar1332));
                    end
                end
              else
                begin
                  if (($signed(reg1338[(1'h0):(1'h0)]) ?
                      $unsigned($signed(reg1268)) : forvar1365[(3'h7):(3'h6)]))
                    begin
                      reg1235 <= (&reg1223);
                      reg1236 <= (!reg1296[(2'h2):(1'h0)]);
                      reg1237 <= {forvar1207};
                      reg1238 <= forvar1239[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg1235 <= (reg1238[(3'h4):(2'h3)] ?
                          reg1187 : ((((8'hba) ? (8'h9f) : reg1265) ?
                                  (reg1223 < reg1358) : (!reg1352)) ?
                              ($unsigned(reg1211) <= forvar1273[(3'h5):(3'h4)]) : $signed((reg1187 ?
                                  reg1243 : forvar1166))));
                      reg1236 <= (reg1338 < $signed($unsigned($signed(reg1330))));
                      reg1237 <= reg1320;
                      reg1238 <= (((8'hb4) ^~ reg1251[(1'h0):(1'h0)]) ?
                          (((reg1180 ?
                              reg1241 : (8'hba)) != {forvar1291}) + forvar1158) : (~&(^~(reg1159 ?
                              reg1220 : forvar1243))));
                    end
                  if ((forvar1210[(3'h4):(2'h2)] ?
                      forvar1162[(3'h6):(3'h5)] : (~&(~^forvar1221[(3'h4):(3'h4)]))))
                    begin
                      reg1239 <= $signed(reg1330);
                      reg1240 <= $unsigned(reg1237);
                      reg1241 <= {reg1347};
                      reg1242 <= reg1321;
                    end
                  else
                    begin
                      reg1239 <= reg1268;
                      reg1240 <= (reg1236 ~^ $unsigned({$unsigned((8'hab))}));
                    end
                  if (reg1218)
                    begin
                      reg1243 <= ($signed((reg1241[(1'h1):(1'h1)] ?
                              (forvar1298 ?
                                  reg1242 : forvar1282) : (forvar1197 ?
                                  forvar1210 : forvar1163))) ?
                          forvar1341[(3'h4):(2'h2)] : $unsigned(($unsigned(forvar1179) ?
                              $signed(reg1260) : reg1167[(4'hb):(2'h2)])));
                      reg1244 <= ($unsigned(reg1246[(4'ha):(3'h5)]) ?
                          $unsigned({$signed(reg1245)}) : (^$unsigned({reg1190})));
                      reg1245 <= wire1147[(1'h1):(1'h0)];
                      reg1246 <= ($unsigned($unsigned((forvar1151 ?
                          reg1259 : reg1269))) & $unsigned((reg1337 & (forvar1202 <= reg1366))));
                    end
                  else
                    begin
                      reg1243 <= (~&forvar1165);
                      reg1244 <= ($unsigned(((-(8'h9c)) ?
                          (!reg1241) : $unsigned(forvar1209))) ^~ $unsigned((8'hac)));
                      reg1245 <= $unsigned(forvar1330);
                    end
                end
            end
          if ((+(+$unsigned($signed(reg1253)))))
            begin
              for (forvar1247 = (1'h0); (forvar1247 < (2'h2)); forvar1247 = (forvar1247 + (1'h1)))
                begin
                  for (forvar1248 = (1'h0); (forvar1248 < (1'h1)); forvar1248 = (forvar1248 + (1'h1)))
                    begin
                      reg1249 <= reg1195[(4'h8):(2'h2)];
                    end
                  for (forvar1250 = (1'h0); (forvar1250 < (2'h3)); forvar1250 = (forvar1250 + (1'h1)))
                    begin
                      reg1251 <= (reg1180[(1'h0):(1'h0)] ?
                          $signed($signed($unsigned(forvar1207))) : (reg1267[(1'h0):(1'h0)] ?
                              ($unsigned(reg1342) * (forvar1310 ?
                                  reg1338 : reg1348)) : forvar1232[(3'h4):(1'h0)]));
                    end
                  for (forvar1252 = (1'h0); (forvar1252 < (2'h2)); forvar1252 = (forvar1252 + (1'h1)))
                    begin
                      reg1253 <= $signed((~^reg1349[(1'h0):(1'h0)]));
                      reg1254 <= $unsigned(reg1211);
                      reg1255 <= reg1149[(2'h3):(1'h1)];
                    end
                  if (((&reg1216) ?
                      wire585 : (({forvar1252} ?
                              wire1147 : reg1276[(1'h1):(1'h1)]) ?
                          $unsigned((forvar1186 ?
                              reg1325 : (8'hb1))) : {$signed(reg1198)})))
                    begin
                      reg1256 <= ((((+reg1184) ?
                          forvar1196 : $unsigned(forvar1167)) | forvar1246[(3'h4):(1'h0)]) * reg1321[(1'h0):(1'h0)]);
                      reg1257 <= reg1291[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1256 <= (reg1150 ?
                          $unsigned(reg1318) : $signed($signed($unsigned(reg1357))));
                      reg1257 <= $unsigned(({$unsigned(reg1291)} ?
                          forvar1314 : $unsigned(((8'hac) > reg1241))));
                    end
                end
            end
          else
            begin
              if (((($unsigned((8'h9e)) ? (~^reg1187) : $unsigned(reg1256)) ?
                      forvar1304 : $signed({reg1352})) ?
                  $unsigned($signed({reg1266})) : ($unsigned({reg1230}) >> {$signed(reg1206)})))
                begin
                  for (forvar1247 = (1'h0); (forvar1247 < (2'h3)); forvar1247 = (forvar1247 + (1'h1)))
                    begin
                      reg1248 <= {$signed((^~(-reg1179)))};
                      reg1249 <= ($signed(((~reg1311) | forvar1167)) ?
                          ({$signed(forvar1306)} > {(~reg1309)}) : ((forvar1310 & $unsigned((8'hb5))) ?
                              ((reg1249 ? wire1145 : forvar1365) ?
                                  reg1256[(4'h9):(4'h8)] : (|reg1240)) : ((reg1314 < reg1168) && $signed((8'h9e)))));
                    end
                  reg1250 <= $unsigned((~|$unsigned($signed(reg1163))));
                  if (($signed(reg1191) ?
                      $signed(reg1328[(3'h4):(1'h0)]) : forvar1153))
                    begin
                      reg1251 <= ($signed(((+(8'hb3)) <= reg1320[(1'h0):(1'h0)])) == reg1178[(4'hf):(4'ha)]);
                      reg1252 <= reg1305;
                      reg1253 <= (reg1258[(1'h1):(1'h0)] ?
                          (((forvar1262 ?
                              reg1232 : reg1357) << forvar1192[(2'h2):(2'h2)]) >> (^~(reg1209 ^ (8'ha3)))) : (8'had));
                      reg1254 <= forvar1168[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1251 <= reg1160;
                      reg1252 <= (forvar1248 && forvar1218[(3'h6):(1'h0)]);
                      reg1253 <= ($signed({(reg1256 ? (8'h9d) : reg1280)}) ?
                          $unsigned(reg1166[(2'h2):(2'h2)]) : $unsigned(wire588));
                    end
                end
              else
                begin
                  if (reg1312)
                    begin
                      reg1247 <= reg1176;
                      reg1248 <= {(~^$unsigned($signed(reg1153)))};
                    end
                  else
                    begin
                      reg1247 <= (|$unsigned(reg1358));
                      reg1248 <= {$signed(forvar1351[(3'h4):(1'h0)])};
                    end
                end
            end
          if ({(^~forvar1158[(1'h1):(1'h0)])})
            begin
              for (forvar1258 = (1'h0); (forvar1258 < (1'h1)); forvar1258 = (forvar1258 + (1'h1)))
                begin
                  for (forvar1259 = (1'h0); (forvar1259 < (1'h1)); forvar1259 = (forvar1259 + (1'h1)))
                    begin
                      reg1260 <= forvar1166[(3'h6):(3'h6)];
                    end
                  for (forvar1261 = (1'h0); (forvar1261 < (2'h2)); forvar1261 = (forvar1261 + (1'h1)))
                    begin
                      reg1262 <= $unsigned(reg1280);
                      reg1263 <= forvar1169;
                      reg1264 <= $signed($signed(reg1187[(1'h0):(1'h0)]));
                      reg1265 <= {((forvar1332[(4'ha):(3'h4)] ^~ $signed(forvar1239)) ?
                              {{reg1314}} : (+$unsigned(reg1154)))};
                    end
                end
              reg1266 <= {$unsigned($signed((reg1343 ? reg1361 : forvar1196)))};
            end
          else
            begin
              reg1258 <= (($unsigned(forvar1306) ?
                      reg1359 : reg1262[(1'h0):(1'h0)]) ?
                  $unsigned((reg1176[(4'hb):(4'h8)] <= {wire585})) : forvar1192[(3'h5):(2'h3)]);
              for (forvar1259 = (1'h0); (forvar1259 < (2'h3)); forvar1259 = (forvar1259 + (1'h1)))
                begin
                  for (forvar1260 = (1'h0); (forvar1260 < (1'h0)); forvar1260 = (forvar1260 + (1'h1)))
                    begin
                      reg1261 <= ($unsigned((forvar1233[(4'h8):(4'h8)] ?
                              reg1315[(1'h1):(1'h0)] : $signed(reg1203))) ?
                          reg1325 : $unsigned(reg1321));
                    end
                  if (((!reg1350[(4'h8):(1'h1)]) ?
                      reg1169[(3'h5):(3'h5)] : $signed({$signed((8'ha0))})))
                    begin
                      reg1262 <= $unsigned(reg1218[(2'h3):(1'h1)]);
                      reg1263 <= (!forvar1233[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1262 <= (8'ha6);
                      reg1263 <= $signed(((forvar1158[(1'h0):(1'h0)] > reg1279[(1'h1):(1'h0)]) ?
                          (^{reg1316}) : $signed((forvar1167 ^ wire590))));
                    end
                  for (forvar1264 = (1'h0); (forvar1264 < (1'h0)); forvar1264 = (forvar1264 + (1'h1)))
                    begin
                      reg1265 <= {$signed(((forvar1241 >> reg1245) ?
                              $signed((8'ha0)) : (forvar1167 ?
                                  forvar1158 : reg1157)))};
                      reg1266 <= (!forvar1252);
                      reg1267 <= reg1242[(4'h8):(1'h0)];
                      reg1268 <= $unsigned($signed(((!reg1161) ?
                          wire586 : reg1222)));
                    end
                  for (forvar1269 = (1'h0); (forvar1269 < (2'h3)); forvar1269 = (forvar1269 + (1'h1)))
                    begin
                      reg1270 <= forvar1162;
                    end
                end
              for (forvar1271 = (1'h0); (forvar1271 < (2'h3)); forvar1271 = (forvar1271 + (1'h1)))
                begin
                  if (((reg1269[(2'h3):(2'h3)] * ($signed(reg1301) + $unsigned(reg1330))) & $signed(reg1187[(2'h2):(2'h2)])))
                    begin
                      reg1272 <= (((+reg1361[(2'h2):(1'h0)]) ?
                              (|reg1327[(3'h7):(3'h7)]) : (~&((8'ha3) ^~ reg1266))) ?
                          (~reg1201) : forvar1157);
                    end
                  else
                    begin
                      reg1272 <= reg1235;
                      reg1273 <= (~&((forvar1168[(4'h9):(1'h0)] ?
                          (|reg1310) : (8'had)) >= (~^$signed(forvar1201))));
                      reg1274 <= $signed(((!(forvar1262 ? reg1193 : (8'hb5))) ?
                          (+(reg1201 ? reg1353 : reg1207)) : ((~&reg1255) ?
                              forvar1161 : reg1231)));
                    end
                  if ($unsigned($signed($unsigned((reg1213 <= forvar1192)))))
                    begin
                      reg1275 <= ($signed((reg1325[(3'h7):(3'h5)] ?
                              (forvar1246 ? reg1359 : reg1203) : forvar1150)) ?
                          $signed(($signed(wire590) ?
                              {reg1159} : $signed(reg1352))) : (^$signed(reg1250)));
                      reg1276 <= (-{$unsigned((8'h9d))});
                      reg1277 <= (+((~&$unsigned(reg1272)) - $unsigned($signed(reg1180))));
                    end
                  else
                    begin
                      reg1275 <= $unsigned(((^(|forvar1154)) ?
                          forvar1269[(2'h3):(1'h1)] : reg1213[(3'h7):(3'h7)]));
                      reg1276 <= $signed($unsigned(((8'hb9) ?
                          reg1231[(2'h3):(2'h3)] : wire1145[(2'h2):(2'h2)])));
                      reg1277 <= $unsigned(($unsigned(reg1327) ?
                          $unsigned(reg1187[(1'h0):(1'h0)]) : $signed((~|(8'ha9)))));
                    end
                  if (((forvar1262[(3'h6):(3'h6)] | $unsigned((forvar1258 & reg1251))) ?
                      (($signed(reg1348) ? $unsigned(reg1338) : (-reg1348)) ?
                          $signed((reg1208 >> forvar1256)) : (-((8'ha7) ?
                              reg1187 : forvar1207))) : (+$unsigned((forvar1265 >>> (8'ha5))))))
                    begin
                      reg1278 <= $signed($unsigned($signed($signed(wire589))));
                      reg1279 <= (-(((reg1248 + reg1278) >>> (~|reg1236)) >= {$signed(reg1245)}));
                    end
                  else
                    begin
                      reg1278 <= $unsigned((reg1361[(1'h0):(1'h0)] ?
                          reg1309 : (-$signed(reg1152))));
                    end
                end
            end
        end
      for (forvar1368 = (1'h0); (forvar1368 < (2'h3)); forvar1368 = (forvar1368 + (1'h1)))
        begin
          if ((($signed((forvar1368 >> (8'hb1))) << $signed($signed((8'ha0)))) <= reg1331))
            begin
              if ((reg1216 >>> ($signed($signed(reg1241)) + (!(forvar1365 & reg1355)))))
                begin
                  reg1369 <= ((forvar1261 ?
                      (((8'hba) ? reg1177 : forvar1209) ?
                          forvar1282[(1'h0):(1'h0)] : (reg1366 <= forvar1238)) : {reg1208}) << ($signed((reg1334 ^ reg1226)) ?
                      ({reg1176} == reg1233[(2'h2):(2'h2)]) : forvar1323[(4'hd):(1'h1)]));
                  if ({forvar1233})
                    begin
                      reg1370 <= reg1227;
                      reg1371 <= $signed({{$unsigned(reg1211)}});
                    end
                  else
                    begin
                      reg1370 <= (forvar1295 || ($signed($signed(forvar1350)) ?
                          (reg1219 ^~ ((8'hb7) ?
                              (8'hb7) : (8'hb8))) : reg1366[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  if (reg1194)
                    begin
                      reg1369 <= {(8'hb0)};
                      reg1370 <= (|forvar1271);
                    end
                  else
                    begin
                      reg1369 <= ($unsigned((~&(forvar1282 < reg1304))) ?
                          (8'haa) : reg1370);
                      reg1370 <= reg1303[(1'h1):(1'h0)];
                      reg1371 <= ($unsigned((+reg1152[(3'h4):(1'h0)])) & reg1318);
                    end
                end
              if ($signed($signed((reg1209 | (|(8'h9c))))))
                begin
                  if ((reg1327[(3'h7):(3'h5)] ?
                      reg1241[(2'h2):(1'h1)] : $unsigned(($signed((8'haf)) ?
                          $unsigned(reg1328) : reg1272[(4'ha):(3'h4)]))))
                    begin
                      reg1372 <= (reg1311 ?
                          (($unsigned((8'hb2)) >>> $signed(forvar1246)) ?
                              $signed($signed(reg1159)) : (-reg1272[(2'h2):(1'h0)])) : $signed($signed((~&forvar1183))));
                      reg1373 <= reg1232[(3'h5):(1'h0)];
                    end
                  else
                    begin
                      reg1372 <= forvar1243;
                    end
                  if (forvar1233)
                    begin
                      reg1374 <= (((|reg1306) ^ ((forvar1152 * forvar1207) ?
                          (reg1213 >>> reg1259) : $unsigned(reg1243))) || ((+((8'hba) ?
                              reg1186 : reg1358)) ?
                          reg1279[(2'h3):(2'h2)] : reg1276));
                      reg1375 <= $unsigned($unsigned(reg1203));
                      reg1376 <= (((8'hb0) & reg1152) >>> (~|reg1185[(1'h0):(1'h0)]));
                      reg1377 <= $unsigned(reg1252);
                    end
                  else
                    begin
                      reg1374 <= (!forvar1207[(2'h2):(1'h1)]);
                      reg1375 <= (((^~wire585) ^~ ((forvar1310 << reg1239) >= (forvar1264 < forvar1207))) || (&(forvar1271 ^ ((8'hba) ?
                          forvar1183 : reg1331))));
                    end
                  for (forvar1378 = (1'h0); (forvar1378 < (1'h0)); forvar1378 = (forvar1378 + (1'h1)))
                    begin
                      reg1379 <= (reg1213[(4'hb):(3'h4)] >> reg1276[(1'h0):(1'h0)]);
                      reg1380 <= (^~reg1196[(1'h0):(1'h0)]);
                    end
                  if ({(&$unsigned($unsigned((8'hba))))})
                    begin
                      reg1381 <= ((~|{(|reg1287)}) >>> {$signed((wire587 ?
                              (8'ha2) : reg1325))});
                      reg1382 <= (~&(^({(8'ha4)} ?
                          (forvar1282 ?
                              reg1261 : reg1369) : reg1199[(2'h2):(2'h2)])));
                      reg1383 <= ((!(~&(~reg1369))) ?
                          reg1185 : ((forvar1210[(1'h0):(1'h0)] <<< ((8'ha7) ?
                              reg1182 : reg1190)) ~^ {(forvar1299 ?
                                  reg1267 : reg1168)}));
                    end
                  else
                    begin
                      reg1381 <= (forvar1328 ?
                          ((forvar1281 ?
                              {reg1232} : $unsigned(reg1174)) && $unsigned(reg1329[(4'h9):(4'h9)])) : {($unsigned((8'hb4)) >> (reg1238 ?
                                  forvar1219 : forvar1334))});
                      reg1382 <= $unsigned((~^$unsigned((forvar1330 ?
                          (8'ha2) : reg1316))));
                      reg1383 <= {$signed(($unsigned(reg1287) >> wire589[(3'h6):(2'h3)]))};
                    end
                end
              else
                begin
                  reg1372 <= ($signed(((!forvar1290) >= $unsigned(reg1342))) ?
                      $signed($signed((^forvar1304))) : $signed($unsigned({reg1375})));
                  for (forvar1373 = (1'h0); (forvar1373 < (2'h2)); forvar1373 = (forvar1373 + (1'h1)))
                    begin
                      reg1374 <= reg1268[(2'h3):(2'h3)];
                    end
                  reg1375 <= reg1248[(1'h1):(1'h0)];
                  if (reg1267)
                    begin
                      reg1376 <= forvar1258;
                      reg1377 <= reg1310[(3'h6):(1'h0)];
                      reg1378 <= (8'hb6);
                    end
                  else
                    begin
                      reg1376 <= ((reg1193 ?
                          $signed(forvar1169[(4'hb):(4'hb)]) : reg1162) ~^ forvar1223);
                      reg1377 <= $signed($signed((reg1214 ?
                          $unsigned(reg1200) : reg1243)));
                      reg1378 <= forvar1238[(2'h2):(2'h2)];
                      reg1379 <= forvar1341[(3'h5):(3'h4)];
                    end
                end
            end
          else
            begin
              reg1369 <= ($unsigned($signed(reg1172[(3'h7):(3'h4)])) ?
                  forvar1295 : (~^(^{forvar1271})));
              for (forvar1370 = (1'h0); (forvar1370 < (1'h0)); forvar1370 = (forvar1370 + (1'h1)))
                begin
                  for (forvar1371 = (1'h0); (forvar1371 < (2'h3)); forvar1371 = (forvar1371 + (1'h1)))
                    begin
                      reg1372 <= (((8'hb4) ? reg1237[(2'h2):(2'h2)] : reg1271) ?
                          {reg1203[(4'hd):(2'h3)]} : ((forvar1246[(3'h5):(1'h1)] && $unsigned(forvar1169)) >> (8'had)));
                      reg1373 <= (|$unsigned($unsigned($unsigned(reg1313))));
                    end
                  reg1374 <= forvar1157;
                end
            end
          if (forvar1219)
            begin
              if ((wire1147 <= reg1178))
                begin
                  for (forvar1384 = (1'h0); (forvar1384 < (2'h3)); forvar1384 = (forvar1384 + (1'h1)))
                    begin
                      reg1385 <= $signed((+((8'hb8) <= $unsigned(reg1154))));
                      reg1386 <= $unsigned(reg1346[(3'h5):(1'h1)]);
                    end
                  if (reg1343[(1'h0):(1'h0)])
                    begin
                      reg1387 <= $unsigned((((forvar1341 ?
                          forvar1158 : forvar1305) >> (forvar1273 < forvar1154)) * $unsigned((forvar1341 ?
                          reg1274 : forvar1247))));
                      reg1388 <= {$unsigned(wire586[(3'h7):(2'h2)])};
                    end
                  else
                    begin
                      reg1387 <= $unsigned((((reg1262 ^ reg1180) ?
                              reg1320[(2'h3):(2'h2)] : $signed(forvar1205)) ?
                          ((reg1222 ? reg1201 : reg1359) ?
                              ((8'ha6) != reg1257) : (-reg1235)) : $signed(reg1315)));
                      reg1388 <= (reg1214[(3'h4):(1'h0)] <= $unsigned($signed((forvar1299 <= forvar1274))));
                      reg1389 <= {$unsigned(reg1348)};
                      reg1390 <= (reg1157 ?
                          (&$unsigned($unsigned(forvar1378))) : $signed(({reg1211} != (wire586 ?
                              (8'ha1) : reg1156))));
                    end
                end
              else
                begin
                  reg1384 <= forvar1351;
                  if ($unsigned($signed(((reg1360 >> reg1385) ?
                      (~reg1381) : (~|reg1166)))))
                    begin
                      reg1385 <= ((8'hb2) ~^ (|reg1323));
                      reg1386 <= ({reg1344[(2'h3):(2'h3)]} ?
                          ($signed((reg1266 ^~ reg1306)) ^ reg1304[(4'ha):(3'h5)]) : $unsigned(($signed((8'hb6)) > $unsigned(reg1204))));
                    end
                  else
                    begin
                      reg1385 <= forvar1161[(4'hb):(3'h4)];
                      reg1386 <= $signed($signed(forvar1152[(2'h3):(2'h3)]));
                    end
                end
            end
          else
            begin
              reg1384 <= ((~reg1313[(3'h5):(1'h0)]) ?
                  {$signed(forvar1334[(1'h0):(1'h0)])} : (&forvar1252));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1391 = (1'h0); (forvar1391 < (2'h3)); forvar1391 = (forvar1391 + (1'h1)))
        begin
          reg1392 <= (forvar1274 ^~ $unsigned((~|$signed(reg1171))));
          for (forvar1393 = (1'h0); (forvar1393 < (2'h3)); forvar1393 = (forvar1393 + (1'h1)))
            begin
              if ({reg1288})
                begin
                  for (forvar1394 = (1'h0); (forvar1394 < (1'h1)); forvar1394 = (forvar1394 + (1'h1)))
                    begin
                      reg1395 <= $signed($unsigned((^~(|reg1243))));
                      reg1396 <= $signed((~{$unsigned(forvar1192)}));
                    end
                  if (reg1364)
                    begin
                      reg1397 <= (8'h9e);
                    end
                  else
                    begin
                      reg1397 <= forvar1212;
                      reg1398 <= $signed($signed((-$signed(reg1158))));
                    end
                end
              else
                begin
                  reg1394 <= (^reg1272[(3'h7):(1'h1)]);
                  for (forvar1395 = (1'h0); (forvar1395 < (2'h3)); forvar1395 = (forvar1395 + (1'h1)))
                    begin
                      reg1396 <= $signed((8'ha5));
                      reg1397 <= $unsigned((~|reg1313));
                      reg1398 <= reg1301;
                    end
                  if ($signed(($signed((reg1262 ? (8'hac) : reg1272)) ?
                      $signed($unsigned(reg1229)) : (~|$signed(reg1370)))))
                    begin
                      reg1399 <= $unsigned($signed(reg1258));
                      reg1400 <= (forvar1351[(1'h1):(1'h0)] ?
                          (!(|reg1370[(2'h2):(2'h2)])) : forvar1239[(1'h1):(1'h0)]);
                      reg1401 <= $unsigned(reg1348[(1'h1):(1'h1)]);
                      reg1402 <= $signed($signed((~|(8'hac))));
                    end
                  else
                    begin
                      reg1399 <= (reg1262[(1'h0):(1'h0)] ?
                          $signed((~|$unsigned(reg1367))) : $unsigned($signed(forvar1188)));
                    end
                  for (forvar1403 = (1'h0); (forvar1403 < (1'h1)); forvar1403 = (forvar1403 + (1'h1)))
                    begin
                      reg1404 <= (^~($unsigned($unsigned(reg1173)) || reg1366));
                      reg1405 <= reg1189;
                      reg1406 <= (~(((-reg1203) < reg1352[(4'hb):(3'h7)]) ?
                          $signed((~&reg1397)) : (&forvar1330)));
                      reg1407 <= ($unsigned($signed((reg1358 ?
                          forvar1166 : forvar1274))) >> {reg1222});
                    end
                end
              for (forvar1408 = (1'h0); (forvar1408 < (1'h0)); forvar1408 = (forvar1408 + (1'h1)))
                begin
                  for (forvar1409 = (1'h0); (forvar1409 < (1'h1)); forvar1409 = (forvar1409 + (1'h1)))
                    begin
                      reg1410 <= (~^reg1351);
                      reg1411 <= ((~(&$unsigned(reg1226))) ?
                          ($signed(reg1205) ?
                              $signed($signed(reg1152)) : ((forvar1192 != reg1377) << (~&reg1378))) : $signed(((^~reg1260) ?
                              $unsigned(forvar1409) : forvar1260)));
                      reg1412 <= (reg1152[(1'h0):(1'h0)] >> $unsigned((^~$unsigned(reg1200))));
                    end
                end
            end
          for (forvar1413 = (1'h0); (forvar1413 < (2'h2)); forvar1413 = (forvar1413 + (1'h1)))
            begin
              for (forvar1414 = (1'h0); (forvar1414 < (1'h0)); forvar1414 = (forvar1414 + (1'h1)))
                begin
                  reg1415 <= ({((~^reg1354) ?
                          {(8'ha8)} : (reg1193 ^~ forvar1299))} == (((reg1166 & reg1396) <= ((8'ha5) ?
                          (8'h9d) : reg1399)) ?
                      ($signed(reg1287) >>> forvar1188) : {$unsigned(reg1247)}));
                  if ((reg1271[(2'h2):(1'h1)] ?
                      (~^(8'hba)) : ((8'ha5) == ((~^reg1254) ^ reg1317))))
                    begin
                      reg1416 <= (~&(~^((^(8'h9f)) ?
                          (reg1297 ^ reg1404) : (^forvar1243))));
                      reg1417 <= (forvar1264 <<< ((|$signed(reg1338)) - $signed((forvar1171 << reg1265))));
                      reg1418 <= (($unsigned((forvar1371 && (8'hb0))) ?
                          $signed((8'hb2)) : ((~|reg1253) ?
                              (reg1174 ? reg1345 : reg1245) : (forvar1149 ?
                                  (8'ha3) : reg1297))) >> ($signed($unsigned(reg1190)) && ($signed(forvar1251) < (reg1220 || forvar1251))));
                    end
                  else
                    begin
                      reg1416 <= ($unsigned($signed(reg1320[(3'h7):(1'h0)])) <= (forvar1159[(2'h2):(1'h1)] != ($signed(forvar1165) ?
                          {forvar1183} : reg1287)));
                      reg1417 <= ((~&((-forvar1264) <= $signed(forvar1243))) == (~|((reg1395 <<< forvar1304) ?
                          (!forvar1232) : (8'hac))));
                    end
                end
              for (forvar1419 = (1'h0); (forvar1419 < (2'h2)); forvar1419 = (forvar1419 + (1'h1)))
                begin
                  if (((({(8'h9c)} | (reg1183 ? (8'ha7) : forvar1281)) ?
                          {reg1378[(1'h0):(1'h0)]} : forvar1370[(2'h2):(1'h1)]) ?
                      ($signed($signed(forvar1269)) ?
                          {$signed(reg1397)} : $unsigned($unsigned(reg1244))) : forvar1265))
                    begin
                      reg1420 <= $unsigned(forvar1252);
                      reg1421 <= $unsigned(($unsigned((reg1306 ?
                          (8'hb9) : forvar1178)) | (~^forvar1305)));
                      reg1422 <= (~&$signed(reg1340));
                      reg1423 <= ({$signed($signed((8'hb9)))} < forvar1393[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg1420 <= $unsigned({($signed(reg1248) ?
                              (~^reg1171) : (forvar1219 ^~ forvar1330))});
                    end
                  for (forvar1424 = (1'h0); (forvar1424 < (1'h0)); forvar1424 = (forvar1424 + (1'h1)))
                    begin
                      reg1425 <= $signed({(~^$unsigned(reg1154))});
                    end
                end
            end
          for (forvar1426 = (1'h0); (forvar1426 < (2'h2)); forvar1426 = (forvar1426 + (1'h1)))
            begin
              reg1427 <= reg1189;
              for (forvar1428 = (1'h0); (forvar1428 < (1'h0)); forvar1428 = (forvar1428 + (1'h1)))
                begin
                  reg1429 <= $signed(forvar1218[(3'h4):(2'h2)]);
                  for (forvar1430 = (1'h0); (forvar1430 < (2'h2)); forvar1430 = (forvar1430 + (1'h1)))
                    begin
                      reg1431 <= $unsigned((&reg1313[(3'h5):(2'h2)]));
                      reg1432 <= reg1400;
                    end
                  for (forvar1433 = (1'h0); (forvar1433 < (2'h3)); forvar1433 = (forvar1433 + (1'h1)))
                    begin
                      reg1434 <= $signed(reg1258[(4'h8):(2'h2)]);
                      reg1435 <= reg1215[(3'h4):(3'h4)];
                    end
                  if (reg1307[(4'hb):(1'h1)])
                    begin
                      reg1436 <= (!reg1420[(4'ha):(1'h1)]);
                    end
                  else
                    begin
                      reg1436 <= {((reg1287 ?
                              (reg1379 <= forvar1272) : (reg1269 - reg1350)) << reg1189[(3'h7):(3'h5)])};
                      reg1437 <= (&((forvar1323[(4'he):(1'h1)] ?
                              $unsigned((8'haf)) : $signed(reg1180)) ?
                          {reg1173} : (8'ha9)));
                    end
                end
              if ((8'h9d))
                begin
                  if ((8'hb0))
                    begin
                      reg1438 <= reg1250[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg1438 <= (($unsigned($signed(reg1350)) <= (reg1227 ^~ {reg1374})) ?
                          (forvar1179[(3'h4):(1'h0)] ?
                              {(~|reg1307)} : forvar1256) : $unsigned({(forvar1158 ~^ reg1239)}));
                      reg1439 <= ((({reg1344} >= {reg1169}) ?
                          $signed($unsigned(reg1216)) : (&$signed(forvar1201))) <= $unsigned($signed((reg1175 * reg1243))));
                      reg1440 <= reg1217[(3'h5):(3'h5)];
                    end
                end
              else
                begin
                  for (forvar1438 = (1'h0); (forvar1438 < (1'h1)); forvar1438 = (forvar1438 + (1'h1)))
                    begin
                      reg1439 <= $unsigned($signed(forvar1384[(3'h5):(2'h3)]));
                      reg1440 <= $signed((forvar1368[(4'ha):(4'h8)] ?
                          {(^~forvar1269)} : $signed(reg1392)));
                      reg1441 <= $signed($signed($unsigned((reg1287 ?
                          reg1162 : reg1326))));
                    end
                end
              reg1442 <= $signed($unsigned(($signed(reg1198) >= (+reg1156))));
            end
        end
      for (forvar1443 = (1'h0); (forvar1443 < (1'h1)); forvar1443 = (forvar1443 + (1'h1)))
        begin
          if ((({reg1371[(2'h2):(1'h0)]} ?
                  ($signed((8'ha4)) - (reg1231 ?
                      reg1210 : reg1429)) : (reg1398[(3'h4):(2'h2)] ?
                      ((8'hb5) ? reg1333 : reg1261) : $unsigned(reg1360))) ?
              (~reg1352[(4'hd):(3'h5)]) : $unsigned($unsigned((reg1330 != reg1249)))))
            begin
              reg1444 <= (8'h9e);
              reg1445 <= $signed(((|forvar1150[(1'h1):(1'h0)]) == (|$signed(reg1347))));
              for (forvar1446 = (1'h0); (forvar1446 < (1'h1)); forvar1446 = (forvar1446 + (1'h1)))
                begin
                  reg1447 <= (reg1370 && (^~forvar1169));
                  for (forvar1448 = (1'h0); (forvar1448 < (2'h3)); forvar1448 = (forvar1448 + (1'h1)))
                    begin
                      reg1449 <= $signed($signed($signed((&reg1372))));
                    end
                  reg1450 <= reg1268[(3'h6):(3'h6)];
                end
            end
          else
            begin
              if ((!(|(~forvar1224))))
                begin
                  if ($unsigned(($unsigned((&forvar1298)) + forvar1226[(1'h1):(1'h0)])))
                    begin
                      reg1444 <= (($unsigned(reg1340[(2'h2):(1'h0)]) ?
                          (((8'hb4) | reg1357) | $signed(forvar1246)) : (^~$signed(reg1418))) && (|reg1371[(2'h2):(2'h2)]));
                      reg1445 <= $unsigned((8'ha7));
                      reg1446 <= {$unsigned(({reg1239} ?
                              (reg1322 << reg1291) : (&reg1360)))};
                      reg1447 <= $unsigned($unsigned($signed({reg1399})));
                    end
                  else
                    begin
                      reg1444 <= $signed({((reg1154 ? reg1195 : (8'ha3)) ?
                              {forvar1247} : (reg1265 ?
                                  forvar1166 : reg1314))});
                      reg1445 <= (({reg1178[(2'h3):(2'h3)]} ?
                              $unsigned((reg1250 ?
                                  reg1259 : reg1181)) : (((8'haf) && reg1247) || reg1334)) ?
                          (reg1389[(3'h4):(1'h1)] ?
                              (8'hb2) : forvar1285) : forvar1232);
                    end
                  if (forvar1243)
                    begin
                      reg1448 <= forvar1153[(4'hf):(2'h3)];
                      reg1449 <= ($signed(reg1264) <= (reg1434 >> $unsigned((reg1216 ?
                          forvar1443 : reg1264))));
                      reg1450 <= $unsigned(((&$signed(reg1339)) ?
                          $unsigned($unsigned(forvar1179)) : (8'hb9)));
                      reg1451 <= forvar1248;
                    end
                  else
                    begin
                      reg1448 <= $signed({$unsigned(reg1356)});
                      reg1449 <= ((^$unsigned((reg1400 ?
                          reg1411 : reg1441))) >>> (~|((reg1334 ~^ reg1150) ?
                          $unsigned(reg1206) : (reg1362 ?
                              forvar1262 : reg1160))));
                      reg1450 <= (!reg1276);
                      reg1451 <= (8'ha1);
                    end
                end
              else
                begin
                  if ((~&forvar1438))
                    begin
                      reg1444 <= $signed({(^~((8'h9d) - reg1311))});
                    end
                  else
                    begin
                      reg1444 <= reg1176[(2'h3):(2'h3)];
                      reg1445 <= reg1210;
                      reg1446 <= (|reg1427[(3'h6):(3'h6)]);
                      reg1447 <= {$unsigned($signed((^reg1304)))};
                    end
                  for (forvar1448 = (1'h0); (forvar1448 < (1'h0)); forvar1448 = (forvar1448 + (1'h1)))
                    begin
                      reg1449 <= {reg1213};
                    end
                  for (forvar1450 = (1'h0); (forvar1450 < (2'h3)); forvar1450 = (forvar1450 + (1'h1)))
                    begin
                      reg1451 <= reg1287[(4'h9):(1'h1)];
                      reg1452 <= forvar1186[(2'h3):(1'h0)];
                      reg1453 <= ({{{reg1318}}} + (($unsigned(forvar1438) ^ $signed(reg1308)) >> ($unsigned(reg1186) == (reg1166 ?
                          reg1256 : reg1213))));
                    end
                  for (forvar1454 = (1'h0); (forvar1454 < (1'h0)); forvar1454 = (forvar1454 + (1'h1)))
                    begin
                      reg1455 <= reg1155[(4'hb):(3'h5)];
                    end
                end
              for (forvar1456 = (1'h0); (forvar1456 < (1'h1)); forvar1456 = (forvar1456 + (1'h1)))
                begin
                  if ({($unsigned(forvar1186[(2'h3):(2'h2)]) ?
                          {$signed(reg1181)} : reg1349[(3'h7):(3'h4)])})
                    begin
                      reg1457 <= $signed(reg1240);
                      reg1458 <= ({$unsigned($unsigned(forvar1363))} ?
                          ($signed($unsigned((8'ha4))) >= $signed((reg1211 & (8'h9c)))) : ($unsigned((forvar1250 << reg1218)) ?
                              (^(reg1314 == reg1291)) : $signed($signed(reg1427))));
                      reg1459 <= ({wire585} ^ ((+$unsigned(forvar1350)) ?
                          wire1145 : forvar1213));
                      reg1460 <= ($signed((((8'h9d) << forvar1262) ?
                          (reg1342 ^ reg1444) : (~^reg1228))) | (^reg1436));
                    end
                  else
                    begin
                      reg1457 <= $signed((reg1340 ?
                          $signed((&reg1236)) : (-$unsigned(forvar1273))));
                    end
                end
              reg1461 <= reg1331[(3'h5):(2'h3)];
              for (forvar1462 = (1'h0); (forvar1462 < (2'h3)); forvar1462 = (forvar1462 + (1'h1)))
                begin
                  for (forvar1463 = (1'h0); (forvar1463 < (1'h0)); forvar1463 = (forvar1463 + (1'h1)))
                    begin
                      reg1464 <= ((~|reg1459[(3'h6):(3'h6)]) ?
                          $signed($signed({reg1377})) : $unsigned(reg1439));
                      reg1465 <= $unsigned($signed((~(!(8'haa)))));
                      reg1466 <= ($unsigned($signed(reg1155)) ?
                          $signed(reg1199[(4'hb):(3'h5)]) : (8'haa));
                      reg1467 <= reg1350[(4'h9):(4'h9)];
                    end
                  reg1468 <= (~^$signed(((8'hb8) ?
                      (forvar1214 - (8'hb5)) : reg1167[(4'hc):(4'h8)])));
                end
            end
          if (((reg1170[(2'h2):(1'h1)] ?
                  forvar1212 : (forvar1256 - (reg1406 <<< (8'ha2)))) ?
              ($unsigned($signed(reg1273)) ?
                  $unsigned({reg1416}) : (((8'ha3) == (8'ha7)) - (^reg1272))) : (^~{forvar1161[(3'h5):(1'h0)]})))
            begin
              for (forvar1469 = (1'h0); (forvar1469 < (1'h0)); forvar1469 = (forvar1469 + (1'h1)))
                begin
                  if (reg1149[(2'h3):(2'h3)])
                    begin
                      reg1470 <= reg1181;
                      reg1471 <= (8'ha1);
                    end
                  else
                    begin
                      reg1470 <= ($unsigned({$unsigned((8'had))}) ?
                          $signed($signed((reg1233 == reg1167))) : reg1314);
                      reg1471 <= reg1154[(2'h3):(1'h0)];
                    end
                  for (forvar1472 = (1'h0); (forvar1472 < (2'h2)); forvar1472 = (forvar1472 + (1'h1)))
                    begin
                      reg1473 <= (8'hb7);
                      reg1474 <= ((forvar1168[(4'ha):(2'h3)] >> forvar1265[(4'hb):(3'h4)]) ?
                          forvar1282[(4'h8):(4'h8)] : (reg1417[(2'h3):(2'h2)] <= $unsigned($signed((8'h9d)))));
                      reg1475 <= ((reg1402 + $unsigned(forvar1273)) ?
                          {$unsigned((reg1241 ~^ forvar1209))} : (!forvar1256[(4'hd):(3'h4)]));
                    end
                  if ({reg1452})
                    begin
                      reg1476 <= (8'hb4);
                      reg1477 <= $unsigned($unsigned(reg1421));
                      reg1478 <= ($signed(((reg1400 ?
                          forvar1282 : reg1337) >= $signed(reg1344))) + reg1314);
                      reg1479 <= reg1239[(4'h9):(1'h1)];
                    end
                  else
                    begin
                      reg1476 <= $signed((8'haf));
                    end
                end
              for (forvar1480 = (1'h0); (forvar1480 < (1'h0)); forvar1480 = (forvar1480 + (1'h1)))
                begin
                  reg1481 <= (^~((reg1404[(1'h0):(1'h0)] ~^ ((8'ha5) ^~ reg1307)) ?
                      ((reg1149 <<< forvar1152) * $unsigned(reg1396)) : (|$signed(wire587))));
                  reg1482 <= ($unsigned((8'hb1)) == forvar1430[(4'he):(3'h7)]);
                end
            end
          else
            begin
              if ((reg1383 & (~(^$unsigned(forvar1409)))))
                begin
                  if (((+forvar1243) + $signed(forvar1443)))
                    begin
                      reg1469 <= (~^$signed(((!reg1418) ^~ (reg1327 ?
                          reg1459 : (8'hb1)))));
                      reg1470 <= (~|(~|(~|(forvar1443 ? reg1259 : reg1466))));
                      reg1471 <= reg1194;
                      reg1472 <= ($unsigned($unsigned((|(8'hb1)))) & reg1242);
                    end
                  else
                    begin
                      reg1469 <= $signed(forvar1179[(4'h8):(4'h8)]);
                      reg1470 <= reg1264;
                    end
                  if (((-reg1189) - (&((reg1174 ~^ (8'hae)) * $signed(reg1366)))))
                    begin
                      reg1473 <= (8'ha8);
                      reg1474 <= (8'ha7);
                    end
                  else
                    begin
                      reg1473 <= reg1209;
                      reg1474 <= $unsigned($signed(((-reg1151) ?
                          (reg1286 ? reg1263 : reg1353) : (reg1161 ?
                              (8'hb5) : wire1145))));
                      reg1475 <= $unsigned({(-(reg1274 || reg1157))});
                      reg1476 <= (8'h9e);
                    end
                  if (($unsigned((forvar1157 && (forvar1183 + reg1287))) ?
                      reg1189 : reg1182))
                    begin
                      reg1477 <= reg1332;
                      reg1478 <= {reg1218[(3'h5):(3'h4)]};
                    end
                  else
                    begin
                      reg1477 <= ($signed($signed($unsigned(forvar1177))) ?
                          (^~reg1293) : reg1383[(1'h1):(1'h0)]);
                      reg1478 <= {forvar1334[(1'h0):(1'h0)]};
                    end
                  for (forvar1479 = (1'h0); (forvar1479 < (1'h1)); forvar1479 = (forvar1479 + (1'h1)))
                    begin
                      reg1480 <= ({$unsigned((&reg1152))} ?
                          $unsigned((-$signed(reg1461))) : (((-reg1273) ?
                                  (forvar1409 ?
                                      forvar1391 : reg1392) : wire1145) ?
                              (8'hb3) : ((reg1400 >> forvar1247) ^ $signed((8'hb7)))));
                      reg1481 <= (^$signed((+reg1312)));
                      reg1482 <= (reg1218[(4'h8):(2'h3)] ?
                          wire586 : (reg1358[(3'h5):(3'h5)] ^ forvar1384));
                      reg1483 <= (^(!(~((8'h9f) >> (8'hb0)))));
                    end
                end
              else
                begin
                  reg1469 <= $unsigned(reg1326[(2'h2):(1'h1)]);
                  if (reg1177)
                    begin
                      reg1470 <= reg1472;
                      reg1471 <= forvar1298;
                    end
                  else
                    begin
                      reg1470 <= $signed((+(-(reg1411 * forvar1156))));
                    end
                  if ((reg1321 <<< ((~&$unsigned(wire588)) ?
                      reg1345 : reg1364)))
                    begin
                      reg1472 <= $signed((reg1468 + {((8'ha9) <= reg1290)}));
                      reg1473 <= {(((forvar1463 - reg1286) ?
                              (forvar1210 || reg1284) : (reg1199 ?
                                  forvar1186 : forvar1371)) <= ($unsigned(reg1251) ?
                              (reg1158 + forvar1354) : (reg1404 ?
                                  (8'hb4) : reg1300)))};
                      reg1474 <= ({$unsigned((&reg1387))} * forvar1424);
                      reg1475 <= (($unsigned($signed((8'had))) ?
                          (!{reg1234}) : (~|reg1304)) < (8'ha5));
                    end
                  else
                    begin
                      reg1472 <= ((($signed(reg1241) < $unsigned(reg1165)) << ((forvar1260 ?
                              reg1231 : reg1476) & (reg1458 <<< wire1145))) ?
                          $signed($unsigned(forvar1196)) : (~^$signed(reg1239[(3'h6):(3'h4)])));
                    end
                  if ($signed(reg1347[(1'h1):(1'h0)]))
                    begin
                      reg1476 <= ($signed($signed($signed((8'haf)))) ?
                          (reg1392 & ((reg1483 == forvar1163) | (reg1196 ?
                              reg1261 : reg1467))) : (^~$signed(((8'ha7) == reg1347))));
                    end
                  else
                    begin
                      reg1476 <= (^($unsigned(forvar1264[(2'h2):(1'h1)]) + {reg1204}));
                      reg1477 <= {($unsigned((-reg1447)) >> $unsigned(reg1400[(3'h7):(2'h2)]))};
                    end
                end
              if (reg1199[(4'hb):(3'h5)])
                begin
                  for (forvar1484 = (1'h0); (forvar1484 < (2'h3)); forvar1484 = (forvar1484 + (1'h1)))
                    begin
                      reg1485 <= reg1162;
                      reg1486 <= $unsigned(((reg1314[(1'h1):(1'h1)] * (reg1302 ?
                              (8'ha7) : forvar1229)) ?
                          {(reg1397 ? reg1284 : forvar1183)} : reg1246));
                      reg1487 <= $unsigned(forvar1480);
                    end
                  for (forvar1488 = (1'h0); (forvar1488 < (2'h2)); forvar1488 = (forvar1488 + (1'h1)))
                    begin
                      reg1489 <= {(|forvar1373)};
                      reg1490 <= reg1381;
                    end
                end
              else
                begin
                  if ((^~reg1208))
                    begin
                      reg1484 <= reg1214[(4'hd):(1'h0)];
                    end
                  else
                    begin
                      reg1484 <= $signed($signed((forvar1201[(3'h6):(2'h3)] <= $signed(forvar1163))));
                    end
                  if ($signed(($signed((reg1340 > reg1154)) << {{reg1173}})))
                    begin
                      reg1485 <= (+(forvar1285[(2'h2):(1'h0)] ?
                          {reg1449[(1'h0):(1'h0)]} : {$signed(reg1400)}));
                      reg1486 <= (($unsigned((reg1229 ?
                          reg1291 : reg1149)) > reg1153[(4'ha):(4'h9)]) && reg1349[(4'he):(4'hc)]);
                    end
                  else
                    begin
                      reg1485 <= (8'hac);
                      reg1486 <= $signed((8'hb5));
                      reg1487 <= reg1449;
                    end
                end
              if (((^{{(8'hb9)}}) < ({{forvar1394}} ?
                  $unsigned((+wire587)) : $signed(reg1325))))
                begin
                  if ((reg1324 < reg1350))
                    begin
                      reg1491 <= {$unsigned(reg1411)};
                      reg1492 <= reg1482[(2'h2):(1'h1)];
                      reg1493 <= (reg1166 ?
                          forvar1168[(3'h7):(2'h2)] : $signed((reg1311 < (reg1189 ?
                              reg1208 : forvar1433))));
                      reg1494 <= $signed(reg1193[(4'h9):(3'h6)]);
                    end
                  else
                    begin
                      reg1491 <= $signed((($unsigned(reg1228) & (reg1306 ?
                          reg1378 : reg1247)) * reg1435));
                      reg1492 <= (forvar1363 ?
                          $signed(((reg1222 & reg1246) ?
                              wire586[(3'h6):(3'h5)] : $unsigned(forvar1148))) : forvar1448);
                      reg1493 <= (&(-$unsigned((&reg1181))));
                    end
                  for (forvar1495 = (1'h0); (forvar1495 < (2'h2)); forvar1495 = (forvar1495 + (1'h1)))
                    begin
                      reg1496 <= reg1479[(1'h0):(1'h0)];
                      reg1497 <= $signed((((&reg1439) ?
                              (forvar1419 ? reg1268 : forvar1394) : ((8'h9e) ?
                                  forvar1212 : (8'hb9))) ?
                          $signed($unsigned(forvar1488)) : $unsigned((-(8'ha7)))));
                      reg1498 <= reg1151[(2'h2):(1'h1)];
                      reg1499 <= $unsigned($signed({(reg1358 ?
                              reg1187 : reg1179)}));
                    end
                  for (forvar1500 = (1'h0); (forvar1500 < (1'h1)); forvar1500 = (forvar1500 + (1'h1)))
                    begin
                      reg1501 <= ({{(^~reg1460)}} >= $signed($signed((^reg1457))));
                    end
                  reg1502 <= (reg1184[(4'he):(3'h5)] + {forvar1246[(2'h2):(2'h2)]});
                end
              else
                begin
                  if ($unsigned(forvar1463))
                    begin
                      reg1491 <= reg1412[(1'h1):(1'h0)];
                      reg1492 <= forvar1314;
                      reg1493 <= (^~(~reg1262[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg1491 <= $signed(forvar1169);
                      reg1492 <= (^~(8'hac));
                      reg1493 <= reg1407;
                    end
                  if ((&(^~reg1231[(4'hd):(1'h0)])))
                    begin
                      reg1494 <= ($unsigned((~^reg1235[(4'hc):(3'h6)])) <= {(8'hb9)});
                      reg1495 <= ($signed(reg1254) <= reg1415[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1494 <= $signed(reg1349);
                      reg1495 <= {(8'ha5)};
                    end
                  for (forvar1496 = (1'h0); (forvar1496 < (1'h1)); forvar1496 = (forvar1496 + (1'h1)))
                    begin
                      reg1497 <= {$unsigned((forvar1438[(4'h9):(2'h3)] >>> $unsigned(reg1352)))};
                      reg1498 <= ((({reg1230} ?
                              (reg1213 ~^ forvar1156) : (reg1348 ?
                                  forvar1446 : reg1196)) ?
                          (reg1502 ?
                              (&reg1171) : $signed(forvar1328)) : $signed((reg1155 <<< forvar1166))) ~^ $signed(forvar1262));
                    end
                end
              if ((8'h9e))
                begin
                  reg1503 <= {forvar1221};
                  for (forvar1504 = (1'h0); (forvar1504 < (1'h1)); forvar1504 = (forvar1504 + (1'h1)))
                    begin
                      reg1505 <= $signed(forvar1409);
                      reg1506 <= (~&reg1243);
                    end
                  if (reg1248)
                    begin
                      reg1507 <= $unsigned($unsigned({$signed(reg1297)}));
                      reg1508 <= $signed(reg1325);
                    end
                  else
                    begin
                      reg1507 <= reg1348;
                    end
                end
              else
                begin
                  if (($unsigned($signed((^~reg1314))) != (forvar1426 ^ ((reg1479 ?
                          forvar1223 : forvar1446) ?
                      (-forvar1484) : (reg1268 > reg1435)))))
                    begin
                      reg1503 <= reg1330;
                      reg1504 <= forvar1153[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1503 <= reg1451[(1'h1):(1'h0)];
                      reg1504 <= (+($unsigned(reg1333) ?
                          (!$unsigned((8'ha5))) : forvar1323));
                      reg1505 <= $signed((((reg1325 == forvar1496) ?
                              forvar1246[(1'h0):(1'h0)] : reg1341[(3'h4):(2'h3)]) ?
                          $signed({reg1422}) : reg1447));
                    end
                  if (forvar1395[(3'h7):(3'h6)])
                    begin
                      reg1506 <= (-(forvar1351 ?
                          ((^forvar1256) >>> $unsigned(reg1336)) : (~$unsigned(reg1405))));
                      reg1507 <= reg1487[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1506 <= $signed($unsigned((!(|reg1448))));
                      reg1507 <= reg1256[(4'h8):(2'h2)];
                    end
                end
            end
        end
    end
  module1509 modinst1736 (.clk(clk), .wire1510(forvar1163), .wire1513(reg1311), .y(wire1735), .wire1512(reg1317), .wire1511(reg1306));
  always
    @(posedge clk) begin
      for (forvar1737 = (1'h0); (forvar1737 < (2'h2)); forvar1737 = (forvar1737 + (1'h1)))
        begin
          reg1738 <= {$signed((forvar1328 ~^ $unsigned(reg1205)))};
          for (forvar1739 = (1'h0); (forvar1739 < (2'h2)); forvar1739 = (forvar1739 + (1'h1)))
            begin
              for (forvar1740 = (1'h0); (forvar1740 < (2'h2)); forvar1740 = (forvar1740 + (1'h1)))
                begin
                  for (forvar1741 = (1'h0); (forvar1741 < (1'h1)); forvar1741 = (forvar1741 + (1'h1)))
                    begin
                      reg1742 <= (^~($signed((~&(8'hb2))) ?
                          reg1200 : $unsigned(reg1439[(1'h1):(1'h0)])));
                      reg1743 <= $signed($signed($unsigned(reg1496[(4'he):(3'h7)])));
                      reg1744 <= $signed((+{(+reg1162)}));
                      reg1745 <= forvar1156[(3'h5):(1'h0)];
                    end
                  for (forvar1746 = (1'h0); (forvar1746 < (1'h0)); forvar1746 = (forvar1746 + (1'h1)))
                    begin
                      reg1747 <= $signed((-$signed(((8'haa) && forvar1348))));
                      reg1748 <= $signed((!$unsigned((~|(8'ha0)))));
                      reg1749 <= $unsigned($signed((~&{reg1297})));
                      reg1750 <= (~|$signed((~&(forvar1462 ?
                          forvar1469 : (8'ha9)))));
                    end
                  if ($unsigned((((forvar1274 >>> reg1750) ^~ $signed(reg1398)) != ($unsigned((8'ha5)) <<< (forvar1298 ?
                      wire589 : (8'ha0))))))
                    begin
                      reg1751 <= (^(^~(8'hb1)));
                      reg1752 <= ({(&(~|reg1187))} != $signed(reg1422));
                      reg1753 <= (reg1328 ?
                          {(|(~|reg1360))} : ((8'h9f) ~^ forvar1251[(3'h6):(1'h1)]));
                    end
                  else
                    begin
                      reg1751 <= ((~|((forvar1363 < (8'hb0)) != $signed(reg1315))) ?
                          (+((&reg1467) >> (8'ha4))) : $signed(reg1229[(1'h1):(1'h0)]));
                    end
                end
            end
          for (forvar1754 = (1'h0); (forvar1754 < (2'h2)); forvar1754 = (forvar1754 + (1'h1)))
            begin
              for (forvar1755 = (1'h0); (forvar1755 < (1'h0)); forvar1755 = (forvar1755 + (1'h1)))
                begin
                  if (reg1461[(1'h0):(1'h0)])
                    begin
                      reg1756 <= reg1332;
                    end
                  else
                    begin
                      reg1756 <= $unsigned((&reg1288[(2'h2):(1'h0)]));
                      reg1757 <= forvar1426[(4'h8):(1'h0)];
                      reg1758 <= (forvar1456 ?
                          ((&wire587) ^ ($signed(reg1201) >>> (reg1437 ?
                              forvar1285 : reg1193))) : $unsigned((|$signed(reg1496))));
                      reg1759 <= $signed($unsigned(forvar1219));
                    end
                  for (forvar1760 = (1'h0); (forvar1760 < (1'h0)); forvar1760 = (forvar1760 + (1'h1)))
                    begin
                      reg1761 <= (({reg1445[(3'h4):(3'h4)]} ?
                          ((~&reg1359) + reg1358[(3'h5):(3'h4)]) : $unsigned(reg1291[(4'ha):(2'h2)])) | ($unsigned(reg1757) ?
                          ((reg1453 & forvar1241) << (reg1353 ?
                              forvar1158 : (8'hb4))) : $signed((^~reg1351))));
                      reg1762 <= (&$signed(forvar1472));
                      reg1763 <= (&(((~&forvar1426) ?
                              (reg1435 && reg1302) : $unsigned(reg1331)) ?
                          ((reg1379 <<< reg1271) ?
                              (forvar1166 ?
                                  (8'haa) : reg1249) : reg1262) : (~^reg1193)));
                      reg1764 <= reg1389;
                    end
                end
              for (forvar1765 = (1'h0); (forvar1765 < (1'h0)); forvar1765 = (forvar1765 + (1'h1)))
                begin
                  if ((reg1199[(4'h9):(3'h4)] ?
                      (reg1247[(2'h3):(1'h1)] ?
                          reg1385[(4'he):(4'hb)] : $signed(forvar1739)) : $unsigned((reg1455 ?
                          (8'hb6) : ((8'hb4) ? reg1346 : reg1172)))))
                    begin
                      reg1766 <= {((~(~|reg1362)) ?
                              (reg1420 < $signed((8'haf))) : ({reg1752} - $unsigned(reg1498)))};
                    end
                  else
                    begin
                      reg1766 <= (~(~^reg1323[(4'h9):(1'h0)]));
                      reg1767 <= (({(forvar1197 ?
                              reg1190 : forvar1151)} ^~ ((reg1467 * forvar1414) >>> (wire588 ^~ reg1246))) ^~ ((((8'ha9) ?
                              forvar1755 : (8'hb4)) != (^(8'hb1))) ?
                          $unsigned((~&reg1297)) : (|((8'ha4) >>> reg1405))));
                    end
                  for (forvar1768 = (1'h0); (forvar1768 < (1'h1)); forvar1768 = (forvar1768 + (1'h1)))
                    begin
                      reg1769 <= $unsigned($signed($unsigned((reg1174 ?
                          forvar1737 : (8'h9f)))));
                      reg1770 <= reg1336[(2'h2):(2'h2)];
                      reg1771 <= reg1251[(2'h3):(1'h0)];
                    end
                end
              for (forvar1772 = (1'h0); (forvar1772 < (2'h3)); forvar1772 = (forvar1772 + (1'h1)))
                begin
                  if ((reg1440 ?
                      forvar1332[(3'h4):(1'h0)] : ({(reg1361 ?
                              forvar1426 : reg1208)} | ((reg1168 ?
                              reg1354 : reg1444) ?
                          reg1248[(2'h2):(1'h1)] : (reg1487 ?
                              reg1265 : reg1161)))))
                    begin
                      reg1773 <= $unsigned($unsigned((8'hb9)));
                    end
                  else
                    begin
                      reg1773 <= (((~forvar1162) << (reg1416 >= (8'hae))) >>> {$signed((reg1339 ?
                              reg1214 : (8'hab)))});
                      reg1774 <= (forvar1183 ?
                          $signed((reg1279[(2'h2):(2'h2)] * $signed(reg1287))) : ({((8'had) ~^ forvar1373)} < {$signed(forvar1306)}));
                      reg1775 <= (+$signed(reg1171[(3'h6):(3'h4)]));
                    end
                  for (forvar1776 = (1'h0); (forvar1776 < (2'h2)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 <= forvar1413;
                      reg1778 <= (reg1193 ?
                          reg1335 : $unsigned($signed((^~(8'haa)))));
                      reg1779 <= reg1273[(2'h2):(1'h0)];
                      reg1780 <= forvar1350;
                    end
                  for (forvar1781 = (1'h0); (forvar1781 < (2'h2)); forvar1781 = (forvar1781 + (1'h1)))
                    begin
                      reg1782 <= ((reg1183[(3'h4):(1'h1)] ?
                              {reg1407} : (^~forvar1384[(3'h5):(3'h4)])) ?
                          $unsigned(($unsigned(reg1377) ?
                              reg1355[(3'h4):(1'h0)] : $signed(reg1377))) : (8'ha4));
                      reg1783 <= ((((&(8'ha4)) ?
                                  (reg1266 ~^ reg1354) : $unsigned((8'hb7))) ?
                              $signed({wire590}) : wire1147) ?
                          (((forvar1269 ?
                              forvar1186 : reg1159) + (reg1232 ~^ reg1197)) <<< reg1402) : forvar1162);
                      reg1784 <= $signed($signed((|$signed(reg1312))));
                      reg1785 <= (reg1382 ?
                          $unsigned(reg1758[(1'h1):(1'h0)]) : ({$unsigned(reg1769)} <= ($signed(reg1780) >>> forvar1419)));
                    end
                  for (forvar1786 = (1'h0); (forvar1786 < (1'h0)); forvar1786 = (forvar1786 + (1'h1)))
                    begin
                      reg1787 <= ((wire590[(1'h0):(1'h0)] ?
                          {(!forvar1250)} : $signed($unsigned(reg1490))) * $signed($signed((reg1243 | reg1334))));
                      reg1788 <= reg1217;
                      reg1789 <= (reg1158[(3'h7):(3'h7)] < $signed(($unsigned(reg1237) ?
                          ((8'h9d) || reg1507) : $signed(reg1784))));
                    end
                end
              for (forvar1790 = (1'h0); (forvar1790 < (2'h2)); forvar1790 = (forvar1790 + (1'h1)))
                begin
                  if ($unsigned((!$unsigned((forvar1291 == reg1747)))))
                    begin
                      reg1791 <= (((reg1350 ?
                              (reg1370 * forvar1285) : $unsigned(forvar1403)) ?
                          $unsigned(reg1215[(1'h1):(1'h0)]) : (~&$unsigned(forvar1209))) + $signed($unsigned({forvar1395})));
                    end
                  else
                    begin
                      reg1791 <= (reg1254 ?
                          reg1751[(2'h3):(2'h2)] : ({(reg1296 <= reg1249)} ?
                              ((~forvar1328) << (8'h9f)) : {(reg1324 ?
                                      reg1475 : (8'hb9))}));
                    end
                  for (forvar1792 = (1'h0); (forvar1792 < (1'h0)); forvar1792 = (forvar1792 + (1'h1)))
                    begin
                      reg1793 <= (reg1421 ^ ((reg1156[(3'h4):(3'h4)] ?
                              $signed(reg1216) : reg1223) ?
                          $unsigned($unsigned(reg1466)) : (8'hb9)));
                      reg1794 <= (&(forvar1472[(2'h2):(1'h1)] ?
                          $unsigned((reg1280 ? reg1158 : reg1446)) : reg1230));
                      reg1795 <= reg1399;
                    end
                  reg1796 <= $signed($signed((!reg1272[(3'h6):(1'h1)])));
                  if ((forvar1306 <= (-forvar1213)))
                    begin
                      reg1797 <= ((8'ha3) | $unsigned((8'had)));
                      reg1798 <= ($unsigned($signed(reg1209[(3'h4):(1'h0)])) == {(8'haa)});
                      reg1799 <= forvar1157;
                      reg1800 <= forvar1239;
                    end
                  else
                    begin
                      reg1797 <= (8'ha9);
                      reg1798 <= {$unsigned(reg1254)};
                      reg1799 <= reg1429;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg1801 <= $unsigned($signed(reg1180[(3'h4):(2'h3)]));
      for (forvar1802 = (1'h0); (forvar1802 < (2'h3)); forvar1802 = (forvar1802 + (1'h1)))
        begin
          if ($signed($signed($signed({(8'ha0)}))))
            begin
              if ($unsigned($unsigned($unsigned({reg1388}))))
                begin
                  reg1803 <= reg1474[(2'h2):(1'h0)];
                end
              else
                begin
                  if (({reg1492} ?
                      (~&(wire585[(2'h3):(2'h3)] & (reg1434 ?
                          reg1150 : reg1343))) : (($signed(forvar1323) ?
                          $unsigned(reg1296) : $unsigned((8'hb4))) >>> forvar1469[(4'hd):(3'h5)])))
                    begin
                      reg1803 <= $signed(reg1249[(1'h1):(1'h1)]);
                      reg1804 <= $unsigned(reg1230);
                    end
                  else
                    begin
                      reg1803 <= reg1378;
                      reg1804 <= reg1480[(3'h4):(3'h4)];
                    end
                  reg1805 <= $signed(reg1465[(3'h7):(3'h5)]);
                  if (reg1357)
                    begin
                      reg1806 <= $signed(((8'h9e) <<< reg1407[(3'h7):(1'h1)]));
                      reg1807 <= (+{(reg1355[(4'ha):(2'h2)] & (reg1204 <= reg1778))});
                      reg1808 <= {((reg1223[(2'h3):(2'h3)] * forvar1393[(3'h5):(3'h5)]) >= (~|$signed(reg1436)))};
                    end
                  else
                    begin
                      reg1806 <= reg1375;
                      reg1807 <= (((^~(8'hb6)) ?
                              forvar1348[(4'hb):(4'h9)] : reg1487) ?
                          ($unsigned((reg1235 ?
                              forvar1496 : reg1230)) != $signed((forvar1219 ?
                              wire1147 : reg1340))) : $signed($signed(reg1222[(3'h7):(1'h1)])));
                      reg1808 <= reg1234[(4'hd):(4'hb)];
                    end
                end
              if ($unsigned($unsigned(((-reg1217) & forvar1430[(2'h2):(1'h0)]))))
                begin
                  for (forvar1809 = (1'h0); (forvar1809 < (1'h1)); forvar1809 = (forvar1809 + (1'h1)))
                    begin
                      reg1810 <= forvar1809;
                      reg1811 <= (~^($unsigned(forvar1162) ^~ $signed((reg1320 >>> reg1193))));
                      reg1812 <= (reg1377 ?
                          reg1472 : $signed(($unsigned(forvar1221) >> {reg1441})));
                    end
                  for (forvar1813 = (1'h0); (forvar1813 < (2'h2)); forvar1813 = (forvar1813 + (1'h1)))
                    begin
                      reg1814 <= $signed({({reg1464} ?
                              $unsigned(reg1445) : $signed(reg1370))});
                      reg1815 <= forvar1290;
                      reg1816 <= (^(($unsigned((8'h9e)) <= reg1392[(1'h1):(1'h1)]) > $unsigned((~forvar1454))));
                      reg1817 <= reg1407;
                    end
                end
              else
                begin
                  for (forvar1809 = (1'h0); (forvar1809 < (2'h2)); forvar1809 = (forvar1809 + (1'h1)))
                    begin
                      reg1810 <= $unsigned($signed(reg1290[(4'ha):(4'ha)]));
                    end
                  if ((reg1464[(3'h4):(1'h1)] - ((|(|reg1338)) ?
                      {(reg1795 || forvar1243)} : ($signed(reg1313) ?
                          (^~reg1487) : (forvar1354 < reg1259)))))
                    begin
                      reg1811 <= reg1800;
                      reg1812 <= (8'hb1);
                    end
                  else
                    begin
                      reg1811 <= ((((^forvar1393) ?
                                  $signed(reg1227) : (reg1372 != reg1496)) ?
                              $unsigned(reg1318[(5'h10):(1'h0)]) : (~&reg1356)) ?
                          reg1238[(3'h5):(2'h3)] : $unsigned({$signed(reg1277)}));
                      reg1812 <= $signed((({forvar1262} ?
                          {reg1771} : $signed(forvar1351)) != (8'hb6)));
                    end
                  if (reg1312)
                    begin
                      reg1813 <= forvar1298;
                      reg1814 <= (8'ha9);
                      reg1815 <= ((~^{$unsigned(reg1369)}) ?
                          reg1767 : reg1769[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg1813 <= $unsigned($signed(reg1375));
                      reg1814 <= $signed($signed((((8'ha7) | reg1271) << {(8'ha3)})));
                      reg1815 <= ($signed((~{reg1473})) * (reg1225 >= forvar1384[(1'h0):(1'h0)]));
                    end
                  for (forvar1816 = (1'h0); (forvar1816 < (1'h1)); forvar1816 = (forvar1816 + (1'h1)))
                    begin
                      reg1817 <= {forvar1177[(1'h0):(1'h0)]};
                      reg1818 <= ({$unsigned(reg1470[(4'ha):(1'h0)])} ?
                          $signed(((forvar1213 - reg1782) ?
                              wire585[(2'h2):(1'h0)] : $unsigned((8'h9f)))) : $signed((reg1232 ?
                              (|reg1193) : (~&(8'ha9)))));
                      reg1819 <= (($unsigned($signed((8'ha1))) ?
                          ($unsigned(reg1301) ^~ reg1165[(4'h8):(3'h7)]) : reg1172) ^ reg1425[(3'h7):(3'h5)]);
                      reg1820 <= $unsigned(forvar1239);
                    end
                end
            end
          else
            begin
              for (forvar1803 = (1'h0); (forvar1803 < (1'h1)); forvar1803 = (forvar1803 + (1'h1)))
                begin
                  if (reg1286[(4'hb):(2'h3)])
                    begin
                      reg1804 <= $signed(((forvar1250[(1'h0):(1'h0)] ?
                          $signed((8'ha2)) : (reg1233 && forvar1323)) >= (reg1291[(1'h0):(1'h0)] != ((8'hac) + (8'hb2)))));
                      reg1805 <= $unsigned(forvar1169);
                      reg1806 <= ((^~{(reg1390 ?
                              reg1182 : reg1184)}) < ($unsigned((^~reg1234)) == reg1266[(4'h9):(3'h5)]));
                    end
                  else
                    begin
                      reg1804 <= (forvar1233 + (-$unsigned($unsigned(reg1478))));
                    end
                end
              for (forvar1807 = (1'h0); (forvar1807 < (1'h0)); forvar1807 = (forvar1807 + (1'h1)))
                begin
                  for (forvar1808 = (1'h0); (forvar1808 < (2'h3)); forvar1808 = (forvar1808 + (1'h1)))
                    begin
                      reg1809 <= reg1442[(2'h2):(1'h0)];
                    end
                end
              reg1810 <= reg1381[(2'h3):(1'h1)];
            end
          for (forvar1821 = (1'h0); (forvar1821 < (1'h0)); forvar1821 = (forvar1821 + (1'h1)))
            begin
              for (forvar1822 = (1'h0); (forvar1822 < (2'h2)); forvar1822 = (forvar1822 + (1'h1)))
                begin
                  reg1823 <= $signed($signed(((+forvar1157) ?
                      (reg1259 * (8'ha6)) : (reg1301 >>> reg1255))));
                end
            end
          reg1824 <= ($unsigned(reg1431[(3'h6):(3'h6)]) * ($unsigned(reg1213[(1'h0):(1'h0)]) ?
              wire1147 : reg1759[(2'h2):(1'h0)]));
          reg1825 <= $signed(forvar1469[(1'h1):(1'h0)]);
        end
    end
  always
    @(posedge clk) begin
      reg1826 <= (!(((~|forvar1755) != (forvar1363 ? reg1816 : reg1357)) ?
          forvar1426 : ($unsigned(reg1508) | reg1787)));
      reg1827 <= ({({reg1410} + {reg1400})} ?
          reg1763[(4'he):(4'hd)] : {$unsigned((&reg1472))});
      if (reg1167)
        begin
          if ($signed(reg1815[(3'h4):(2'h2)]))
            begin
              if (reg1180)
                begin
                  reg1828 <= reg1287[(1'h1):(1'h0)];
                  if ((-reg1176))
                    begin
                      reg1829 <= (8'hac);
                      reg1830 <= $signed(($unsigned(reg1389) * (^~forvar1207)));
                    end
                  else
                    begin
                      reg1829 <= $signed($unsigned(($unsigned(reg1779) ?
                          $unsigned(forvar1807) : reg1759[(1'h1):(1'h0)])));
                    end
                  for (forvar1831 = (1'h0); (forvar1831 < (2'h3)); forvar1831 = (forvar1831 + (1'h1)))
                    begin
                      reg1832 <= ((reg1379[(4'hb):(2'h3)] <= (+(forvar1226 ?
                          (8'hb0) : reg1276))) >> (^~$signed((reg1745 ?
                          reg1418 : reg1265))));
                      reg1833 <= $signed($unsigned(((reg1824 ?
                              reg1487 : wire590) ?
                          (+forvar1251) : forvar1394[(4'h9):(4'h8)])));
                      reg1834 <= (~&({(forvar1281 ? forvar1168 : reg1232)} ?
                          reg1233[(1'h0):(1'h0)] : $unsigned(reg1417[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  if (forvar1419[(3'h7):(2'h3)])
                    begin
                      reg1828 <= $unsigned(($signed($unsigned(reg1168)) ~^ reg1187[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg1828 <= (forvar1479 ?
                          reg1434[(4'he):(4'hc)] : (~^((8'h9c) ?
                              {forvar1469} : (reg1457 == (8'hb9)))));
                      reg1829 <= (^~($signed((-forvar1306)) ?
                          ((reg1246 ? (8'haf) : reg1369) ?
                              forvar1816 : $signed(reg1369)) : $signed((forvar1394 == reg1163))));
                      reg1830 <= (~|{(reg1471 ? (+reg1217) : forvar1149)});
                      reg1831 <= {$signed((forvar1149 ?
                              (!(8'ha4)) : ((8'had) ? (8'ha9) : forvar1196)))};
                    end
                end
              reg1835 <= $unsigned((!((reg1320 ? reg1464 : reg1315) ?
                  forvar1370 : $signed(reg1228))));
              for (forvar1836 = (1'h0); (forvar1836 < (2'h2)); forvar1836 = (forvar1836 + (1'h1)))
                begin
                  for (forvar1837 = (1'h0); (forvar1837 < (1'h0)); forvar1837 = (forvar1837 + (1'h1)))
                    begin
                      reg1838 <= ({(~|(reg1380 ^~ reg1271))} ?
                          (!(~&reg1195[(4'h9):(1'h1)])) : (reg1829 | $unsigned($unsigned(reg1438))));
                    end
                end
              reg1839 <= $unsigned({reg1229});
            end
          else
            begin
              for (forvar1828 = (1'h0); (forvar1828 < (1'h0)); forvar1828 = (forvar1828 + (1'h1)))
                begin
                  reg1829 <= (+$signed(($unsigned(reg1227) ?
                      $signed(reg1354) : (~^forvar1210))));
                  for (forvar1830 = (1'h0); (forvar1830 < (2'h3)); forvar1830 = (forvar1830 + (1'h1)))
                    begin
                      reg1831 <= $unsigned(($signed(((8'h9c) ?
                              (8'ha1) : (8'hb7))) ?
                          reg1489 : (~^forvar1214)));
                      reg1832 <= $signed($unsigned(forvar1792[(1'h1):(1'h0)]));
                      reg1833 <= (8'haf);
                      reg1834 <= reg1789;
                    end
                  for (forvar1835 = (1'h0); (forvar1835 < (2'h2)); forvar1835 = (forvar1835 + (1'h1)))
                    begin
                      reg1836 <= $signed((^~$unsigned({reg1257})));
                      reg1837 <= (~&(^~$unsigned(reg1494)));
                      reg1838 <= (&({(!forvar1496)} == (reg1431[(3'h5):(1'h1)] - reg1189[(2'h2):(1'h1)])));
                    end
                end
              if ((8'haf))
                begin
                  reg1839 <= reg1411[(4'ha):(3'h5)];
                end
              else
                begin
                  for (forvar1839 = (1'h0); (forvar1839 < (2'h2)); forvar1839 = (forvar1839 + (1'h1)))
                    begin
                      reg1840 <= reg1785[(3'h4):(2'h2)];
                      reg1841 <= $unsigned((8'hb3));
                      reg1842 <= (^~reg1485[(2'h2):(1'h1)]);
                    end
                end
            end
        end
      else
        begin
          if ($unsigned($unsigned({forvar1414[(1'h1):(1'h0)]})))
            begin
              for (forvar1828 = (1'h0); (forvar1828 < (2'h3)); forvar1828 = (forvar1828 + (1'h1)))
                begin
                  reg1829 <= reg1190;
                end
              for (forvar1830 = (1'h0); (forvar1830 < (1'h1)); forvar1830 = (forvar1830 + (1'h1)))
                begin
                  for (forvar1831 = (1'h0); (forvar1831 < (2'h3)); forvar1831 = (forvar1831 + (1'h1)))
                    begin
                      reg1832 <= reg1212[(3'h5):(2'h3)];
                      reg1833 <= $signed((($signed((8'ha8)) ?
                              $unsigned(reg1448) : (|reg1242)) ?
                          $unsigned((|reg1401)) : ((reg1189 ?
                                  (8'ha3) : reg1493) ?
                              (8'ha0) : forvar1790)));
                      reg1834 <= reg1244;
                    end
                  if (((($unsigned(reg1482) ? {reg1309} : (reg1809 + reg1390)) ?
                      $unsigned(forvar1807) : {reg1808[(1'h0):(1'h0)]}) > ((|(^~forvar1504)) - ($unsigned(reg1369) & {forvar1157}))))
                    begin
                      reg1835 <= (reg1364[(1'h0):(1'h0)] || $signed((^~reg1229[(2'h2):(1'h1)])));
                      reg1836 <= $unsigned($unsigned((((8'h9d) ?
                          (8'had) : reg1405) * reg1825)));
                      reg1837 <= $signed((((|reg1157) >>> {(8'ha8)}) ?
                          (^~reg1381[(3'h5):(1'h0)]) : {$unsigned(forvar1161)}));
                    end
                  else
                    begin
                      reg1835 <= reg1355;
                      reg1836 <= (~&reg1229);
                      reg1837 <= $signed(reg1249[(3'h4):(2'h2)]);
                      reg1838 <= reg1177;
                    end
                  reg1839 <= forvar1212;
                  for (forvar1840 = (1'h0); (forvar1840 < (2'h2)); forvar1840 = (forvar1840 + (1'h1)))
                    begin
                      reg1841 <= (({(forvar1202 > reg1174)} & ((|reg1423) && reg1478[(4'hd):(2'h2)])) ?
                          reg1484[(1'h0):(1'h0)] : reg1163[(1'h1):(1'h0)]);
                      reg1842 <= (!($signed(reg1376) ? reg1397 : reg1227));
                      reg1843 <= $unsigned({$unsigned($signed(reg1262))});
                    end
                end
              if ((~$unsigned((forvar1330 ?
                  (~|reg1828) : (reg1216 ? reg1435 : (8'hb1))))))
                begin
                  for (forvar1844 = (1'h0); (forvar1844 < (2'h2)); forvar1844 = (forvar1844 + (1'h1)))
                    begin
                      reg1845 <= {({$unsigned(forvar1500)} < reg1219)};
                      reg1846 <= forvar1807[(3'h7):(2'h3)];
                    end
                end
              else
                begin
                  if ($unsigned(forvar1480[(2'h3):(1'h0)]))
                    begin
                      reg1844 <= $unsigned($unsigned($signed($signed(forvar1223))));
                      reg1845 <= (-reg1154[(1'h1):(1'h0)]);
                      reg1846 <= ($signed($unsigned((forvar1161 == reg1260))) < reg1345);
                    end
                  else
                    begin
                      reg1844 <= (reg1233[(2'h2):(1'h1)] < (&{(forvar1480 <= reg1308)}));
                    end
                  reg1847 <= reg1823;
                  if ($signed(reg1243[(1'h1):(1'h0)]))
                    begin
                      reg1848 <= (forvar1167[(3'h4):(1'h0)] <<< reg1459);
                      reg1849 <= $unsigned($unsigned(forvar1239[(4'ha):(4'h9)]));
                    end
                  else
                    begin
                      reg1848 <= $unsigned({((reg1196 | reg1823) | (+reg1849))});
                      reg1849 <= $signed(reg1470);
                      reg1850 <= ((((^reg1349) >>> (~|reg1457)) != {(reg1794 >> reg1480)}) >= (|(reg1458[(3'h4):(1'h1)] * reg1766)));
                    end
                end
            end
          else
            begin
              for (forvar1828 = (1'h0); (forvar1828 < (1'h0)); forvar1828 = (forvar1828 + (1'h1)))
                begin
                  if ({(^$signed(reg1370[(2'h3):(2'h3)]))})
                    begin
                      reg1829 <= (+reg1209[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1829 <= $signed($signed(({forvar1337} ?
                          $signed(forvar1290) : forvar1463[(3'h5):(2'h2)])));
                      reg1830 <= {$unsigned($unsigned((reg1154 ?
                              forvar1822 : reg1178)))};
                      reg1831 <= $signed({$unsigned(((8'ha6) < reg1481))});
                    end
                  reg1832 <= reg1219;
                  for (forvar1833 = (1'h0); (forvar1833 < (1'h0)); forvar1833 = (forvar1833 + (1'h1)))
                    begin
                      reg1834 <= $unsigned(reg1321);
                      reg1835 <= (forvar1450 ?
                          {(reg1749[(1'h1):(1'h1)] ?
                                  reg1406[(1'h0):(1'h0)] : (~|reg1369))} : $unsigned(($signed(reg1323) ?
                              forvar1772 : reg1497)));
                      reg1836 <= reg1247;
                    end
                  for (forvar1837 = (1'h0); (forvar1837 < (1'h0)); forvar1837 = (forvar1837 + (1'h1)))
                    begin
                      reg1838 <= ($unsigned(reg1489) ?
                          ($unsigned(reg1788) ^~ ($unsigned((8'ha2)) ?
                              (reg1327 + reg1169) : $unsigned(reg1303))) : (!(reg1757[(1'h1):(1'h0)] <<< (8'hb4))));
                    end
                end
              if (($signed({{reg1816}}) > $unsigned((~|(forvar1214 ?
                  reg1199 : forvar1265)))))
                begin
                  for (forvar1839 = (1'h0); (forvar1839 < (1'h0)); forvar1839 = (forvar1839 + (1'h1)))
                    begin
                      reg1840 <= $unsigned(($signed((&forvar1305)) && ((-reg1421) << reg1225[(3'h5):(1'h1)])));
                      reg1841 <= reg1340;
                      reg1842 <= (!(~&(reg1820[(4'h8):(2'h3)] < $unsigned(forvar1186))));
                    end
                  if (reg1388[(2'h3):(1'h0)])
                    begin
                      reg1843 <= (($signed(((8'hba) ? forvar1169 : (8'hb7))) ?
                          (reg1831 ?
                              reg1421[(1'h1):(1'h0)] : (8'ha4)) : ((~reg1183) | $signed(reg1389))) - $unsigned($unsigned(reg1445)));
                      reg1844 <= $unsigned($signed((8'ha5)));
                      reg1845 <= (~|{($signed(reg1342) + wire586[(4'h8):(1'h1)])});
                      reg1846 <= $signed($unsigned((reg1412[(2'h2):(2'h2)] ?
                          $unsigned(forvar1251) : reg1267)));
                    end
                  else
                    begin
                      reg1843 <= ($unsigned((~^(forvar1334 >>> reg1767))) <<< reg1816);
                      reg1844 <= reg1340[(1'h0):(1'h0)];
                      reg1845 <= reg1824[(4'h8):(3'h7)];
                    end
                  if (forvar1786)
                    begin
                      reg1847 <= $signed(reg1399[(1'h0):(1'h0)]);
                      reg1848 <= (forvar1285 ?
                          $unsigned(((~reg1367) >> $unsigned((8'haa)))) : reg1484);
                      reg1849 <= (~^((|$signed(reg1457)) ?
                          (reg1815[(2'h2):(1'h0)] ?
                              $unsigned(reg1205) : $unsigned((8'hb4))) : ($signed((8'had)) ?
                              (^~forvar1463) : $signed(reg1216))));
                    end
                  else
                    begin
                      reg1847 <= (forvar1781[(1'h0):(1'h0)] ?
                          (&{(forvar1831 | reg1324)}) : $signed({(reg1229 ?
                                  (8'hae) : reg1752)}));
                      reg1848 <= (^$signed(reg1162));
                      reg1849 <= ($unsigned(reg1274) ~^ $signed(forvar1179[(1'h0):(1'h0)]));
                      reg1850 <= ((~&forvar1231[(2'h2):(2'h2)]) ?
                          $unsigned(forvar1231[(1'h1):(1'h1)]) : ({(8'hab)} ?
                              forvar1394 : {reg1301[(4'hc):(3'h5)]}));
                    end
                end
              else
                begin
                  if (reg1194)
                    begin
                      reg1839 <= $unsigned(reg1157);
                    end
                  else
                    begin
                      reg1839 <= forvar1741[(3'h5):(2'h3)];
                      reg1840 <= $signed(reg1795[(1'h0):(1'h0)]);
                    end
                  reg1841 <= $signed($unsigned(reg1475));
                  reg1842 <= $unsigned(reg1274[(2'h3):(1'h0)]);
                  reg1843 <= reg1831;
                end
            end
          for (forvar1851 = (1'h0); (forvar1851 < (2'h2)); forvar1851 = (forvar1851 + (1'h1)))
            begin
              reg1852 <= reg1339;
              for (forvar1853 = (1'h0); (forvar1853 < (2'h3)); forvar1853 = (forvar1853 + (1'h1)))
                begin
                  if ({(((^~reg1292) ?
                          (forvar1384 ? forvar1426 : reg1825) : ((8'hac) ?
                              forvar1433 : reg1767)) == {((8'h9d) & reg1280)})})
                    begin
                      reg1854 <= ((wire587[(4'hc):(4'h8)] <<< forvar1430) >>> $signed((&(^~reg1347))));
                      reg1855 <= reg1297;
                      reg1856 <= (8'h9f);
                      reg1857 <= $unsigned(forvar1180);
                    end
                  else
                    begin
                      reg1854 <= (|(($unsigned(reg1157) ?
                          (-reg1276) : reg1847[(2'h3):(2'h3)]) >>> (&(reg1195 >> reg1785))));
                      reg1855 <= reg1437;
                    end
                  if ($signed((|reg1218[(2'h2):(2'h2)])))
                    begin
                      reg1858 <= {($unsigned((reg1502 ?
                              forvar1224 : reg1857)) >> ((reg1197 < reg1303) ?
                              (reg1778 == forvar1330) : (reg1177 & reg1183)))};
                      reg1859 <= ((8'ha2) <= (({forvar1259} ?
                          (reg1294 && forvar1472) : $unsigned(forvar1232)) >> reg1473[(3'h6):(1'h0)]));
                    end
                  else
                    begin
                      reg1858 <= $signed(((-forvar1228[(1'h1):(1'h1)]) ?
                          {forvar1809[(2'h2):(1'h1)]} : ((reg1289 + forvar1261) ?
                              {reg1806} : $unsigned((8'hb0)))));
                    end
                  if ($signed($unsigned(reg1275[(1'h1):(1'h0)])))
                    begin
                      reg1860 <= {reg1149[(3'h6):(3'h6)]};
                      reg1861 <= reg1474;
                      reg1862 <= (reg1742[(3'h5):(1'h0)] ?
                          {((forvar1414 ^~ reg1358) ?
                                  $unsigned((8'hb3)) : forvar1772[(1'h0):(1'h0)])} : reg1189[(3'h7):(2'h2)]);
                    end
                  else
                    begin
                      reg1860 <= ((wire1145 ?
                          {(reg1859 > forvar1792)} : (reg1337 <<< reg1793[(4'hc):(4'h9)])) - $unsigned(reg1465[(1'h0):(1'h0)]));
                    end
                end
              if (forvar1157)
                begin
                  if ($signed((~|reg1306[(4'h8):(2'h3)])))
                    begin
                      reg1863 <= (({((8'hae) || (8'had))} ?
                          $signed((^~forvar1171)) : (+(forvar1256 ?
                              (8'hb8) : reg1369))) && forvar1229);
                    end
                  else
                    begin
                      reg1863 <= (8'ha5);
                      reg1864 <= ($unsigned((((8'ha6) == reg1838) > $unsigned(reg1400))) && $unsigned(($signed((8'hac)) ?
                          forvar1269 : (~reg1378))));
                      reg1865 <= $signed($signed($signed($unsigned(reg1201))));
                      reg1866 <= forvar1840[(3'h7):(2'h3)];
                    end
                  reg1867 <= reg1249[(4'h8):(3'h6)];
                  reg1868 <= {{reg1177}};
                end
              else
                begin
                  for (forvar1863 = (1'h0); (forvar1863 < (1'h1)); forvar1863 = (forvar1863 + (1'h1)))
                    begin
                      reg1864 <= $signed($unsigned($unsigned(forvar1836[(3'h4):(2'h3)])));
                      reg1865 <= (^((reg1469[(2'h2):(1'h1)] >= ((8'hba) << forvar1450)) << $signed($signed(reg1353))));
                      reg1866 <= forvar1409;
                    end
                end
              for (forvar1869 = (1'h0); (forvar1869 < (2'h3)); forvar1869 = (forvar1869 + (1'h1)))
                begin
                  for (forvar1870 = (1'h0); (forvar1870 < (2'h2)); forvar1870 = (forvar1870 + (1'h1)))
                    begin
                      reg1871 <= {$signed($unsigned((~|forvar1246)))};
                    end
                  for (forvar1872 = (1'h0); (forvar1872 < (1'h0)); forvar1872 = (forvar1872 + (1'h1)))
                    begin
                      reg1873 <= (~^(~$unsigned({reg1301})));
                    end
                  for (forvar1874 = (1'h0); (forvar1874 < (2'h3)); forvar1874 = (forvar1874 + (1'h1)))
                    begin
                      reg1875 <= (~^$signed(((8'hb8) <<< (&reg1507))));
                    end
                  reg1876 <= $unsigned(reg1168);
                end
            end
          for (forvar1877 = (1'h0); (forvar1877 < (2'h3)); forvar1877 = (forvar1877 + (1'h1)))
            begin
              for (forvar1878 = (1'h0); (forvar1878 < (2'h3)); forvar1878 = (forvar1878 + (1'h1)))
                begin
                  for (forvar1879 = (1'h0); (forvar1879 < (1'h1)); forvar1879 = (forvar1879 + (1'h1)))
                    begin
                      reg1880 <= ({{$signed(reg1818)}} ?
                          ($unsigned((-(8'hba))) >>> $signed($unsigned(reg1336))) : (forvar1878[(3'h5):(1'h1)] <= (~forvar1863)));
                      reg1881 <= (reg1153 && forvar1391);
                      reg1882 <= reg1775;
                      reg1883 <= (~^reg1344[(3'h7):(2'h3)]);
                    end
                  for (forvar1884 = (1'h0); (forvar1884 < (1'h0)); forvar1884 = (forvar1884 + (1'h1)))
                    begin
                      reg1885 <= ($unsigned($signed($signed(reg1388))) ?
                          (((reg1813 <<< forvar1354) && reg1239) && (forvar1271[(2'h3):(2'h3)] ?
                              $unsigned((8'ha4)) : $unsigned(reg1346))) : ($unsigned($unsigned(forvar1414)) > ($signed((8'ha6)) <<< (reg1157 << reg1412))));
                      reg1886 <= reg1800[(1'h0):(1'h0)];
                      reg1887 <= ((((reg1215 ?
                              reg1209 : reg1833) | reg1239[(3'h5):(1'h1)]) ?
                          ((reg1864 > reg1169) ?
                              ((8'hb2) ?
                                  (8'hb3) : (8'hb4)) : {forvar1872}) : reg1820[(3'h7):(3'h7)]) & (8'ha7));
                      reg1888 <= (-$signed(($signed(reg1348) ?
                          {reg1437} : (reg1451 != reg1458))));
                    end
                  for (forvar1889 = (1'h0); (forvar1889 < (1'h1)); forvar1889 = (forvar1889 + (1'h1)))
                    begin
                      reg1890 <= (reg1775 + $signed(reg1201));
                    end
                end
              for (forvar1891 = (1'h0); (forvar1891 < (2'h2)); forvar1891 = (forvar1891 + (1'h1)))
                begin
                  reg1892 <= (reg1887 ?
                      $unsigned((~|(8'hb1))) : ({reg1186[(3'h4):(2'h3)]} == $unsigned(reg1800)));
                  if (reg1842[(2'h2):(1'h1)])
                    begin
                      reg1893 <= ((forvar1394[(3'h4):(2'h2)] <<< (((8'ha5) ?
                              forvar1201 : forvar1306) > $signed(reg1829))) ?
                          ($signed(reg1265) >= (-(8'hb8))) : $signed((^~(!reg1448))));
                    end
                  else
                    begin
                      reg1893 <= forvar1247;
                    end
                  if (forvar1443)
                    begin
                      reg1894 <= reg1455[(2'h2):(1'h1)];
                      reg1895 <= $unsigned((($signed(reg1170) ?
                              (~^reg1469) : (reg1243 != reg1504)) ?
                          forvar1273[(4'ha):(4'h8)] : (((8'hb4) << (8'ha7)) <<< forvar1186[(2'h2):(1'h0)])));
                      reg1896 <= $signed($signed({(!(8'hb9))}));
                    end
                  else
                    begin
                      reg1894 <= ($unsigned($signed(reg1749)) ?
                          ($signed($unsigned(reg1886)) || (reg1446 * (&(8'had)))) : (((~|reg1785) ?
                                  forvar1844[(3'h5):(3'h4)] : reg1481) ?
                              (8'hb5) : (~|$unsigned((8'hb3)))));
                      reg1895 <= reg1751;
                      reg1896 <= $signed((forvar1314[(3'h6):(3'h4)] != reg1795));
                    end
                  reg1897 <= reg1211[(3'h6):(1'h0)];
                end
              for (forvar1898 = (1'h0); (forvar1898 < (2'h3)); forvar1898 = (forvar1898 + (1'h1)))
                begin
                  if (reg1434[(4'h8):(4'h8)])
                    begin
                      reg1899 <= ($signed((forvar1298[(1'h0):(1'h0)] & (reg1452 >> forvar1354))) ?
                          $unsigned($signed(reg1200[(3'h6):(3'h4)])) : (reg1244[(2'h2):(1'h0)] | ({reg1421} < $signed(reg1389))));
                      reg1900 <= reg1886;
                    end
                  else
                    begin
                      reg1899 <= ($unsigned($signed({reg1346})) ?
                          $signed(forvar1746[(2'h2):(1'h0)]) : reg1442);
                      reg1900 <= reg1863[(1'h1):(1'h1)];
                      reg1901 <= ($signed($unsigned(reg1168)) * reg1881);
                      reg1902 <= $signed(((wire590[(3'h6):(2'h3)] ?
                          reg1893[(2'h3):(1'h0)] : reg1227[(2'h2):(2'h2)]) ^ forvar1889));
                    end
                  reg1903 <= (+reg1373);
                  if (reg1270)
                    begin
                      reg1904 <= reg1388[(3'h4):(2'h2)];
                      reg1905 <= ((reg1460 - $unsigned($signed(reg1823))) <<< (({reg1902} ?
                              (forvar1878 ^ reg1833) : $signed((8'h9c))) ?
                          (|$unsigned(wire1145)) : forvar1201[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg1904 <= forvar1755;
                      reg1905 <= reg1196[(2'h3):(1'h1)];
                      reg1906 <= ($signed($signed(reg1252)) ?
                          reg1436[(4'h8):(1'h1)] : $signed({(forvar1469 ?
                                  (8'ha8) : reg1436)}));
                      reg1907 <= $signed(($signed((reg1241 & forvar1809)) | reg1859[(3'h6):(2'h3)]));
                    end
                  if (reg1404)
                    begin
                      reg1908 <= forvar1760;
                      reg1909 <= reg1397;
                      reg1910 <= ($signed(reg1155[(1'h1):(1'h1)]) > ((8'haa) == ($signed((8'hb6)) >= (reg1307 - reg1174))));
                    end
                  else
                    begin
                      reg1908 <= {($signed((+(8'hb7))) >> $signed($unsigned(reg1471)))};
                      reg1909 <= $unsigned((((forvar1163 || reg1384) ?
                          (8'hb6) : {(8'hac)}) | $signed((reg1329 ?
                          reg1823 : reg1327))));
                    end
                end
              for (forvar1911 = (1'h0); (forvar1911 < (1'h1)); forvar1911 = (forvar1911 + (1'h1)))
                begin
                  reg1912 <= $unsigned($signed(forvar1737[(1'h0):(1'h0)]));
                  reg1913 <= (reg1799[(2'h2):(1'h1)] > reg1378);
                end
            end
          for (forvar1914 = (1'h0); (forvar1914 < (1'h0)); forvar1914 = (forvar1914 + (1'h1)))
            begin
              for (forvar1915 = (1'h0); (forvar1915 < (1'h0)); forvar1915 = (forvar1915 + (1'h1)))
                begin
                  for (forvar1916 = (1'h0); (forvar1916 < (2'h2)); forvar1916 = (forvar1916 + (1'h1)))
                    begin
                      reg1917 <= (-$unsigned(((forvar1408 ? reg1490 : (8'haf)) ?
                          (8'hb5) : {reg1206})));
                      reg1918 <= $unsigned(((((8'hba) <<< forvar1741) ?
                          (reg1269 * (8'ha4)) : (|reg1241)) < reg1834[(1'h0):(1'h0)]));
                    end
                  if ($signed($unsigned($unsigned(reg1797))))
                    begin
                      reg1919 <= $unsigned((&forvar1151));
                      reg1920 <= (8'h9c);
                      reg1921 <= forvar1426;
                    end
                  else
                    begin
                      reg1919 <= $signed({forvar1836[(4'h8):(4'h8)]});
                      reg1920 <= $unsigned((8'hb2));
                    end
                end
            end
        end
    end
  assign wire1922 = $unsigned((~|forvar1438));
  module1923 modinst2668 (.clk(clk), .y(wire2667), .wire1925(reg1255), .wire1924(reg1283), .wire1926(reg1203), .wire1927(forvar1165), .wire1928(reg1767));
  assign wire2669 = (-reg1322);
  assign wire2670 = ($unsigned((reg1331[(4'h8):(3'h4)] && forvar1446)) > reg1215[(3'h5):(2'h2)]);
  assign wire2671 = (~^{(8'ha3)});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module287  (y, clk, wire292, wire291, wire290, wire289, wire288);
  output wire [(32'hd6a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire292;
  input wire signed [(4'hb):(1'h0)] wire291;
  input wire signed [(5'h10):(1'h0)] wire290;
  input wire signed [(4'ha):(1'h0)] wire289;
  input wire [(4'h8):(1'h0)] wire288;
  wire [(4'ha):(1'h0)] wire580;
  wire [(4'hf):(1'h0)] wire579;
  wire [(4'ha):(1'h0)] wire578;
  wire signed [(5'h10):(1'h0)] wire577;
  reg [(2'h2):(1'h0)] reg576 = (1'h0);
  reg [(4'hf):(1'h0)] reg575 = (1'h0);
  reg [(3'h5):(1'h0)] reg574 = (1'h0);
  reg [(5'h10):(1'h0)] forvar573 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar572 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg571 = (1'h0);
  reg [(4'h8):(1'h0)] reg570 = (1'h0);
  reg [(2'h3):(1'h0)] reg569 = (1'h0);
  reg [(4'hc):(1'h0)] reg568 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar567 = (1'h0);
  reg [(3'h4):(1'h0)] reg563 = (1'h0);
  reg [(4'he):(1'h0)] reg562 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar558 = (1'h0);
  reg [(4'hd):(1'h0)] forvar556 = (1'h0);
  reg [(2'h3):(1'h0)] forvar555 = (1'h0);
  reg [(4'hb):(1'h0)] forvar549 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg567 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg566 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg565 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg564 = (1'h0);
  reg [(4'h8):(1'h0)] forvar563 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar562 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg561 = (1'h0);
  reg [(3'h5):(1'h0)] reg560 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg559 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg558 = (1'h0);
  reg [(3'h7):(1'h0)] forvar554 = (1'h0);
  reg [(4'ha):(1'h0)] forvar552 = (1'h0);
  reg [(2'h3):(1'h0)] reg544 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg543 = (1'h0);
  reg [(4'hb):(1'h0)] reg542 = (1'h0);
  reg [(4'hd):(1'h0)] forvar541 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar508 = (1'h0);
  reg [(3'h7):(1'h0)] reg538 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar537 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar529 = (1'h0);
  reg [(2'h3):(1'h0)] forvar527 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg525 = (1'h0);
  reg [(3'h5):(1'h0)] forvar524 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar523 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg522 = (1'h0);
  reg [(3'h4):(1'h0)] reg520 = (1'h0);
  reg [(2'h2):(1'h0)] reg517 = (1'h0);
  reg [(3'h7):(1'h0)] forvar514 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar512 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg509 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg557 = (1'h0);
  reg [(5'h10):(1'h0)] reg556 = (1'h0);
  reg [(2'h2):(1'h0)] reg555 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg554 = (1'h0);
  reg [(5'h10):(1'h0)] reg553 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg552 = (1'h0);
  reg [(4'ha):(1'h0)] reg551 = (1'h0);
  reg signed [(4'he):(1'h0)] reg550 = (1'h0);
  reg [(4'he):(1'h0)] reg549 = (1'h0);
  reg [(5'h10):(1'h0)] reg548 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg547 = (1'h0);
  reg [(4'hd):(1'h0)] reg546 = (1'h0);
  reg [(3'h5):(1'h0)] reg545 = (1'h0);
  reg [(5'h10):(1'h0)] forvar544 = (1'h0);
  reg [(2'h2):(1'h0)] forvar543 = (1'h0);
  reg [(2'h2):(1'h0)] forvar542 = (1'h0);
  reg [(4'hb):(1'h0)] reg541 = (1'h0);
  reg [(2'h2):(1'h0)] reg540 = (1'h0);
  reg [(3'h5):(1'h0)] reg539 = (1'h0);
  reg [(5'h10):(1'h0)] forvar538 = (1'h0);
  reg [(2'h2):(1'h0)] reg534 = (1'h0);
  reg [(4'hc):(1'h0)] reg537 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar536 = (1'h0);
  reg [(4'hd):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar534 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar533 = (1'h0);
  reg [(4'h9):(1'h0)] reg532 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg531 = (1'h0);
  reg [(3'h5):(1'h0)] reg530 = (1'h0);
  reg [(3'h6):(1'h0)] reg529 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg528 = (1'h0);
  reg [(4'hb):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg526 = (1'h0);
  reg [(4'h9):(1'h0)] forvar525 = (1'h0);
  reg [(2'h3):(1'h0)] reg524 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg523 = (1'h0);
  reg [(5'h10):(1'h0)] forvar522 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg521 = (1'h0);
  reg [(3'h5):(1'h0)] forvar520 = (1'h0);
  reg [(4'hc):(1'h0)] reg511 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg519 = (1'h0);
  reg [(3'h5):(1'h0)] reg518 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar517 = (1'h0);
  reg [(3'h5):(1'h0)] reg516 = (1'h0);
  reg [(4'h9):(1'h0)] reg515 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg514 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg513 = (1'h0);
  reg [(4'h9):(1'h0)] reg512 = (1'h0);
  reg [(5'h10):(1'h0)] forvar511 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg510 = (1'h0);
  reg [(5'h10):(1'h0)] forvar509 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg508 = (1'h0);
  reg [(4'hd):(1'h0)] reg507 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar489 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar481 = (1'h0);
  reg [(2'h2):(1'h0)] reg479 = (1'h0);
  reg [(3'h4):(1'h0)] forvar473 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar471 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg506 = (1'h0);
  reg [(3'h7):(1'h0)] reg505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg504 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar503 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg502 = (1'h0);
  reg [(4'hb):(1'h0)] forvar501 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg493 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar492 = (1'h0);
  reg signed [(4'he):(1'h0)] reg500 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg499 = (1'h0);
  reg [(2'h2):(1'h0)] reg498 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg497 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg496 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg495 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg494 = (1'h0);
  reg [(4'hd):(1'h0)] forvar493 = (1'h0);
  reg [(4'ha):(1'h0)] reg491 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar470 = (1'h0);
  reg [(3'h4):(1'h0)] forvar467 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar485 = (1'h0);
  reg [(4'hd):(1'h0)] reg484 = (1'h0);
  reg [(4'he):(1'h0)] forvar483 = (1'h0);
  reg [(3'h6):(1'h0)] forvar482 = (1'h0);
  reg [(3'h7):(1'h0)] reg480 = (1'h0);
  reg signed [(4'he):(1'h0)] reg477 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar468 = (1'h0);
  reg [(4'hd):(1'h0)] reg492 = (1'h0);
  reg [(4'he):(1'h0)] forvar491 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg490 = (1'h0);
  reg [(2'h3):(1'h0)] reg489 = (1'h0);
  reg [(3'h5):(1'h0)] reg488 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg487 = (1'h0);
  reg [(3'h5):(1'h0)] reg486 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg485 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar484 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg483 = (1'h0);
  reg signed [(4'he):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg481 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar480 = (1'h0);
  reg [(2'h2):(1'h0)] forvar479 = (1'h0);
  reg [(4'he):(1'h0)] forvar472 = (1'h0);
  reg [(5'h10):(1'h0)] forvar469 = (1'h0);
  reg [(3'h6):(1'h0)] reg478 = (1'h0);
  reg [(4'h9):(1'h0)] forvar477 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg476 = (1'h0);
  reg [(3'h7):(1'h0)] reg475 = (1'h0);
  reg [(4'hf):(1'h0)] reg474 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg473 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg472 = (1'h0);
  reg [(4'hd):(1'h0)] reg471 = (1'h0);
  reg [(4'h9):(1'h0)] reg470 = (1'h0);
  reg [(4'hd):(1'h0)] reg469 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg468 = (1'h0);
  reg [(3'h7):(1'h0)] reg467 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg466 = (1'h0);
  reg [(4'he):(1'h0)] reg465 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg464 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg463 = (1'h0);
  reg [(4'hc):(1'h0)] forvar462 = (1'h0);
  reg [(5'h10):(1'h0)] reg461 = (1'h0);
  reg [(4'hc):(1'h0)] forvar459 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg456 = (1'h0);
  reg [(3'h7):(1'h0)] reg460 = (1'h0);
  reg [(2'h2):(1'h0)] reg459 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg458 = (1'h0);
  reg [(4'hc):(1'h0)] reg457 = (1'h0);
  reg [(4'hf):(1'h0)] forvar456 = (1'h0);
  reg [(5'h10):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar454 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg445 = (1'h0);
  reg [(5'h10):(1'h0)] reg444 = (1'h0);
  reg [(4'hc):(1'h0)] forvar443 = (1'h0);
  reg [(3'h6):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar452 = (1'h0);
  reg [(4'hf):(1'h0)] reg451 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg450 = (1'h0);
  reg [(5'h10):(1'h0)] reg449 = (1'h0);
  reg [(4'ha):(1'h0)] reg448 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar447 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg446 = (1'h0);
  reg [(3'h4):(1'h0)] forvar445 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar444 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg443 = (1'h0);
  reg [(4'hd):(1'h0)] forvar442 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg441 = (1'h0);
  reg [(4'hf):(1'h0)] reg440 = (1'h0);
  reg [(3'h7):(1'h0)] reg439 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg438 = (1'h0);
  reg [(3'h5):(1'h0)] forvar437 = (1'h0);
  reg [(4'h8):(1'h0)] reg436 = (1'h0);
  reg [(4'ha):(1'h0)] reg435 = (1'h0);
  reg [(4'hb):(1'h0)] reg434 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar433 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg432 = (1'h0);
  reg [(2'h2):(1'h0)] forvar430 = (1'h0);
  reg [(4'h9):(1'h0)] forvar421 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg419 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg414 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg413 = (1'h0);
  reg [(4'hf):(1'h0)] reg431 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg430 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg429 = (1'h0);
  reg [(4'hf):(1'h0)] reg428 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar427 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg424 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg422 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg427 = (1'h0);
  reg [(4'hf):(1'h0)] reg426 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg425 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar424 = (1'h0);
  reg [(4'h9):(1'h0)] reg423 = (1'h0);
  reg [(3'h6):(1'h0)] forvar422 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg421 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg420 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar419 = (1'h0);
  reg [(4'hb):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg417 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg416 = (1'h0);
  reg [(4'hb):(1'h0)] reg415 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar414 = (1'h0);
  reg [(5'h10):(1'h0)] forvar413 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar404 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg403 = (1'h0);
  reg [(4'hc):(1'h0)] reg407 = (1'h0);
  reg [(3'h5):(1'h0)] reg406 = (1'h0);
  reg [(4'h8):(1'h0)] forvar405 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar399 = (1'h0);
  reg [(4'hb):(1'h0)] forvar391 = (1'h0);
  reg [(4'h9):(1'h0)] reg396 = (1'h0);
  reg [(2'h3):(1'h0)] forvar379 = (1'h0);
  reg [(3'h6):(1'h0)] reg386 = (1'h0);
  reg [(2'h2):(1'h0)] reg385 = (1'h0);
  reg [(3'h5):(1'h0)] forvar382 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg381 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar378 = (1'h0);
  reg signed [(4'he):(1'h0)] reg376 = (1'h0);
  reg [(4'h8):(1'h0)] reg412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg411 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg410 = (1'h0);
  reg [(4'hf):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg408 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar407 = (1'h0);
  reg [(4'he):(1'h0)] forvar406 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg405 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg404 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar403 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg402 = (1'h0);
  reg [(5'h10):(1'h0)] reg401 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar400 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg399 = (1'h0);
  reg [(3'h4):(1'h0)] reg398 = (1'h0);
  reg [(3'h7):(1'h0)] forvar397 = (1'h0);
  reg [(2'h2):(1'h0)] forvar396 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg395 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg394 = (1'h0);
  reg [(4'hf):(1'h0)] reg393 = (1'h0);
  reg [(5'h10):(1'h0)] reg392 = (1'h0);
  reg [(3'h6):(1'h0)] reg391 = (1'h0);
  reg [(3'h7):(1'h0)] reg390 = (1'h0);
  reg [(2'h3):(1'h0)] reg389 = (1'h0);
  reg [(3'h4):(1'h0)] reg388 = (1'h0);
  reg [(4'hf):(1'h0)] reg387 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar386 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar385 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg383 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg382 = (1'h0);
  reg [(5'h10):(1'h0)] forvar381 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg379 = (1'h0);
  reg [(3'h6):(1'h0)] reg378 = (1'h0);
  reg [(5'h10):(1'h0)] forvar377 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar376 = (1'h0);
  reg [(3'h4):(1'h0)] reg375 = (1'h0);
  reg [(4'h9):(1'h0)] reg374 = (1'h0);
  reg [(4'he):(1'h0)] forvar373 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg372 = (1'h0);
  reg [(4'hc):(1'h0)] reg371 = (1'h0);
  reg [(4'he):(1'h0)] reg370 = (1'h0);
  reg [(4'h8):(1'h0)] forvar369 = (1'h0);
  reg [(5'h10):(1'h0)] reg368 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg367 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg366 = (1'h0);
  reg [(4'h8):(1'h0)] forvar365 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar364 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar363 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg362 = (1'h0);
  reg [(5'h10):(1'h0)] reg361 = (1'h0);
  reg [(4'hc):(1'h0)] reg360 = (1'h0);
  reg [(4'hc):(1'h0)] forvar359 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg358 = (1'h0);
  reg [(4'hf):(1'h0)] reg357 = (1'h0);
  reg [(3'h4):(1'h0)] forvar353 = (1'h0);
  reg [(4'he):(1'h0)] reg352 = (1'h0);
  reg [(3'h5):(1'h0)] forvar351 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg347 = (1'h0);
  reg [(4'hc):(1'h0)] reg356 = (1'h0);
  reg [(4'hd):(1'h0)] reg355 = (1'h0);
  reg [(3'h5):(1'h0)] reg354 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg353 = (1'h0);
  reg [(4'he):(1'h0)] forvar352 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg351 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg350 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg348 = (1'h0);
  reg [(4'hd):(1'h0)] forvar347 = (1'h0);
  reg [(4'he):(1'h0)] reg346 = (1'h0);
  reg [(4'hc):(1'h0)] reg344 = (1'h0);
  reg [(4'ha):(1'h0)] forvar342 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg341 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg345 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar344 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg342 = (1'h0);
  reg [(4'hf):(1'h0)] forvar341 = (1'h0);
  reg [(2'h2):(1'h0)] reg340 = (1'h0);
  reg [(4'h8):(1'h0)] reg339 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg338 = (1'h0);
  reg [(3'h6):(1'h0)] forvar337 = (1'h0);
  reg [(3'h5):(1'h0)] forvar336 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg325 = (1'h0);
  reg [(3'h7):(1'h0)] reg335 = (1'h0);
  reg [(3'h7):(1'h0)] reg334 = (1'h0);
  reg signed [(4'he):(1'h0)] reg333 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg332 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg331 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar329 = (1'h0);
  reg [(3'h6):(1'h0)] reg328 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg326 = (1'h0);
  reg [(4'hb):(1'h0)] forvar325 = (1'h0);
  reg [(5'h10):(1'h0)] reg324 = (1'h0);
  reg [(4'hd):(1'h0)] reg323 = (1'h0);
  reg [(3'h7):(1'h0)] reg322 = (1'h0);
  reg [(2'h2):(1'h0)] reg321 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar320 = (1'h0);
  reg [(4'ha):(1'h0)] reg319 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg318 = (1'h0);
  reg [(2'h3):(1'h0)] reg317 = (1'h0);
  reg [(3'h6):(1'h0)] reg316 = (1'h0);
  reg [(3'h5):(1'h0)] forvar315 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg314 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar313 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg312 = (1'h0);
  reg [(4'he):(1'h0)] reg311 = (1'h0);
  reg [(3'h5):(1'h0)] reg310 = (1'h0);
  reg [(2'h3):(1'h0)] reg309 = (1'h0);
  reg [(2'h2):(1'h0)] forvar308 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar306 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg305 = (1'h0);
  reg [(3'h4):(1'h0)] reg304 = (1'h0);
  reg signed [(4'he):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg302 = (1'h0);
  reg [(4'h8):(1'h0)] reg301 = (1'h0);
  reg [(4'hf):(1'h0)] reg300 = (1'h0);
  reg [(2'h2):(1'h0)] reg299 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg298 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg297 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar296 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg296 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar295 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar294 = (1'h0);
  wire [(4'he):(1'h0)] wire293;
  assign y = {wire580,
                 wire579,
                 wire578,
                 wire577,
                 reg576,
                 reg575,
                 reg574,
                 forvar573,
                 forvar572,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 forvar567,
                 reg563,
                 reg562,
                 forvar558,
                 forvar556,
                 forvar555,
                 forvar549,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 forvar563,
                 forvar562,
                 reg561,
                 reg560,
                 reg559,
                 reg558,
                 forvar554,
                 forvar552,
                 reg544,
                 reg543,
                 reg542,
                 forvar541,
                 forvar508,
                 reg538,
                 forvar537,
                 forvar529,
                 forvar527,
                 reg525,
                 forvar524,
                 forvar523,
                 reg522,
                 reg520,
                 reg517,
                 forvar514,
                 forvar512,
                 reg509,
                 reg557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 forvar544,
                 forvar543,
                 forvar542,
                 reg541,
                 reg540,
                 reg539,
                 forvar538,
                 reg534,
                 reg537,
                 forvar536,
                 reg535,
                 forvar534,
                 forvar533,
                 reg532,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 forvar525,
                 reg524,
                 reg523,
                 forvar522,
                 reg521,
                 forvar520,
                 reg511,
                 reg519,
                 reg518,
                 forvar517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 forvar511,
                 reg510,
                 forvar509,
                 reg508,
                 reg507,
                 forvar489,
                 forvar481,
                 reg479,
                 forvar473,
                 forvar471,
                 reg506,
                 reg505,
                 reg504,
                 forvar503,
                 reg502,
                 forvar501,
                 reg493,
                 forvar492,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 forvar493,
                 reg491,
                 forvar470,
                 forvar467,
                 forvar485,
                 reg484,
                 forvar483,
                 forvar482,
                 reg480,
                 reg477,
                 forvar468,
                 reg492,
                 forvar491,
                 reg490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 forvar484,
                 reg483,
                 reg482,
                 reg481,
                 forvar480,
                 forvar479,
                 forvar472,
                 forvar469,
                 reg478,
                 forvar477,
                 reg476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 forvar462,
                 reg461,
                 forvar459,
                 reg456,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 forvar456,
                 reg455,
                 forvar454,
                 reg445,
                 reg444,
                 forvar443,
                 reg453,
                 forvar452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 forvar447,
                 reg446,
                 forvar445,
                 forvar444,
                 reg443,
                 forvar442,
                 reg441,
                 reg440,
                 reg439,
                 reg438,
                 forvar437,
                 reg436,
                 reg435,
                 reg434,
                 forvar433,
                 reg432,
                 forvar430,
                 forvar421,
                 reg419,
                 reg414,
                 reg413,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 forvar427,
                 reg424,
                 reg422,
                 reg427,
                 reg426,
                 reg425,
                 forvar424,
                 reg423,
                 forvar422,
                 reg421,
                 reg420,
                 forvar419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 forvar414,
                 forvar413,
                 forvar404,
                 reg403,
                 reg407,
                 reg406,
                 forvar405,
                 forvar399,
                 forvar391,
                 reg396,
                 forvar379,
                 reg386,
                 reg385,
                 forvar382,
                 reg381,
                 forvar378,
                 reg376,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 forvar407,
                 forvar406,
                 reg405,
                 reg404,
                 forvar403,
                 reg402,
                 reg401,
                 forvar400,
                 reg399,
                 reg398,
                 forvar397,
                 forvar396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 forvar386,
                 forvar385,
                 reg384,
                 reg383,
                 reg382,
                 forvar381,
                 reg380,
                 reg379,
                 reg378,
                 forvar377,
                 forvar376,
                 reg375,
                 reg374,
                 forvar373,
                 reg372,
                 reg371,
                 reg370,
                 forvar369,
                 reg368,
                 reg367,
                 reg366,
                 forvar365,
                 forvar364,
                 forvar363,
                 reg362,
                 reg361,
                 reg360,
                 forvar359,
                 reg358,
                 reg357,
                 forvar353,
                 reg352,
                 forvar351,
                 reg347,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 forvar352,
                 reg351,
                 reg350,
                 reg349,
                 reg348,
                 forvar347,
                 reg346,
                 reg344,
                 forvar342,
                 reg341,
                 reg345,
                 forvar344,
                 reg343,
                 reg342,
                 forvar341,
                 reg340,
                 reg339,
                 reg338,
                 forvar337,
                 forvar336,
                 reg325,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 reg330,
                 forvar329,
                 reg328,
                 reg327,
                 reg326,
                 forvar325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 forvar320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 forvar315,
                 reg314,
                 forvar313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 forvar308,
                 reg307,
                 forvar306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 forvar296,
                 reg296,
                 forvar295,
                 forvar294,
                 wire293,
                 (1'h0)};
  assign wire293 = {(((~&wire291) || (wire291 ?
                           wire289 : wire290)) | $signed((&(8'haa))))};
  always
    @(posedge clk) begin
      for (forvar294 = (1'h0); (forvar294 < (2'h2)); forvar294 = (forvar294 + (1'h1)))
        begin
          if ({(8'ha3)})
            begin
              if (({(~^(wire291 | forvar294))} || wire293))
                begin
                  for (forvar295 = (1'h0); (forvar295 < (1'h1)); forvar295 = (forvar295 + (1'h1)))
                    begin
                      reg296 <= (8'haa);
                    end
                end
              else
                begin
                  for (forvar295 = (1'h0); (forvar295 < (2'h2)); forvar295 = (forvar295 + (1'h1)))
                    begin
                      reg296 <= reg296;
                    end
                end
            end
          else
            begin
              for (forvar295 = (1'h0); (forvar295 < (1'h0)); forvar295 = (forvar295 + (1'h1)))
                begin
                  for (forvar296 = (1'h0); (forvar296 < (2'h2)); forvar296 = (forvar296 + (1'h1)))
                    begin
                      reg297 <= ($unsigned($signed(wire289)) ^~ {{((8'hac) <= (8'h9c))}});
                      reg298 <= $signed((-forvar294[(2'h2):(2'h2)]));
                    end
                  if (wire289[(1'h0):(1'h0)])
                    begin
                      reg299 <= reg298[(2'h3):(2'h3)];
                      reg300 <= $unsigned((reg297[(3'h4):(1'h1)] * ((reg296 <= forvar294) <= (8'ha2))));
                      reg301 <= $signed(reg298);
                    end
                  else
                    begin
                      reg299 <= (~^($unsigned($unsigned(forvar294)) << (reg296 ?
                          reg300 : forvar294[(4'h9):(3'h7)])));
                      reg300 <= ((!{$signed(wire288)}) ? (!reg299) : forvar296);
                      reg301 <= $signed($signed((^~reg297[(1'h1):(1'h0)])));
                    end
                end
              if (($signed($signed($unsigned(wire290))) ^~ wire288))
                begin
                  if (reg300)
                    begin
                      reg302 <= wire292;
                      reg303 <= {reg298};
                      reg304 <= (8'h9e);
                      reg305 <= forvar294;
                    end
                  else
                    begin
                      reg302 <= $signed(((|(^~wire290)) ?
                          $signed(forvar294) : ((~|reg305) ?
                              reg297[(1'h0):(1'h0)] : $signed(wire293))));
                    end
                  for (forvar306 = (1'h0); (forvar306 < (2'h3)); forvar306 = (forvar306 + (1'h1)))
                    begin
                      reg307 <= (($unsigned((^reg305)) ?
                          wire291[(2'h3):(2'h3)] : (&((8'ha2) > wire288))) >>> $unsigned($unsigned(reg303)));
                    end
                end
              else
                begin
                  if ($unsigned(($unsigned(wire288[(1'h1):(1'h1)]) >= (~^wire289[(3'h7):(3'h6)]))))
                    begin
                      reg302 <= reg301[(3'h7):(2'h3)];
                      reg303 <= $signed((^wire288[(3'h4):(2'h2)]));
                      reg304 <= (($signed((!(8'hb5))) - (8'ha3)) ?
                          {($signed(reg296) ?
                                  (8'hb4) : wire291)} : ({$signed((8'hac))} ?
                              reg301[(1'h1):(1'h0)] : ((reg300 ^~ forvar295) ?
                                  $unsigned(reg303) : forvar294)));
                    end
                  else
                    begin
                      reg302 <= {forvar294[(4'h9):(3'h7)]};
                      reg303 <= wire293[(4'he):(4'hc)];
                    end
                end
              for (forvar308 = (1'h0); (forvar308 < (2'h3)); forvar308 = (forvar308 + (1'h1)))
                begin
                  if (($signed((|$signed(reg298))) == (!($unsigned(wire293) ?
                      forvar295 : forvar296))))
                    begin
                      reg309 <= $unsigned(reg296[(4'hd):(1'h0)]);
                      reg310 <= {{(^{wire293})}};
                    end
                  else
                    begin
                      reg309 <= {((~&(^(8'haf))) <= forvar294[(1'h1):(1'h0)])};
                      reg310 <= ((forvar308[(1'h0):(1'h0)] || $unsigned($signed(wire288))) ^~ ($signed(reg298) || (+((8'had) ?
                          (8'hb8) : forvar308))));
                      reg311 <= $signed(({(~forvar296)} ~^ $signed(reg300[(4'hd):(1'h0)])));
                      reg312 <= $signed({$unsigned((+reg304))});
                    end
                  for (forvar313 = (1'h0); (forvar313 < (2'h3)); forvar313 = (forvar313 + (1'h1)))
                    begin
                      reg314 <= (^~reg297[(3'h6):(3'h4)]);
                    end
                  for (forvar315 = (1'h0); (forvar315 < (1'h0)); forvar315 = (forvar315 + (1'h1)))
                    begin
                      reg316 <= {reg296};
                      reg317 <= {$unsigned((8'ha5))};
                      reg318 <= $unsigned(wire289);
                      reg319 <= (~$unsigned($unsigned((~&wire289))));
                    end
                  for (forvar320 = (1'h0); (forvar320 < (2'h2)); forvar320 = (forvar320 + (1'h1)))
                    begin
                      reg321 <= $unsigned(($signed(reg303) ?
                          reg318 : $unsigned($unsigned(reg302))));
                      reg322 <= reg299;
                      reg323 <= $signed((($unsigned(forvar320) ?
                              {reg303} : $unsigned(reg299)) ?
                          reg302[(2'h3):(1'h0)] : reg321[(2'h2):(1'h1)]));
                      reg324 <= forvar315[(2'h3):(2'h3)];
                    end
                end
              if ((~|(((8'ha4) ?
                  reg314[(2'h3):(2'h3)] : $unsigned(forvar308)) + reg309[(1'h0):(1'h0)])))
                begin
                  for (forvar325 = (1'h0); (forvar325 < (1'h1)); forvar325 = (forvar325 + (1'h1)))
                    begin
                      reg326 <= (wire291 & {(8'ha0)});
                      reg327 <= reg299;
                      reg328 <= $signed(wire292[(4'h8):(2'h3)]);
                    end
                  for (forvar329 = (1'h0); (forvar329 < (2'h3)); forvar329 = (forvar329 + (1'h1)))
                    begin
                      reg330 <= $signed(reg304);
                      reg331 <= (8'hae);
                      reg332 <= forvar295;
                    end
                  if ((reg318 ^~ $unsigned($signed($unsigned((8'h9c))))))
                    begin
                      reg333 <= $signed(($unsigned(reg323[(3'h4):(1'h0)]) ?
                          $signed({(8'h9d)}) : reg305[(1'h0):(1'h0)]));
                      reg334 <= (|{$signed($unsigned((8'hae)))});
                      reg335 <= ($unsigned((~&wire291[(4'ha):(3'h6)])) ?
                          (((wire289 <<< wire290) ?
                              (wire293 ^~ forvar313) : {wire288}) * (~&reg314[(1'h1):(1'h0)])) : (^~$unsigned({reg322})));
                    end
                  else
                    begin
                      reg333 <= forvar325[(3'h5):(1'h0)];
                      reg334 <= (!$signed($unsigned($unsigned(reg333))));
                      reg335 <= forvar296[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  if (((((!reg334) ?
                      forvar306[(3'h4):(3'h4)] : (reg327 ~^ reg309)) ^ forvar320[(1'h1):(1'h1)]) + $signed((~&$unsigned(forvar320)))))
                    begin
                      reg325 <= $unsigned(reg301[(3'h5):(1'h1)]);
                      reg326 <= reg334[(3'h7):(3'h4)];
                      reg327 <= ((8'hae) > reg333);
                      reg328 <= $signed((+forvar295[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg325 <= forvar308;
                      reg326 <= $signed(reg298);
                    end
                  for (forvar329 = (1'h0); (forvar329 < (1'h0)); forvar329 = (forvar329 + (1'h1)))
                    begin
                      reg330 <= reg317;
                    end
                end
            end
          for (forvar336 = (1'h0); (forvar336 < (1'h0)); forvar336 = (forvar336 + (1'h1)))
            begin
              if (((({reg301} ?
                  forvar306 : $signed(wire292)) >= $unsigned(reg334[(1'h0):(1'h0)])) >>> reg305[(1'h0):(1'h0)]))
                begin
                  for (forvar337 = (1'h0); (forvar337 < (1'h1)); forvar337 = (forvar337 + (1'h1)))
                    begin
                      reg338 <= (&(&{(~&reg316)}));
                      reg339 <= wire288[(4'h8):(3'h5)];
                      reg340 <= reg338;
                    end
                  for (forvar341 = (1'h0); (forvar341 < (1'h1)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= (&(((reg318 * forvar306) ?
                              (8'ha0) : (~|reg317)) ?
                          $unsigned(wire290[(2'h2):(2'h2)]) : $signed(reg316[(1'h0):(1'h0)])));
                    end
                  reg343 <= (-((+(~reg298)) ? {(~^reg331)} : {reg342}));
                  for (forvar344 = (1'h0); (forvar344 < (2'h2)); forvar344 = (forvar344 + (1'h1)))
                    begin
                      reg345 <= {(((reg309 ?
                              reg309 : reg326) - reg332) ^~ $unsigned((wire288 && forvar306)))};
                    end
                end
              else
                begin
                  for (forvar337 = (1'h0); (forvar337 < (1'h1)); forvar337 = (forvar337 + (1'h1)))
                    begin
                      reg338 <= (&forvar341[(4'hc):(4'h9)]);
                      reg339 <= (reg319[(1'h0):(1'h0)] - reg297);
                      reg340 <= (&$signed(({reg303} ?
                          (forvar306 < forvar313) : $unsigned(reg302))));
                      reg341 <= (~&(-((~wire293) ?
                          (reg345 <= forvar294) : $signed(forvar308))));
                    end
                  for (forvar342 = (1'h0); (forvar342 < (1'h0)); forvar342 = (forvar342 + (1'h1)))
                    begin
                      reg343 <= (^(^~$unsigned((reg303 ? forvar294 : reg342))));
                    end
                  if ($unsigned(reg312))
                    begin
                      reg344 <= (~$signed(((&reg338) ?
                          $unsigned(reg317) : reg343[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg344 <= wire291;
                      reg345 <= $unsigned($unsigned((~^(8'hb1))));
                      reg346 <= (^$unsigned((&$signed(forvar329))));
                    end
                end
            end
          if ($signed(wire292))
            begin
              for (forvar347 = (1'h0); (forvar347 < (1'h0)); forvar347 = (forvar347 + (1'h1)))
                begin
                  if (reg296[(4'h8):(3'h6)])
                    begin
                      reg348 <= $unsigned(forvar336);
                      reg349 <= (~(+$signed(reg297)));
                      reg350 <= ($unsigned(reg307[(3'h7):(1'h1)]) ?
                          (^reg338[(2'h3):(1'h0)]) : reg314[(2'h3):(1'h0)]);
                      reg351 <= ($unsigned(wire288) - reg311[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg348 <= forvar294;
                    end
                  for (forvar352 = (1'h0); (forvar352 < (2'h2)); forvar352 = (forvar352 + (1'h1)))
                    begin
                      reg353 <= $signed(reg332);
                      reg354 <= (^reg331);
                      reg355 <= reg339;
                    end
                  reg356 <= reg297[(2'h3):(2'h3)];
                end
            end
          else
            begin
              if ({(&(~^(!reg318)))})
                begin
                  if (($unsigned((8'h9f)) ?
                      ($signed($signed(reg316)) ^ $unsigned(((8'h9e) ?
                          reg299 : reg334))) : reg298[(4'h9):(3'h6)]))
                    begin
                      reg347 <= $unsigned((!wire293[(3'h5):(3'h4)]));
                      reg348 <= (~({{(8'had)}} <<< ($signed(forvar336) ^ (reg304 ?
                          (8'ha4) : (8'h9f)))));
                      reg349 <= reg335;
                      reg350 <= ($unsigned(reg335[(1'h0):(1'h0)]) >= (^{forvar308[(1'h0):(1'h0)]}));
                    end
                  else
                    begin
                      reg347 <= (|(reg347 ?
                          ((reg318 >> reg345) > ((8'ha3) ?
                              forvar320 : (8'ha8))) : ($unsigned(reg307) & reg319)));
                      reg348 <= (((((8'hae) >>> forvar341) <<< {reg345}) ?
                              $unsigned((^reg338)) : ($signed(forvar337) != $signed(reg333))) ?
                          reg347 : $signed($signed((+forvar315))));
                      reg349 <= (forvar313 ?
                          ((forvar341 ?
                              (-reg351) : forvar320) >> $signed(reg348)) : (&$unsigned(((8'hb0) ?
                              wire292 : forvar306))));
                      reg350 <= (^((&$signed(reg312)) ^ $signed({reg356})));
                    end
                  for (forvar351 = (1'h0); (forvar351 < (2'h3)); forvar351 = (forvar351 + (1'h1)))
                    begin
                      reg352 <= reg332;
                    end
                  for (forvar353 = (1'h0); (forvar353 < (2'h2)); forvar353 = (forvar353 + (1'h1)))
                    begin
                      reg354 <= $unsigned($signed((&(forvar313 ~^ reg316))));
                    end
                  if (($unsigned(forvar353) ?
                      {(~&(forvar352 ? reg330 : forvar353))} : reg332))
                    begin
                      reg355 <= (~&(((forvar329 ? (8'hac) : reg332) ?
                          ((8'ha4) && forvar315) : $unsigned(reg349)) >> $unsigned(reg327[(4'he):(4'he)])));
                    end
                  else
                    begin
                      reg355 <= reg311[(1'h0):(1'h0)];
                      reg356 <= $unsigned(reg335);
                      reg357 <= ((^~wire293) ?
                          (reg326[(3'h6):(1'h0)] ?
                              reg309[(2'h2):(1'h1)] : ((&reg319) ?
                                  {(8'ha1)} : reg355[(3'h7):(3'h4)])) : reg317);
                      reg358 <= (~{$unsigned($signed(reg335))});
                    end
                end
              else
                begin
                  reg347 <= (((reg334[(3'h6):(3'h4)] ~^ (reg302 - reg310)) ?
                          ($unsigned(reg300) ^~ (reg324 ?
                              reg353 : reg299)) : $signed((&reg342))) ?
                      $signed($signed($unsigned(reg353))) : (forvar336[(2'h3):(2'h2)] ?
                          $signed((reg350 ?
                              reg317 : reg346)) : reg333[(1'h1):(1'h0)]));
                  reg348 <= $unsigned(forvar342[(2'h3):(2'h2)]);
                end
              for (forvar359 = (1'h0); (forvar359 < (2'h3)); forvar359 = (forvar359 + (1'h1)))
                begin
                  if ($unsigned($signed(forvar295)))
                    begin
                      reg360 <= (~|$unsigned(reg340[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg360 <= $signed(reg325[(3'h4):(1'h0)]);
                      reg361 <= (~|$unsigned(forvar329));
                      reg362 <= (|({(&reg309)} ?
                          ((reg335 >>> wire288) ?
                              $unsigned(forvar342) : $signed(reg305)) : $unsigned((reg300 ?
                              (8'h9d) : wire290))));
                    end
                end
            end
          for (forvar363 = (1'h0); (forvar363 < (2'h2)); forvar363 = (forvar363 + (1'h1)))
            begin
              for (forvar364 = (1'h0); (forvar364 < (1'h0)); forvar364 = (forvar364 + (1'h1)))
                begin
                  for (forvar365 = (1'h0); (forvar365 < (1'h1)); forvar365 = (forvar365 + (1'h1)))
                    begin
                      reg366 <= ($unsigned((~(forvar352 <<< wire292))) >>> ((reg311 ?
                              (^~reg303) : (reg327 ^~ reg330)) ?
                          (reg342[(4'he):(3'h7)] ?
                              {reg301} : (reg348 ?
                                  forvar359 : forvar329)) : {(reg354 < reg362)}));
                      reg367 <= (((8'hb9) ?
                          $signed((forvar329 ?
                              (8'had) : reg327)) : (reg296[(4'he):(3'h5)] ?
                              reg333 : $unsigned(reg352))) == $signed(reg331));
                      reg368 <= $unsigned(reg299);
                    end
                  for (forvar369 = (1'h0); (forvar369 < (1'h1)); forvar369 = (forvar369 + (1'h1)))
                    begin
                      reg370 <= (8'ha8);
                      reg371 <= (!forvar341);
                    end
                  reg372 <= $signed({$unsigned((forvar296 >>> reg355))});
                  for (forvar373 = (1'h0); (forvar373 < (2'h3)); forvar373 = (forvar373 + (1'h1)))
                    begin
                      reg374 <= {forvar336[(3'h4):(2'h3)]};
                      reg375 <= reg344;
                    end
                end
            end
        end
      if (reg338)
        begin
          for (forvar376 = (1'h0); (forvar376 < (2'h3)); forvar376 = (forvar376 + (1'h1)))
            begin
              for (forvar377 = (1'h0); (forvar377 < (2'h3)); forvar377 = (forvar377 + (1'h1)))
                begin
                  if (reg302)
                    begin
                      reg378 <= (^((8'hb6) ?
                          reg367[(2'h2):(2'h2)] : $signed(reg305[(3'h6):(3'h5)])));
                      reg379 <= (&$signed(({reg319} - {reg346})));
                      reg380 <= (&(+$unsigned($signed(reg345))));
                    end
                  else
                    begin
                      reg378 <= forvar320[(1'h1):(1'h0)];
                    end
                  for (forvar381 = (1'h0); (forvar381 < (2'h3)); forvar381 = (forvar381 + (1'h1)))
                    begin
                      reg382 <= reg357[(2'h3):(2'h3)];
                      reg383 <= ((^~(~(reg361 ?
                          (8'hb2) : forvar377))) ^ $unsigned($unsigned(((8'hab) <<< reg316))));
                      reg384 <= (({(reg378 ?
                                  (8'hb2) : reg330)} >= (~^(forvar364 ?
                              forvar381 : reg338))) ?
                          wire288 : ($signed($unsigned(reg333)) > $unsigned($unsigned(forvar359))));
                    end
                end
              for (forvar385 = (1'h0); (forvar385 < (2'h2)); forvar385 = (forvar385 + (1'h1)))
                begin
                  for (forvar386 = (1'h0); (forvar386 < (2'h2)); forvar386 = (forvar386 + (1'h1)))
                    begin
                      reg387 <= $signed($signed(reg355[(2'h3):(2'h2)]));
                      reg388 <= (&(($signed((8'hb8)) ^ $signed(forvar351)) ?
                          reg312 : {reg346}));
                    end
                  if (((-{reg382}) ?
                      forvar325[(2'h3):(1'h0)] : {((reg346 >= reg298) ?
                              (reg322 ?
                                  (8'h9f) : reg319) : (reg316 >> (8'ha1)))}))
                    begin
                      reg389 <= forvar295;
                      reg390 <= reg356[(4'hb):(3'h7)];
                      reg391 <= ($unsigned($signed($unsigned(reg312))) ?
                          $unsigned(($signed((8'h9c)) ?
                              (~|reg298) : $signed(reg300))) : $unsigned(($signed(reg319) | $unsigned(forvar336))));
                      reg392 <= (reg314[(4'h8):(3'h7)] ?
                          (-($unsigned(forvar385) ?
                              (reg383 >> (8'hb8)) : (reg378 ?
                                  forvar363 : reg311))) : {{forvar329}});
                    end
                  else
                    begin
                      reg389 <= (((^~$unsigned(reg352)) ?
                              wire293 : $signed((forvar351 ?
                                  forvar353 : reg351))) ?
                          forvar313 : reg304[(2'h2):(1'h1)]);
                      reg390 <= ((-forvar341[(4'hc):(4'h8)]) >>> $signed(wire293[(1'h1):(1'h0)]));
                      reg391 <= {$unsigned($signed($signed(reg340)))};
                      reg392 <= wire293;
                    end
                  reg393 <= $unsigned(reg298[(4'h8):(3'h4)]);
                  if (($unsigned(((|reg296) == $signed((8'hb6)))) >> {reg296[(4'h8):(3'h6)]}))
                    begin
                      reg394 <= ((~^((!reg302) ^ (reg378 ? reg296 : reg353))) ?
                          wire289[(3'h6):(1'h1)] : reg390);
                    end
                  else
                    begin
                      reg394 <= ($signed(reg335) ?
                          (~&reg299) : reg345[(1'h0):(1'h0)]);
                      reg395 <= ($unsigned($signed((reg319 >>> reg333))) ?
                          forvar341 : (|((reg345 ?
                              forvar295 : reg322) ^ $signed(reg380))));
                    end
                end
            end
          for (forvar396 = (1'h0); (forvar396 < (2'h3)); forvar396 = (forvar396 + (1'h1)))
            begin
              for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
                begin
                  if ($unsigned(($unsigned(reg316) != $unsigned(forvar315))))
                    begin
                      reg398 <= (~&reg303);
                    end
                  else
                    begin
                      reg398 <= $signed(forvar385[(3'h5):(1'h1)]);
                      reg399 <= reg310[(3'h5):(3'h5)];
                    end
                  for (forvar400 = (1'h0); (forvar400 < (1'h0)); forvar400 = (forvar400 + (1'h1)))
                    begin
                      reg401 <= reg398;
                      reg402 <= $unsigned($unsigned(((wire290 != reg338) ?
                          reg345 : (forvar308 >>> (8'hb6)))));
                    end
                  for (forvar403 = (1'h0); (forvar403 < (1'h0)); forvar403 = (forvar403 + (1'h1)))
                    begin
                      reg404 <= (^~(~&$signed(((8'hb9) ? reg333 : forvar315))));
                      reg405 <= ($unsigned((~reg305)) <<< ((&{reg303}) ?
                          ($unsigned(reg309) >> ((8'h9e) ?
                              reg297 : (8'had))) : $signed({reg352})));
                    end
                end
              for (forvar406 = (1'h0); (forvar406 < (1'h1)); forvar406 = (forvar406 + (1'h1)))
                begin
                  for (forvar407 = (1'h0); (forvar407 < (2'h3)); forvar407 = (forvar407 + (1'h1)))
                    begin
                      reg408 <= $signed({(reg328[(2'h3):(2'h2)] <= reg345)});
                      reg409 <= $unsigned((~&(reg332[(3'h6):(3'h5)] < {reg389})));
                      reg410 <= reg354;
                      reg411 <= {(reg340 <= (!(^~reg331)))};
                    end
                end
            end
          reg412 <= reg374[(2'h2):(1'h0)];
        end
      else
        begin
          reg376 <= reg357;
          for (forvar377 = (1'h0); (forvar377 < (2'h2)); forvar377 = (forvar377 + (1'h1)))
            begin
              if ((~($signed((-reg323)) ?
                  {(8'ha3)} : $unsigned($unsigned(reg384)))))
                begin
                  for (forvar378 = (1'h0); (forvar378 < (2'h2)); forvar378 = (forvar378 + (1'h1)))
                    begin
                      reg379 <= $unsigned(((!(reg353 ? reg409 : reg347)) ?
                          $signed($signed(reg298)) : (!reg372)));
                      reg380 <= ($unsigned(((reg314 > forvar364) >= forvar353[(3'h4):(3'h4)])) >> (8'hb7));
                      reg381 <= $unsigned($signed($unsigned((reg362 ?
                          reg383 : reg335))));
                    end
                  for (forvar382 = (1'h0); (forvar382 < (2'h2)); forvar382 = (forvar382 + (1'h1)))
                    begin
                      reg383 <= (~^$signed((|forvar400[(3'h6):(3'h6)])));
                      reg384 <= reg402[(2'h3):(2'h2)];
                      reg385 <= (((~(^~(8'ha0))) ?
                          reg366[(3'h5):(1'h0)] : (forvar377[(2'h3):(1'h0)] < $unsigned(reg350))) - (reg384[(3'h5):(1'h0)] ?
                          forvar382 : reg317[(2'h3):(1'h0)]));
                    end
                  reg386 <= $unsigned((forvar377 && (+(forvar378 ?
                      reg303 : reg303))));
                  if ((~($signed($unsigned(forvar381)) ?
                      (reg338 < {wire290}) : wire290)))
                    begin
                      reg387 <= ((reg332[(3'h5):(3'h5)] ?
                          reg379 : reg376[(4'h9):(4'h8)]) ~^ ((^~$signed(forvar315)) ?
                          $signed($unsigned(forvar397)) : (~&(~&forvar347))));
                      reg388 <= (8'hb6);
                      reg389 <= (^~$unsigned($signed(reg330)));
                      reg390 <= reg316[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg387 <= $unsigned(($unsigned((~|reg345)) ?
                          ($unsigned(forvar386) >> $signed(reg304)) : $signed($signed(wire293))));
                      reg388 <= $signed($unsigned((|$signed(reg389))));
                      reg389 <= ($unsigned($unsigned(((8'ha5) || (8'ha9)))) < $unsigned(((reg374 >>> reg394) ?
                          reg343 : (reg311 - forvar342))));
                    end
                end
              else
                begin
                  reg378 <= $signed({$unsigned(((8'ha1) | wire292))});
                  for (forvar379 = (1'h0); (forvar379 < (1'h1)); forvar379 = (forvar379 + (1'h1)))
                    begin
                      reg380 <= ($signed(reg372[(1'h1):(1'h1)]) ?
                          {reg404} : reg361[(4'h8):(4'h8)]);
                      reg381 <= (|forvar351[(1'h0):(1'h0)]);
                    end
                  if ($signed((~|{$unsigned(forvar406)})))
                    begin
                      reg382 <= reg353[(1'h1):(1'h1)];
                      reg383 <= $signed(reg331[(3'h5):(3'h5)]);
                      reg384 <= (~|$signed(((reg411 | reg309) ~^ reg327)));
                      reg385 <= (!reg409);
                    end
                  else
                    begin
                      reg382 <= {forvar306};
                      reg383 <= reg409;
                      reg384 <= reg296;
                    end
                  if (((reg311 ?
                          ((reg375 ? forvar344 : forvar369) ?
                              (reg348 == forvar342) : forvar344) : ((reg310 < reg370) ?
                              ((8'ha4) ?
                                  reg307 : forvar359) : $unsigned(forvar385))) ?
                      ((~&reg383) ?
                          forvar353 : reg327) : ($unsigned($signed(reg382)) ?
                          reg412[(1'h1):(1'h1)] : ($unsigned(forvar351) ?
                              reg402 : $unsigned(forvar353)))))
                    begin
                      reg386 <= $signed($unsigned((&reg348[(2'h3):(1'h1)])));
                      reg387 <= ((!(reg331 != $signed(reg322))) ~^ reg393[(4'hf):(4'hd)]);
                    end
                  else
                    begin
                      reg386 <= ((((~|reg304) ?
                              (forvar386 ~^ forvar369) : $unsigned(reg410)) >> (^~$signed(reg372))) ?
                          reg372[(2'h2):(1'h0)] : (reg357 >> $unsigned((wire289 >= reg350))));
                    end
                end
              if ($unsigned(reg301[(3'h6):(1'h0)]))
                begin
                  if ({reg344[(4'h9):(3'h5)]})
                    begin
                      reg391 <= (+(reg404 ?
                          {(forvar381 || forvar400)} : $signed($signed(forvar397))));
                      reg392 <= reg360;
                      reg393 <= ($signed(forvar325[(3'h6):(3'h5)]) ?
                          $unsigned($unsigned($unsigned(forvar373))) : $unsigned(forvar381));
                    end
                  else
                    begin
                      reg391 <= $signed(reg370[(4'hb):(3'h5)]);
                    end
                  if (reg334[(3'h7):(1'h0)])
                    begin
                      reg394 <= ($unsigned((~^(reg332 || (8'haa)))) <<< reg372);
                    end
                  else
                    begin
                      reg394 <= $unsigned({reg331});
                      reg395 <= $signed(forvar306);
                      reg396 <= reg393[(3'h7):(2'h2)];
                    end
                  for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
                    begin
                      reg398 <= reg386;
                    end
                end
              else
                begin
                  for (forvar391 = (1'h0); (forvar391 < (2'h3)); forvar391 = (forvar391 + (1'h1)))
                    begin
                      reg392 <= (^~reg311[(2'h3):(2'h3)]);
                      reg393 <= reg374[(3'h6):(1'h0)];
                    end
                end
              for (forvar399 = (1'h0); (forvar399 < (1'h1)); forvar399 = (forvar399 + (1'h1)))
                begin
                  for (forvar400 = (1'h0); (forvar400 < (1'h0)); forvar400 = (forvar400 + (1'h1)))
                    begin
                      reg401 <= reg317;
                      reg402 <= reg370;
                    end
                end
              if (((8'ha3) < $unsigned(reg348[(2'h3):(1'h1)])))
                begin
                  for (forvar403 = (1'h0); (forvar403 < (2'h3)); forvar403 = (forvar403 + (1'h1)))
                    begin
                      reg404 <= $signed($signed(forvar377[(3'h7):(3'h4)]));
                    end
                  for (forvar405 = (1'h0); (forvar405 < (1'h1)); forvar405 = (forvar405 + (1'h1)))
                    begin
                      reg406 <= $signed(reg358);
                      reg407 <= ((((reg401 ?
                                  forvar308 : forvar306) | $signed(reg395)) ?
                              forvar353 : (|$unsigned(forvar396))) ?
                          ((~^(reg392 ?
                              (8'h9f) : forvar369)) != forvar342) : (8'hb1));
                      reg408 <= $signed((8'hb6));
                    end
                end
              else
                begin
                  reg403 <= wire290;
                  for (forvar404 = (1'h0); (forvar404 < (2'h2)); forvar404 = (forvar404 + (1'h1)))
                    begin
                      reg405 <= (8'h9f);
                      reg406 <= reg296;
                      reg407 <= forvar376[(1'h0):(1'h0)];
                      reg408 <= $signed($unsigned(forvar369));
                    end
                  if (reg325[(2'h2):(1'h0)])
                    begin
                      reg409 <= ({((+(8'haf)) ?
                                  reg376[(4'ha):(3'h5)] : $signed(reg374))} ?
                          (^~((reg395 ?
                              (8'haa) : reg405) ~^ (reg381 <= forvar325))) : {(~&(forvar315 != reg346))});
                    end
                  else
                    begin
                      reg409 <= ((forvar295 ?
                          reg332 : (~^reg297[(2'h2):(2'h2)])) && (-(forvar406[(2'h2):(2'h2)] ?
                          wire289[(3'h5):(2'h2)] : (forvar405 ~^ reg410))));
                      reg410 <= (($signed($unsigned(reg347)) ?
                              forvar378[(2'h3):(2'h2)] : reg392) ?
                          (forvar308 >>> ($unsigned(forvar377) | reg357)) : ({(~(8'hab))} <= {forvar336}));
                      reg411 <= (reg387[(4'hc):(4'hc)] ?
                          {{reg390}} : ($unsigned(reg378[(1'h0):(1'h0)]) ?
                              (8'hb5) : $unsigned(forvar365)));
                    end
                  reg412 <= (forvar306 ?
                      ($unsigned($signed(wire288)) >= reg389[(1'h0):(1'h0)]) : (($unsigned(forvar377) ?
                              {reg325} : $signed(reg333)) ?
                          wire291 : ((8'ha7) >> $unsigned(reg326))));
                end
            end
          if ($unsigned(($unsigned((forvar376 ? reg393 : reg297)) ?
              ($unsigned(reg386) ? {forvar397} : reg299) : ($unsigned((8'hb0)) ?
                  $unsigned(reg351) : reg399))))
            begin
              for (forvar413 = (1'h0); (forvar413 < (1'h0)); forvar413 = (forvar413 + (1'h1)))
                begin
                  for (forvar414 = (1'h0); (forvar414 < (1'h1)); forvar414 = (forvar414 + (1'h1)))
                    begin
                      reg415 <= reg368[(4'h8):(1'h0)];
                      reg416 <= reg356;
                    end
                  reg417 <= (-((&forvar399) ~^ $signed((&(8'hb8)))));
                  if ($unsigned((wire289[(3'h6):(3'h5)] <<< reg378)))
                    begin
                      reg418 <= reg354[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg418 <= forvar381[(3'h7):(2'h2)];
                    end
                end
              if (reg406)
                begin
                  for (forvar419 = (1'h0); (forvar419 < (1'h1)); forvar419 = (forvar419 + (1'h1)))
                    begin
                      reg420 <= (&$signed((^reg367[(2'h3):(1'h1)])));
                      reg421 <= $signed({((&(8'hb5)) ?
                              (+reg330) : $signed((8'haa)))});
                    end
                  for (forvar422 = (1'h0); (forvar422 < (1'h0)); forvar422 = (forvar422 + (1'h1)))
                    begin
                      reg423 <= (!$signed($unsigned((^~forvar396))));
                    end
                  for (forvar424 = (1'h0); (forvar424 < (2'h2)); forvar424 = (forvar424 + (1'h1)))
                    begin
                      reg425 <= reg301;
                      reg426 <= {(($unsigned(forvar341) ?
                                  reg323 : $signed(forvar399)) ?
                              (!(+reg411)) : $unsigned((^reg412)))};
                      reg427 <= (|($unsigned((reg314 * reg303)) >= (reg322[(1'h1):(1'h1)] || ((8'haa) ?
                          reg411 : (8'hb0)))));
                    end
                end
              else
                begin
                  for (forvar419 = (1'h0); (forvar419 < (2'h2)); forvar419 = (forvar419 + (1'h1)))
                    begin
                      reg420 <= $signed(forvar400);
                      reg421 <= reg342;
                      reg422 <= $signed(forvar385);
                      reg423 <= ($unsigned((&((8'h9d) ? reg345 : reg420))) ?
                          $unsigned($signed($signed(forvar352))) : ($unsigned((+forvar373)) > (&(reg379 + (8'h9f)))));
                    end
                  if (wire292[(3'h6):(2'h2)])
                    begin
                      reg424 <= ({(reg325 >= {forvar391})} ?
                          reg307 : $unsigned((forvar391[(3'h6):(1'h1)] ?
                              $signed((8'hb8)) : (reg423 ? reg311 : reg366))));
                      reg425 <= (reg410 ?
                          reg325[(2'h2):(1'h1)] : $unsigned(({forvar315} ?
                              $signed(forvar352) : forvar378[(1'h1):(1'h0)])));
                      reg426 <= reg417;
                    end
                  else
                    begin
                      reg424 <= $signed(reg310);
                    end
                  for (forvar427 = (1'h0); (forvar427 < (1'h0)); forvar427 = (forvar427 + (1'h1)))
                    begin
                      reg428 <= (reg360[(3'h4):(3'h4)] ?
                          $unsigned(reg388) : (~((reg408 ?
                              forvar386 : reg383) >>> {forvar294})));
                      reg429 <= reg391[(3'h4):(2'h3)];
                      reg430 <= forvar400;
                      reg431 <= (~&{((reg332 ?
                              reg326 : forvar369) >> $signed(reg376))});
                    end
                end
            end
          else
            begin
              if (($signed((reg366 == forvar306)) <= (~$signed(forvar379[(2'h3):(2'h2)]))))
                begin
                  if ($unsigned($unsigned($signed({(8'h9f)}))))
                    begin
                      reg413 <= ((~&forvar352[(1'h0):(1'h0)]) ?
                          (reg405[(2'h2):(1'h0)] != forvar329) : reg321[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg413 <= $signed($signed(forvar399));
                      reg414 <= $unsigned($signed(reg348[(2'h3):(2'h3)]));
                      reg415 <= reg388[(1'h0):(1'h0)];
                      reg416 <= $unsigned({($signed(forvar403) >>> $signed((8'haf)))});
                    end
                  if (reg298)
                    begin
                      reg417 <= ($signed(reg344) & ($signed({reg426}) ?
                          reg362[(3'h4):(1'h0)] : ((-reg398) >>> {reg401})));
                      reg418 <= (($signed((reg385 ^ reg334)) || forvar352[(1'h0):(1'h0)]) ~^ ((~{forvar359}) ?
                          (~(~^reg356)) : (8'ha0)));
                    end
                  else
                    begin
                      reg417 <= {(reg416[(3'h4):(1'h1)] << ($signed(forvar378) ?
                              (reg414 ?
                                  forvar365 : reg366) : (reg339 < reg326)))};
                      reg418 <= reg421[(4'hc):(1'h0)];
                      reg419 <= ({((forvar397 ? reg314 : (8'ha8)) ?
                              $signed(forvar403) : {reg361})} - reg402[(2'h3):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar413 = (1'h0); (forvar413 < (2'h2)); forvar413 = (forvar413 + (1'h1)))
                    begin
                      reg414 <= (reg307 ?
                          $signed(((reg318 ?
                              (8'ha6) : reg405) ~^ $signed(reg302))) : (($unsigned(reg345) ?
                              (reg387 != reg333) : $signed(reg345)) | reg325));
                      reg415 <= ((~|$unsigned($signed(reg331))) ?
                          (((forvar313 == reg348) || $unsigned(reg388)) >> reg389) : reg322);
                      reg416 <= reg322[(3'h7):(3'h5)];
                    end
                end
              reg420 <= reg425[(1'h1):(1'h0)];
              if ($unsigned(forvar315))
                begin
                  reg421 <= $unsigned($unsigned((-(wire293 ?
                      reg360 : reg389))));
                end
              else
                begin
                  for (forvar421 = (1'h0); (forvar421 < (2'h3)); forvar421 = (forvar421 + (1'h1)))
                    begin
                      reg422 <= forvar347;
                      reg423 <= $unsigned(reg423[(1'h0):(1'h0)]);
                      reg424 <= (^~reg347);
                      reg425 <= ((reg322 ?
                              ((reg380 <= forvar336) - reg396) : reg354[(1'h0):(1'h0)]) ?
                          ($unsigned((+reg303)) == forvar379) : {$unsigned({reg378})});
                    end
                  if ((8'hb1))
                    begin
                      reg426 <= forvar344;
                      reg427 <= ($signed((!forvar351[(3'h4):(1'h1)])) < ($signed((forvar329 != reg415)) ?
                          reg404 : ($signed(reg415) * (reg384 ?
                              reg386 : reg419))));
                      reg428 <= (~&((reg386[(2'h3):(2'h2)] ?
                              $signed(reg378) : (-reg346)) ?
                          reg314[(1'h0):(1'h0)] : reg408[(2'h3):(1'h0)]));
                      reg429 <= ((((reg314 && reg362) ?
                          reg428[(4'he):(3'h5)] : reg351) ~^ ((-forvar386) ^~ (reg370 ?
                          reg331 : reg382))) * $signed($unsigned($signed(forvar396))));
                    end
                  else
                    begin
                      reg426 <= wire292[(3'h5):(2'h3)];
                    end
                  for (forvar430 = (1'h0); (forvar430 < (1'h1)); forvar430 = (forvar430 + (1'h1)))
                    begin
                      reg431 <= ($unsigned($unsigned($unsigned(reg298))) & forvar353);
                      reg432 <= reg342;
                    end
                end
              for (forvar433 = (1'h0); (forvar433 < (1'h0)); forvar433 = (forvar433 + (1'h1)))
                begin
                  if (($signed($signed((reg296 > reg406))) >>> $signed((8'h9c))))
                    begin
                      reg434 <= $unsigned(($signed(reg389[(1'h1):(1'h1)]) ?
                          $signed(forvar337) : $signed({forvar336})));
                      reg435 <= reg413[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg434 <= (($unsigned((reg346 - forvar373)) & forvar325) * $unsigned({(reg332 ?
                              reg303 : reg299)}));
                      reg435 <= (reg395 ?
                          ((reg430 ?
                              reg382[(4'ha):(4'h8)] : forvar365) ^~ (forvar315[(3'h4):(2'h3)] ?
                              {(8'hb3)} : reg341)) : reg428);
                      reg436 <= reg356;
                    end
                end
            end
        end
      for (forvar437 = (1'h0); (forvar437 < (2'h3)); forvar437 = (forvar437 + (1'h1)))
        begin
          reg438 <= (|reg360);
          reg439 <= $signed($signed({(^reg438)}));
          reg440 <= forvar306;
        end
    end
  always
    @(posedge clk) begin
      reg441 <= ($signed(forvar397) ^~ (reg374[(1'h0):(1'h0)] | reg349[(2'h2):(2'h2)]));
      for (forvar442 = (1'h0); (forvar442 < (1'h1)); forvar442 = (forvar442 + (1'h1)))
        begin
          if (reg321[(1'h0):(1'h0)])
            begin
              reg443 <= (~^reg354);
              for (forvar444 = (1'h0); (forvar444 < (1'h0)); forvar444 = (forvar444 + (1'h1)))
                begin
                  for (forvar445 = (1'h0); (forvar445 < (2'h3)); forvar445 = (forvar445 + (1'h1)))
                    begin
                      reg446 <= (8'hb4);
                    end
                  for (forvar447 = (1'h0); (forvar447 < (2'h3)); forvar447 = (forvar447 + (1'h1)))
                    begin
                      reg448 <= $signed(((((8'hb3) <<< reg419) | (forvar377 ?
                              reg310 : reg342)) ?
                          $signed((~&reg296)) : $signed(reg322[(3'h6):(1'h0)])));
                      reg449 <= $signed((^~$signed({(8'h9d)})));
                      reg450 <= (^~(8'h9e));
                      reg451 <= (+$signed(((reg385 ? reg423 : reg304) ?
                          reg338[(4'ha):(4'ha)] : $unsigned((8'ha3)))));
                    end
                  for (forvar452 = (1'h0); (forvar452 < (1'h1)); forvar452 = (forvar452 + (1'h1)))
                    begin
                      reg453 <= (reg372[(3'h6):(3'h6)] ?
                          (($signed(reg432) ?
                              ((8'haa) + reg378) : (forvar364 >= forvar422)) ^ {(-reg391)}) : {(+{(8'hb3)})});
                    end
                end
            end
          else
            begin
              for (forvar443 = (1'h0); (forvar443 < (2'h2)); forvar443 = (forvar443 + (1'h1)))
                begin
                  if ($signed($signed((8'hae))))
                    begin
                      reg444 <= reg438;
                      reg445 <= forvar391[(4'h8):(2'h2)];
                      reg446 <= reg375;
                    end
                  else
                    begin
                      reg444 <= ($signed((~&reg417)) ?
                          reg356 : $unsigned($signed((^reg368))));
                      reg445 <= reg378[(2'h2):(2'h2)];
                      reg446 <= (&reg388[(2'h2):(1'h0)]);
                    end
                end
            end
          for (forvar454 = (1'h0); (forvar454 < (2'h3)); forvar454 = (forvar454 + (1'h1)))
            begin
              reg455 <= (~{$unsigned($unsigned(reg379))});
              if (reg371)
                begin
                  for (forvar456 = (1'h0); (forvar456 < (2'h2)); forvar456 = (forvar456 + (1'h1)))
                    begin
                      reg457 <= reg353;
                      reg458 <= reg419[(3'h4):(2'h2)];
                      reg459 <= forvar351[(2'h3):(1'h0)];
                    end
                  reg460 <= (^$unsigned(($signed(forvar369) || $unsigned((8'ha6)))));
                end
              else
                begin
                  if (forvar353[(2'h2):(1'h1)])
                    begin
                      reg456 <= (reg312 ?
                          forvar452[(3'h7):(2'h2)] : (($unsigned(reg352) ?
                              reg460[(1'h1):(1'h1)] : (reg430 ?
                                  wire291 : reg357)) != (~&forvar400)));
                      reg457 <= ({reg451} ?
                          reg339[(3'h6):(3'h4)] : (reg321[(2'h2):(1'h0)] - (^$signed(forvar427))));
                      reg458 <= reg307;
                    end
                  else
                    begin
                      reg456 <= reg404;
                      reg457 <= ((reg460 || (reg446[(3'h7):(1'h0)] & {(8'hb4)})) >= {reg387[(4'hc):(1'h0)]});
                    end
                  for (forvar459 = (1'h0); (forvar459 < (2'h3)); forvar459 = (forvar459 + (1'h1)))
                    begin
                      reg460 <= (((reg388 ^ reg436[(3'h7):(2'h2)]) & $unsigned((reg394 ?
                              reg414 : forvar407))) ?
                          reg296 : {$unsigned($unsigned(reg322))});
                      reg461 <= $unsigned($unsigned(($signed((8'hb0)) ~^ ((8'hb9) >> reg393))));
                    end
                  for (forvar462 = (1'h0); (forvar462 < (2'h3)); forvar462 = (forvar462 + (1'h1)))
                    begin
                      reg463 <= {(-$unsigned($unsigned(forvar396)))};
                      reg464 <= (~|$signed((8'hb4)));
                      reg465 <= ((reg422[(3'h6):(3'h5)] ?
                              forvar400[(3'h6):(2'h2)] : (reg440[(2'h2):(1'h1)] >= (8'h9f))) ?
                          ((&(8'hae)) ?
                              wire293[(4'hc):(4'hb)] : reg428) : reg453[(1'h0):(1'h0)]);
                      reg466 <= (~(&$unsigned((reg353 ? reg332 : forvar353))));
                    end
                end
            end
        end
      if (reg304[(3'h4):(1'h1)])
        begin
          reg467 <= (^({reg419[(4'h9):(3'h7)]} ?
              $signed($signed(reg340)) : $signed(reg457[(3'h7):(3'h4)])));
          if (forvar422[(1'h1):(1'h1)])
            begin
              reg468 <= reg376[(4'hc):(3'h7)];
              if (reg446)
                begin
                  if ((^~({(forvar352 >= forvar397)} ?
                      reg453[(1'h0):(1'h0)] : ((|forvar381) ~^ $unsigned(reg355)))))
                    begin
                      reg469 <= (forvar382[(3'h4):(2'h3)] == (~(forvar454 ?
                          (reg457 * reg412) : forvar462[(4'hc):(4'ha)])));
                      reg470 <= $signed({($unsigned((8'ha3)) | {reg404})});
                      reg471 <= $unsigned((~&reg324));
                    end
                  else
                    begin
                      reg469 <= forvar325[(3'h4):(1'h1)];
                      reg470 <= wire289;
                      reg471 <= {reg335[(3'h6):(3'h5)]};
                      reg472 <= $signed($unsigned((((8'ha0) ? reg357 : reg459) ?
                          (reg333 ^ forvar363) : $unsigned(reg343))));
                    end
                  if ((~^reg341))
                    begin
                      reg473 <= forvar315;
                      reg474 <= reg391;
                      reg475 <= $signed((((reg333 && reg412) + (+reg382)) & (8'h9d)));
                      reg476 <= (($unsigned($unsigned(forvar422)) < ({(8'hb8)} ?
                          ((8'ha7) ?
                              reg466 : reg391) : reg391[(2'h3):(2'h3)])) > (((forvar365 ^ reg469) || $unsigned(reg357)) ?
                          {{(8'hb2)}} : (^~(reg413 ? reg418 : forvar462))));
                    end
                  else
                    begin
                      reg473 <= $signed(({reg411} >= reg312[(1'h0):(1'h0)]));
                    end
                  for (forvar477 = (1'h0); (forvar477 < (2'h3)); forvar477 = (forvar477 + (1'h1)))
                    begin
                      reg478 <= (({$unsigned((8'hb6))} ?
                              (|$signed(reg402)) : reg394) ?
                          (~&(|$unsigned(reg371))) : (reg391 > forvar294));
                    end
                end
              else
                begin
                  for (forvar469 = (1'h0); (forvar469 < (2'h3)); forvar469 = (forvar469 + (1'h1)))
                    begin
                      reg470 <= reg311;
                      reg471 <= $unsigned($signed($signed($signed(reg297))));
                    end
                  for (forvar472 = (1'h0); (forvar472 < (1'h1)); forvar472 = (forvar472 + (1'h1)))
                    begin
                      reg473 <= {((forvar452[(4'hb):(4'ha)] ?
                                  {reg339} : (reg338 <<< forvar337)) ?
                              reg444[(4'h8):(4'h8)] : forvar443[(1'h0):(1'h0)])};
                    end
                end
              for (forvar479 = (1'h0); (forvar479 < (2'h2)); forvar479 = (forvar479 + (1'h1)))
                begin
                  for (forvar480 = (1'h0); (forvar480 < (1'h0)); forvar480 = (forvar480 + (1'h1)))
                    begin
                      reg481 <= (reg327[(4'ha):(4'ha)] ?
                          $unsigned(forvar456[(4'hc):(4'ha)]) : (forvar391[(4'ha):(3'h5)] ?
                              (!(-reg384)) : $unsigned($unsigned(reg298))));
                      reg482 <= ($unsigned(wire293[(3'h7):(2'h3)]) * (reg385[(2'h2):(1'h1)] | (!$unsigned(reg362))));
                      reg483 <= reg375;
                    end
                  for (forvar484 = (1'h0); (forvar484 < (2'h2)); forvar484 = (forvar484 + (1'h1)))
                    begin
                      reg485 <= $unsigned($signed((((8'hb6) ?
                              reg399 : forvar296) ?
                          (reg449 >>> (8'h9f)) : reg472[(2'h3):(2'h2)])));
                      reg486 <= (($unsigned($signed((8'ha0))) <= $unsigned(reg471[(3'h5):(1'h0)])) ?
                          {{forvar320[(1'h1):(1'h1)]}} : $unsigned((forvar452 & (forvar406 >= reg467))));
                    end
                  if (reg463)
                    begin
                      reg487 <= {(reg453 <= reg342[(1'h0):(1'h0)])};
                      reg488 <= $unsigned((-reg343));
                      reg489 <= $signed({(reg389 <= forvar365[(3'h6):(3'h6)])});
                      reg490 <= $signed((-($signed(forvar386) != (forvar295 ?
                          reg444 : forvar306))));
                    end
                  else
                    begin
                      reg487 <= reg304[(1'h0):(1'h0)];
                      reg488 <= (forvar430 ?
                          ((reg414 == forvar445[(2'h3):(1'h0)]) ?
                              reg303[(2'h2):(2'h2)] : {$signed(reg348)}) : $signed(forvar480));
                      reg489 <= (~^$unsigned((!(~reg328))));
                      reg490 <= ($signed(((~^(8'hb3)) >> (+(8'hb4)))) ?
                          forvar296 : (~((reg323 ?
                              (8'ha8) : reg453) | (|forvar413))));
                    end
                end
              for (forvar491 = (1'h0); (forvar491 < (2'h3)); forvar491 = (forvar491 + (1'h1)))
                begin
                  reg492 <= reg463[(3'h4):(2'h2)];
                end
            end
          else
            begin
              for (forvar468 = (1'h0); (forvar468 < (2'h2)); forvar468 = (forvar468 + (1'h1)))
                begin
                  if ($unsigned(reg393[(2'h2):(2'h2)]))
                    begin
                      reg469 <= (~^$unsigned(forvar405[(3'h6):(1'h0)]));
                      reg470 <= (reg398[(1'h0):(1'h0)] ?
                          forvar433[(3'h4):(3'h4)] : ((((8'hb5) >= reg490) ?
                                  {(8'ha1)} : $unsigned(forvar296)) ?
                              reg460 : (^~reg413[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg469 <= (~^($signed((reg490 + forvar359)) <= (^(reg435 >>> reg392))));
                      reg470 <= ($signed((reg324 ?
                          {reg332} : $unsigned(forvar352))) ~^ (({(8'hb4)} ^ (reg382 == forvar444)) <= $unsigned($unsigned(reg420))));
                      reg471 <= reg423;
                      reg472 <= $signed(reg305);
                    end
                  if (($signed(reg399[(5'h10):(4'hc)]) ?
                      reg298 : (^forvar351[(2'h2):(1'h0)])))
                    begin
                      reg473 <= forvar454;
                      reg474 <= forvar422[(3'h6):(1'h0)];
                      reg475 <= $signed(forvar405[(1'h1):(1'h0)]);
                      reg476 <= (!($signed((reg489 >= (8'ha9))) ?
                          {forvar376[(2'h2):(1'h1)]} : (~|forvar459)));
                    end
                  else
                    begin
                      reg473 <= ($unsigned((~|reg356)) ?
                          wire289[(4'ha):(2'h3)] : reg435[(3'h6):(3'h4)]);
                    end
                  if ($unsigned(reg471))
                    begin
                      reg477 <= (-reg319[(1'h0):(1'h0)]);
                      reg478 <= forvar479;
                    end
                  else
                    begin
                      reg477 <= reg374;
                      reg478 <= ($signed($signed((~forvar454))) ?
                          {reg361[(4'hc):(3'h4)]} : ($unsigned((forvar386 - reg366)) - reg489));
                    end
                  for (forvar479 = (1'h0); (forvar479 < (1'h1)); forvar479 = (forvar479 + (1'h1)))
                    begin
                      reg480 <= forvar341[(4'hb):(3'h5)];
                      reg481 <= (reg344 > $signed(reg316));
                    end
                end
              for (forvar482 = (1'h0); (forvar482 < (2'h3)); forvar482 = (forvar482 + (1'h1)))
                begin
                  for (forvar483 = (1'h0); (forvar483 < (2'h3)); forvar483 = (forvar483 + (1'h1)))
                    begin
                      reg484 <= forvar369[(3'h4):(1'h0)];
                    end
                  for (forvar485 = (1'h0); (forvar485 < (2'h3)); forvar485 = (forvar485 + (1'h1)))
                    begin
                      reg486 <= $unsigned(reg478);
                      reg487 <= forvar491[(2'h3):(2'h2)];
                    end
                end
            end
        end
      else
        begin
          for (forvar467 = (1'h0); (forvar467 < (1'h1)); forvar467 = (forvar467 + (1'h1)))
            begin
              reg468 <= reg299;
              reg469 <= reg487[(2'h2):(1'h1)];
            end
          if ((8'hb2))
            begin
              for (forvar470 = (1'h0); (forvar470 < (2'h3)); forvar470 = (forvar470 + (1'h1)))
                begin
                  if (((8'ha6) ?
                      (forvar454 ~^ forvar477[(4'h9):(3'h5)]) : reg385[(2'h2):(2'h2)]))
                    begin
                      reg471 <= (((~|(reg461 ? forvar472 : reg310)) ?
                              $signed(reg314) : {$unsigned(reg411)}) ?
                          $signed(reg418[(3'h5):(2'h2)]) : ((forvar382[(2'h3):(2'h2)] ?
                              (reg432 ?
                                  reg383 : reg340) : reg356) + forvar399[(2'h3):(1'h1)]));
                      reg472 <= {reg417};
                      reg473 <= $signed($signed(wire290[(4'hf):(3'h6)]));
                      reg474 <= forvar419;
                    end
                  else
                    begin
                      reg471 <= $unsigned($signed($signed((reg316 <= (8'hab)))));
                      reg472 <= $unsigned(reg305);
                    end
                  if (forvar363)
                    begin
                      reg475 <= (-{reg411[(1'h1):(1'h1)]});
                      reg476 <= reg325[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg475 <= ($signed((reg307[(3'h7):(3'h4)] ^~ forvar483[(3'h4):(2'h2)])) ~^ (8'ha9));
                      reg476 <= forvar469[(1'h1):(1'h0)];
                      reg477 <= {($signed($signed(forvar341)) << {(~reg410)})};
                      reg478 <= reg449[(4'ha):(2'h3)];
                    end
                  for (forvar479 = (1'h0); (forvar479 < (2'h3)); forvar479 = (forvar479 + (1'h1)))
                    begin
                      reg480 <= $unsigned(reg482[(4'he):(4'hd)]);
                      reg481 <= (((&(forvar480 ? forvar462 : reg375)) ?
                              (-(forvar353 ?
                                  reg357 : (8'hb4))) : $unsigned((reg367 ?
                                  (8'haa) : reg482))) ?
                          $signed($unsigned(forvar422[(3'h4):(2'h2)])) : ($unsigned($signed(reg450)) ?
                              (&reg360[(1'h0):(1'h0)]) : ($signed((8'ha1)) ?
                                  {wire291} : {reg480})));
                    end
                end
              if (($signed((reg317[(1'h0):(1'h0)] ? (&forvar462) : {reg356})) ?
                  reg470[(4'h8):(2'h3)] : $signed(forvar386)))
                begin
                  for (forvar482 = (1'h0); (forvar482 < (1'h1)); forvar482 = (forvar482 + (1'h1)))
                    begin
                      reg483 <= (~^(!$unsigned((8'ha4))));
                      reg484 <= $unsigned((8'h9c));
                      reg485 <= (^~$unsigned((^~$signed(reg395))));
                    end
                  if (reg484)
                    begin
                      reg486 <= $unsigned(((reg304[(2'h2):(1'h1)] ?
                          (&reg370) : forvar443) && reg352[(4'he):(4'hb)]));
                      reg487 <= (reg339[(2'h2):(2'h2)] ?
                          $unsigned(reg343[(3'h4):(2'h3)]) : (~^({reg484} ?
                              (forvar477 ?
                                  reg426 : forvar480) : (forvar364 ^~ reg341))));
                      reg488 <= (~&reg472[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg486 <= reg484;
                      reg487 <= forvar413[(4'hf):(2'h2)];
                      reg488 <= (~(forvar483[(2'h2):(1'h0)] ?
                          forvar479[(1'h0):(1'h0)] : $signed((~&reg349))));
                      reg489 <= reg417;
                    end
                  if (((reg358[(1'h0):(1'h0)] - $unsigned($signed(forvar344))) ?
                      ({$unsigned(forvar467)} ?
                          (-reg489[(1'h1):(1'h1)]) : ((reg394 ?
                              reg456 : reg465) | (!reg404))) : forvar403[(3'h6):(3'h6)]))
                    begin
                      reg490 <= {(^((+forvar352) != $unsigned(forvar414)))};
                    end
                  else
                    begin
                      reg490 <= (($unsigned(forvar407) >>> $signed(forvar480)) || forvar359[(4'ha):(3'h5)]);
                    end
                  reg491 <= reg415;
                end
              else
                begin
                  for (forvar482 = (1'h0); (forvar482 < (2'h3)); forvar482 = (forvar482 + (1'h1)))
                    begin
                      reg483 <= $signed((8'hb9));
                    end
                end
              if ((forvar353 ?
                  (~|({reg314} ?
                      reg312[(2'h3):(1'h1)] : {reg420})) : ($unsigned(reg384[(4'h8):(1'h1)]) ?
                      ((reg448 < reg426) <<< reg391) : $signed($unsigned(reg403)))))
                begin
                  reg492 <= (-reg311[(1'h1):(1'h0)]);
                  for (forvar493 = (1'h0); (forvar493 < (1'h0)); forvar493 = (forvar493 + (1'h1)))
                    begin
                      reg494 <= (reg407 + {($unsigned(reg345) >= $unsigned((8'ha3)))});
                    end
                  if ((+$signed(forvar320)))
                    begin
                      reg495 <= (8'ha0);
                      reg496 <= (((|reg330) >> $signed($signed(reg362))) * reg436[(2'h3):(2'h2)]);
                      reg497 <= (&(|forvar482));
                    end
                  else
                    begin
                      reg495 <= (reg411[(1'h1):(1'h0)] <= (reg411[(1'h1):(1'h0)] ?
                          (reg371[(4'h8):(2'h3)] - reg396) : {(forvar470 <<< reg388)}));
                      reg496 <= reg327[(4'hd):(3'h4)];
                      reg497 <= forvar373;
                      reg498 <= (forvar378 ?
                          forvar472[(4'hc):(4'h8)] : (8'hb5));
                    end
                  if (reg368[(2'h3):(2'h3)])
                    begin
                      reg499 <= reg460[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg499 <= ((+(~^$signed(reg299))) ?
                          (~|reg379[(2'h2):(1'h0)]) : ((reg498 ?
                              $unsigned(reg469) : $unsigned(forvar378)) <= $unsigned(((8'hb5) <= forvar396))));
                      reg500 <= $signed($signed(forvar320[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar492 = (1'h0); (forvar492 < (1'h0)); forvar492 = (forvar492 + (1'h1)))
                    begin
                      reg493 <= (~|({reg344} & (reg471[(3'h7):(2'h3)] + reg492)));
                      reg494 <= $signed(forvar433[(3'h5):(1'h1)]);
                      reg495 <= reg391;
                    end
                  if ($unsigned($unsigned((|(reg360 <<< (8'hba))))))
                    begin
                      reg496 <= (^~(reg425 ?
                          ((reg366 ? forvar468 : (8'hae)) ?
                              (forvar382 ?
                                  reg358 : forvar493) : {(8'ha2)}) : reg381[(2'h3):(1'h1)]));
                      reg497 <= (8'h9c);
                      reg498 <= $signed((^$unsigned(((8'haf) ?
                          wire292 : reg414))));
                      reg499 <= $signed($unsigned((8'hb2)));
                    end
                  else
                    begin
                      reg496 <= {$signed(reg398[(1'h0):(1'h0)])};
                      reg497 <= reg461;
                      reg498 <= (-(($signed(forvar491) ?
                              $signed(reg375) : $signed((8'hb7))) ?
                          forvar421[(3'h6):(2'h3)] : {$signed((8'ha2))}));
                      reg499 <= {$signed((reg416[(2'h3):(2'h3)] && (~|reg328)))};
                    end
                end
              for (forvar501 = (1'h0); (forvar501 < (2'h3)); forvar501 = (forvar501 + (1'h1)))
                begin
                  reg502 <= (forvar421[(2'h2):(2'h2)] ?
                      reg300 : wire288[(2'h2):(1'h0)]);
                  for (forvar503 = (1'h0); (forvar503 < (1'h0)); forvar503 = (forvar503 + (1'h1)))
                    begin
                      reg504 <= reg390;
                      reg505 <= ({forvar424} ?
                          ((&forvar364) ?
                              $unsigned(reg314[(3'h4):(1'h1)]) : $unsigned(forvar407[(2'h3):(2'h2)])) : $signed(reg432));
                      reg506 <= forvar296;
                    end
                end
            end
          else
            begin
              for (forvar470 = (1'h0); (forvar470 < (1'h1)); forvar470 = (forvar470 + (1'h1)))
                begin
                  for (forvar471 = (1'h0); (forvar471 < (2'h3)); forvar471 = (forvar471 + (1'h1)))
                    begin
                      reg472 <= $signed($signed((^{reg383})));
                    end
                end
              if ($signed((^~forvar353[(1'h0):(1'h0)])))
                begin
                  for (forvar473 = (1'h0); (forvar473 < (2'h2)); forvar473 = (forvar473 + (1'h1)))
                    begin
                      reg474 <= reg476[(2'h2):(2'h2)];
                      reg475 <= {{reg375}};
                    end
                  if (reg324[(1'h1):(1'h1)])
                    begin
                      reg476 <= reg357;
                      reg477 <= {((+{forvar456}) ~^ reg388[(2'h3):(1'h0)])};
                    end
                  else
                    begin
                      reg476 <= (8'ha9);
                      reg477 <= $unsigned(reg353[(1'h1):(1'h0)]);
                      reg478 <= reg465;
                    end
                  reg479 <= reg446;
                end
              else
                begin
                  for (forvar473 = (1'h0); (forvar473 < (2'h3)); forvar473 = (forvar473 + (1'h1)))
                    begin
                      reg474 <= forvar294[(1'h1):(1'h1)];
                    end
                end
              reg480 <= (($signed({reg341}) ?
                  $signed($unsigned(reg341)) : (reg493 ?
                      $signed(forvar373) : (8'ha2))) >>> reg439[(3'h4):(2'h3)]);
              if ((8'ha3))
                begin
                  for (forvar481 = (1'h0); (forvar481 < (1'h1)); forvar481 = (forvar481 + (1'h1)))
                    begin
                      reg482 <= ({{(~&reg502)}} > (+(~|(~^(8'hb6)))));
                      reg483 <= (~$signed($unsigned((8'ha9))));
                      reg484 <= $signed(($signed(reg492) | (forvar491 ?
                          $signed((8'hb9)) : forvar462[(1'h1):(1'h1)])));
                    end
                  for (forvar485 = (1'h0); (forvar485 < (1'h0)); forvar485 = (forvar485 + (1'h1)))
                    begin
                      reg486 <= ((8'ha7) ?
                          $unsigned(((reg367 ?
                              reg314 : reg325) || (8'hab))) : (~^$unsigned($unsigned((8'ha5)))));
                      reg487 <= (forvar295[(3'h4):(1'h1)] ~^ reg404);
                      reg488 <= ($unsigned(reg419) <<< $signed(forvar396[(2'h2):(2'h2)]));
                    end
                end
              else
                begin
                  if (({$unsigned(reg347)} >= (8'hb7)))
                    begin
                      reg481 <= forvar381[(1'h0):(1'h0)];
                      reg482 <= (reg311 <= $unsigned({forvar427}));
                      reg483 <= reg378[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg481 <= ((($unsigned(reg298) ?
                          (+(8'hb6)) : $signed(reg401)) <<< $signed((forvar295 ^~ reg383))) <<< ((((8'hba) | reg341) ?
                          (reg460 | (8'hba)) : forvar427) == ((reg344 ^~ reg430) <= (~|(8'hb8)))));
                      reg482 <= (forvar480[(2'h3):(1'h0)] ?
                          (!($unsigned((8'hb6)) ?
                              (forvar405 + reg349) : (forvar491 - reg497))) : $unsigned((reg312 ?
                              (forvar491 < reg399) : $signed(reg468))));
                    end
                  for (forvar484 = (1'h0); (forvar484 < (1'h0)); forvar484 = (forvar484 + (1'h1)))
                    begin
                      reg485 <= $signed($signed(((forvar382 & reg500) ?
                          $unsigned(forvar493) : $signed(reg497))));
                      reg486 <= $signed((~&reg506[(3'h7):(1'h1)]));
                      reg487 <= $signed($unsigned(reg296));
                      reg488 <= $signed((+(|{reg339})));
                    end
                  for (forvar489 = (1'h0); (forvar489 < (2'h2)); forvar489 = (forvar489 + (1'h1)))
                    begin
                      reg490 <= ($unsigned(((&reg341) ?
                              {reg457} : $signed(forvar462))) ?
                          (reg398[(3'h4):(1'h0)] && {reg353}) : $signed((!forvar406[(3'h6):(3'h6)])));
                    end
                end
            end
          reg507 <= (8'ha7);
        end
      if ($signed(({(~^reg464)} ?
          (8'hb3) : $unsigned((forvar480 << forvar306)))))
        begin
          reg508 <= forvar421[(2'h2):(2'h2)];
          for (forvar509 = (1'h0); (forvar509 < (2'h3)); forvar509 = (forvar509 + (1'h1)))
            begin
              if (reg403)
                begin
                  reg510 <= forvar503;
                  for (forvar511 = (1'h0); (forvar511 < (2'h2)); forvar511 = (forvar511 + (1'h1)))
                    begin
                      reg512 <= {$signed((|reg480))};
                    end
                  if ($unsigned((|(+(8'hb5)))))
                    begin
                      reg513 <= {{reg412}};
                    end
                  else
                    begin
                      reg513 <= {$unsigned($signed($signed(reg505)))};
                      reg514 <= (!$signed((~|((8'h9e) ? (8'hba) : reg492))));
                      reg515 <= (reg407[(4'h8):(4'h8)] ?
                          reg508[(3'h5):(1'h0)] : reg354);
                      reg516 <= reg461;
                    end
                  for (forvar517 = (1'h0); (forvar517 < (1'h1)); forvar517 = (forvar517 + (1'h1)))
                    begin
                      reg518 <= (reg380 - reg375);
                      reg519 <= $unsigned((~^(8'hb1)));
                    end
                end
              else
                begin
                  reg510 <= $unsigned((forvar456[(2'h3):(1'h0)] ~^ ((forvar363 ?
                          reg489 : reg302) ?
                      (reg453 ? reg441 : forvar421) : reg464)));
                  reg511 <= (^~$unsigned((((8'had) ? reg358 : reg334) ?
                      $signed(reg328) : (forvar484 ? reg483 : wire289))));
                end
              if ($signed($signed(reg297)))
                begin
                  for (forvar520 = (1'h0); (forvar520 < (1'h1)); forvar520 = (forvar520 + (1'h1)))
                    begin
                      reg521 <= (forvar365[(2'h3):(1'h1)] ?
                          $unsigned($signed((reg408 ?
                              reg476 : forvar479))) : $signed((|(forvar477 >> reg362))));
                    end
                  for (forvar522 = (1'h0); (forvar522 < (1'h1)); forvar522 = (forvar522 + (1'h1)))
                    begin
                      reg523 <= {(^~(^~reg470))};
                      reg524 <= ({reg408[(1'h1):(1'h0)]} >= (|$signed($signed(forvar483))));
                    end
                  for (forvar525 = (1'h0); (forvar525 < (2'h3)); forvar525 = (forvar525 + (1'h1)))
                    begin
                      reg526 <= (forvar347 + $signed(forvar485[(2'h2):(1'h1)]));
                      reg527 <= reg352;
                      reg528 <= ($signed(reg468[(4'h8):(1'h0)]) ?
                          reg430 : {reg338});
                    end
                  if (reg481[(4'ha):(3'h7)])
                    begin
                      reg529 <= (~|(($unsigned(reg458) ?
                              (&reg491) : ((8'ha7) ? forvar503 : (8'hac))) ?
                          ({reg389} + {(8'h9e)}) : reg460[(3'h6):(3'h5)]));
                      reg530 <= ($signed((~((8'ha2) ?
                          (8'ha8) : forvar414))) ~^ $signed($signed(reg302[(2'h3):(2'h2)])));
                      reg531 <= (({(reg391 ? reg473 : reg307)} ?
                          (reg372 > (&reg334)) : $signed((~^reg334))) == $signed((-forvar427[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg529 <= forvar325;
                      reg530 <= (reg494[(3'h6):(2'h3)] ?
                          $signed(forvar525[(4'h9):(3'h7)]) : (8'hb5));
                      reg531 <= $signed((forvar296[(1'h0):(1'h0)] ?
                          ($signed(reg477) ?
                              (8'hb6) : reg466[(1'h1):(1'h1)]) : (reg381[(4'ha):(2'h2)] << (forvar329 ?
                              (8'hab) : reg358))));
                    end
                end
              else
                begin
                  for (forvar520 = (1'h0); (forvar520 < (1'h1)); forvar520 = (forvar520 + (1'h1)))
                    begin
                      reg521 <= (~$unsigned($unsigned($unsigned(reg496))));
                    end
                  for (forvar522 = (1'h0); (forvar522 < (1'h1)); forvar522 = (forvar522 + (1'h1)))
                    begin
                      reg523 <= reg450[(2'h3):(2'h2)];
                      reg524 <= (((((8'h9d) ?
                                  forvar520 : forvar365) ^~ (forvar485 && forvar501)) ?
                              forvar442[(1'h0):(1'h0)] : ($unsigned(reg314) | forvar313[(3'h7):(2'h3)])) ?
                          reg367[(1'h1):(1'h1)] : (+reg514));
                    end
                end
              reg532 <= $signed(reg386[(3'h5):(1'h1)]);
            end
          for (forvar533 = (1'h0); (forvar533 < (2'h3)); forvar533 = (forvar533 + (1'h1)))
            begin
              if (reg351[(1'h1):(1'h0)])
                begin
                  for (forvar534 = (1'h0); (forvar534 < (1'h1)); forvar534 = (forvar534 + (1'h1)))
                    begin
                      reg535 <= reg421;
                    end
                  for (forvar536 = (1'h0); (forvar536 < (2'h3)); forvar536 = (forvar536 + (1'h1)))
                    begin
                      reg537 <= (forvar381[(3'h4):(3'h4)] ?
                          (^~{$signed(reg347)}) : ((forvar509[(4'h8):(4'h8)] + (~^reg302)) >= reg316));
                    end
                end
              else
                begin
                  reg534 <= reg416[(4'h9):(3'h7)];
                  reg535 <= (reg444 ?
                      forvar489 : ($signed((reg429 && reg486)) ?
                          reg422[(1'h0):(1'h0)] : (~forvar403)));
                end
              if (($signed(forvar503[(1'h1):(1'h1)]) || $unsigned($signed($unsigned(forvar308)))))
                begin
                  for (forvar538 = (1'h0); (forvar538 < (1'h0)); forvar538 = (forvar538 + (1'h1)))
                    begin
                      reg539 <= $signed($signed($unsigned((reg507 ?
                          reg532 : forvar481))));
                      reg540 <= (^~reg456[(2'h3):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar538 = (1'h0); (forvar538 < (1'h0)); forvar538 = (forvar538 + (1'h1)))
                    begin
                      reg539 <= reg314[(1'h0):(1'h0)];
                      reg540 <= $unsigned((&((reg531 <<< reg490) >>> (~|reg368))));
                      reg541 <= reg423;
                    end
                end
            end
          for (forvar542 = (1'h0); (forvar542 < (1'h0)); forvar542 = (forvar542 + (1'h1)))
            begin
              for (forvar543 = (1'h0); (forvar543 < (1'h1)); forvar543 = (forvar543 + (1'h1)))
                begin
                  for (forvar544 = (1'h0); (forvar544 < (2'h3)); forvar544 = (forvar544 + (1'h1)))
                    begin
                      reg545 <= $signed(($unsigned({forvar363}) ?
                          ($unsigned(reg349) ?
                              (+reg439) : reg384[(2'h3):(1'h1)]) : $signed($signed(reg322))));
                      reg546 <= $signed(reg360);
                      reg547 <= reg441;
                      reg548 <= {(&$unsigned($unsigned(reg325)))};
                    end
                  if (((^{$signed(reg340)}) ?
                      reg507[(3'h7):(3'h4)] : forvar427))
                    begin
                      reg549 <= $signed($unsigned(forvar536));
                      reg550 <= $signed($signed($signed((reg335 ?
                          reg330 : reg500))));
                      reg551 <= reg399;
                      reg552 <= {forvar534};
                    end
                  else
                    begin
                      reg549 <= (8'hb0);
                      reg550 <= ($signed(((reg361 == reg406) ^ (reg495 <= (8'hb5)))) ?
                          ($signed(reg391) < $signed({forvar336})) : $unsigned((forvar342[(4'h9):(4'h9)] || reg545[(1'h1):(1'h1)])));
                    end
                  if ((+reg469[(4'h8):(4'h8)]))
                    begin
                      reg553 <= (reg407 ?
                          (((reg489 <= forvar493) << $signed(reg379)) ?
                              (reg434 ~^ (^reg551)) : (&reg448[(2'h3):(1'h0)])) : $unsigned(((^~forvar414) ?
                              $unsigned(reg335) : forvar536)));
                      reg554 <= forvar313[(2'h3):(1'h0)];
                      reg555 <= (reg519 ?
                          reg360[(1'h1):(1'h0)] : forvar344[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg553 <= (({reg339} >> (|(~|reg372))) ?
                          forvar351 : {$unsigned(reg529[(1'h1):(1'h0)])});
                      reg554 <= {((~^reg330) >>> reg401)};
                      reg555 <= {reg328};
                      reg556 <= ((forvar468[(4'h8):(3'h4)] == (reg409 <<< $signed(reg528))) ^~ $unsigned(reg441));
                    end
                end
              reg557 <= $signed((|{(forvar379 > (8'hab))}));
            end
        end
      else
        begin
          if ($unsigned(reg327))
            begin
              if ($signed((8'haa)))
                begin
                  if ((reg556[(1'h1):(1'h1)] ^ $unsigned(((~wire292) ?
                      $signed((8'h9f)) : reg414[(2'h3):(2'h3)]))))
                    begin
                      reg508 <= (($unsigned((reg494 ?
                          reg384 : (8'hb1))) && (reg296 && $signed((8'ha3)))) <<< reg326);
                    end
                  else
                    begin
                      reg508 <= {reg540[(1'h0):(1'h0)]};
                    end
                end
              else
                begin
                  if (reg420)
                    begin
                      reg508 <= {((|reg540[(1'h1):(1'h0)]) ?
                              $signed({reg376}) : $unsigned(reg420))};
                      reg509 <= {({reg353} ^~ $signed((forvar503 ~^ reg361)))};
                      reg510 <= ($unsigned(((forvar447 + reg500) ?
                          (reg539 + reg449) : (&forvar353))) << (forvar400 ?
                          (^(reg556 ?
                              (8'hb1) : (8'ha8))) : {(forvar543 && (8'hb3))}));
                    end
                  else
                    begin
                      reg508 <= (((reg488 != (!(8'h9f))) ?
                          ((reg393 ?
                              reg518 : forvar294) == (forvar341 <= forvar533)) : reg356[(3'h7):(3'h4)]) <= ($signed({(8'hb3)}) != ($unsigned(reg334) & $unsigned(forvar456))));
                    end
                end
              for (forvar511 = (1'h0); (forvar511 < (2'h2)); forvar511 = (forvar511 + (1'h1)))
                begin
                  for (forvar512 = (1'h0); (forvar512 < (2'h2)); forvar512 = (forvar512 + (1'h1)))
                    begin
                      reg513 <= $signed((~&(reg300[(4'he):(4'h9)] ?
                          reg391[(1'h1):(1'h0)] : {reg321})));
                    end
                  for (forvar514 = (1'h0); (forvar514 < (2'h3)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= $unsigned((~&reg456[(3'h4):(2'h2)]));
                    end
                  if (((~|(^{reg449})) ^ reg376))
                    begin
                      reg516 <= (8'hac);
                      reg517 <= reg356;
                      reg518 <= {(&reg553)};
                    end
                  else
                    begin
                      reg516 <= $signed((forvar525[(2'h3):(1'h0)] > (~^{forvar482})));
                      reg517 <= forvar313[(1'h1):(1'h0)];
                      reg518 <= $unsigned($signed(reg317));
                      reg519 <= (reg488[(2'h2):(1'h1)] && ({reg344[(3'h5):(3'h4)]} <<< $signed((reg459 ?
                          forvar404 : wire291))));
                    end
                  if (reg399[(1'h1):(1'h1)])
                    begin
                      reg520 <= $unsigned((reg425 != reg394));
                      reg521 <= (((~reg458[(2'h3):(2'h3)]) | $unsigned($signed(forvar443))) ?
                          ({(8'hb2)} ?
                              $unsigned($signed(forvar296)) : $signed((reg466 ?
                                  forvar396 : forvar376))) : reg409);
                      reg522 <= reg491;
                    end
                  else
                    begin
                      reg520 <= forvar543[(1'h0):(1'h0)];
                      reg521 <= (((reg407 ?
                              (reg463 << reg382) : reg556) * reg408) ?
                          $signed(forvar351) : (^~(~$signed((8'ha3)))));
                      reg522 <= ((8'hb4) >> $unsigned((~(forvar385 ?
                          reg405 : reg302))));
                    end
                end
              for (forvar523 = (1'h0); (forvar523 < (2'h3)); forvar523 = (forvar523 + (1'h1)))
                begin
                  for (forvar524 = (1'h0); (forvar524 < (2'h2)); forvar524 = (forvar524 + (1'h1)))
                    begin
                      reg525 <= ($unsigned(reg357[(4'h8):(1'h0)]) >>> wire288);
                      reg526 <= (+(reg551[(4'h8):(1'h0)] ?
                          ((reg488 ? (8'haf) : reg524) ?
                              (8'hac) : (~&reg441)) : (reg343[(1'h1):(1'h0)] <<< (~&reg403))));
                    end
                  for (forvar527 = (1'h0); (forvar527 < (2'h2)); forvar527 = (forvar527 + (1'h1)))
                    begin
                      reg528 <= {(~|$unsigned($unsigned(reg352)))};
                    end
                  for (forvar529 = (1'h0); (forvar529 < (2'h3)); forvar529 = (forvar529 + (1'h1)))
                    begin
                      reg530 <= ((^$signed($unsigned(reg355))) >> ((~&$signed(forvar378)) ~^ reg525));
                      reg531 <= (8'hac);
                      reg532 <= {reg441};
                    end
                  for (forvar533 = (1'h0); (forvar533 < (1'h1)); forvar533 = (forvar533 + (1'h1)))
                    begin
                      reg534 <= $signed(($unsigned((~reg410)) ?
                          reg347[(3'h6):(2'h3)] : (8'haa)));
                      reg535 <= (reg341[(1'h1):(1'h0)] ?
                          reg535 : reg347[(3'h4):(2'h3)]);
                    end
                end
              for (forvar536 = (1'h0); (forvar536 < (2'h3)); forvar536 = (forvar536 + (1'h1)))
                begin
                  for (forvar537 = (1'h0); (forvar537 < (1'h0)); forvar537 = (forvar537 + (1'h1)))
                    begin
                      reg538 <= (8'hb4);
                      reg539 <= forvar501;
                      reg540 <= (((^$signed((8'hb3))) >>> reg525) != ((~|(reg468 ?
                          (8'hba) : reg445)) && reg537[(2'h2):(2'h2)]));
                    end
                end
            end
          else
            begin
              if ((({reg309} ?
                  ($unsigned((8'hac)) == (|reg506)) : $signed($signed(reg522))) - forvar365))
                begin
                  for (forvar508 = (1'h0); (forvar508 < (1'h1)); forvar508 = (forvar508 + (1'h1)))
                    begin
                      reg509 <= (forvar320[(2'h2):(2'h2)] <= $unsigned($unsigned($signed(forvar514))));
                    end
                  if ((reg497[(4'hf):(3'h6)] >= $signed(((reg487 ?
                      reg527 : forvar493) < {reg372}))))
                    begin
                      reg510 <= (8'h9e);
                      reg511 <= reg438[(1'h1):(1'h0)];
                      reg512 <= $signed($signed(((forvar381 ?
                          reg493 : (8'h9d)) << (!forvar534))));
                    end
                  else
                    begin
                      reg510 <= $signed(reg316[(3'h5):(1'h0)]);
                      reg511 <= $signed(({(reg459 + reg495)} | $signed(reg335)));
                    end
                  if ($signed(reg554))
                    begin
                      reg513 <= ((reg435 || forvar489) - ({((8'ha3) && reg468)} <= $signed((reg460 ?
                          reg459 : forvar308))));
                      reg514 <= (&(~^($unsigned(reg362) >> $unsigned(wire290))));
                    end
                  else
                    begin
                      reg513 <= (~^$unsigned($unsigned($unsigned((8'hb7)))));
                      reg514 <= (|forvar483);
                      reg515 <= $unsigned(reg493);
                    end
                end
              else
                begin
                  if ((~&(~&(reg451[(4'hc):(1'h1)] ?
                      reg449[(4'he):(4'hc)] : $unsigned((8'hab))))))
                    begin
                      reg508 <= (8'ha4);
                      reg509 <= (forvar527 & reg380);
                      reg510 <= $signed((((reg478 ?
                          reg382 : reg366) - $unsigned(forvar379)) == ({forvar406} ?
                          $unsigned(reg468) : reg556[(3'h5):(3'h5)])));
                    end
                  else
                    begin
                      reg508 <= ((forvar373[(4'hd):(2'h2)] ?
                              (~(&reg496)) : reg429) ?
                          (8'hb1) : reg351[(2'h3):(2'h2)]);
                      reg509 <= reg409[(2'h2):(1'h1)];
                      reg510 <= ($unsigned($signed((forvar489 ~^ reg423))) ?
                          ($signed((forvar369 <= (8'ha0))) ?
                              forvar462 : ($unsigned(reg362) >= forvar459[(4'ha):(4'h8)])) : ((forvar489 <= (~&reg344)) ?
                              (reg483 ?
                                  $signed(reg528) : (~|(8'hb7))) : $unsigned($unsigned(reg356))));
                    end
                  for (forvar511 = (1'h0); (forvar511 < (1'h1)); forvar511 = (forvar511 + (1'h1)))
                    begin
                      reg512 <= forvar405[(4'h8):(2'h3)];
                      reg513 <= $unsigned(($signed($unsigned(reg402)) >>> reg326));
                    end
                  for (forvar514 = (1'h0); (forvar514 < (2'h2)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= (reg445[(1'h1):(1'h0)] ?
                          reg399 : (forvar413[(3'h7):(2'h2)] + $signed((~&reg444))));
                      reg516 <= {{reg340}};
                    end
                end
              for (forvar517 = (1'h0); (forvar517 < (2'h2)); forvar517 = (forvar517 + (1'h1)))
                begin
                  if ({wire292[(1'h1):(1'h1)]})
                    begin
                      reg518 <= $unsigned(reg516);
                    end
                  else
                    begin
                      reg518 <= forvar369[(1'h1):(1'h1)];
                      reg519 <= $signed($unsigned(((^~wire289) <= $signed(forvar529))));
                      reg520 <= ({forvar336} + forvar406[(3'h4):(1'h1)]);
                    end
                  reg521 <= (8'hb3);
                  for (forvar522 = (1'h0); (forvar522 < (2'h3)); forvar522 = (forvar522 + (1'h1)))
                    begin
                      reg523 <= ($unsigned({((8'hba) >> reg416)}) ?
                          (forvar483 ?
                              (reg352 == reg307[(1'h0):(1'h0)]) : $signed($unsigned(reg418))) : {(reg314 != (reg531 ?
                                  (8'hb6) : reg403))});
                    end
                end
            end
          if ($signed((-reg332)))
            begin
              for (forvar541 = (1'h0); (forvar541 < (1'h1)); forvar541 = (forvar541 + (1'h1)))
                begin
                  if ($unsigned($unsigned($signed(forvar433))))
                    begin
                      reg542 <= ({reg473[(2'h3):(1'h0)]} || reg415[(2'h3):(2'h2)]);
                      reg543 <= ($signed($unsigned((^forvar294))) ?
                          $unsigned(forvar482) : {reg509});
                    end
                  else
                    begin
                      reg542 <= (+forvar473[(1'h1):(1'h1)]);
                      reg543 <= (({(forvar508 - forvar485)} ?
                              forvar442[(1'h1):(1'h1)] : ({forvar413} >= reg529)) ?
                          (~|$unsigned($signed(forvar378))) : reg482);
                      reg544 <= {$unsigned(reg386)};
                      reg545 <= reg402;
                    end
                  if ($unsigned($unsigned($unsigned(reg516[(3'h4):(1'h0)]))))
                    begin
                      reg546 <= $signed((forvar520[(2'h3):(2'h3)] | reg434));
                      reg547 <= forvar509;
                    end
                  else
                    begin
                      reg546 <= reg426[(4'hb):(1'h1)];
                      reg547 <= ({reg375} + forvar442[(4'hc):(2'h2)]);
                      reg548 <= forvar359[(4'ha):(1'h1)];
                      reg549 <= reg548[(5'h10):(4'ha)];
                    end
                  if (reg468[(4'h8):(4'h8)])
                    begin
                      reg550 <= (&$signed({reg493[(1'h1):(1'h0)]}));
                      reg551 <= (((+(reg351 ?
                          reg311 : reg389)) || (~&{reg492})) & ((8'hb1) ?
                          $unsigned(reg385[(1'h0):(1'h0)]) : $unsigned((forvar517 >> reg375))));
                    end
                  else
                    begin
                      reg550 <= reg525;
                    end
                end
              for (forvar552 = (1'h0); (forvar552 < (2'h2)); forvar552 = (forvar552 + (1'h1)))
                begin
                  reg553 <= reg403;
                  for (forvar554 = (1'h0); (forvar554 < (2'h2)); forvar554 = (forvar554 + (1'h1)))
                    begin
                      reg555 <= $signed(reg411);
                    end
                  if ($signed(forvar493[(2'h2):(1'h0)]))
                    begin
                      reg556 <= ({(~^(reg330 ? reg493 : reg343))} ?
                          $signed($signed(reg460[(3'h5):(1'h1)])) : forvar517[(4'h8):(1'h1)]);
                      reg557 <= ((reg544 | (~$unsigned(reg487))) ?
                          forvar527[(2'h2):(2'h2)] : (8'hb8));
                      reg558 <= ((+(forvar467 << $unsigned(forvar529))) == reg330[(3'h6):(3'h6)]);
                      reg559 <= (forvar359 ?
                          ((8'hb7) ?
                              $unsigned({forvar485}) : $signed((reg491 ?
                                  reg368 : (8'hba)))) : (forvar482 ?
                              reg461[(2'h3):(1'h1)] : ((reg398 * reg383) ?
                                  (reg552 ?
                                      forvar400 : forvar472) : $signed(reg298))));
                    end
                  else
                    begin
                      reg556 <= $unsigned(reg357);
                    end
                  reg560 <= $unsigned(((~(8'ha7)) ?
                      {(~|reg431)} : $signed({reg307})));
                end
              reg561 <= ((~($signed((8'hb4)) ?
                      $unsigned(forvar364) : forvar492[(1'h0):(1'h0)])) ?
                  $signed((^~(reg487 << reg525))) : ($unsigned((reg355 || (8'had))) ?
                      $unsigned((reg559 ^ forvar544)) : $unsigned(forvar534)));
              for (forvar562 = (1'h0); (forvar562 < (2'h3)); forvar562 = (forvar562 + (1'h1)))
                begin
                  for (forvar563 = (1'h0); (forvar563 < (2'h2)); forvar563 = (forvar563 + (1'h1)))
                    begin
                      reg564 <= ((+reg314[(3'h5):(2'h2)]) ?
                          $unsigned($signed((forvar406 < forvar479))) : $unsigned($signed((reg486 ?
                              reg345 : (8'hac)))));
                      reg565 <= $signed((~|({reg535} - (reg441 == forvar512))));
                      reg566 <= forvar396;
                    end
                  reg567 <= (~^reg471[(3'h7):(2'h2)]);
                end
            end
          else
            begin
              if (((|$unsigned(reg550[(1'h0):(1'h0)])) + (^$signed((reg441 == (8'h9e))))))
                begin
                  for (forvar541 = (1'h0); (forvar541 < (2'h2)); forvar541 = (forvar541 + (1'h1)))
                    begin
                      reg542 <= (reg414 ?
                          (forvar503 ?
                              (!((8'ha3) ? (8'h9d) : (8'h9e))) : ((forvar554 ?
                                  forvar421 : forvar351) ^~ (!reg401))) : reg296);
                      reg543 <= ((reg457[(4'h9):(1'h0)] != (^~(~reg476))) != reg314[(1'h0):(1'h0)]);
                    end
                  for (forvar544 = (1'h0); (forvar544 < (1'h0)); forvar544 = (forvar544 + (1'h1)))
                    begin
                      reg545 <= $unsigned(((&reg441[(4'h8):(1'h1)]) | forvar482));
                    end
                end
              else
                begin
                  if ((+(((|(8'h9f)) ?
                          (forvar329 ~^ reg547) : $unsigned((8'haa))) ?
                      reg502 : forvar508[(2'h3):(2'h2)])))
                    begin
                      reg541 <= (~&(((~|forvar517) ^~ (reg298 ?
                          (8'hb8) : reg386)) * ((!reg496) ?
                          reg350[(2'h2):(1'h1)] : $signed(reg560))));
                      reg542 <= reg439[(3'h4):(1'h0)];
                      reg543 <= $unsigned(forvar537[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg541 <= (($unsigned((forvar482 ? reg300 : reg326)) ?
                              $signed(((8'h9c) << (8'hb1))) : $unsigned(((8'ha1) <<< (8'ha3)))) ?
                          {reg390[(3'h6):(1'h0)]} : wire289);
                      reg542 <= reg358[(2'h2):(1'h1)];
                      reg543 <= ((((reg466 ?
                              reg565 : reg358) == $unsigned(reg432)) ^ reg484) ?
                          reg361[(3'h5):(3'h4)] : $signed(((~^reg344) ?
                              reg438 : $unsigned(forvar422))));
                    end
                  for (forvar544 = (1'h0); (forvar544 < (2'h2)); forvar544 = (forvar544 + (1'h1)))
                    begin
                      reg545 <= (({forvar419} ~^ $signed((&reg478))) <<< wire292[(1'h1):(1'h1)]);
                      reg546 <= $unsigned((reg531 < reg466[(1'h0):(1'h0)]));
                      reg547 <= $signed((~$signed(reg545)));
                      reg548 <= $unsigned((($signed(forvar407) || (reg542 - reg565)) ?
                          $signed((reg297 ?
                              (8'hb0) : wire292)) : reg368[(5'h10):(4'hf)]));
                    end
                  for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
                    begin
                      reg550 <= ((~|((^~reg438) - ((8'haf) ?
                          reg495 : reg408))) << ($signed($signed((8'hab))) ?
                          (~&(~(8'hb6))) : $signed({reg530})));
                      reg551 <= $unsigned($unsigned(forvar542[(1'h0):(1'h0)]));
                    end
                  if ({reg567[(3'h7):(2'h2)]})
                    begin
                      reg552 <= (((~|(^~reg413)) || {{reg323}}) - reg319);
                      reg553 <= forvar501[(4'h8):(1'h0)];
                      reg554 <= $unsigned(($signed($unsigned(reg318)) < (^{reg439})));
                    end
                  else
                    begin
                      reg552 <= {(reg483[(2'h2):(2'h2)] ?
                              (reg326 == (forvar437 ?
                                  reg504 : forvar437)) : reg548[(3'h7):(3'h4)])};
                    end
                end
              for (forvar555 = (1'h0); (forvar555 < (2'h3)); forvar555 = (forvar555 + (1'h1)))
                begin
                  for (forvar556 = (1'h0); (forvar556 < (1'h0)); forvar556 = (forvar556 + (1'h1)))
                    begin
                      reg557 <= ((~^forvar424) ?
                          (((~^(8'hb9)) ?
                                  (forvar520 ?
                                      forvar523 : forvar556) : {(8'hb6)}) ?
                              $unsigned($signed(forvar452)) : (~|forvar477)) : ($signed((~forvar508)) ?
                              $signed((~reg443)) : (forvar556 ?
                                  {reg500} : reg352[(4'h8):(2'h2)])));
                    end
                end
              for (forvar558 = (1'h0); (forvar558 < (2'h2)); forvar558 = (forvar558 + (1'h1)))
                begin
                  if (reg383)
                    begin
                      reg559 <= (^(reg560[(3'h5):(2'h2)] && $signed((reg561 > (8'h9c)))));
                      reg560 <= forvar386[(4'h9):(3'h5)];
                      reg561 <= $unsigned((~$signed(reg350)));
                    end
                  else
                    begin
                      reg559 <= {$signed((!(+reg339)))};
                      reg560 <= ((~^(reg361[(3'h4):(2'h3)] <= (reg405 >>> reg522))) > reg475[(3'h7):(1'h1)]);
                      reg561 <= forvar537;
                    end
                  reg562 <= $unsigned(($signed($unsigned(reg376)) ^ (~^forvar413[(3'h5):(2'h3)])));
                  if ((((-$unsigned((8'hb6))) ?
                      reg374 : (!$signed((8'ha5)))) << (+((^~forvar481) ?
                      reg354 : (reg469 ? reg387 : (8'haa))))))
                    begin
                      reg563 <= reg410;
                    end
                  else
                    begin
                      reg563 <= reg494;
                      reg564 <= reg331[(2'h3):(2'h3)];
                      reg565 <= (~(8'hb6));
                      reg566 <= $signed((((!reg461) - (+forvar509)) ?
                          (~forvar468) : {(forvar454 < reg558)}));
                    end
                  for (forvar567 = (1'h0); (forvar567 < (1'h0)); forvar567 = (forvar567 + (1'h1)))
                    begin
                      reg568 <= reg469;
                      reg569 <= {reg470[(1'h1):(1'h1)]};
                      reg570 <= reg393[(4'he):(4'hc)];
                      reg571 <= (^~forvar543[(1'h0):(1'h0)]);
                    end
                end
            end
          for (forvar572 = (1'h0); (forvar572 < (2'h3)); forvar572 = (forvar572 + (1'h1)))
            begin
              for (forvar573 = (1'h0); (forvar573 < (2'h3)); forvar573 = (forvar573 + (1'h1)))
                begin
                  if ($unsigned($unsigned(forvar562[(2'h2):(2'h2)])))
                    begin
                      reg574 <= reg486;
                      reg575 <= (!$unsigned(forvar472));
                    end
                  else
                    begin
                      reg574 <= $unsigned($unsigned($signed((reg426 ?
                          reg356 : reg388))));
                      reg575 <= ($unsigned(reg384[(2'h2):(2'h2)]) ~^ $unsigned(($unsigned(reg408) + $unsigned(reg338))));
                      reg576 <= (-reg500[(3'h4):(2'h2)]);
                    end
                end
            end
        end
    end
  assign wire577 = ({reg494[(4'h8):(3'h7)]} ?
                       reg358[(4'h8):(4'h8)] : ($unsigned(reg300) ?
                           $unsigned((reg309 != forvar315)) : reg569[(2'h3):(2'h3)]));
  assign wire578 = (-(8'hb9));
  assign wire579 = (reg405 <= (^((reg343 ?
                       (8'hac) : reg564) > $signed(forvar543))));
  assign wire580 = (($signed((reg464 ? reg478 : (8'hb2))) ? reg440 : (8'hb6)) ?
                       reg521 : $unsigned((~(&forvar379))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module227
#(parameter param284 = (!(~(((8'hb2) ? (8'haf) : (8'hb7)) >> (^~(8'hb5))))))
(y, clk, wire231, wire230, wire229, wire228);
  output wire [(32'h1ff):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire231;
  input wire [(2'h3):(1'h0)] wire230;
  input wire signed [(3'h7):(1'h0)] wire229;
  input wire signed [(4'hb):(1'h0)] wire228;
  wire signed [(4'h8):(1'h0)] wire283;
  wire [(4'hf):(1'h0)] wire282;
  wire signed [(2'h2):(1'h0)] wire281;
  wire [(2'h2):(1'h0)] wire280;
  wire [(4'he):(1'h0)] wire279;
  wire signed [(3'h7):(1'h0)] wire278;
  wire [(5'h10):(1'h0)] wire277;
  reg signed [(4'h8):(1'h0)] reg276 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg258 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar257 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar252 = (1'h0);
  reg [(4'he):(1'h0)] reg256 = (1'h0);
  reg [(2'h2):(1'h0)] reg251 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg275 = (1'h0);
  reg [(4'ha):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg272 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar271 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg270 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar269 = (1'h0);
  reg [(4'h9):(1'h0)] reg268 = (1'h0);
  reg [(4'h8):(1'h0)] reg267 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg266 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg265 = (1'h0);
  reg [(4'h8):(1'h0)] forvar264 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg263 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg262 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg261 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg260 = (1'h0);
  reg [(4'hb):(1'h0)] reg259 = (1'h0);
  reg [(4'h9):(1'h0)] forvar258 = (1'h0);
  reg [(3'h5):(1'h0)] reg257 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar256 = (1'h0);
  reg [(3'h5):(1'h0)] reg255 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg254 = (1'h0);
  reg [(2'h3):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg252 = (1'h0);
  reg [(4'hb):(1'h0)] forvar251 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar250 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg241 = (1'h0);
  reg [(3'h4):(1'h0)] forvar240 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar234 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg249 = (1'h0);
  reg [(3'h7):(1'h0)] reg248 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg247 = (1'h0);
  reg [(4'hc):(1'h0)] reg246 = (1'h0);
  reg [(4'h9):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg244 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg243 = (1'h0);
  reg [(4'h8):(1'h0)] reg242 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar241 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg240 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg239 = (1'h0);
  reg [(2'h3):(1'h0)] reg238 = (1'h0);
  reg [(4'h8):(1'h0)] reg237 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg236 = (1'h0);
  reg [(3'h5):(1'h0)] forvar235 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg235 = (1'h0);
  reg signed [(4'he):(1'h0)] reg234 = (1'h0);
  wire [(3'h7):(1'h0)] wire233;
  wire [(3'h4):(1'h0)] wire232;
  assign y = {wire283,
                 wire282,
                 wire281,
                 wire280,
                 wire279,
                 wire278,
                 wire277,
                 reg276,
                 reg258,
                 forvar257,
                 forvar252,
                 reg256,
                 reg251,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 forvar271,
                 reg270,
                 forvar269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 forvar264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 forvar258,
                 reg257,
                 forvar256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 forvar251,
                 forvar250,
                 reg241,
                 forvar240,
                 forvar234,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 forvar241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 forvar235,
                 reg235,
                 reg234,
                 wire233,
                 wire232,
                 (1'h0)};
  assign wire232 = ({($signed(wire231) ~^ wire229[(2'h2):(2'h2)])} | (((wire229 == (8'ha0)) < wire230[(1'h0):(1'h0)]) ?
                       {(wire230 > wire231)} : wire228[(4'h8):(2'h3)]));
  assign wire233 = wire231[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      if ((wire228 ? wire232[(3'h4):(2'h2)] : wire229))
        begin
          reg234 <= ($unsigned($unsigned(wire231[(1'h0):(1'h0)])) ?
              {$unsigned((wire232 | wire228))} : (({wire229} && $unsigned(wire233)) > (+$signed(wire230))));
          if (wire233)
            begin
              reg235 <= {(wire229[(3'h4):(1'h0)] ~^ ((wire232 ?
                      wire232 : wire228) <<< $signed(wire230)))};
            end
          else
            begin
              for (forvar235 = (1'h0); (forvar235 < (2'h2)); forvar235 = (forvar235 + (1'h1)))
                begin
                  reg236 <= ((8'hb2) >>> wire229[(1'h0):(1'h0)]);
                  if (reg236)
                    begin
                      reg237 <= $signed(wire230);
                      reg238 <= (!reg235[(1'h1):(1'h0)]);
                      reg239 <= (($signed((reg234 ? reg238 : reg234)) ?
                          ({wire231} ?
                              (^~(8'hb3)) : (reg234 ?
                                  (8'hba) : reg234)) : {$unsigned(reg236)}) ^~ (|reg234[(1'h1):(1'h1)]));
                      reg240 <= reg236;
                    end
                  else
                    begin
                      reg237 <= $unsigned((forvar235 ?
                          (^(wire232 ^~ reg238)) : ($unsigned(wire231) - (wire231 ?
                              (8'hb8) : wire231))));
                      reg238 <= (~&wire230[(1'h1):(1'h1)]);
                      reg239 <= reg236;
                    end
                  for (forvar241 = (1'h0); (forvar241 < (2'h2)); forvar241 = (forvar241 + (1'h1)))
                    begin
                      reg242 <= (($unsigned((reg235 ? wire228 : (8'hb0))) ?
                              ({(8'hb4)} <<< (reg240 <<< forvar235)) : wire228) ?
                          $unsigned((-wire232[(2'h2):(1'h0)])) : ((-$signed(reg234)) ?
                              {(+reg240)} : wire230[(2'h2):(1'h0)]));
                      reg243 <= wire232[(3'h4):(1'h1)];
                      reg244 <= (8'hb7);
                    end
                  if ($signed($signed(((reg244 ?
                      reg239 : wire229) <= {(8'ha1)}))))
                    begin
                      reg245 <= $signed(wire230);
                      reg246 <= $unsigned($unsigned(((!reg242) ?
                          (wire233 * (8'ha2)) : $unsigned(forvar235))));
                      reg247 <= $signed(reg243[(3'h4):(1'h0)]);
                      reg248 <= $signed({wire233[(1'h1):(1'h1)]});
                    end
                  else
                    begin
                      reg245 <= (((reg234[(3'h6):(3'h4)] + $unsigned(wire230)) - (reg235[(1'h0):(1'h0)] ?
                              (reg239 ? reg240 : reg247) : (|wire232))) ?
                          $unsigned(((~(8'hb7)) ?
                              $unsigned((8'hb3)) : (forvar235 ?
                                  reg247 : reg247))) : (&((reg235 ?
                                  wire233 : reg239) ?
                              (reg245 ^~ reg242) : {wire232})));
                      reg246 <= (|$unsigned(reg248));
                    end
                end
            end
          reg249 <= ({forvar241[(3'h4):(1'h0)]} >= wire233);
        end
      else
        begin
          if ($unsigned({({reg244} ? (!reg245) : $unsigned((8'hb1)))}))
            begin
              if (reg243[(1'h1):(1'h0)])
                begin
                  if (($unsigned($signed($signed(wire231))) << $unsigned((^{wire229}))))
                    begin
                      reg234 <= $unsigned(((((8'ha8) ? wire229 : reg249) ?
                              (forvar241 | wire228) : {wire233}) ?
                          {(wire229 == (8'hb1))} : {wire230[(1'h0):(1'h0)]}));
                      reg235 <= (-{$signed((wire231 ? (8'haa) : reg235))});
                      reg236 <= $signed($unsigned({$signed(reg234)}));
                      reg237 <= (wire230 ?
                          reg236[(2'h2):(2'h2)] : ((((8'ha2) ?
                                  reg249 : reg236) >> (&(8'ha0))) ?
                              wire229 : (reg238[(1'h0):(1'h0)] ?
                                  ((8'hb7) && (8'hb8)) : (wire230 ?
                                      reg236 : reg238))));
                    end
                  else
                    begin
                      reg234 <= ((8'ha1) ?
                          (8'ha6) : (((wire233 < reg242) & wire228) ?
                              $unsigned((reg244 <<< forvar241)) : {reg235}));
                    end
                end
              else
                begin
                  for (forvar234 = (1'h0); (forvar234 < (2'h3)); forvar234 = (forvar234 + (1'h1)))
                    begin
                      reg235 <= ($unsigned(reg240) >> reg249[(2'h2):(1'h0)]);
                    end
                end
              reg238 <= reg248;
              reg239 <= {wire233};
            end
          else
            begin
              for (forvar234 = (1'h0); (forvar234 < (2'h3)); forvar234 = (forvar234 + (1'h1)))
                begin
                  reg235 <= (($signed(wire231) ~^ (^(-wire233))) ?
                      $unsigned(reg242) : {($signed(forvar241) ?
                              (wire228 ^ reg249) : $signed(reg243))});
                  if (((8'ha2) ?
                      $signed($signed($signed(reg235))) : $unsigned(reg236[(1'h0):(1'h0)])))
                    begin
                      reg236 <= reg246[(4'h8):(1'h1)];
                      reg237 <= wire231;
                      reg238 <= (~^(!{$signed(reg244)}));
                    end
                  else
                    begin
                      reg236 <= reg235[(1'h1):(1'h0)];
                      reg237 <= $signed(reg236);
                      reg238 <= (-reg234[(1'h0):(1'h0)]);
                    end
                end
              reg239 <= ((~^((^reg248) ?
                      (wire233 ? wire232 : reg242) : (reg240 ?
                          reg247 : wire230))) ?
                  (reg249 ?
                      $signed((reg236 ?
                          wire232 : (8'ha4))) : $unsigned(reg246[(2'h3):(2'h2)])) : reg247);
              if ((~|$unsigned($signed(wire231[(3'h4):(1'h0)]))))
                begin
                  reg240 <= reg246[(1'h1):(1'h0)];
                end
              else
                begin
                  for (forvar240 = (1'h0); (forvar240 < (1'h1)); forvar240 = (forvar240 + (1'h1)))
                    begin
                      reg241 <= wire228;
                    end
                  if (($unsigned(((!reg242) ?
                          (reg236 ? reg247 : reg246) : reg243)) ?
                      (((wire230 + reg243) ?
                          (+wire232) : reg241[(1'h0):(1'h0)]) >= reg237) : (reg240[(1'h1):(1'h0)] <= (^~reg244))))
                    begin
                      reg242 <= (^~$unsigned({(~&(8'ha5))}));
                      reg243 <= forvar240;
                    end
                  else
                    begin
                      reg242 <= {(reg240[(3'h5):(2'h3)] ? reg249 : reg244)};
                      reg243 <= (~^((^reg239[(3'h5):(2'h3)]) ?
                          (reg246 < $signed((8'hac))) : (reg241 ?
                              $unsigned(reg242) : (reg246 ?
                                  reg242 : wire229))));
                      reg244 <= (({$signed(reg243)} ?
                          (wire229 <<< (reg244 == (8'ha7))) : reg238[(2'h3):(1'h1)]) <= ({$unsigned((8'hb1))} ?
                          wire232[(2'h2):(1'h0)] : $signed(((8'hab) << wire233))));
                    end
                end
            end
        end
      for (forvar250 = (1'h0); (forvar250 < (2'h2)); forvar250 = (forvar250 + (1'h1)))
        begin
          if ($signed($unsigned($unsigned((+reg244)))))
            begin
              for (forvar251 = (1'h0); (forvar251 < (1'h1)); forvar251 = (forvar251 + (1'h1)))
                begin
                  reg252 <= forvar240[(2'h2):(2'h2)];
                end
              if (reg239)
                begin
                  if ((({(forvar234 ^~ wire228)} < $signed(reg246)) != (reg247 ?
                      ({reg234} ?
                          (reg249 ? reg238 : forvar240) : (reg240 ?
                              forvar250 : wire230)) : ({forvar241} ?
                          (&reg248) : (reg242 && reg249)))))
                    begin
                      reg253 <= forvar250;
                    end
                  else
                    begin
                      reg253 <= $unsigned((((forvar234 ?
                          reg247 : reg245) * (reg245 ?
                          reg252 : reg239)) ^ reg238[(2'h2):(1'h0)]));
                      reg254 <= reg236[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  if ($unsigned((8'had)))
                    begin
                      reg253 <= (~&{$unsigned(reg237)});
                      reg254 <= ({((+(8'ha5)) & reg236)} > $unsigned(forvar234));
                    end
                  else
                    begin
                      reg253 <= ($unsigned(wire229) <<< {$signed(reg237[(4'h8):(2'h3)])});
                      reg254 <= $signed($unsigned(forvar250[(3'h4):(3'h4)]));
                      reg255 <= reg234[(4'he):(4'ha)];
                    end
                  for (forvar256 = (1'h0); (forvar256 < (2'h3)); forvar256 = (forvar256 + (1'h1)))
                    begin
                      reg257 <= $unsigned(reg240[(4'ha):(1'h0)]);
                    end
                end
              for (forvar258 = (1'h0); (forvar258 < (1'h1)); forvar258 = (forvar258 + (1'h1)))
                begin
                  reg259 <= $unsigned(reg243[(1'h0):(1'h0)]);
                  reg260 <= ((^~((reg241 ?
                      reg254 : (8'ha7)) || forvar241[(4'h8):(3'h5)])) & $unsigned($signed($signed(reg244))));
                  if (reg237[(3'h4):(2'h3)])
                    begin
                      reg261 <= (~^(!$unsigned({(8'hb6)})));
                    end
                  else
                    begin
                      reg261 <= (~$signed($unsigned((forvar256 == (8'ha5)))));
                      reg262 <= ($signed({forvar234}) ~^ (~|($signed(reg237) ^ ((8'hb6) ?
                          reg234 : forvar240))));
                    end
                  reg263 <= (~^reg257[(1'h1):(1'h1)]);
                end
              for (forvar264 = (1'h0); (forvar264 < (1'h0)); forvar264 = (forvar264 + (1'h1)))
                begin
                  if ($unsigned((reg246 && $unsigned(reg238[(2'h2):(2'h2)]))))
                    begin
                      reg265 <= {reg260[(3'h5):(3'h5)]};
                      reg266 <= ({$unsigned((reg241 >> forvar240))} <= ((|(reg244 > reg252)) >= reg238));
                      reg267 <= (~^{$unsigned(reg243[(1'h0):(1'h0)])});
                      reg268 <= wire230[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg265 <= ($unsigned(reg268[(4'h8):(3'h4)]) ?
                          reg260[(3'h5):(3'h4)] : wire229);
                      reg266 <= ((reg255 > $signed((reg260 ?
                          wire230 : reg265))) >> $unsigned((reg243[(3'h4):(3'h4)] * (reg268 ?
                          reg267 : wire231))));
                      reg267 <= $signed((&((forvar264 ?
                          forvar241 : forvar241) * (reg260 ?
                          reg262 : reg246))));
                    end
                  for (forvar269 = (1'h0); (forvar269 < (2'h3)); forvar269 = (forvar269 + (1'h1)))
                    begin
                      reg270 <= $unsigned($unsigned((forvar264 ?
                          reg239 : (wire230 ^~ reg241))));
                    end
                  for (forvar271 = (1'h0); (forvar271 < (1'h1)); forvar271 = (forvar271 + (1'h1)))
                    begin
                      reg272 <= (($signed((reg235 ?
                              (8'ha4) : reg249)) && $signed($unsigned((8'hb2)))) ?
                          (^(reg234[(4'he):(4'h8)] ^ (reg263 ?
                              reg255 : reg248))) : {($signed(forvar256) ?
                                  (&reg235) : wire228[(3'h7):(3'h7)])});
                      reg273 <= forvar234[(1'h1):(1'h0)];
                      reg274 <= $signed(forvar264[(2'h2):(1'h0)]);
                      reg275 <= forvar264;
                    end
                end
            end
          else
            begin
              reg251 <= {$signed(reg275[(1'h1):(1'h1)])};
              if ((|$unsigned(reg243[(2'h3):(2'h3)])))
                begin
                  reg252 <= $unsigned(forvar241[(1'h1):(1'h0)]);
                  reg253 <= (($unsigned($signed(reg275)) == $signed((&(8'ha0)))) + $signed($unsigned($signed(reg257))));
                  if ((reg241[(2'h2):(2'h2)] ?
                      ((|(wire230 ?
                          (8'hb5) : forvar241)) | (~^reg234[(1'h0):(1'h0)])) : $signed(({(8'hac)} ?
                          $unsigned(reg251) : $signed(reg236)))))
                    begin
                      reg254 <= {(-(reg239 >> {forvar256}))};
                    end
                  else
                    begin
                      reg254 <= (reg238 ?
                          (wire233[(2'h2):(2'h2)] & (~(reg241 ?
                              reg254 : reg255))) : reg245[(3'h7):(1'h1)]);
                      reg255 <= $unsigned((($signed(reg257) >> reg251) ~^ {(reg253 ?
                              (8'hac) : reg255)}));
                      reg256 <= (-reg273[(2'h3):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar252 = (1'h0); (forvar252 < (1'h1)); forvar252 = (forvar252 + (1'h1)))
                    begin
                      reg253 <= $signed($signed(((reg251 <= reg272) ?
                          $unsigned(forvar251) : reg262[(4'h9):(3'h6)])));
                    end
                  if (reg244)
                    begin
                      reg254 <= (reg246[(3'h4):(2'h2)] >= (~$signed({reg246})));
                      reg255 <= (^forvar251);
                    end
                  else
                    begin
                      reg254 <= $signed((wire230[(2'h2):(1'h0)] * reg241));
                    end
                  reg256 <= $unsigned((~|reg243));
                  for (forvar257 = (1'h0); (forvar257 < (2'h2)); forvar257 = (forvar257 + (1'h1)))
                    begin
                      reg258 <= reg263[(4'hb):(3'h7)];
                      reg259 <= $unsigned(($signed((reg247 ?
                              reg274 : wire232)) ?
                          (-reg275[(3'h7):(3'h4)]) : ((forvar256 && reg270) ?
                              (^~forvar256) : reg256)));
                    end
                end
            end
          reg276 <= $signed((^($signed(wire230) <= (!reg246))));
        end
    end
  assign wire277 = $unsigned(reg256[(2'h2):(1'h0)]);
  assign wire278 = ({reg245[(4'h9):(2'h2)]} ~^ forvar264);
  assign wire279 = {{reg247[(2'h2):(1'h0)]}};
  assign wire280 = $signed(($unsigned($unsigned(reg256)) - ($signed(forvar251) ?
                       {reg259} : (|reg259))));
  assign wire281 = (8'had);
  assign wire282 = reg246[(4'h8):(3'h4)];
  assign wire283 = (reg244[(2'h3):(1'h1)] ?
                       (wire233 ^ reg270) : (~|reg254[(1'h1):(1'h1)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1923  (y, clk, wire1928, wire1927, wire1926, wire1925, wire1924);
  output wire [(32'h1f4f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h8):(1'h0)] wire1928;
  input wire signed [(4'ha):(1'h0)] wire1927;
  input wire signed [(3'h5):(1'h0)] wire1926;
  input wire signed [(3'h5):(1'h0)] wire1925;
  input wire [(3'h7):(1'h0)] wire1924;
  wire [(2'h2):(1'h0)] wire2666;
  wire [(2'h3):(1'h0)] wire2665;
  wire [(4'h9):(1'h0)] wire2664;
  wire signed [(3'h6):(1'h0)] wire2663;
  wire signed [(4'h9):(1'h0)] wire2662;
  wire [(3'h5):(1'h0)] wire2661;
  wire signed [(3'h7):(1'h0)] wire2660;
  reg [(3'h5):(1'h0)] reg2659 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2658 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2657 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2656 = (1'h0);
  reg [(4'h9):(1'h0)] reg2655 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2654 = (1'h0);
  reg [(4'hd):(1'h0)] reg2653 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2652 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2651 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2639 = (1'h0);
  reg [(3'h4):(1'h0)] reg2650 = (1'h0);
  reg [(3'h4):(1'h0)] reg2649 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2648 = (1'h0);
  reg [(4'hd):(1'h0)] reg2647 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2646 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2645 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2644 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2643 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2642 = (1'h0);
  reg [(5'h10):(1'h0)] reg2641 = (1'h0);
  reg [(3'h5):(1'h0)] reg2640 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2639 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2638 = (1'h0);
  reg [(4'hd):(1'h0)] reg2630 = (1'h0);
  reg [(3'h7):(1'h0)] reg2637 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2636 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2635 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2634 = (1'h0);
  reg [(4'he):(1'h0)] reg2633 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2632 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2631 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2630 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2629 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2628 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2627 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2626 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2625 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2624 = (1'h0);
  reg [(3'h6):(1'h0)] reg2623 = (1'h0);
  reg [(3'h7):(1'h0)] reg2622 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2621 = (1'h0);
  reg [(3'h5):(1'h0)] reg2620 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2618 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2619 = (1'h0);
  reg [(3'h4):(1'h0)] reg2618 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2617 = (1'h0);
  reg [(4'hf):(1'h0)] reg2616 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2613 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2615 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2614 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2613 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2612 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2611 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2610 = (1'h0);
  reg [(3'h5):(1'h0)] reg2609 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2608 = (1'h0);
  reg [(5'h10):(1'h0)] reg2607 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2606 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2605 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2604 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2603 = (1'h0);
  reg [(4'hd):(1'h0)] reg2602 = (1'h0);
  reg [(5'h10):(1'h0)] reg2601 = (1'h0);
  reg [(4'hb):(1'h0)] reg2600 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2599 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2598 = (1'h0);
  reg [(4'hf):(1'h0)] reg2597 = (1'h0);
  reg [(4'hc):(1'h0)] reg2596 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2595 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2594 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2593 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2592 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2591 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2589 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2587 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2586 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2585 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2584 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2583 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2578 = (1'h0);
  reg [(3'h5):(1'h0)] reg2575 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2590 = (1'h0);
  reg [(4'hf):(1'h0)] reg2589 = (1'h0);
  reg [(3'h4):(1'h0)] reg2588 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2587 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2586 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2585 = (1'h0);
  reg [(4'hd):(1'h0)] reg2584 = (1'h0);
  reg [(3'h4):(1'h0)] reg2581 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2577 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2576 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2583 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2582 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2581 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2580 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2579 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2578 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2577 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2576 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2575 = (1'h0);
  reg [(4'h9):(1'h0)] reg2574 = (1'h0);
  reg [(5'h10):(1'h0)] reg2573 = (1'h0);
  reg [(2'h2):(1'h0)] reg2572 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2571 = (1'h0);
  reg [(2'h2):(1'h0)] reg2570 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2569 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2568 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2567 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2566 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2565 = (1'h0);
  reg [(4'hb):(1'h0)] reg2564 = (1'h0);
  reg [(2'h2):(1'h0)] reg2563 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2562 = (1'h0);
  reg [(4'he):(1'h0)] reg2561 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2560 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2559 = (1'h0);
  reg [(4'hc):(1'h0)] reg2558 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2557 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2556 = (1'h0);
  reg [(4'hf):(1'h0)] reg2555 = (1'h0);
  reg [(2'h3):(1'h0)] reg2554 = (1'h0);
  reg [(3'h4):(1'h0)] reg2553 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2552 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2551 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2550 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2539 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2549 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2548 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2547 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2546 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2545 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2544 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2543 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2542 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2541 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2540 = (1'h0);
  reg [(4'hb):(1'h0)] reg2539 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2538 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2537 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2536 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2531 = (1'h0);
  reg [(5'h10):(1'h0)] reg2528 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2527 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2536 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2535 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2534 = (1'h0);
  reg [(3'h5):(1'h0)] reg2533 = (1'h0);
  reg [(4'he):(1'h0)] reg2532 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2531 = (1'h0);
  reg [(4'hc):(1'h0)] reg2530 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2529 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2528 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2527 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2526 = (1'h0);
  reg [(4'he):(1'h0)] reg2523 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2519 = (1'h0);
  reg [(2'h3):(1'h0)] reg2518 = (1'h0);
  reg [(3'h7):(1'h0)] reg2525 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2524 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2523 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2522 = (1'h0);
  reg [(2'h2):(1'h0)] reg2521 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2520 = (1'h0);
  reg [(3'h5):(1'h0)] reg2519 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2518 = (1'h0);
  reg [(3'h5):(1'h0)] reg2517 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2516 = (1'h0);
  reg [(4'hd):(1'h0)] reg2515 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2514 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2513 = (1'h0);
  reg [(4'ha):(1'h0)] reg2512 = (1'h0);
  reg [(3'h4):(1'h0)] reg2476 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2475 = (1'h0);
  reg [(2'h2):(1'h0)] reg2472 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2471 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2467 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2511 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2510 = (1'h0);
  reg [(4'hd):(1'h0)] reg2509 = (1'h0);
  reg [(2'h2):(1'h0)] reg2508 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2507 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2506 = (1'h0);
  reg [(5'h10):(1'h0)] reg2505 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2504 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2503 = (1'h0);
  reg [(2'h2):(1'h0)] reg2502 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2501 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2500 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2499 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2498 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2497 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2496 = (1'h0);
  reg [(3'h6):(1'h0)] reg2495 = (1'h0);
  reg [(4'hf):(1'h0)] reg2494 = (1'h0);
  reg [(4'h9):(1'h0)] reg2493 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2492 = (1'h0);
  reg [(4'ha):(1'h0)] reg2491 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2489 = (1'h0);
  reg [(3'h5):(1'h0)] reg2487 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2490 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2489 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2488 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2487 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2486 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2485 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2484 = (1'h0);
  reg [(4'h8):(1'h0)] reg2483 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2482 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2481 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2480 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2479 = (1'h0);
  reg [(3'h4):(1'h0)] reg2478 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2477 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2476 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2475 = (1'h0);
  reg [(4'hf):(1'h0)] reg2474 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2473 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2472 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2471 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2470 = (1'h0);
  reg [(4'hd):(1'h0)] reg2469 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2468 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2467 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2466 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire2465;
  reg signed [(2'h2):(1'h0)] reg2464 = (1'h0);
  reg [(2'h3):(1'h0)] reg2463 = (1'h0);
  reg [(4'hb):(1'h0)] reg2462 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2461 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2460 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2459 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2458 = (1'h0);
  reg [(5'h10):(1'h0)] reg2457 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2456 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2451 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2448 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2446 = (1'h0);
  reg [(4'he):(1'h0)] forvar2440 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2450 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2441 = (1'h0);
  reg [(2'h3):(1'h0)] reg2456 = (1'h0);
  reg [(4'hb):(1'h0)] reg2455 = (1'h0);
  reg [(5'h10):(1'h0)] reg2454 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2453 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2452 = (1'h0);
  reg [(5'h10):(1'h0)] reg2451 = (1'h0);
  reg [(5'h10):(1'h0)] reg2450 = (1'h0);
  reg [(4'ha):(1'h0)] reg2449 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2448 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2447 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2446 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2445 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2444 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2443 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2442 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2441 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2440 = (1'h0);
  reg [(4'h9):(1'h0)] reg2439 = (1'h0);
  reg [(5'h10):(1'h0)] reg2436 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2434 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2432 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2431 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2430 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2426 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2425 = (1'h0);
  reg [(3'h4):(1'h0)] reg2413 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2410 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2407 = (1'h0);
  reg [(4'h8):(1'h0)] reg2395 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2402 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2399 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2394 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2392 = (1'h0);
  reg [(2'h2):(1'h0)] reg2387 = (1'h0);
  reg [(4'h9):(1'h0)] reg2383 = (1'h0);
  reg [(4'hf):(1'h0)] reg2438 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2414 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2428 = (1'h0);
  reg [(4'hb):(1'h0)] reg2437 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2436 = (1'h0);
  reg [(3'h5):(1'h0)] reg2435 = (1'h0);
  reg [(4'h9):(1'h0)] reg2434 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2433 = (1'h0);
  reg [(2'h3):(1'h0)] reg2432 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2431 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2430 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2429 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2428 = (1'h0);
  reg [(4'h9):(1'h0)] reg2427 = (1'h0);
  reg [(2'h2):(1'h0)] reg2426 = (1'h0);
  reg [(3'h5):(1'h0)] reg2425 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2422 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2420 = (1'h0);
  reg [(4'h8):(1'h0)] reg2418 = (1'h0);
  reg [(3'h7):(1'h0)] reg2416 = (1'h0);
  reg [(4'hb):(1'h0)] reg2424 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2423 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2422 = (1'h0);
  reg [(5'h10):(1'h0)] reg2421 = (1'h0);
  reg [(2'h2):(1'h0)] reg2420 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2419 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2418 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2417 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2416 = (1'h0);
  reg [(4'h8):(1'h0)] reg2415 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2414 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2413 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2409 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2404 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2412 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2411 = (1'h0);
  reg [(3'h7):(1'h0)] reg2410 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2409 = (1'h0);
  reg [(3'h6):(1'h0)] reg2408 = (1'h0);
  reg [(4'hf):(1'h0)] reg2407 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2406 = (1'h0);
  reg [(4'hc):(1'h0)] reg2405 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2404 = (1'h0);
  reg [(4'hb):(1'h0)] reg2403 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2402 = (1'h0);
  reg [(2'h3):(1'h0)] reg2401 = (1'h0);
  reg [(2'h3):(1'h0)] reg2400 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2399 = (1'h0);
  reg [(5'h10):(1'h0)] reg2398 = (1'h0);
  reg [(2'h3):(1'h0)] reg2397 = (1'h0);
  reg [(4'h9):(1'h0)] reg2396 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2395 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2394 = (1'h0);
  reg [(3'h7):(1'h0)] reg2393 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2392 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2391 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2390 = (1'h0);
  reg [(4'ha):(1'h0)] reg2389 = (1'h0);
  reg [(4'hb):(1'h0)] reg2388 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2387 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2386 = (1'h0);
  reg [(3'h5):(1'h0)] reg2385 = (1'h0);
  reg [(2'h2):(1'h0)] reg2384 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2383 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2382 = (1'h0);
  reg [(4'h9):(1'h0)] reg2373 = (1'h0);
  reg [(4'he):(1'h0)] forvar2371 = (1'h0);
  reg [(4'h9):(1'h0)] reg2381 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2380 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2379 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2370 = (1'h0);
  reg [(3'h5):(1'h0)] reg2378 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2377 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2376 = (1'h0);
  reg [(3'h5):(1'h0)] reg2375 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2374 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2373 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2372 = (1'h0);
  reg [(3'h6):(1'h0)] reg2371 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2370 = (1'h0);
  reg [(4'h9):(1'h0)] reg2369 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2368 = (1'h0);
  reg [(3'h5):(1'h0)] reg2367 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2366 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2365 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2364 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2363 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2362 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2361 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2352 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2351 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2349 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2348 = (1'h0);
  reg [(4'hc):(1'h0)] reg2346 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2359 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2357 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2355 = (1'h0);
  reg [(2'h3):(1'h0)] reg2354 = (1'h0);
  reg [(4'hf):(1'h0)] reg2360 = (1'h0);
  reg [(4'he):(1'h0)] reg2359 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2358 = (1'h0);
  reg [(3'h7):(1'h0)] reg2357 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2356 = (1'h0);
  reg [(3'h6):(1'h0)] reg2355 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2354 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2353 = (1'h0);
  reg [(4'he):(1'h0)] reg2352 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2351 = (1'h0);
  reg [(3'h7):(1'h0)] reg2350 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2349 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2348 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2347 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2346 = (1'h0);
  reg [(4'h8):(1'h0)] reg2345 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2344 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2343 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2339 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2335 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2342 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2341 = (1'h0);
  reg [(3'h6):(1'h0)] reg2340 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2339 = (1'h0);
  reg [(4'hf):(1'h0)] reg2338 = (1'h0);
  reg [(3'h4):(1'h0)] reg2337 = (1'h0);
  reg [(3'h7):(1'h0)] reg2336 = (1'h0);
  reg [(4'hf):(1'h0)] reg2335 = (1'h0);
  reg [(3'h7):(1'h0)] reg2334 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2333 = (1'h0);
  reg [(4'hf):(1'h0)] reg2332 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2331 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2330 = (1'h0);
  reg [(4'he):(1'h0)] reg2329 = (1'h0);
  reg [(4'hc):(1'h0)] reg2328 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2327 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2326 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2325 = (1'h0);
  reg [(4'ha):(1'h0)] reg2324 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2323 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2322 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2321 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2320 = (1'h0);
  reg [(4'h8):(1'h0)] reg2319 = (1'h0);
  reg [(3'h6):(1'h0)] reg2318 = (1'h0);
  reg [(4'ha):(1'h0)] reg2317 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2316 = (1'h0);
  reg [(4'hb):(1'h0)] reg2315 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2314 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2313 = (1'h0);
  reg [(4'hc):(1'h0)] reg2312 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2311 = (1'h0);
  reg [(2'h3):(1'h0)] reg2310 = (1'h0);
  reg [(4'he):(1'h0)] reg2309 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2308 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2307 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2306 = (1'h0);
  reg [(3'h7):(1'h0)] reg2305 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2304 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2303 = (1'h0);
  reg [(4'he):(1'h0)] forvar2301 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2283 = (1'h0);
  reg [(4'ha):(1'h0)] reg2276 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2296 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2293 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2289 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2287 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2285 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2282 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2280 = (1'h0);
  reg [(3'h5):(1'h0)] reg2279 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2275 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2302 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2298 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2295 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2290 = (1'h0);
  reg [(4'ha):(1'h0)] reg2301 = (1'h0);
  reg [(5'h10):(1'h0)] reg2300 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2299 = (1'h0);
  reg [(4'hd):(1'h0)] reg2298 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2297 = (1'h0);
  reg [(4'h9):(1'h0)] reg2296 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2295 = (1'h0);
  reg [(3'h7):(1'h0)] reg2294 = (1'h0);
  reg [(4'hf):(1'h0)] reg2293 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2292 = (1'h0);
  reg [(5'h10):(1'h0)] reg2291 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2290 = (1'h0);
  reg [(5'h10):(1'h0)] reg2289 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2288 = (1'h0);
  reg [(4'ha):(1'h0)] reg2287 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2286 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2285 = (1'h0);
  reg [(4'h8):(1'h0)] reg2284 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2283 = (1'h0);
  reg [(4'hf):(1'h0)] reg2282 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2281 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2280 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2279 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2278 = (1'h0);
  reg [(4'h8):(1'h0)] reg2277 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2276 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2275 = (1'h0);
  reg [(4'hf):(1'h0)] reg2274 = (1'h0);
  reg [(4'he):(1'h0)] reg2273 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2270 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2272 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2271 = (1'h0);
  reg [(3'h5):(1'h0)] reg2270 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2269 = (1'h0);
  reg [(4'ha):(1'h0)] reg2269 = (1'h0);
  reg [(2'h3):(1'h0)] reg2268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2267 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2266 = (1'h0);
  reg [(4'he):(1'h0)] reg2265 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2264 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2263 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2262 = (1'h0);
  reg [(2'h3):(1'h0)] reg2261 = (1'h0);
  reg [(3'h5):(1'h0)] reg2260 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2259 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2257 = (1'h0);
  reg [(3'h4):(1'h0)] reg2256 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2255 = (1'h0);
  reg [(2'h2):(1'h0)] reg2254 = (1'h0);
  reg [(4'he):(1'h0)] reg2253 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2252 = (1'h0);
  reg [(4'hd):(1'h0)] reg2251 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2250 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2249 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2248 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2247 = (1'h0);
  reg [(4'h8):(1'h0)] reg2246 = (1'h0);
  reg [(2'h3):(1'h0)] reg2245 = (1'h0);
  reg [(2'h3):(1'h0)] reg2244 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2243 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2242 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2241 = (1'h0);
  reg [(4'h9):(1'h0)] reg2240 = (1'h0);
  reg [(4'he):(1'h0)] reg2239 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2238 = (1'h0);
  reg [(4'h8):(1'h0)] reg2237 = (1'h0);
  reg [(3'h6):(1'h0)] reg2236 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2235 = (1'h0);
  reg [(4'hd):(1'h0)] reg2234 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2233 = (1'h0);
  reg [(2'h2):(1'h0)] reg2232 = (1'h0);
  reg [(3'h7):(1'h0)] reg2231 = (1'h0);
  reg [(3'h7):(1'h0)] reg2230 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2229 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2228 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2164 = (1'h0);
  reg [(4'hb):(1'h0)] reg2227 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2226 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2225 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2224 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2220 = (1'h0);
  reg [(3'h5):(1'h0)] reg2223 = (1'h0);
  reg [(4'h8):(1'h0)] reg2222 = (1'h0);
  reg [(2'h3):(1'h0)] reg2221 = (1'h0);
  reg [(4'h8):(1'h0)] reg2220 = (1'h0);
  reg [(5'h10):(1'h0)] reg2219 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2218 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2217 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2216 = (1'h0);
  reg [(3'h7):(1'h0)] reg2215 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2214 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2213 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2212 = (1'h0);
  reg [(4'hc):(1'h0)] reg2211 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2210 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2209 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2208 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2205 = (1'h0);
  reg [(4'h9):(1'h0)] reg2201 = (1'h0);
  reg [(3'h6):(1'h0)] reg2207 = (1'h0);
  reg [(4'he):(1'h0)] reg2206 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2205 = (1'h0);
  reg [(2'h3):(1'h0)] reg2204 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2203 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2202 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2201 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2200 = (1'h0);
  reg [(2'h3):(1'h0)] reg2199 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2198 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2197 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2196 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2195 = (1'h0);
  reg [(3'h6):(1'h0)] reg2194 = (1'h0);
  reg [(4'he):(1'h0)] reg2193 = (1'h0);
  reg [(4'hb):(1'h0)] reg2192 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2191 = (1'h0);
  reg [(4'h8):(1'h0)] reg2190 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2189 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2187 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2182 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2179 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2177 = (1'h0);
  reg [(4'hc):(1'h0)] reg2174 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2173 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2172 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2168 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2167 = (1'h0);
  reg [(5'h10):(1'h0)] reg2166 = (1'h0);
  reg [(3'h5):(1'h0)] reg2163 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2162 = (1'h0);
  reg [(3'h4):(1'h0)] reg2188 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2187 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2186 = (1'h0);
  reg [(2'h3):(1'h0)] reg2185 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2183 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2182 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2181 = (1'h0);
  reg [(4'h8):(1'h0)] reg2180 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2179 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2178 = (1'h0);
  reg [(4'hd):(1'h0)] reg2177 = (1'h0);
  reg [(3'h7):(1'h0)] reg2176 = (1'h0);
  reg [(4'he):(1'h0)] reg2175 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2174 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2173 = (1'h0);
  reg [(4'h9):(1'h0)] reg2172 = (1'h0);
  reg [(4'h8):(1'h0)] reg2171 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2170 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2169 = (1'h0);
  reg [(3'h6):(1'h0)] reg2168 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2167 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2166 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2165 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2164 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2163 = (1'h0);
  reg [(3'h5):(1'h0)] reg2162 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2161 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2160 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2159 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2158 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2157 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2156 = (1'h0);
  reg [(4'hf):(1'h0)] reg2155 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2154 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2153 = (1'h0);
  reg [(3'h5):(1'h0)] reg2152 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2151 = (1'h0);
  reg [(4'hc):(1'h0)] reg2150 = (1'h0);
  reg [(4'h8):(1'h0)] reg2149 = (1'h0);
  reg [(4'hf):(1'h0)] reg2148 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2147 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2146 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2145 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2144 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2143 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2142 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2141 = (1'h0);
  reg [(3'h5):(1'h0)] reg2140 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2139 = (1'h0);
  reg [(3'h5):(1'h0)] reg2138 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2137 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2136 = (1'h0);
  reg [(3'h5):(1'h0)] reg2135 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2134 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2133 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2132 = (1'h0);
  reg [(4'h9):(1'h0)] reg2128 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2127 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2126 = (1'h0);
  reg [(4'hb):(1'h0)] reg2131 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2130 = (1'h0);
  reg [(3'h4):(1'h0)] reg2129 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2128 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2127 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2126 = (1'h0);
  reg [(3'h7):(1'h0)] reg2119 = (1'h0);
  reg [(3'h4):(1'h0)] reg2125 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2124 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2123 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2122 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2121 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2120 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2119 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2118 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2117 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2116 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2115 = (1'h0);
  reg [(4'he):(1'h0)] reg2114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2113 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2112 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2111 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2103 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2102 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2110 = (1'h0);
  reg [(4'hd):(1'h0)] reg2109 = (1'h0);
  reg [(2'h3):(1'h0)] reg2108 = (1'h0);
  reg [(4'ha):(1'h0)] reg2107 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2106 = (1'h0);
  reg [(2'h3):(1'h0)] reg2105 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2104 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2103 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2102 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2101 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2100 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2099 = (1'h0);
  reg [(4'hd):(1'h0)] reg2098 = (1'h0);
  reg [(4'h8):(1'h0)] reg2097 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2096 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2095 = (1'h0);
  reg [(2'h2):(1'h0)] reg2094 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2093 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2091 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2086 = (1'h0);
  reg [(3'h7):(1'h0)] reg2084 = (1'h0);
  reg [(4'hc):(1'h0)] reg2092 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2091 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2090 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2089 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2088 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2087 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2086 = (1'h0);
  reg [(3'h7):(1'h0)] reg2085 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2084 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2083 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2082 = (1'h0);
  reg [(4'hd):(1'h0)] reg2081 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2058 = (1'h0);
  reg [(4'hf):(1'h0)] reg2053 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2052 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2051 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2050 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2047 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2080 = (1'h0);
  reg [(4'hc):(1'h0)] reg2079 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2078 = (1'h0);
  reg [(4'h8):(1'h0)] reg2077 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2076 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2075 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2074 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2073 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2072 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2071 = (1'h0);
  reg [(4'hd):(1'h0)] reg2070 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2069 = (1'h0);
  reg [(3'h6):(1'h0)] reg2068 = (1'h0);
  reg [(2'h2):(1'h0)] reg2067 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2066 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2065 = (1'h0);
  reg [(3'h4):(1'h0)] reg2064 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2063 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2062 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2061 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2060 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2059 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2058 = (1'h0);
  reg [(5'h10):(1'h0)] reg2057 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2056 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2055 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2054 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2053 = (1'h0);
  reg [(4'he):(1'h0)] forvar2052 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2051 = (1'h0);
  reg [(4'hb):(1'h0)] reg2050 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2049 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2048 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2047 = (1'h0);
  reg [(4'h9):(1'h0)] reg2046 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2041 = (1'h0);
  reg [(3'h6):(1'h0)] reg2045 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2044 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2043 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2042 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2041 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2040 = (1'h0);
  reg [(3'h5):(1'h0)] reg2035 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2039 = (1'h0);
  reg [(3'h7):(1'h0)] reg2038 = (1'h0);
  reg [(4'h8):(1'h0)] reg2037 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2036 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2035 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2025 = (1'h0);
  reg [(3'h6):(1'h0)] reg2034 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2033 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2032 = (1'h0);
  reg [(4'ha):(1'h0)] reg2031 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2030 = (1'h0);
  reg [(4'h9):(1'h0)] reg2029 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2028 = (1'h0);
  reg [(2'h3):(1'h0)] reg2027 = (1'h0);
  reg [(4'hb):(1'h0)] reg2026 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2025 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2024 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2023 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2022 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2020 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2015 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2013 = (1'h0);
  reg [(4'h8):(1'h0)] reg2011 = (1'h0);
  reg [(4'h8):(1'h0)] reg2021 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2020 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2019 = (1'h0);
  reg [(5'h10):(1'h0)] reg2018 = (1'h0);
  reg [(2'h2):(1'h0)] reg2017 = (1'h0);
  reg [(3'h5):(1'h0)] reg2016 = (1'h0);
  reg [(4'hf):(1'h0)] reg2015 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2014 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2013 = (1'h0);
  reg [(3'h5):(1'h0)] reg2012 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2011 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2010 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2009 = (1'h0);
  reg [(4'he):(1'h0)] forvar2001 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2008 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2007 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2006 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2005 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2004 = (1'h0);
  reg [(2'h3):(1'h0)] reg2003 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2002 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2001 = (1'h0);
  reg [(2'h3):(1'h0)] reg2000 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1999 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1998 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1980 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1974 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1976 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1971 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1970 = (1'h0);
  reg [(4'hd):(1'h0)] reg1997 = (1'h0);
  reg [(4'hb):(1'h0)] reg1996 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1995 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1991 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1994 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1993 = (1'h0);
  reg [(4'hc):(1'h0)] reg1992 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1991 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1983 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1990 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1989 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1988 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1987 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1986 = (1'h0);
  reg [(2'h3):(1'h0)] reg1985 = (1'h0);
  reg [(4'hc):(1'h0)] reg1984 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1983 = (1'h0);
  reg [(5'h10):(1'h0)] reg1982 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1981 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1980 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1979 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1978 = (1'h0);
  reg [(3'h5):(1'h0)] reg1977 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1976 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1967 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1975 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1974 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1973 = (1'h0);
  reg [(3'h6):(1'h0)] reg1972 = (1'h0);
  reg [(5'h10):(1'h0)] reg1971 = (1'h0);
  reg [(4'hc):(1'h0)] reg1970 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1969 = (1'h0);
  reg [(4'hd):(1'h0)] reg1968 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1967 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1966 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1965 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1963 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1962 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1964 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1963 = (1'h0);
  reg [(4'hf):(1'h0)] reg1962 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1961 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1960 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1959 = (1'h0);
  reg [(3'h6):(1'h0)] reg1958 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1957 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1956 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1955 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1954 = (1'h0);
  reg [(4'h8):(1'h0)] reg1953 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1952 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1948 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1947 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1951 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1950 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1949 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1948 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1947 = (1'h0);
  reg [(4'h8):(1'h0)] reg1946 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1941 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1939 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1936 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1945 = (1'h0);
  reg [(4'he):(1'h0)] reg1944 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1943 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1942 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1941 = (1'h0);
  reg [(4'hf):(1'h0)] reg1938 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1934 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1933 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1931 = (1'h0);
  reg [(2'h3):(1'h0)] reg1940 = (1'h0);
  reg [(3'h4):(1'h0)] reg1939 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1938 = (1'h0);
  reg [(4'h9):(1'h0)] reg1937 = (1'h0);
  reg [(3'h5):(1'h0)] reg1936 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1935 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1934 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1933 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1932 = (1'h0);
  reg [(3'h7):(1'h0)] reg1931 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1930 = (1'h0);
  reg [(5'h10):(1'h0)] reg1929 = (1'h0);
  assign y = {wire2666,
                 wire2665,
                 wire2664,
                 wire2663,
                 wire2662,
                 wire2661,
                 wire2660,
                 reg2659,
                 forvar2658,
                 reg2657,
                 reg2656,
                 reg2655,
                 forvar2654,
                 reg2653,
                 reg2652,
                 forvar2651,
                 reg2639,
                 reg2650,
                 reg2649,
                 reg2648,
                 reg2647,
                 forvar2646,
                 reg2645,
                 reg2644,
                 reg2643,
                 reg2642,
                 reg2641,
                 reg2640,
                 forvar2639,
                 forvar2638,
                 reg2630,
                 reg2637,
                 reg2636,
                 reg2635,
                 reg2634,
                 reg2633,
                 reg2632,
                 reg2631,
                 forvar2630,
                 reg2629,
                 forvar2628,
                 reg2627,
                 reg2626,
                 reg2625,
                 forvar2624,
                 reg2623,
                 reg2622,
                 reg2621,
                 reg2620,
                 forvar2618,
                 reg2619,
                 reg2618,
                 reg2617,
                 reg2616,
                 reg2613,
                 reg2615,
                 reg2614,
                 forvar2613,
                 forvar2612,
                 reg2611,
                 reg2610,
                 reg2609,
                 reg2608,
                 reg2607,
                 forvar2606,
                 forvar2605,
                 forvar2604,
                 forvar2603,
                 reg2602,
                 reg2601,
                 reg2600,
                 reg2599,
                 reg2598,
                 reg2597,
                 reg2596,
                 reg2595,
                 forvar2594,
                 reg2593,
                 reg2592,
                 reg2591,
                 forvar2589,
                 forvar2587,
                 reg2586,
                 forvar2585,
                 forvar2584,
                 forvar2583,
                 forvar2578,
                 reg2575,
                 reg2590,
                 reg2589,
                 reg2588,
                 reg2587,
                 forvar2586,
                 reg2585,
                 reg2584,
                 reg2581,
                 forvar2577,
                 reg2576,
                 reg2583,
                 reg2582,
                 forvar2581,
                 reg2580,
                 reg2579,
                 reg2578,
                 reg2577,
                 forvar2576,
                 forvar2575,
                 reg2574,
                 reg2573,
                 reg2572,
                 reg2571,
                 reg2570,
                 reg2569,
                 reg2568,
                 reg2567,
                 reg2566,
                 reg2565,
                 reg2564,
                 reg2563,
                 forvar2562,
                 reg2561,
                 reg2560,
                 reg2559,
                 reg2558,
                 reg2557,
                 forvar2556,
                 reg2555,
                 reg2554,
                 reg2553,
                 reg2552,
                 forvar2551,
                 forvar2550,
                 forvar2539,
                 reg2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2545,
                 reg2544,
                 forvar2543,
                 reg2542,
                 reg2541,
                 reg2540,
                 reg2539,
                 reg2538,
                 reg2537,
                 forvar2536,
                 reg2531,
                 reg2528,
                 forvar2527,
                 reg2536,
                 reg2535,
                 reg2534,
                 reg2533,
                 reg2532,
                 forvar2531,
                 reg2530,
                 reg2529,
                 forvar2528,
                 reg2527,
                 forvar2526,
                 reg2523,
                 forvar2519,
                 reg2518,
                 reg2525,
                 reg2524,
                 forvar2523,
                 reg2522,
                 reg2521,
                 reg2520,
                 reg2519,
                 forvar2518,
                 reg2517,
                 reg2516,
                 reg2515,
                 forvar2514,
                 forvar2513,
                 reg2512,
                 reg2476,
                 reg2475,
                 reg2472,
                 forvar2471,
                 reg2467,
                 reg2511,
                 forvar2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 forvar2506,
                 reg2505,
                 reg2504,
                 reg2503,
                 reg2502,
                 forvar2501,
                 reg2500,
                 reg2499,
                 reg2498,
                 forvar2497,
                 forvar2496,
                 reg2495,
                 reg2494,
                 reg2493,
                 reg2492,
                 reg2491,
                 forvar2489,
                 reg2487,
                 reg2490,
                 reg2489,
                 reg2488,
                 forvar2487,
                 reg2486,
                 reg2485,
                 forvar2484,
                 reg2483,
                 forvar2482,
                 reg2481,
                 reg2480,
                 forvar2479,
                 reg2478,
                 reg2477,
                 forvar2476,
                 forvar2475,
                 reg2474,
                 reg2473,
                 forvar2472,
                 reg2471,
                 reg2470,
                 reg2469,
                 reg2468,
                 forvar2467,
                 forvar2466,
                 wire2465,
                 reg2464,
                 reg2463,
                 reg2462,
                 forvar2461,
                 reg2460,
                 reg2459,
                 reg2458,
                 reg2457,
                 forvar2456,
                 forvar2451,
                 forvar2448,
                 forvar2446,
                 forvar2440,
                 forvar2450,
                 forvar2441,
                 reg2456,
                 reg2455,
                 reg2454,
                 reg2453,
                 reg2452,
                 reg2451,
                 reg2450,
                 reg2449,
                 reg2448,
                 reg2447,
                 reg2446,
                 reg2445,
                 reg2444,
                 reg2443,
                 reg2442,
                 reg2441,
                 reg2440,
                 reg2439,
                 reg2436,
                 forvar2434,
                 forvar2432,
                 forvar2431,
                 reg2430,
                 forvar2426,
                 forvar2425,
                 reg2413,
                 forvar2410,
                 forvar2407,
                 reg2395,
                 forvar2402,
                 reg2399,
                 reg2394,
                 reg2392,
                 reg2387,
                 reg2383,
                 reg2438,
                 forvar2414,
                 forvar2428,
                 reg2437,
                 forvar2436,
                 reg2435,
                 reg2434,
                 reg2433,
                 reg2432,
                 reg2431,
                 forvar2430,
                 reg2429,
                 reg2428,
                 reg2427,
                 reg2426,
                 reg2425,
                 reg2422,
                 forvar2420,
                 reg2418,
                 reg2416,
                 reg2424,
                 reg2423,
                 forvar2422,
                 reg2421,
                 reg2420,
                 reg2419,
                 forvar2418,
                 reg2417,
                 forvar2416,
                 reg2415,
                 reg2414,
                 forvar2413,
                 forvar2409,
                 forvar2404,
                 reg2412,
                 reg2411,
                 reg2410,
                 reg2409,
                 reg2408,
                 reg2407,
                 reg2406,
                 reg2405,
                 reg2404,
                 reg2403,
                 reg2402,
                 reg2401,
                 reg2400,
                 forvar2399,
                 reg2398,
                 reg2397,
                 reg2396,
                 forvar2395,
                 forvar2394,
                 reg2393,
                 forvar2392,
                 reg2391,
                 reg2390,
                 reg2389,
                 reg2388,
                 forvar2387,
                 forvar2386,
                 reg2385,
                 reg2384,
                 forvar2383,
                 forvar2382,
                 reg2373,
                 forvar2371,
                 reg2381,
                 reg2380,
                 forvar2379,
                 forvar2370,
                 reg2378,
                 reg2377,
                 reg2376,
                 reg2375,
                 reg2374,
                 forvar2373,
                 reg2372,
                 reg2371,
                 reg2370,
                 reg2369,
                 forvar2368,
                 reg2367,
                 reg2366,
                 reg2365,
                 forvar2364,
                 forvar2363,
                 forvar2362,
                 forvar2361,
                 forvar2352,
                 forvar2351,
                 forvar2349,
                 forvar2348,
                 reg2346,
                 forvar2359,
                 forvar2357,
                 forvar2355,
                 reg2354,
                 reg2360,
                 reg2359,
                 reg2358,
                 reg2357,
                 reg2356,
                 reg2355,
                 forvar2354,
                 reg2353,
                 reg2352,
                 reg2351,
                 reg2350,
                 reg2349,
                 reg2348,
                 reg2347,
                 forvar2346,
                 reg2345,
                 reg2344,
                 reg2343,
                 reg2339,
                 forvar2335,
                 reg2342,
                 reg2341,
                 reg2340,
                 forvar2339,
                 reg2338,
                 reg2337,
                 reg2336,
                 reg2335,
                 reg2334,
                 reg2333,
                 reg2332,
                 reg2331,
                 forvar2330,
                 reg2329,
                 reg2328,
                 reg2327,
                 reg2326,
                 forvar2325,
                 reg2324,
                 forvar2323,
                 forvar2322,
                 forvar2321,
                 reg2320,
                 reg2319,
                 reg2318,
                 reg2317,
                 forvar2316,
                 reg2315,
                 reg2314,
                 forvar2313,
                 reg2312,
                 forvar2311,
                 reg2310,
                 reg2309,
                 reg2308,
                 reg2307,
                 reg2306,
                 reg2305,
                 reg2304,
                 forvar2303,
                 forvar2301,
                 forvar2283,
                 reg2276,
                 forvar2296,
                 forvar2293,
                 forvar2289,
                 forvar2287,
                 reg2285,
                 forvar2282,
                 reg2280,
                 reg2279,
                 forvar2275,
                 reg2302,
                 forvar2298,
                 reg2295,
                 reg2290,
                 reg2301,
                 reg2300,
                 reg2299,
                 reg2298,
                 reg2297,
                 reg2296,
                 forvar2295,
                 reg2294,
                 reg2293,
                 reg2292,
                 reg2291,
                 forvar2290,
                 reg2289,
                 reg2288,
                 reg2287,
                 reg2286,
                 forvar2285,
                 reg2284,
                 reg2283,
                 reg2282,
                 forvar2281,
                 forvar2280,
                 forvar2279,
                 reg2278,
                 reg2277,
                 forvar2276,
                 reg2275,
                 reg2274,
                 reg2273,
                 forvar2270,
                 reg2272,
                 reg2271,
                 reg2270,
                 forvar2269,
                 reg2269,
                 reg2268,
                 reg2267,
                 reg2266,
                 reg2265,
                 forvar2264,
                 forvar2263,
                 reg2262,
                 reg2261,
                 reg2260,
                 reg2259,
                 reg2258,
                 reg2257,
                 reg2256,
                 forvar2255,
                 reg2254,
                 reg2253,
                 reg2252,
                 reg2251,
                 forvar2250,
                 reg2249,
                 forvar2248,
                 forvar2247,
                 reg2246,
                 reg2245,
                 reg2244,
                 forvar2243,
                 reg2242,
                 reg2241,
                 reg2240,
                 reg2239,
                 forvar2238,
                 reg2237,
                 reg2236,
                 reg2235,
                 reg2234,
                 reg2233,
                 reg2232,
                 reg2231,
                 reg2230,
                 forvar2229,
                 forvar2228,
                 reg2164,
                 reg2227,
                 reg2226,
                 reg2225,
                 reg2224,
                 forvar2220,
                 reg2223,
                 reg2222,
                 reg2221,
                 reg2220,
                 reg2219,
                 reg2218,
                 reg2217,
                 reg2216,
                 reg2215,
                 reg2214,
                 forvar2213,
                 forvar2212,
                 reg2211,
                 forvar2210,
                 reg2209,
                 forvar2208,
                 forvar2205,
                 reg2201,
                 reg2207,
                 reg2206,
                 reg2205,
                 reg2204,
                 reg2203,
                 reg2202,
                 forvar2201,
                 reg2200,
                 reg2199,
                 reg2198,
                 reg2197,
                 forvar2196,
                 reg2195,
                 reg2194,
                 reg2193,
                 reg2192,
                 reg2191,
                 reg2190,
                 reg2189,
                 forvar2187,
                 forvar2182,
                 reg2179,
                 forvar2177,
                 reg2174,
                 reg2173,
                 forvar2172,
                 forvar2168,
                 forvar2167,
                 reg2166,
                 reg2163,
                 forvar2162,
                 reg2188,
                 reg2187,
                 reg2186,
                 reg2185,
                 reg2184,
                 reg2183,
                 reg2182,
                 reg2181,
                 reg2180,
                 forvar2179,
                 reg2178,
                 reg2177,
                 reg2176,
                 reg2175,
                 forvar2174,
                 forvar2173,
                 reg2172,
                 reg2171,
                 reg2170,
                 reg2169,
                 reg2168,
                 reg2167,
                 forvar2166,
                 reg2165,
                 forvar2164,
                 forvar2163,
                 reg2162,
                 reg2161,
                 reg2160,
                 reg2159,
                 reg2158,
                 forvar2157,
                 reg2156,
                 reg2155,
                 reg2154,
                 forvar2153,
                 reg2152,
                 reg2151,
                 reg2150,
                 reg2149,
                 reg2148,
                 reg2147,
                 reg2146,
                 forvar2145,
                 forvar2144,
                 forvar2143,
                 reg2142,
                 reg2141,
                 reg2140,
                 reg2139,
                 reg2138,
                 reg2137,
                 forvar2136,
                 reg2135,
                 reg2134,
                 forvar2133,
                 forvar2132,
                 reg2128,
                 forvar2127,
                 reg2126,
                 reg2131,
                 reg2130,
                 reg2129,
                 forvar2128,
                 reg2127,
                 forvar2126,
                 reg2119,
                 reg2125,
                 forvar2124,
                 reg2123,
                 forvar2122,
                 reg2121,
                 reg2120,
                 forvar2119,
                 reg2118,
                 reg2117,
                 forvar2116,
                 forvar2115,
                 reg2114,
                 reg2113,
                 reg2112,
                 forvar2111,
                 forvar2103,
                 reg2102,
                 reg2110,
                 reg2109,
                 reg2108,
                 reg2107,
                 forvar2106,
                 reg2105,
                 reg2104,
                 reg2103,
                 forvar2102,
                 reg2101,
                 forvar2100,
                 reg2099,
                 reg2098,
                 reg2097,
                 forvar2096,
                 forvar2095,
                 reg2094,
                 reg2093,
                 reg2091,
                 forvar2086,
                 reg2084,
                 reg2092,
                 forvar2091,
                 reg2090,
                 reg2089,
                 reg2088,
                 reg2087,
                 reg2086,
                 reg2085,
                 forvar2084,
                 forvar2083,
                 forvar2082,
                 reg2081,
                 reg2058,
                 reg2053,
                 reg2052,
                 reg2051,
                 forvar2050,
                 reg2047,
                 reg2080,
                 reg2079,
                 forvar2078,
                 reg2077,
                 reg2076,
                 forvar2075,
                 reg2074,
                 reg2073,
                 reg2072,
                 reg2071,
                 reg2070,
                 reg2069,
                 reg2068,
                 reg2067,
                 forvar2066,
                 forvar2065,
                 reg2064,
                 reg2063,
                 forvar2062,
                 reg2061,
                 reg2060,
                 reg2059,
                 forvar2058,
                 reg2057,
                 reg2056,
                 reg2055,
                 reg2054,
                 forvar2053,
                 forvar2052,
                 forvar2051,
                 reg2050,
                 forvar2049,
                 forvar2048,
                 forvar2047,
                 reg2046,
                 forvar2041,
                 reg2045,
                 reg2044,
                 reg2043,
                 reg2042,
                 reg2041,
                 forvar2040,
                 reg2035,
                 reg2039,
                 reg2038,
                 reg2037,
                 reg2036,
                 forvar2035,
                 forvar2025,
                 reg2034,
                 forvar2033,
                 reg2032,
                 reg2031,
                 forvar2030,
                 reg2029,
                 forvar2028,
                 reg2027,
                 reg2026,
                 reg2025,
                 reg2024,
                 forvar2023,
                 forvar2022,
                 reg2020,
                 forvar2015,
                 reg2013,
                 reg2011,
                 reg2021,
                 forvar2020,
                 reg2019,
                 reg2018,
                 reg2017,
                 reg2016,
                 reg2015,
                 reg2014,
                 forvar2013,
                 reg2012,
                 forvar2011,
                 reg2010,
                 reg2009,
                 forvar2001,
                 reg2008,
                 forvar2007,
                 reg2006,
                 reg2005,
                 forvar2004,
                 reg2003,
                 reg2002,
                 reg2001,
                 reg2000,
                 forvar1999,
                 forvar1998,
                 forvar1980,
                 forvar1974,
                 reg1976,
                 forvar1971,
                 forvar1970,
                 reg1997,
                 reg1996,
                 reg1995,
                 reg1991,
                 reg1994,
                 reg1993,
                 reg1992,
                 forvar1991,
                 forvar1983,
                 reg1990,
                 reg1989,
                 reg1988,
                 reg1987,
                 reg1986,
                 reg1985,
                 reg1984,
                 reg1983,
                 reg1982,
                 reg1981,
                 reg1980,
                 reg1979,
                 reg1978,
                 reg1977,
                 forvar1976,
                 reg1967,
                 reg1975,
                 reg1974,
                 reg1973,
                 reg1972,
                 reg1971,
                 reg1970,
                 reg1969,
                 reg1968,
                 forvar1967,
                 reg1966,
                 reg1965,
                 reg1963,
                 forvar1962,
                 reg1964,
                 forvar1963,
                 reg1962,
                 reg1961,
                 reg1960,
                 forvar1959,
                 reg1958,
                 reg1957,
                 forvar1956,
                 reg1955,
                 reg1954,
                 reg1953,
                 reg1952,
                 reg1948,
                 forvar1947,
                 reg1951,
                 reg1950,
                 reg1949,
                 forvar1948,
                 reg1947,
                 reg1946,
                 reg1941,
                 forvar1939,
                 forvar1936,
                 reg1945,
                 reg1944,
                 forvar1943,
                 reg1942,
                 forvar1941,
                 reg1938,
                 reg1934,
                 forvar1933,
                 forvar1931,
                 reg1940,
                 reg1939,
                 forvar1938,
                 reg1937,
                 reg1936,
                 reg1935,
                 forvar1934,
                 reg1933,
                 reg1932,
                 reg1931,
                 forvar1930,
                 reg1929,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1929 <= (wire1928[(3'h7):(3'h5)] ^~ {wire1924[(1'h0):(1'h0)]});
    end
  always
    @(posedge clk) begin
      for (forvar1930 = (1'h0); (forvar1930 < (2'h2)); forvar1930 = (forvar1930 + (1'h1)))
        begin
          if ((8'ha0))
            begin
              if ((wire1925[(3'h4):(2'h2)] || (wire1925 ?
                  {reg1929[(1'h0):(1'h0)]} : ((wire1927 ? wire1927 : wire1927) ?
                      {wire1925} : wire1927))))
                begin
                  if ({($unsigned((8'haf)) < ((reg1929 ? forvar1930 : (8'hb1)) ?
                          (~|(8'h9f)) : {wire1927}))})
                    begin
                      reg1931 <= wire1928;
                      reg1932 <= reg1929[(4'hd):(1'h0)];
                      reg1933 <= $unsigned($signed((reg1931[(2'h3):(2'h3)] ?
                          wire1926[(2'h3):(2'h3)] : {wire1927})));
                    end
                  else
                    begin
                      reg1931 <= wire1928[(1'h1):(1'h1)];
                      reg1932 <= ({$unsigned((wire1927 ~^ reg1931))} ?
                          ($signed(((8'h9f) ? wire1928 : wire1926)) ?
                              $unsigned($unsigned(wire1928)) : ((8'hac) ?
                                  {reg1931} : (~&wire1924))) : wire1928[(2'h3):(2'h2)]);
                    end
                  for (forvar1934 = (1'h0); (forvar1934 < (1'h0)); forvar1934 = (forvar1934 + (1'h1)))
                    begin
                      reg1935 <= wire1926;
                    end
                  if (($signed(($signed(wire1924) >= (reg1932 + wire1924))) ?
                      reg1932[(3'h7):(2'h3)] : $signed(((reg1932 | wire1927) ?
                          (^~reg1933) : (wire1926 ? reg1933 : wire1927)))))
                    begin
                      reg1936 <= (reg1935 ?
                          (reg1931 ?
                              $unsigned(forvar1934) : ($unsigned((8'hae)) ?
                                  {reg1932} : wire1925)) : $signed($unsigned((8'hb0))));
                      reg1937 <= {$unsigned($unsigned(reg1936))};
                    end
                  else
                    begin
                      reg1936 <= reg1935;
                      reg1937 <= forvar1930;
                    end
                  for (forvar1938 = (1'h0); (forvar1938 < (2'h3)); forvar1938 = (forvar1938 + (1'h1)))
                    begin
                      reg1939 <= (+(({wire1925} ?
                              (~|wire1924) : reg1935[(1'h1):(1'h0)]) ?
                          $unsigned(wire1927) : $signed($signed(reg1932))));
                      reg1940 <= reg1932[(3'h5):(3'h5)];
                    end
                end
              else
                begin
                  for (forvar1931 = (1'h0); (forvar1931 < (2'h3)); forvar1931 = (forvar1931 + (1'h1)))
                    begin
                      reg1932 <= ((~$signed(reg1935)) ?
                          $unsigned(reg1932) : $signed(reg1933));
                    end
                  for (forvar1933 = (1'h0); (forvar1933 < (1'h1)); forvar1933 = (forvar1933 + (1'h1)))
                    begin
                      reg1934 <= reg1929[(4'hb):(3'h7)];
                      reg1935 <= (+(+(reg1940 >> $signed(reg1939))));
                    end
                  if ((~&wire1928))
                    begin
                      reg1936 <= {$unsigned($unsigned($signed(forvar1934)))};
                      reg1937 <= (&forvar1933[(1'h1):(1'h1)]);
                      reg1938 <= $unsigned((|((reg1939 ?
                          (8'hb0) : reg1929) >= (forvar1938 || (8'h9c)))));
                      reg1939 <= $signed(reg1939);
                    end
                  else
                    begin
                      reg1936 <= $signed($unsigned({$signed(wire1925)}));
                      reg1937 <= (-(8'hb9));
                      reg1938 <= ((8'h9e) << reg1934[(4'ha):(2'h2)]);
                      reg1939 <= reg1933[(1'h1):(1'h0)];
                    end
                end
              for (forvar1941 = (1'h0); (forvar1941 < (1'h0)); forvar1941 = (forvar1941 + (1'h1)))
                begin
                  if ((((8'ha6) <= reg1931) >> reg1937))
                    begin
                      reg1942 <= ((~^$signed(((8'hae) ?
                          wire1924 : reg1935))) > {((-forvar1938) >>> (forvar1933 << wire1928))});
                    end
                  else
                    begin
                      reg1942 <= (+$unsigned($signed((wire1926 <<< forvar1931))));
                    end
                  for (forvar1943 = (1'h0); (forvar1943 < (2'h3)); forvar1943 = (forvar1943 + (1'h1)))
                    begin
                      reg1944 <= reg1937;
                      reg1945 <= ($unsigned((^~$signed(forvar1941))) ?
                          {((reg1933 <= reg1929) > {wire1924})} : $signed($signed(reg1931)));
                    end
                end
            end
          else
            begin
              for (forvar1931 = (1'h0); (forvar1931 < (1'h0)); forvar1931 = (forvar1931 + (1'h1)))
                begin
                  if (((forvar1943[(2'h3):(2'h3)] ?
                          $unsigned(reg1936) : (+$unsigned(reg1940))) ?
                      (((forvar1938 ? reg1939 : reg1944) ^~ (reg1937 ?
                              reg1934 : (8'ha6))) ?
                          (wire1926[(2'h2):(1'h0)] ?
                              ((8'haf) && reg1931) : $unsigned(reg1936)) : $unsigned((~^wire1924))) : (-$signed($signed(forvar1938)))))
                    begin
                      reg1932 <= reg1937;
                      reg1933 <= $signed(reg1929[(3'h7):(1'h0)]);
                      reg1934 <= wire1926[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg1932 <= reg1929[(3'h6):(1'h0)];
                      reg1933 <= ({(reg1939 ?
                              $unsigned(forvar1934) : {wire1925})} && (~reg1933[(1'h0):(1'h0)]));
                      reg1934 <= {($signed(((8'ha7) ?
                              reg1931 : reg1929)) & $unsigned((forvar1933 - (8'ha9))))};
                    end
                  reg1935 <= forvar1933[(4'h9):(1'h1)];
                  for (forvar1936 = (1'h0); (forvar1936 < (2'h3)); forvar1936 = (forvar1936 + (1'h1)))
                    begin
                      reg1937 <= (($unsigned($unsigned(forvar1943)) < {$signed(wire1924)}) ?
                          (~$unsigned((reg1942 ?
                              wire1928 : reg1929))) : ((8'hb4) > {(wire1926 ?
                                  (8'ha9) : (8'had))}));
                    end
                end
              for (forvar1938 = (1'h0); (forvar1938 < (2'h3)); forvar1938 = (forvar1938 + (1'h1)))
                begin
                  for (forvar1939 = (1'h0); (forvar1939 < (1'h1)); forvar1939 = (forvar1939 + (1'h1)))
                    begin
                      reg1940 <= ($signed(($unsigned(reg1944) && (-forvar1938))) ?
                          (^reg1931) : reg1944);
                      reg1941 <= (-wire1924[(3'h5):(3'h4)]);
                      reg1942 <= wire1928[(3'h4):(1'h1)];
                    end
                  for (forvar1943 = (1'h0); (forvar1943 < (1'h0)); forvar1943 = (forvar1943 + (1'h1)))
                    begin
                      reg1944 <= ((^(~|(^~reg1944))) ?
                          ((reg1936[(3'h5):(3'h4)] + (forvar1938 ?
                                  (8'hac) : (8'h9c))) ?
                              $unsigned($unsigned(reg1942)) : $signed($signed(forvar1936))) : ((~&(8'h9c)) > forvar1930[(3'h6):(1'h0)]));
                      reg1945 <= wire1924;
                      reg1946 <= reg1945;
                    end
                end
              if ((forvar1930[(4'ha):(3'h5)] | forvar1938[(1'h0):(1'h0)]))
                begin
                  reg1947 <= $signed(reg1934[(4'hc):(3'h7)]);
                  for (forvar1948 = (1'h0); (forvar1948 < (1'h0)); forvar1948 = (forvar1948 + (1'h1)))
                    begin
                      reg1949 <= (8'hb0);
                      reg1950 <= ($unsigned((~&(|(8'had)))) & reg1947);
                      reg1951 <= wire1925;
                    end
                end
              else
                begin
                  for (forvar1947 = (1'h0); (forvar1947 < (2'h2)); forvar1947 = (forvar1947 + (1'h1)))
                    begin
                      reg1948 <= $signed((8'hb9));
                      reg1949 <= reg1950[(4'h8):(3'h5)];
                      reg1950 <= {(wire1928 ^~ $signed(reg1945))};
                      reg1951 <= ((&(reg1951[(4'h8):(3'h4)] >> (reg1933 != reg1933))) ?
                          (8'had) : (~|((!reg1949) ?
                              $signed((8'hba)) : {reg1933})));
                    end
                  if (reg1949[(1'h1):(1'h1)])
                    begin
                      reg1952 <= (($unsigned($unsigned(forvar1934)) ?
                          (&$signed(forvar1947)) : (((8'ha7) ?
                              reg1932 : reg1951) >>> reg1942[(1'h0):(1'h0)])) ^ $signed((-reg1938[(4'h9):(3'h5)])));
                    end
                  else
                    begin
                      reg1952 <= {((^reg1932) << (reg1946[(1'h1):(1'h0)] + $signed(reg1952)))};
                      reg1953 <= (reg1937 <= (forvar1939 ?
                          ($unsigned(reg1932) ?
                              reg1932[(3'h5):(3'h4)] : (~|reg1931)) : (^~(forvar1941 ?
                              forvar1930 : reg1936))));
                      reg1954 <= ((((forvar1938 ?
                              reg1936 : forvar1931) != $unsigned(wire1927)) ?
                          $signed((wire1927 ?
                              (8'h9f) : reg1934)) : reg1934[(3'h6):(3'h6)]) < reg1942[(2'h3):(2'h3)]);
                      reg1955 <= $signed($signed($unsigned($signed(forvar1934))));
                    end
                  for (forvar1956 = (1'h0); (forvar1956 < (2'h2)); forvar1956 = (forvar1956 + (1'h1)))
                    begin
                      reg1957 <= $signed((wire1928 - forvar1947[(2'h3):(2'h3)]));
                      reg1958 <= {$unsigned($unsigned($signed(reg1940)))};
                    end
                end
              if ({($signed((wire1925 >>> (8'ha9))) ?
                      reg1934[(4'h8):(1'h1)] : $signed(((8'hb9) <= reg1933)))})
                begin
                  for (forvar1959 = (1'h0); (forvar1959 < (2'h2)); forvar1959 = (forvar1959 + (1'h1)))
                    begin
                      reg1960 <= (((reg1950[(3'h6):(1'h1)] << reg1935) ?
                          reg1931 : ((+reg1949) ?
                              (reg1948 ? reg1932 : forvar1948) : ((8'hb3) ?
                                  (8'ha5) : wire1924))) << $unsigned($signed($unsigned(reg1941))));
                    end
                  reg1961 <= $signed(((reg1952[(3'h7):(1'h0)] ^ (^~reg1936)) ?
                      reg1931[(3'h5):(3'h5)] : $signed($signed(reg1958))));
                  reg1962 <= ($unsigned((reg1941 ?
                          $unsigned(reg1938) : $signed(reg1935))) ?
                      reg1934[(3'h7):(3'h6)] : ({forvar1938[(1'h1):(1'h0)]} << ($signed(wire1928) >> {reg1957})));
                  for (forvar1963 = (1'h0); (forvar1963 < (2'h2)); forvar1963 = (forvar1963 + (1'h1)))
                    begin
                      reg1964 <= $signed({$signed((reg1941 ?
                              (8'hb4) : reg1941))});
                    end
                end
              else
                begin
                  for (forvar1959 = (1'h0); (forvar1959 < (2'h2)); forvar1959 = (forvar1959 + (1'h1)))
                    begin
                      reg1960 <= $signed((~&$unsigned(reg1937[(1'h0):(1'h0)])));
                      reg1961 <= reg1950;
                    end
                  for (forvar1962 = (1'h0); (forvar1962 < (1'h0)); forvar1962 = (forvar1962 + (1'h1)))
                    begin
                      reg1963 <= forvar1956;
                      reg1964 <= {{reg1955[(3'h4):(1'h0)]}};
                      reg1965 <= reg1955[(3'h6):(3'h4)];
                    end
                  reg1966 <= reg1954;
                end
            end
          if ($unsigned(reg1960))
            begin
              if (reg1963)
                begin
                  for (forvar1967 = (1'h0); (forvar1967 < (2'h3)); forvar1967 = (forvar1967 + (1'h1)))
                    begin
                      reg1968 <= ($unsigned(forvar1956) ?
                          (reg1935[(2'h3):(1'h1)] ^~ ({reg1939} ?
                              {(8'ha7)} : ((8'had) && reg1951))) : $signed(((reg1935 ^ reg1952) ?
                              (~reg1944) : $unsigned(reg1932))));
                      reg1969 <= reg1938;
                    end
                  if ($unsigned(((reg1968 ?
                      $signed(reg1960) : (~^reg1953)) - forvar1948[(1'h1):(1'h0)])))
                    begin
                      reg1970 <= reg1940[(2'h2):(1'h1)];
                      reg1971 <= reg1949[(1'h0):(1'h0)];
                      reg1972 <= $unsigned(reg1945[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1970 <= $signed($unsigned((forvar1947[(1'h0):(1'h0)] <<< (reg1964 <= reg1968))));
                      reg1971 <= (~^((~&{(8'h9c)}) ?
                          $signed((^forvar1948)) : $unsigned((forvar1963 | reg1950))));
                      reg1972 <= reg1932[(2'h3):(2'h3)];
                    end
                  if (forvar1947[(2'h3):(2'h3)])
                    begin
                      reg1973 <= $unsigned((8'h9e));
                      reg1974 <= wire1928[(4'h8):(2'h2)];
                      reg1975 <= $signed($unsigned({forvar1943[(1'h0):(1'h0)]}));
                    end
                  else
                    begin
                      reg1973 <= ((^~{(reg1972 ?
                              reg1961 : forvar1947)}) > (!forvar1948[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  reg1967 <= reg1953;
                end
              if (((reg1972 ?
                  reg1970[(1'h1):(1'h1)] : reg1929) == (|{(reg1939 || forvar1934)})))
                begin
                  for (forvar1976 = (1'h0); (forvar1976 < (2'h3)); forvar1976 = (forvar1976 + (1'h1)))
                    begin
                      reg1977 <= reg1973;
                      reg1978 <= $unsigned(forvar1962);
                      reg1979 <= (^~($unsigned((!reg1958)) != (^wire1927[(4'ha):(2'h3)])));
                    end
                  if (($unsigned($unsigned($signed(reg1944))) & (((wire1926 ?
                      reg1951 : wire1924) - ((8'h9d) & reg1951)) | reg1948)))
                    begin
                      reg1980 <= forvar1947[(3'h4):(1'h0)];
                      reg1981 <= $signed(((8'h9f) > $signed(((8'hac) ?
                          forvar1930 : forvar1938))));
                      reg1982 <= reg1937[(4'h9):(3'h6)];
                      reg1983 <= {reg1975[(2'h2):(1'h0)]};
                    end
                  else
                    begin
                      reg1980 <= $signed(forvar1943[(3'h4):(2'h3)]);
                      reg1981 <= (+$unsigned($unsigned((reg1967 < reg1980))));
                      reg1982 <= $unsigned($signed($signed((forvar1936 - reg1961))));
                      reg1983 <= (~&$unsigned(forvar1962));
                    end
                  if ($unsigned((~|(^(reg1937 ? reg1945 : reg1939)))))
                    begin
                      reg1984 <= ({(~^(^~(8'ha8)))} <<< $signed($unsigned((8'ha5))));
                      reg1985 <= ((!reg1970) ?
                          {reg1934[(3'h7):(3'h4)]} : (^~((^(8'ha1)) ?
                              reg1937 : $unsigned(reg1945))));
                      reg1986 <= {(~&$signed((~&reg1934)))};
                      reg1987 <= forvar1963;
                    end
                  else
                    begin
                      reg1984 <= ((~reg1949) ?
                          (~^reg1944[(3'h5):(1'h0)]) : (8'ha6));
                      reg1985 <= (!(~|((reg1960 - forvar1963) ?
                          reg1962 : (^~reg1952))));
                      reg1986 <= $signed($unsigned((((8'hb3) ?
                              reg1942 : reg1985) ?
                          $unsigned(reg1933) : wire1927[(1'h1):(1'h1)])));
                    end
                  if ((^(8'hb9)))
                    begin
                      reg1988 <= forvar1931;
                      reg1989 <= (reg1934[(4'ha):(3'h4)] ?
                          $signed(($unsigned(reg1979) | {(8'ha3)})) : wire1924[(3'h7):(2'h3)]);
                      reg1990 <= (&(reg1969 >= reg1931));
                    end
                  else
                    begin
                      reg1988 <= $signed((wire1924 ?
                          (forvar1963 ?
                              $signed(reg1942) : $unsigned(reg1929)) : $signed((forvar1931 ?
                              forvar1943 : forvar1956))));
                      reg1989 <= $signed(({$signed(reg1940)} ?
                          (~|$unsigned(wire1926)) : (reg1939[(1'h0):(1'h0)] ?
                              reg1937[(3'h7):(2'h2)] : reg1929)));
                      reg1990 <= (~reg1989[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar1976 = (1'h0); (forvar1976 < (1'h1)); forvar1976 = (forvar1976 + (1'h1)))
                    begin
                      reg1977 <= ({$unsigned((~^reg1988))} ?
                          (forvar1962[(3'h5):(1'h0)] >> (~^reg1974[(2'h3):(1'h0)])) : (-(|$signed(reg1951))));
                      reg1978 <= reg1960[(4'h8):(1'h0)];
                    end
                  if (reg1958)
                    begin
                      reg1979 <= wire1928;
                      reg1980 <= $signed(forvar1963);
                      reg1981 <= $unsigned($signed(reg1952));
                      reg1982 <= ($signed($unsigned($signed((8'hab)))) != $signed(forvar1967[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1979 <= $unsigned((wire1926[(3'h5):(2'h3)] ?
                          $signed((reg1979 >>> reg1988)) : (|(!forvar1967))));
                      reg1980 <= $unsigned(($signed(forvar1976) ?
                          reg1953 : (forvar1963 ?
                              $unsigned((8'hb2)) : reg1963[(4'h9):(4'h9)])));
                      reg1981 <= (&((reg1985 - (8'ha1)) ?
                          ($signed(reg1937) && {reg1974}) : (~forvar1939[(1'h0):(1'h0)])));
                      reg1982 <= forvar1938;
                    end
                  for (forvar1983 = (1'h0); (forvar1983 < (2'h3)); forvar1983 = (forvar1983 + (1'h1)))
                    begin
                      reg1984 <= $signed(wire1924);
                      reg1985 <= $unsigned($unsigned(reg1942[(4'h8):(1'h1)]));
                    end
                end
              if (reg1967[(3'h7):(2'h2)])
                begin
                  for (forvar1991 = (1'h0); (forvar1991 < (2'h2)); forvar1991 = (forvar1991 + (1'h1)))
                    begin
                      reg1992 <= (!$signed((^~reg1985)));
                      reg1993 <= ($unsigned($unsigned(forvar1976)) & $unsigned(((reg1989 ?
                              reg1971 : reg1971) ?
                          ((8'haf) != forvar1963) : reg1973)));
                      reg1994 <= ((8'ha4) < $unsigned((-(|reg1937))));
                    end
                end
              else
                begin
                  if (($signed((+(~&reg1941))) - $signed($signed(reg1974))))
                    begin
                      reg1991 <= $signed($unsigned($signed(((8'h9c) ?
                          reg1960 : reg1941))));
                    end
                  else
                    begin
                      reg1991 <= ($unsigned((~^forvar1931[(1'h0):(1'h0)])) ?
                          ($signed((reg1986 ?
                              reg1971 : reg1971)) | {$signed(reg1970)}) : (&((~^reg1933) >= reg1958)));
                      reg1992 <= $signed($signed(((~(8'hb0)) || reg1977)));
                    end
                  if (reg1975[(2'h3):(1'h1)])
                    begin
                      reg1993 <= (8'ha7);
                    end
                  else
                    begin
                      reg1993 <= (~(^($unsigned(reg1962) ?
                          $signed((8'hb0)) : (|(8'hab)))));
                      reg1994 <= wire1925[(2'h3):(2'h3)];
                    end
                  if (reg1961[(3'h7):(3'h5)])
                    begin
                      reg1995 <= {$unsigned(reg1946[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg1995 <= $unsigned((^~((&reg1988) == {forvar1948})));
                      reg1996 <= (-$unsigned(reg1957));
                      reg1997 <= $unsigned($signed(((-(8'hb6)) >> reg1991)));
                    end
                end
            end
          else
            begin
              if ({reg1978})
                begin
                  if (((forvar1959[(2'h3):(1'h1)] <<< $signed($unsigned((8'hb2)))) + (-$signed($unsigned((8'haf))))))
                    begin
                      reg1967 <= forvar1948;
                      reg1968 <= {$unsigned((((8'hb9) ^~ reg1971) == $signed(wire1925)))};
                      reg1969 <= $signed((((reg1938 >> reg1934) ~^ (~forvar1948)) ?
                          $unsigned(((8'hb1) || forvar1933)) : (reg1969 ?
                              {reg1933} : (|reg1931))));
                    end
                  else
                    begin
                      reg1967 <= $signed((reg1971 ?
                          $unsigned((reg1997 ^~ reg1951)) : ((reg1987 ?
                              reg1953 : forvar1959) - forvar1956)));
                    end
                  for (forvar1970 = (1'h0); (forvar1970 < (1'h0)); forvar1970 = (forvar1970 + (1'h1)))
                    begin
                      reg1971 <= reg1952;
                    end
                end
              else
                begin
                  for (forvar1967 = (1'h0); (forvar1967 < (2'h2)); forvar1967 = (forvar1967 + (1'h1)))
                    begin
                      reg1968 <= forvar1933;
                      reg1969 <= $unsigned($signed((reg1964 && (reg1994 <= forvar1963))));
                    end
                  reg1970 <= $signed($signed($signed(reg1963[(3'h7):(1'h1)])));
                  for (forvar1971 = (1'h0); (forvar1971 < (1'h0)); forvar1971 = (forvar1971 + (1'h1)))
                    begin
                      reg1972 <= (!($signed((reg1996 ?
                          reg1974 : reg1929)) & reg1986[(3'h6):(3'h5)]));
                      reg1973 <= (|$signed(reg1974[(3'h6):(3'h6)]));
                    end
                end
              if ((~|(reg1935 <= forvar1948[(3'h5):(1'h1)])))
                begin
                  if ($signed((-$unsigned($unsigned(reg1993)))))
                    begin
                      reg1974 <= forvar1948[(1'h0):(1'h0)];
                      reg1975 <= ($unsigned((reg1985[(2'h2):(2'h2)] ?
                              reg1931[(3'h5):(2'h2)] : $unsigned(forvar1933))) ?
                          (reg1942 ?
                              (+$unsigned(reg1971)) : (((8'ha5) ?
                                  reg1946 : (8'ha0)) & (!reg1969))) : $signed(((8'hae) ?
                              (forvar1983 + reg1981) : $signed(reg1949))));
                    end
                  else
                    begin
                      reg1974 <= (8'hb8);
                      reg1975 <= (+reg1942[(3'h6):(3'h6)]);
                    end
                  reg1976 <= (reg1982 != ($unsigned((|(8'hac))) ?
                      (^$unsigned(reg1950)) : (((8'h9d) >>> reg1967) ?
                          (-reg1963) : (reg1984 < reg1950))));
                  reg1977 <= reg1953[(4'h8):(3'h4)];
                end
              else
                begin
                  for (forvar1974 = (1'h0); (forvar1974 < (2'h3)); forvar1974 = (forvar1974 + (1'h1)))
                    begin
                      reg1975 <= reg1961;
                      reg1976 <= ($signed($unsigned((8'had))) - {$unsigned(reg1988)});
                      reg1977 <= {($signed((8'hb3)) != $signed((!reg1995)))};
                      reg1978 <= reg1991[(3'h5):(2'h3)];
                    end
                  reg1979 <= (^~(8'hb5));
                  for (forvar1980 = (1'h0); (forvar1980 < (2'h3)); forvar1980 = (forvar1980 + (1'h1)))
                    begin
                      reg1981 <= (^{(~&$signed(forvar1931))});
                      reg1982 <= reg1957;
                      reg1983 <= $signed($unsigned($signed(reg1969)));
                      reg1984 <= $signed(({(8'hb9)} || ($signed(reg1970) - reg1987[(3'h6):(2'h3)])));
                    end
                end
            end
        end
      for (forvar1998 = (1'h0); (forvar1998 < (2'h3)); forvar1998 = (forvar1998 + (1'h1)))
        begin
          for (forvar1999 = (1'h0); (forvar1999 < (2'h2)); forvar1999 = (forvar1999 + (1'h1)))
            begin
              if ((-(forvar1991 ? {reg1953} : wire1927[(4'h8):(2'h2)])))
                begin
                  if ((~{(8'ha4)}))
                    begin
                      reg2000 <= (~&(({reg1984} ?
                          $signed(forvar1934) : reg1936[(1'h1):(1'h1)]) & reg1954));
                      reg2001 <= reg1967;
                      reg2002 <= {$signed(((reg1991 ?
                              forvar1956 : reg1974) != (|reg1971)))};
                    end
                  else
                    begin
                      reg2000 <= (reg1970 == $signed(reg2000[(2'h3):(2'h2)]));
                    end
                  reg2003 <= (~|((!$unsigned(reg1949)) + reg1957[(3'h6):(1'h1)]));
                  for (forvar2004 = (1'h0); (forvar2004 < (2'h2)); forvar2004 = (forvar2004 + (1'h1)))
                    begin
                      reg2005 <= (~|(((^forvar1934) ?
                          {(8'ha6)} : $unsigned((8'ha1))) >> $unsigned((8'hab))));
                      reg2006 <= $unsigned($unsigned((forvar1991 << $signed(reg1951))));
                    end
                  for (forvar2007 = (1'h0); (forvar2007 < (2'h2)); forvar2007 = (forvar2007 + (1'h1)))
                    begin
                      reg2008 <= $signed(((!(reg1991 ?
                          forvar1938 : (8'ha6))) <<< reg1971));
                    end
                end
              else
                begin
                  reg2000 <= $signed({(~reg1950[(4'hb):(3'h5)])});
                  for (forvar2001 = (1'h0); (forvar2001 < (1'h1)); forvar2001 = (forvar2001 + (1'h1)))
                    begin
                      reg2002 <= $unsigned(reg1988[(4'h8):(3'h4)]);
                      reg2003 <= $signed((reg2008 ?
                          $signed((&reg1965)) : ($unsigned(forvar1941) | {reg1997})));
                    end
                  for (forvar2004 = (1'h0); (forvar2004 < (1'h0)); forvar2004 = (forvar2004 + (1'h1)))
                    begin
                      reg2005 <= ($signed((|(reg1967 - wire1924))) ?
                          $unsigned(reg1960[(3'h6):(1'h0)]) : ($unsigned(reg1938) ?
                              ((forvar1967 ? reg1977 : forvar1980) ?
                                  reg2005[(1'h1):(1'h1)] : $signed(reg1967)) : (8'had)));
                      reg2006 <= {((!(reg1951 <= reg1936)) ?
                              reg1972 : ($unsigned(reg1940) << (^~wire1924)))};
                    end
                  for (forvar2007 = (1'h0); (forvar2007 < (1'h0)); forvar2007 = (forvar2007 + (1'h1)))
                    begin
                      reg2008 <= (reg1941 ?
                          (forvar2007 | $unsigned($unsigned(reg1990))) : ($unsigned((reg1972 && forvar1941)) | reg1964));
                      reg2009 <= reg1967;
                      reg2010 <= $signed((reg1958 - $unsigned(((8'hb8) ?
                          reg1947 : reg2008))));
                    end
                end
              if ($signed(reg1952[(4'h9):(4'h9)]))
                begin
                  for (forvar2011 = (1'h0); (forvar2011 < (2'h3)); forvar2011 = (forvar2011 + (1'h1)))
                    begin
                      reg2012 <= reg2000;
                    end
                  for (forvar2013 = (1'h0); (forvar2013 < (1'h1)); forvar2013 = (forvar2013 + (1'h1)))
                    begin
                      reg2014 <= (((~&((8'hb1) ? reg1950 : reg1967)) ?
                              reg1970 : forvar1948) ?
                          $signed($unsigned(reg1970)) : reg1946[(3'h6):(1'h0)]);
                      reg2015 <= $unsigned((^~reg1970));
                    end
                  if (reg1957[(2'h2):(1'h0)])
                    begin
                      reg2016 <= ({(reg1991[(3'h6):(2'h2)] ?
                                  (reg1969 ? reg1945 : reg1955) : (forvar1959 ?
                                      reg2002 : reg1933))} ?
                          {$signed((~&reg1951))} : (+{reg1929[(4'h9):(4'h8)]}));
                      reg2017 <= ($unsigned((reg1940[(2'h2):(2'h2)] ?
                          $unsigned(reg1944) : (forvar2007 ?
                              reg1964 : reg1958))) >> $signed((reg1950[(4'hd):(4'ha)] > (forvar2001 + wire1928))));
                      reg2018 <= $signed($unsigned(reg1932));
                      reg2019 <= $signed(forvar1938);
                    end
                  else
                    begin
                      reg2016 <= ($signed((-$signed(reg1960))) ?
                          (((|reg1952) ?
                                  reg1974[(3'h4):(2'h3)] : $signed(reg1964)) ?
                              $signed(reg2015[(1'h1):(1'h0)]) : ((forvar1967 != reg1973) ^~ reg2005[(4'he):(3'h6)])) : $unsigned($signed((~&reg1986))));
                      reg2017 <= $signed($signed($signed(reg1989[(3'h4):(1'h1)])));
                    end
                  for (forvar2020 = (1'h0); (forvar2020 < (1'h1)); forvar2020 = (forvar2020 + (1'h1)))
                    begin
                      reg2021 <= {reg1978[(3'h6):(2'h3)]};
                    end
                end
              else
                begin
                  if (reg1936)
                    begin
                      reg2011 <= (-{$unsigned($signed(reg2008))});
                      reg2012 <= $unsigned(reg1993[(1'h1):(1'h1)]);
                      reg2013 <= $signed($signed((8'hb4)));
                      reg2014 <= $unsigned((!reg2018[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg2011 <= $unsigned((reg1990 < forvar1963[(4'h9):(3'h7)]));
                      reg2012 <= $unsigned(reg1932[(3'h7):(3'h4)]);
                      reg2013 <= (~|reg1960);
                    end
                  for (forvar2015 = (1'h0); (forvar2015 < (1'h0)); forvar2015 = (forvar2015 + (1'h1)))
                    begin
                      reg2016 <= (reg1941 ?
                          ($signed($unsigned(reg1938)) ?
                              (!(reg1982 ^~ forvar1998)) : ($signed(reg1945) ?
                                  ((8'had) ? reg1950 : forvar2020) : (reg1937 ?
                                      reg1997 : reg1948))) : $unsigned(($signed(reg1953) << (8'ha7))));
                      reg2017 <= reg1984[(2'h3):(2'h3)];
                    end
                  if ($unsigned($signed(((reg1986 != reg1953) ?
                      reg1982[(4'hc):(4'hc)] : forvar1943[(1'h0):(1'h0)]))))
                    begin
                      reg2018 <= reg1945;
                      reg2019 <= (-forvar1976[(2'h2):(1'h1)]);
                      reg2020 <= reg2002;
                      reg2021 <= $signed($unsigned({$signed((8'hb8))}));
                    end
                  else
                    begin
                      reg2018 <= ($signed($unsigned(reg1962[(2'h2):(2'h2)])) << $unsigned(forvar1936));
                      reg2019 <= (^$signed(reg1951[(3'h7):(2'h3)]));
                      reg2020 <= ((reg1969 ?
                          $signed($unsigned(forvar1999)) : ($unsigned((8'hae)) ?
                              reg1947 : (reg1949 + reg1946))) ^~ $signed(forvar2004[(1'h1):(1'h1)]));
                    end
                end
            end
          for (forvar2022 = (1'h0); (forvar2022 < (2'h3)); forvar2022 = (forvar2022 + (1'h1)))
            begin
              if (($unsigned({reg1964}) ?
                  ($unsigned((|reg1989)) | ((forvar2020 == forvar2020) ?
                      $unsigned(reg1970) : (wire1924 ?
                          forvar1938 : forvar1998))) : reg1981))
                begin
                  for (forvar2023 = (1'h0); (forvar2023 < (1'h1)); forvar2023 = (forvar2023 + (1'h1)))
                    begin
                      reg2024 <= (~&({(reg1957 ?
                              (8'hb6) : (8'ha5))} && $unsigned($signed(reg1979))));
                      reg2025 <= (reg1931[(2'h3):(2'h2)] ?
                          ((~^forvar1976) > reg1967) : (($unsigned(reg1947) - (^forvar1931)) <= (+(reg1990 | (8'haa)))));
                      reg2026 <= reg2008[(3'h7):(3'h4)];
                      reg2027 <= (reg2018 ~^ reg2025[(4'h9):(3'h6)]);
                    end
                  for (forvar2028 = (1'h0); (forvar2028 < (2'h2)); forvar2028 = (forvar2028 + (1'h1)))
                    begin
                      reg2029 <= $unsigned($unsigned(((reg1981 ?
                              forvar1980 : (8'h9e)) ?
                          $signed((8'hba)) : (&forvar1956))));
                    end
                  for (forvar2030 = (1'h0); (forvar2030 < (1'h1)); forvar2030 = (forvar2030 + (1'h1)))
                    begin
                      reg2031 <= reg1960[(4'hd):(2'h3)];
                      reg2032 <= reg2029;
                    end
                  for (forvar2033 = (1'h0); (forvar2033 < (2'h3)); forvar2033 = (forvar2033 + (1'h1)))
                    begin
                      reg2034 <= (8'ha8);
                    end
                end
              else
                begin
                  for (forvar2023 = (1'h0); (forvar2023 < (1'h0)); forvar2023 = (forvar2023 + (1'h1)))
                    begin
                      reg2024 <= reg2025[(3'h4):(3'h4)];
                    end
                  for (forvar2025 = (1'h0); (forvar2025 < (2'h2)); forvar2025 = (forvar2025 + (1'h1)))
                    begin
                      reg2026 <= reg2026;
                    end
                end
              if (forvar2011[(3'h5):(3'h5)])
                begin
                  for (forvar2035 = (1'h0); (forvar2035 < (2'h3)); forvar2035 = (forvar2035 + (1'h1)))
                    begin
                      reg2036 <= ($signed({$signed(reg1967)}) * reg1986[(2'h2):(2'h2)]);
                    end
                  if ($signed(((~|$unsigned(wire1924)) ?
                      {$signed((8'h9e))} : reg1960)))
                    begin
                      reg2037 <= (({((8'hb4) || (8'hb7))} ?
                              forvar1948[(1'h0):(1'h0)] : $unsigned((reg2005 ?
                                  forvar2025 : (8'hb0)))) ?
                          $signed(reg2031) : forvar1930[(3'h6):(3'h5)]);
                      reg2038 <= reg2026[(2'h2):(2'h2)];
                      reg2039 <= ($signed(((reg1935 ?
                              (8'ha4) : (8'haa)) ~^ (forvar2025 ?
                              reg2006 : reg1966))) ?
                          reg1979 : $signed(reg1994[(3'h4):(3'h4)]));
                    end
                  else
                    begin
                      reg2037 <= forvar2007;
                    end
                end
              else
                begin
                  reg2035 <= $signed($unsigned($unsigned($unsigned(forvar1959))));
                  if ($unsigned((^~({(8'hb7)} ?
                      forvar1934[(1'h0):(1'h0)] : $unsigned(reg1981)))))
                    begin
                      reg2036 <= forvar2001;
                    end
                  else
                    begin
                      reg2036 <= ($unsigned(reg2003) ?
                          $unsigned($unsigned({reg1935})) : $signed($signed({reg1978})));
                    end
                end
            end
          for (forvar2040 = (1'h0); (forvar2040 < (2'h3)); forvar2040 = (forvar2040 + (1'h1)))
            begin
              if (($unsigned($signed((reg1968 ?
                  reg1987 : forvar2013))) << (reg1980 * ((forvar2025 >>> reg1992) && $signed((8'h9f))))))
                begin
                  if (({$unsigned((reg1985 >= reg1978))} ? (8'hb7) : {reg1991}))
                    begin
                      reg2041 <= reg1970[(4'hb):(4'hb)];
                      reg2042 <= reg2001;
                      reg2043 <= reg1979[(4'h9):(1'h0)];
                      reg2044 <= reg1960;
                    end
                  else
                    begin
                      reg2041 <= reg2012;
                      reg2042 <= reg1963;
                      reg2043 <= reg1931[(2'h2):(2'h2)];
                    end
                  reg2045 <= forvar1999[(2'h3):(2'h3)];
                end
              else
                begin
                  for (forvar2041 = (1'h0); (forvar2041 < (1'h0)); forvar2041 = (forvar2041 + (1'h1)))
                    begin
                      reg2042 <= (~^$unsigned(forvar1991[(1'h1):(1'h0)]));
                      reg2043 <= reg1953[(3'h7):(3'h4)];
                    end
                end
              reg2046 <= reg2034[(1'h1):(1'h0)];
            end
        end
      if (reg1978)
        begin
          for (forvar2047 = (1'h0); (forvar2047 < (1'h0)); forvar2047 = (forvar2047 + (1'h1)))
            begin
              for (forvar2048 = (1'h0); (forvar2048 < (2'h2)); forvar2048 = (forvar2048 + (1'h1)))
                begin
                  for (forvar2049 = (1'h0); (forvar2049 < (2'h3)); forvar2049 = (forvar2049 + (1'h1)))
                    begin
                      reg2050 <= forvar1999[(1'h1):(1'h1)];
                    end
                end
            end
          for (forvar2051 = (1'h0); (forvar2051 < (1'h0)); forvar2051 = (forvar2051 + (1'h1)))
            begin
              for (forvar2052 = (1'h0); (forvar2052 < (2'h3)); forvar2052 = (forvar2052 + (1'h1)))
                begin
                  for (forvar2053 = (1'h0); (forvar2053 < (2'h3)); forvar2053 = (forvar2053 + (1'h1)))
                    begin
                      reg2054 <= ((reg1974 - reg1971) <<< (~^(&reg1970)));
                      reg2055 <= (|$unsigned(({(8'ha4)} != (8'ha3))));
                      reg2056 <= reg2037[(4'h8):(3'h4)];
                      reg2057 <= {$signed(reg1965)};
                    end
                  for (forvar2058 = (1'h0); (forvar2058 < (1'h0)); forvar2058 = (forvar2058 + (1'h1)))
                    begin
                      reg2059 <= reg2055;
                    end
                  if (($unsigned(((reg2013 ?
                      (8'ha0) : reg2027) <= {forvar2013})) - {({wire1927} < (reg2012 ?
                          reg2026 : reg1997))}))
                    begin
                      reg2060 <= reg2005[(3'h6):(3'h4)];
                      reg2061 <= (|($unsigned((~(8'hb9))) == (forvar2051[(1'h1):(1'h1)] ?
                          $unsigned(reg2005) : (reg2003 ?
                              forvar2022 : reg1984))));
                    end
                  else
                    begin
                      reg2060 <= $unsigned(reg1936);
                      reg2061 <= ($unsigned((~(forvar1930 ?
                          reg2036 : forvar1959))) < ((^reg1954) ?
                          (^~{forvar2035}) : reg1958[(3'h5):(3'h5)]));
                    end
                  for (forvar2062 = (1'h0); (forvar2062 < (1'h1)); forvar2062 = (forvar2062 + (1'h1)))
                    begin
                      reg2063 <= $unsigned((reg2015[(4'hd):(3'h7)] ?
                          ({reg1958} ?
                              {reg1938} : reg2059) : ($unsigned((8'hab)) <= (reg2002 ?
                              reg1954 : reg2045))));
                      reg2064 <= reg2020[(3'h7):(1'h0)];
                    end
                end
            end
          for (forvar2065 = (1'h0); (forvar2065 < (1'h1)); forvar2065 = (forvar2065 + (1'h1)))
            begin
              for (forvar2066 = (1'h0); (forvar2066 < (2'h2)); forvar2066 = (forvar2066 + (1'h1)))
                begin
                  if (((($unsigned(reg2003) << (^~reg2039)) ?
                      reg2013[(2'h2):(1'h1)] : reg1997[(4'hd):(1'h1)]) ~^ $signed((~forvar2066))))
                    begin
                      reg2067 <= $signed(((8'ha2) ?
                          ($unsigned(forvar1939) ?
                              (reg2000 > reg1969) : wire1925) : ({(8'ha8)} ?
                              (reg1937 ?
                                  (8'h9d) : reg1993) : $unsigned(reg1962))));
                      reg2068 <= $unsigned(($signed((^~forvar1939)) ?
                          $unsigned($signed(reg1990)) : $signed(forvar1939[(4'h9):(3'h7)])));
                      reg2069 <= ($signed(reg2003[(2'h2):(1'h1)]) ?
                          $unsigned($unsigned(reg1974)) : (^~((forvar2001 == forvar1930) ?
                              forvar1971[(1'h1):(1'h1)] : $unsigned(reg2020))));
                    end
                  else
                    begin
                      reg2067 <= {(8'ha0)};
                      reg2068 <= ((reg2006 & (((8'ha3) ?
                              reg1984 : reg1960) << $signed(forvar1943))) ?
                          reg1961[(1'h1):(1'h1)] : (~&reg1955));
                      reg2069 <= ({((^forvar1943) || (~forvar1941))} >> (8'ha1));
                      reg2070 <= $signed($signed({((8'hb9) > forvar1980)}));
                    end
                  if ($signed((+forvar2023)))
                    begin
                      reg2071 <= (!((~&reg1992) ?
                          forvar1998[(3'h6):(1'h1)] : (^~reg1933)));
                      reg2072 <= reg1933;
                      reg2073 <= $signed(forvar2065[(3'h4):(2'h3)]);
                      reg2074 <= reg2070;
                    end
                  else
                    begin
                      reg2071 <= $signed(($signed((forvar1976 ~^ reg1953)) ?
                          ($signed(forvar1948) ?
                              reg2057 : (forvar1983 ?
                                  reg2067 : forvar2047)) : $unsigned((forvar2040 ?
                              reg2059 : wire1927))));
                      reg2072 <= $unsigned(($signed($signed(reg1951)) ?
                          $unsigned(reg2059) : (reg1962 - (&reg2018))));
                      reg2073 <= {(&($unsigned(forvar1962) ?
                              (forvar1971 ?
                                  reg2025 : forvar2015) : (reg2016 && forvar1930)))};
                    end
                  for (forvar2075 = (1'h0); (forvar2075 < (2'h2)); forvar2075 = (forvar2075 + (1'h1)))
                    begin
                      reg2076 <= $signed({forvar2011});
                      reg2077 <= (({{reg1938}} > reg1929[(5'h10):(4'hd)]) >>> $unsigned((-(^~(8'ha4)))));
                    end
                  for (forvar2078 = (1'h0); (forvar2078 < (1'h0)); forvar2078 = (forvar2078 + (1'h1)))
                    begin
                      reg2079 <= (^reg2055[(2'h2):(2'h2)]);
                    end
                end
              reg2080 <= (+forvar2065);
            end
        end
      else
        begin
          reg2047 <= $unsigned($signed($unsigned((wire1924 ?
              forvar1930 : forvar2053))));
          for (forvar2048 = (1'h0); (forvar2048 < (2'h2)); forvar2048 = (forvar2048 + (1'h1)))
            begin
              for (forvar2049 = (1'h0); (forvar2049 < (1'h0)); forvar2049 = (forvar2049 + (1'h1)))
                begin
                  for (forvar2050 = (1'h0); (forvar2050 < (2'h2)); forvar2050 = (forvar2050 + (1'h1)))
                    begin
                      reg2051 <= ($unsigned((~&((8'h9d) ?
                          reg1936 : forvar2041))) >> (reg1984 ?
                          $unsigned((~^forvar1971)) : ($unsigned(reg1988) ^~ forvar1980)));
                      reg2052 <= {{($signed(forvar1970) & (-reg2041))}};
                      reg2053 <= ((8'ha0) == $unsigned(reg1971[(1'h1):(1'h0)]));
                    end
                  if ($signed((($signed(reg2009) ?
                          $unsigned(reg1953) : (reg1966 ? reg1991 : (8'ha4))) ?
                      (~(forvar1930 ?
                          reg1934 : (8'hb6))) : $signed($unsigned(reg2055)))))
                    begin
                      reg2054 <= reg2047;
                      reg2055 <= ((^$signed({reg1948})) ?
                          (forvar1999 > (8'had)) : forvar1967[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg2054 <= (forvar1934[(1'h0):(1'h0)] ?
                          {(((8'ha3) >> reg2003) <= (~forvar1933))} : reg2015[(1'h0):(1'h0)]);
                      reg2055 <= reg1978;
                      reg2056 <= forvar2066[(1'h0):(1'h0)];
                      reg2057 <= $signed($signed($signed($unsigned(reg2031))));
                    end
                end
              reg2058 <= $unsigned(forvar2035[(3'h5):(2'h2)]);
            end
        end
      reg2081 <= {(&reg1972)};
    end
  always
    @(posedge clk) begin
      for (forvar2082 = (1'h0); (forvar2082 < (1'h0)); forvar2082 = (forvar2082 + (1'h1)))
        begin
          for (forvar2083 = (1'h0); (forvar2083 < (2'h2)); forvar2083 = (forvar2083 + (1'h1)))
            begin
              if (($signed((~|(reg1932 ? reg1955 : reg1947))) ?
                  $unsigned($unsigned($unsigned((8'ha1)))) : (&(-((8'hb3) >= reg1978)))))
                begin
                  for (forvar2084 = (1'h0); (forvar2084 < (2'h3)); forvar2084 = (forvar2084 + (1'h1)))
                    begin
                      reg2085 <= {$signed($signed(reg1944))};
                      reg2086 <= reg2034[(1'h0):(1'h0)];
                      reg2087 <= {(reg2038 ? (~&$signed(reg2003)) : reg2056)};
                    end
                  if ($unsigned(reg2019))
                    begin
                      reg2088 <= wire1928;
                    end
                  else
                    begin
                      reg2088 <= forvar2030[(4'ha):(4'h9)];
                      reg2089 <= $unsigned((reg1991[(2'h3):(1'h0)] ?
                          ((reg1951 ^~ reg2045) ?
                              (wire1925 ?
                                  reg2018 : (8'ha7)) : {reg1996}) : forvar2075[(2'h3):(2'h3)]));
                      reg2090 <= (reg1955[(4'hf):(4'ha)] < (8'hba));
                    end
                  for (forvar2091 = (1'h0); (forvar2091 < (2'h2)); forvar2091 = (forvar2091 + (1'h1)))
                    begin
                      reg2092 <= (~$unsigned(($unsigned(reg2047) <= (reg2051 ?
                          reg1977 : reg1940))));
                    end
                end
              else
                begin
                  if ($unsigned((reg2003 ^ $signed({forvar2051}))))
                    begin
                      reg2084 <= ($signed($unsigned($unsigned(reg2008))) ?
                          ($unsigned((!reg1985)) > ($signed(reg1940) << (8'ha3))) : (+$signed(reg1929[(3'h7):(2'h2)])));
                      reg2085 <= $unsigned((($unsigned(reg2034) << {reg2085}) ?
                          ($signed(reg2006) ?
                              {reg2085} : reg1982[(4'h8):(3'h4)]) : reg1938[(3'h7):(2'h2)]));
                    end
                  else
                    begin
                      reg2084 <= $unsigned(reg2045);
                      reg2085 <= $signed(reg2061);
                    end
                  for (forvar2086 = (1'h0); (forvar2086 < (2'h2)); forvar2086 = (forvar2086 + (1'h1)))
                    begin
                      reg2087 <= (($signed((forvar2086 ?
                              forvar1971 : (8'hb6))) >>> (((8'ha3) ?
                                  reg1963 : reg1949) ?
                              $unsigned(reg2085) : {(8'ha6)})) ?
                          $signed(((wire1925 ?
                              reg2092 : (8'hb2)) <= (reg1971 - (8'hba)))) : reg1944);
                      reg2088 <= ({$unsigned(reg2045)} ?
                          $unsigned(reg2059) : (8'ha6));
                    end
                  if (reg2032)
                    begin
                      reg2089 <= (-($unsigned({forvar2030}) > reg2056));
                      reg2090 <= (~reg1978[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg2089 <= forvar2051[(4'hc):(4'hb)];
                      reg2090 <= forvar2041;
                    end
                  if ($unsigned(reg2054[(2'h2):(1'h1)]))
                    begin
                      reg2091 <= {{reg2005[(4'hd):(2'h3)]}};
                      reg2092 <= ((~^(^~reg1975)) && $signed((-(reg2085 > reg2051))));
                      reg2093 <= forvar2048;
                      reg2094 <= $unsigned(reg2052[(3'h6):(3'h5)]);
                    end
                  else
                    begin
                      reg2091 <= reg2053[(4'hb):(4'h8)];
                    end
                end
              for (forvar2095 = (1'h0); (forvar2095 < (1'h1)); forvar2095 = (forvar2095 + (1'h1)))
                begin
                  for (forvar2096 = (1'h0); (forvar2096 < (1'h1)); forvar2096 = (forvar2096 + (1'h1)))
                    begin
                      reg2097 <= $unsigned(forvar1936[(1'h0):(1'h0)]);
                    end
                  reg2098 <= ($signed(reg2029) << ({forvar2015[(3'h4):(2'h3)]} ?
                      reg2046[(1'h0):(1'h0)] : $signed((reg2087 != (8'hb3)))));
                  reg2099 <= forvar1980[(1'h1):(1'h1)];
                end
            end
          for (forvar2100 = (1'h0); (forvar2100 < (2'h3)); forvar2100 = (forvar2100 + (1'h1)))
            begin
              if ({reg2024[(2'h3):(2'h2)]})
                begin
                  reg2101 <= reg1939;
                  for (forvar2102 = (1'h0); (forvar2102 < (1'h0)); forvar2102 = (forvar2102 + (1'h1)))
                    begin
                      reg2103 <= {(reg2086[(1'h0):(1'h0)] != (~{reg1939}))};
                      reg2104 <= $signed($signed($signed($signed(forvar2078))));
                      reg2105 <= ($unsigned(((~reg1961) > (~|reg2010))) != (^~$unsigned((forvar1983 ?
                          (8'h9f) : forvar2052))));
                    end
                  for (forvar2106 = (1'h0); (forvar2106 < (1'h0)); forvar2106 = (forvar2106 + (1'h1)))
                    begin
                      reg2107 <= forvar2102[(1'h1):(1'h0)];
                      reg2108 <= (reg2041[(4'ha):(2'h3)] ?
                          $signed(reg2087[(1'h1):(1'h0)]) : (reg1931 ?
                              (|(~|reg2036)) : reg2070));
                      reg2109 <= $unsigned($signed($unsigned((-reg1989))));
                    end
                  reg2110 <= (-(~&$signed((8'hb2))));
                end
              else
                begin
                  reg2101 <= {reg2092[(4'hb):(3'h7)]};
                  reg2102 <= ($signed($signed((^(8'h9c)))) ^~ reg2097);
                  for (forvar2103 = (1'h0); (forvar2103 < (2'h3)); forvar2103 = (forvar2103 + (1'h1)))
                    begin
                      reg2104 <= (~^(reg1984[(1'h1):(1'h1)] ?
                          $unsigned((^(8'hab))) : (^~reg2050[(4'hb):(1'h0)])));
                      reg2105 <= ((|$unsigned(((8'hb4) < reg2021))) >= $signed(wire1925[(2'h3):(1'h1)]));
                    end
                end
              for (forvar2111 = (1'h0); (forvar2111 < (1'h0)); forvar2111 = (forvar2111 + (1'h1)))
                begin
                  reg2112 <= (~|reg2010);
                  if ({(reg1982 && {$signed(reg1960)})})
                    begin
                      reg2113 <= $unsigned((!reg2076[(4'hc):(2'h3)]));
                    end
                  else
                    begin
                      reg2113 <= ($unsigned({$unsigned(reg1995)}) ^ (forvar1971 ?
                          $unsigned($signed(reg1981)) : forvar1931));
                    end
                  reg2114 <= (8'ha2);
                end
            end
          for (forvar2115 = (1'h0); (forvar2115 < (2'h2)); forvar2115 = (forvar2115 + (1'h1)))
            begin
              if ($signed($unsigned($unsigned(reg2013[(3'h4):(1'h1)]))))
                begin
                  for (forvar2116 = (1'h0); (forvar2116 < (1'h1)); forvar2116 = (forvar2116 + (1'h1)))
                    begin
                      reg2117 <= reg1946[(3'h5):(3'h4)];
                      reg2118 <= forvar2023;
                    end
                  for (forvar2119 = (1'h0); (forvar2119 < (1'h1)); forvar2119 = (forvar2119 + (1'h1)))
                    begin
                      reg2120 <= forvar2015[(3'h6):(1'h1)];
                      reg2121 <= reg1974;
                    end
                  for (forvar2122 = (1'h0); (forvar2122 < (2'h2)); forvar2122 = (forvar2122 + (1'h1)))
                    begin
                      reg2123 <= reg2113;
                    end
                  for (forvar2124 = (1'h0); (forvar2124 < (2'h2)); forvar2124 = (forvar2124 + (1'h1)))
                    begin
                      reg2125 <= reg2063;
                    end
                end
              else
                begin
                  for (forvar2116 = (1'h0); (forvar2116 < (2'h2)); forvar2116 = (forvar2116 + (1'h1)))
                    begin
                      reg2117 <= (^~{((8'hab) < (forvar2122 ?
                              reg2070 : forvar2066))});
                      reg2118 <= (|((reg2105[(2'h3):(2'h2)] ~^ (^wire1927)) | forvar2115));
                      reg2119 <= $signed(((reg2063 ?
                          $signed((8'hb6)) : $unsigned(reg2027)) < ($signed((8'hb9)) ?
                          (reg2071 ?
                              forvar1956 : forvar1943) : $signed((8'h9c)))));
                      reg2120 <= $unsigned((|(8'hac)));
                    end
                end
              if ((8'hae))
                begin
                  for (forvar2126 = (1'h0); (forvar2126 < (1'h0)); forvar2126 = (forvar2126 + (1'h1)))
                    begin
                      reg2127 <= reg2125;
                    end
                  for (forvar2128 = (1'h0); (forvar2128 < (2'h3)); forvar2128 = (forvar2128 + (1'h1)))
                    begin
                      reg2129 <= reg1951;
                      reg2130 <= {(reg2094 ?
                              (!(reg1932 ?
                                  forvar2030 : forvar2013)) : reg1993)};
                      reg2131 <= reg1958[(3'h6):(3'h5)];
                    end
                end
              else
                begin
                  reg2126 <= ((~&forvar1962[(3'h6):(3'h6)]) ?
                      {$signed($signed(reg1929))} : reg1952);
                  for (forvar2127 = (1'h0); (forvar2127 < (2'h2)); forvar2127 = (forvar2127 + (1'h1)))
                    begin
                      reg2128 <= (+reg2069[(2'h2):(1'h0)]);
                    end
                  if ((+reg2113[(2'h2):(1'h1)]))
                    begin
                      reg2129 <= (~($signed(reg2094) ?
                          $signed($signed((8'ha1))) : ($unsigned(reg2054) ?
                              (reg2092 * reg1977) : {reg2129})));
                      reg2130 <= $unsigned((reg2125[(1'h1):(1'h1)] ?
                          forvar1998 : forvar1970));
                      reg2131 <= (($signed({reg1981}) | (reg2056[(1'h1):(1'h1)] ?
                              (reg2103 ? forvar2035 : reg2080) : (forvar2100 ?
                                  reg2032 : forvar1967))) ?
                          (((reg1937 << forvar1980) ?
                                  $unsigned(forvar2025) : reg2114) ?
                              reg2047[(1'h1):(1'h0)] : (forvar2048[(2'h2):(1'h1)] ?
                                  ((8'ha0) ?
                                      reg1937 : forvar2011) : (-reg2127))) : $unsigned($unsigned($unsigned((8'hb9)))));
                    end
                  else
                    begin
                      reg2129 <= ($signed(forvar2128) + forvar2013[(3'h5):(3'h4)]);
                    end
                end
              for (forvar2132 = (1'h0); (forvar2132 < (1'h0)); forvar2132 = (forvar2132 + (1'h1)))
                begin
                  for (forvar2133 = (1'h0); (forvar2133 < (2'h3)); forvar2133 = (forvar2133 + (1'h1)))
                    begin
                      reg2134 <= (-(~|($unsigned(reg2126) ?
                          (reg2109 > reg2029) : reg2069)));
                      reg2135 <= (reg2121 ? reg2126 : (+{$signed((8'hb4))}));
                    end
                  for (forvar2136 = (1'h0); (forvar2136 < (1'h1)); forvar2136 = (forvar2136 + (1'h1)))
                    begin
                      reg2137 <= reg2002[(3'h6):(3'h5)];
                      reg2138 <= reg2012;
                    end
                  if ($unsigned(reg2088))
                    begin
                      reg2139 <= forvar1962;
                      reg2140 <= $unsigned((forvar2128 ?
                          $signed((^reg2102)) : (reg2137 ?
                              $signed((8'hb4)) : (&wire1924))));
                      reg2141 <= $unsigned(reg2026[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg2139 <= $signed($signed(forvar2001));
                      reg2140 <= $unsigned($signed($signed((8'hab))));
                      reg2141 <= forvar2116;
                    end
                  reg2142 <= (^~forvar1976[(2'h2):(2'h2)]);
                end
            end
        end
      if ($signed($unsigned(($unsigned(reg2059) ? reg1971 : $signed((8'hb2))))))
        begin
          for (forvar2143 = (1'h0); (forvar2143 < (1'h0)); forvar2143 = (forvar2143 + (1'h1)))
            begin
              for (forvar2144 = (1'h0); (forvar2144 < (2'h2)); forvar2144 = (forvar2144 + (1'h1)))
                begin
                  for (forvar2145 = (1'h0); (forvar2145 < (1'h1)); forvar2145 = (forvar2145 + (1'h1)))
                    begin
                      reg2146 <= $unsigned((({reg1977} ?
                              reg2071[(1'h0):(1'h0)] : (-forvar2001)) ?
                          (8'h9f) : (((8'ha3) ? reg2036 : reg1961) ?
                              $signed(forvar2040) : (forvar2030 == reg1985))));
                      reg2147 <= (8'ha6);
                      reg2148 <= (^~$unsigned(reg2009[(4'h9):(2'h2)]));
                    end
                  if ($unsigned($unsigned((!$unsigned(forvar1934)))))
                    begin
                      reg2149 <= reg2107;
                      reg2150 <= reg1983;
                      reg2151 <= (&(reg2041[(3'h5):(1'h0)] >>> (((8'hb6) ^~ reg2025) ?
                          (~^reg2001) : (!reg1947))));
                      reg2152 <= ($unsigned($unsigned((8'hb5))) > $signed((8'hb6)));
                    end
                  else
                    begin
                      reg2149 <= (reg2069 >= ($signed(forvar1939[(3'h4):(2'h3)]) || ((|reg2089) * (forvar2015 ?
                          forvar2095 : reg2038))));
                      reg2150 <= forvar2052[(4'hd):(4'hd)];
                      reg2151 <= (reg2098 ?
                          $unsigned(((+reg2020) ?
                              {reg2053} : reg1983[(2'h2):(1'h0)])) : $unsigned((~&(forvar2133 ^~ reg1981))));
                      reg2152 <= (reg2130[(1'h1):(1'h1)] ?
                          $signed((~|{forvar1980})) : $signed(reg2005[(4'hc):(1'h0)]));
                    end
                  for (forvar2153 = (1'h0); (forvar2153 < (1'h1)); forvar2153 = (forvar2153 + (1'h1)))
                    begin
                      reg2154 <= (8'hb0);
                      reg2155 <= {((reg2118[(1'h0):(1'h0)] ?
                                  reg2056 : $signed(reg1989)) ?
                              reg1963 : (+{forvar2127}))};
                      reg2156 <= ({$signed((wire1924 ?
                              forvar2132 : reg1980))} | ((!{reg2079}) == {(reg2034 ?
                              forvar1936 : reg2151)}));
                    end
                  for (forvar2157 = (1'h0); (forvar2157 < (1'h0)); forvar2157 = (forvar2157 + (1'h1)))
                    begin
                      reg2158 <= (8'ha4);
                      reg2159 <= ((8'ha9) - $signed($unsigned((^forvar2035))));
                      reg2160 <= $unsigned(reg1975[(1'h0):(1'h0)]);
                    end
                end
              reg2161 <= reg2108[(1'h1):(1'h1)];
            end
        end
      else
        begin
          for (forvar2143 = (1'h0); (forvar2143 < (2'h2)); forvar2143 = (forvar2143 + (1'h1)))
            begin
              for (forvar2144 = (1'h0); (forvar2144 < (2'h3)); forvar2144 = (forvar2144 + (1'h1)))
                begin
                  for (forvar2145 = (1'h0); (forvar2145 < (1'h0)); forvar2145 = (forvar2145 + (1'h1)))
                    begin
                      reg2146 <= (forvar2078[(2'h3):(1'h0)] == {$signed(reg2120[(4'h9):(1'h1)])});
                    end
                  reg2147 <= (^$unsigned(reg1936[(1'h0):(1'h0)]));
                end
            end
        end
      if ((reg1990[(2'h3):(1'h0)] != (^~($signed(forvar2040) || reg2130[(2'h2):(2'h2)]))))
        begin
          if (($signed(reg2131) << $unsigned(($unsigned((8'hb7)) ?
              reg2128 : reg2141[(4'hc):(2'h3)]))))
            begin
              reg2162 <= ((forvar2133 ^ (&{reg1967})) ?
                  ($unsigned(forvar2052[(4'ha):(1'h1)]) ?
                      reg1931[(2'h2):(1'h0)] : ({reg1982} >>> (~reg2117))) : (8'ha8));
              for (forvar2163 = (1'h0); (forvar2163 < (2'h3)); forvar2163 = (forvar2163 + (1'h1)))
                begin
                  for (forvar2164 = (1'h0); (forvar2164 < (2'h2)); forvar2164 = (forvar2164 + (1'h1)))
                    begin
                      reg2165 <= $unsigned($unsigned((reg1954[(3'h5):(2'h2)] ?
                          ((8'hb5) ~^ forvar2011) : {reg2138})));
                    end
                  for (forvar2166 = (1'h0); (forvar2166 < (1'h0)); forvar2166 = (forvar2166 + (1'h1)))
                    begin
                      reg2167 <= (($signed({reg2085}) >> (~^((8'ha7) == forvar2115))) ?
                          $signed($unsigned(forvar2119[(1'h1):(1'h0)])) : $unsigned((forvar1967 ?
                              reg2025 : $unsigned((8'hba)))));
                      reg2168 <= reg2069;
                      reg2169 <= ($signed($unsigned($signed((8'ha4)))) && reg2000);
                    end
                  if (($signed(reg2010) ?
                      ({$signed(forvar1963)} >= {forvar2015[(3'h6):(3'h6)]}) : ($unsigned(((8'hb3) - reg2067)) ~^ reg2020)))
                    begin
                      reg2170 <= reg1961;
                      reg2171 <= {(((reg2063 ? reg2091 : reg1987) ?
                                  (|forvar1948) : forvar1947) ?
                              ($signed(reg1978) == (reg2118 ?
                                  forvar2163 : reg2086)) : {$signed(forvar2163)})};
                    end
                  else
                    begin
                      reg2170 <= $signed($unsigned((~|$unsigned((8'hb5)))));
                    end
                  reg2172 <= (((-(forvar2013 ?
                      (8'ha2) : reg2161)) - reg2058[(2'h3):(1'h0)]) ~^ ((-reg2036[(1'h1):(1'h0)]) ?
                      (^~reg1961[(1'h1):(1'h1)]) : ((forvar1939 ?
                          reg2027 : forvar2049) <<< (forvar1947 ^~ forvar1963))));
                end
              for (forvar2173 = (1'h0); (forvar2173 < (1'h1)); forvar2173 = (forvar2173 + (1'h1)))
                begin
                  for (forvar2174 = (1'h0); (forvar2174 < (1'h1)); forvar2174 = (forvar2174 + (1'h1)))
                    begin
                      reg2175 <= (reg2099[(3'h6):(3'h4)] < (forvar2004 ?
                          {reg1993[(1'h0):(1'h0)]} : ((&forvar1947) ?
                              forvar2051[(4'hb):(1'h1)] : (reg1966 ?
                                  reg1932 : (8'hab)))));
                      reg2176 <= reg2021;
                      reg2177 <= {(-(reg1940 <= wire1926))};
                      reg2178 <= ($signed(forvar2136) & $signed((~|(-forvar2084))));
                    end
                  for (forvar2179 = (1'h0); (forvar2179 < (2'h3)); forvar2179 = (forvar2179 + (1'h1)))
                    begin
                      reg2180 <= reg1933;
                      reg2181 <= (($signed((8'hb5)) ?
                          reg2045[(3'h5):(1'h1)] : $signed(reg2073[(3'h4):(3'h4)])) > reg1942[(4'h8):(3'h7)]);
                      reg2182 <= $signed({((~|(8'ha5)) - (~^forvar2157))});
                      reg2183 <= reg2176;
                    end
                  if ((-($unsigned((reg2051 ?
                      (8'ha0) : forvar2102)) >> {$unsigned(reg2071)})))
                    begin
                      reg2184 <= reg2042;
                      reg2185 <= reg1965[(4'h9):(1'h0)];
                      reg2186 <= $unsigned({(~^(~&reg2020))});
                      reg2187 <= $signed((((forvar1934 ? (8'hb6) : wire1924) ?
                              $signed(forvar2007) : $unsigned(forvar2133)) ?
                          {reg2142} : ($unsigned(forvar2100) ^ {reg1935})));
                    end
                  else
                    begin
                      reg2184 <= ($signed($signed($unsigned(reg2130))) ?
                          (^$signed($unsigned((8'haa)))) : (8'had));
                      reg2185 <= reg2154[(2'h3):(1'h0)];
                      reg2186 <= reg1978[(4'h9):(3'h4)];
                      reg2187 <= forvar1930[(3'h5):(3'h5)];
                    end
                  reg2188 <= $signed(reg2051[(3'h4):(3'h4)]);
                end
            end
          else
            begin
              for (forvar2162 = (1'h0); (forvar2162 < (1'h1)); forvar2162 = (forvar2162 + (1'h1)))
                begin
                  reg2163 <= (~|$unsigned((~|reg2125[(1'h1):(1'h1)])));
                  for (forvar2164 = (1'h0); (forvar2164 < (1'h1)); forvar2164 = (forvar2164 + (1'h1)))
                    begin
                      reg2165 <= $signed((8'haf));
                      reg2166 <= $signed(forvar1948[(3'h6):(3'h6)]);
                    end
                end
              for (forvar2167 = (1'h0); (forvar2167 < (2'h2)); forvar2167 = (forvar2167 + (1'h1)))
                begin
                  for (forvar2168 = (1'h0); (forvar2168 < (2'h3)); forvar2168 = (forvar2168 + (1'h1)))
                    begin
                      reg2169 <= ((8'ha5) ?
                          $unsigned(((reg2131 && reg2085) == (reg2110 == reg2079))) : (reg2027 ?
                              $signed((-forvar2051)) : forvar2052[(4'h9):(3'h6)]));
                      reg2170 <= {(8'hb2)};
                    end
                  reg2171 <= $unsigned(reg1982[(1'h0):(1'h0)]);
                  for (forvar2172 = (1'h0); (forvar2172 < (2'h3)); forvar2172 = (forvar2172 + (1'h1)))
                    begin
                      reg2173 <= reg1988;
                      reg2174 <= ((((8'h9e) ?
                              $unsigned(reg2156) : reg1934[(2'h3):(2'h2)]) + reg2038[(2'h3):(2'h2)]) ?
                          $unsigned((~&reg2026[(1'h1):(1'h1)])) : $unsigned({(reg2076 ?
                                  forvar2083 : forvar1934)}));
                      reg2175 <= $unsigned(reg2097[(1'h1):(1'h0)]);
                      reg2176 <= forvar2062;
                    end
                  for (forvar2177 = (1'h0); (forvar2177 < (2'h3)); forvar2177 = (forvar2177 + (1'h1)))
                    begin
                      reg2178 <= (&(reg2005 ?
                          ((reg2102 ? forvar1948 : forvar2132) ?
                              {(8'h9c)} : reg2034) : $unsigned((reg1964 <<< reg2064))));
                      reg2179 <= reg2005[(1'h1):(1'h1)];
                      reg2180 <= forvar1939;
                      reg2181 <= $unsigned(reg1944);
                    end
                end
              if ($unsigned($unsigned(reg2089)))
                begin
                  reg2182 <= reg2042;
                  if ($unsigned({$signed(((8'hae) >>> reg1948))}))
                    begin
                      reg2183 <= $unsigned({$unsigned(forvar2082[(1'h0):(1'h0)])});
                      reg2184 <= $unsigned((reg2018[(4'he):(4'ha)] || ((reg2008 ?
                              (8'hb3) : reg2011) ?
                          (&reg1932) : (forvar2111 == reg2107))));
                    end
                  else
                    begin
                      reg2183 <= (reg1929[(4'hd):(4'h8)] ?
                          (reg2118[(1'h1):(1'h0)] >= $signed((|reg2148))) : {(~|reg2041[(3'h6):(1'h0)])});
                      reg2184 <= $unsigned($signed((reg2019[(2'h2):(2'h2)] ?
                          $unsigned(reg2104) : $unsigned(reg2165))));
                      reg2185 <= ($unsigned(($signed(forvar2048) != (forvar2128 ^ (8'ha8)))) ~^ (8'h9e));
                    end
                  reg2186 <= ($signed((!reg2176[(1'h0):(1'h0)])) ?
                      $unsigned((!((8'ha5) ? reg1953 : reg2086))) : (8'ha1));
                  reg2187 <= ((reg2103 || ($unsigned(reg2109) != $unsigned((8'ha6)))) >> $signed((reg1946 ?
                      reg2185[(1'h0):(1'h0)] : (reg2055 ?
                          forvar2058 : (8'hae)))));
                end
              else
                begin
                  for (forvar2182 = (1'h0); (forvar2182 < (2'h3)); forvar2182 = (forvar2182 + (1'h1)))
                    begin
                      reg2183 <= reg1953[(3'h4):(1'h0)];
                      reg2184 <= $signed((-$unsigned(((8'ha6) ^ reg1996))));
                      reg2185 <= $unsigned($signed((&(reg2080 & reg1940))));
                      reg2186 <= reg2088;
                    end
                  for (forvar2187 = (1'h0); (forvar2187 < (2'h3)); forvar2187 = (forvar2187 + (1'h1)))
                    begin
                      reg2188 <= $signed((+$signed((forvar1959 + reg2057))));
                      reg2189 <= {{((reg2053 >> reg2185) ?
                                  $signed(reg2162) : (~|reg1997))}};
                      reg2190 <= $unsigned({(wire1925 ?
                              (|reg2024) : (reg2126 + reg2067))});
                      reg2191 <= $signed({reg2156});
                    end
                  if (({reg1978[(4'ha):(3'h5)]} && ($signed(reg1954) > (-forvar2086[(3'h6):(3'h5)]))))
                    begin
                      reg2192 <= ($signed($unsigned((wire1924 - forvar2022))) < ($unsigned((reg1942 ?
                          reg2129 : reg2113)) | $signed(reg2008)));
                      reg2193 <= (({reg2127[(1'h0):(1'h0)]} ?
                              {(|(8'hb9))} : $unsigned(reg2051)) ?
                          (reg1929[(5'h10):(2'h2)] ?
                              (forvar2182[(2'h2):(1'h0)] ?
                                  forvar1930[(3'h6):(1'h0)] : $signed(reg2101)) : reg2152) : reg2110[(1'h0):(1'h0)]);
                      reg2194 <= ($signed(reg2031) ? reg1967 : forvar2096);
                      reg2195 <= (~&($signed($signed(reg1994)) << reg1983[(2'h3):(2'h3)]));
                    end
                  else
                    begin
                      reg2192 <= $unsigned(reg2089);
                      reg2193 <= $unsigned((-forvar2066));
                      reg2194 <= (reg1957 ?
                          reg1992[(1'h0):(1'h0)] : $unsigned({(reg2064 + reg2031)}));
                    end
                  for (forvar2196 = (1'h0); (forvar2196 < (2'h2)); forvar2196 = (forvar2196 + (1'h1)))
                    begin
                      reg2197 <= $signed($signed((reg2104 ?
                          (reg1997 ? reg2168 : reg2071) : reg2076)));
                      reg2198 <= $unsigned((~&$unsigned($unsigned(reg2093))));
                      reg2199 <= reg2113[(3'h7):(3'h7)];
                      reg2200 <= forvar2001[(2'h2):(1'h0)];
                    end
                end
              if (reg2118)
                begin
                  for (forvar2201 = (1'h0); (forvar2201 < (1'h1)); forvar2201 = (forvar2201 + (1'h1)))
                    begin
                      reg2202 <= ($unsigned($signed((forvar1983 >>> forvar1983))) + (&$unsigned($unsigned(reg2005))));
                      reg2203 <= wire1925;
                    end
                  if (($signed($signed((|reg2174))) << reg2029))
                    begin
                      reg2204 <= {(reg2068 >= ((reg1948 > reg2150) - (forvar2065 ^ reg2061)))};
                      reg2205 <= forvar2058[(3'h7):(2'h3)];
                      reg2206 <= forvar2115[(4'ha):(3'h5)];
                      reg2207 <= $unsigned({reg2160[(1'h1):(1'h0)]});
                    end
                  else
                    begin
                      reg2204 <= (((forvar2051[(4'hd):(2'h2)] ?
                                  (reg2059 ? reg1950 : reg2099) : forvar1934) ?
                              $signed((reg2038 ^~ (8'hb5))) : $signed((forvar2115 ?
                                  reg2054 : forvar2095))) ?
                          forvar2136[(1'h1):(1'h0)] : reg2019[(4'h8):(1'h0)]);
                      reg2205 <= $unsigned(($signed(reg2150[(1'h1):(1'h1)]) >>> reg1997[(4'ha):(4'h8)]));
                    end
                end
              else
                begin
                  reg2201 <= ($unsigned(reg2206) ?
                      (&$signed(forvar2168)) : $signed((+forvar2174)));
                  if (reg2172[(2'h2):(2'h2)])
                    begin
                      reg2202 <= ($signed(reg1954) >> {$unsigned((^~reg2163))});
                      reg2203 <= (reg1944 ^~ (^~($signed(reg2079) <= (reg2176 ?
                          forvar2065 : forvar1963))));
                      reg2204 <= reg1964;
                    end
                  else
                    begin
                      reg2202 <= (^~(($signed(reg2167) ?
                          (-reg2149) : (reg2055 ?
                              (8'haf) : reg2142)) >> {reg1953}));
                    end
                  for (forvar2205 = (1'h0); (forvar2205 < (2'h3)); forvar2205 = (forvar2205 + (1'h1)))
                    begin
                      reg2206 <= {reg2074};
                      reg2207 <= ($unsigned(((reg2101 <<< forvar2167) & forvar2065)) ?
                          (reg1985 ?
                              {forvar2172[(2'h3):(2'h3)]} : $unsigned(forvar1943)) : $signed(((~|reg2047) ?
                              ((8'hac) == forvar2075) : $unsigned(reg2141))));
                    end
                  for (forvar2208 = (1'h0); (forvar2208 < (2'h3)); forvar2208 = (forvar2208 + (1'h1)))
                    begin
                      reg2209 <= ($unsigned(({reg2073} << $signed(reg2138))) ^ ({reg2018[(5'h10):(4'hb)]} ?
                          {(|wire1928)} : reg1939));
                    end
                end
            end
          for (forvar2210 = (1'h0); (forvar2210 < (2'h3)); forvar2210 = (forvar2210 + (1'h1)))
            begin
              reg2211 <= (|$unsigned($signed((reg2058 ?
                  (8'hb4) : forvar2030))));
              for (forvar2212 = (1'h0); (forvar2212 < (1'h0)); forvar2212 = (forvar2212 + (1'h1)))
                begin
                  for (forvar2213 = (1'h0); (forvar2213 < (1'h0)); forvar2213 = (forvar2213 + (1'h1)))
                    begin
                      reg2214 <= reg2104[(3'h4):(2'h2)];
                      reg2215 <= $unsigned({{$unsigned((8'ha7))}});
                    end
                  if (forvar2153[(3'h5):(1'h0)])
                    begin
                      reg2216 <= reg2141[(3'h4):(2'h3)];
                      reg2217 <= (((^~(8'ha4)) ?
                          $signed($unsigned(reg2174)) : $signed($signed(wire1924))) + $signed(((reg2014 ?
                              forvar1963 : reg1983) ?
                          (+reg1937) : (&reg2076))));
                      reg2218 <= {((8'h9f) ?
                              reg1972[(1'h1):(1'h0)] : (+$signed(forvar1938)))};
                    end
                  else
                    begin
                      reg2216 <= {reg2003[(2'h2):(1'h0)]};
                      reg2217 <= {reg2085[(1'h0):(1'h0)]};
                      reg2218 <= $unsigned({((forvar2051 ? (8'ha8) : reg2109) ?
                              $unsigned(reg2002) : forvar2177[(2'h3):(2'h3)])});
                    end
                  reg2219 <= (reg2128[(4'h8):(3'h6)] & (($unsigned(reg2121) ?
                          (forvar1936 ?
                              forvar1971 : reg2215) : (reg2001 >> forvar2172)) ?
                      $unsigned($signed(reg2031)) : ((reg2024 ~^ forvar2030) ?
                          forvar2035 : wire1928)));
                end
              if ($unsigned(forvar2065))
                begin
                  if ({$unsigned(($unsigned(reg1975) >>> {reg2172}))})
                    begin
                      reg2220 <= forvar2164[(3'h6):(2'h3)];
                      reg2221 <= forvar2127[(2'h3):(1'h0)];
                      reg2222 <= (^($unsigned($unsigned(reg1976)) ?
                          ({reg1983} ?
                              forvar2187[(3'h7):(3'h6)] : {(8'ha1)}) : ($signed(reg2027) ?
                              (reg2101 > reg2163) : reg2074[(3'h4):(3'h4)])));
                      reg2223 <= (~forvar2086);
                    end
                  else
                    begin
                      reg2220 <= $signed((reg1983[(3'h4):(2'h3)] ?
                          $unsigned($unsigned(reg2112)) : (+reg2172[(4'h9):(1'h0)])));
                      reg2221 <= reg2085;
                      reg2222 <= $unsigned((8'h9e));
                      reg2223 <= ($signed(reg2016[(2'h3):(1'h1)]) && $signed(reg2043[(2'h2):(1'h1)]));
                    end
                end
              else
                begin
                  for (forvar2220 = (1'h0); (forvar2220 < (1'h0)); forvar2220 = (forvar2220 + (1'h1)))
                    begin
                      reg2221 <= ((8'h9d) ^~ (reg1964 << (^~(reg2011 ?
                          forvar2065 : reg2223))));
                      reg2222 <= $unsigned(($signed(reg2079) ?
                          (reg2152 ?
                              $signed(reg2223) : (forvar2119 ?
                                  (8'ha6) : reg2093)) : {(~|(8'haf))}));
                      reg2223 <= ((forvar2048[(1'h0):(1'h0)] ?
                          ($signed(forvar2013) ?
                              (reg1946 == (8'hb1)) : (reg2198 >= reg1952)) : reg2084) ~^ reg2179[(1'h1):(1'h1)]);
                      reg2224 <= (reg2097[(1'h0):(1'h0)] ?
                          (((reg1978 == forvar2033) * {reg2181}) ?
                              $signed((reg2005 ?
                                  forvar2040 : reg1958)) : (^~$signed(reg2034))) : (!{$unsigned(forvar1976)}));
                    end
                  if (reg1990[(1'h0):(1'h0)])
                    begin
                      reg2225 <= $unsigned((((^forvar1938) ?
                              reg1958[(1'h0):(1'h0)] : reg2039) ?
                          $signed($unsigned(reg2072)) : ((reg2080 ?
                                  (8'hb8) : reg2014) ?
                              (!forvar2004) : (|forvar2145))));
                    end
                  else
                    begin
                      reg2225 <= (($signed((~^reg2217)) | (!(reg2182 ~^ forvar2001))) ?
                          $unsigned(((forvar1947 < (8'ha5)) ?
                              $unsigned(forvar2004) : (~forvar2177))) : (&((reg2003 ?
                                  reg1950 : reg2202) ?
                              $signed(reg1941) : $signed(reg2045))));
                    end
                end
              reg2226 <= forvar1991[(1'h1):(1'h1)];
            end
          reg2227 <= reg2034;
        end
      else
        begin
          reg2162 <= {$unsigned(($signed(reg2187) ?
                  reg1937 : reg2057[(4'h9):(1'h1)]))};
          if ($signed(reg2009[(4'hb):(4'hb)]))
            begin
              if (reg1954[(2'h2):(1'h1)])
                begin
                  if ((8'ha7))
                    begin
                      reg2163 <= forvar2053;
                      reg2164 <= (reg2032[(1'h0):(1'h0)] ?
                          (^~forvar2025[(2'h2):(2'h2)]) : reg2025);
                      reg2165 <= forvar2013;
                      reg2166 <= reg2169;
                    end
                  else
                    begin
                      reg2163 <= (|($unsigned((reg2192 ~^ reg2061)) > $signed($unsigned(forvar2095))));
                    end
                end
              else
                begin
                  if ((($unsigned((+reg1964)) ?
                      $unsigned($signed(reg2152)) : reg2054) ^ $signed($signed(reg2134))))
                    begin
                      reg2163 <= (forvar1941 <<< (8'ha3));
                    end
                  else
                    begin
                      reg2163 <= (($unsigned($signed(reg2099)) ?
                              reg2046 : ((reg2039 ^~ reg2099) & (reg1980 ^~ (8'h9f)))) ?
                          {reg2059} : reg2205);
                      reg2164 <= (^~reg2223[(2'h2):(2'h2)]);
                      reg2165 <= (reg2221 ^ ((~((8'ha4) <<< reg2047)) ?
                          $unsigned(reg1976) : reg2163[(1'h0):(1'h0)]));
                      reg2166 <= reg2123[(1'h0):(1'h0)];
                    end
                  reg2167 <= $unsigned({$signed(reg2037[(3'h5):(2'h3)])});
                  if (($signed(($unsigned(reg2090) ?
                          (forvar2163 == forvar2103) : {reg2064})) ?
                      (((reg2223 ?
                              reg2139 : reg1963) >= forvar2075[(2'h3):(2'h3)]) ?
                          {{reg2171}} : reg2114) : $signed($unsigned(forvar2196))))
                    begin
                      reg2168 <= ($signed($signed($signed(reg2094))) > forvar2144[(2'h2):(1'h1)]);
                      reg2169 <= (~^reg1988[(3'h5):(3'h4)]);
                      reg2170 <= reg2119[(1'h0):(1'h0)];
                      reg2171 <= $unsigned((reg2156 ?
                          ((reg1963 < reg2051) ?
                              (reg2114 || reg2218) : reg2088) : ($signed(reg2165) ?
                              (reg2031 == reg1932) : $signed((8'ha0)))));
                    end
                  else
                    begin
                      reg2168 <= ((8'hb3) ? {(8'ha9)} : $signed((8'hb4)));
                      reg2169 <= ($unsigned($signed(reg2036[(1'h1):(1'h0)])) ?
                          forvar2174[(4'hb):(1'h0)] : ($unsigned((reg2185 + forvar2096)) <<< ((reg2169 ?
                                  reg1940 : reg2123) ?
                              ((8'hae) ?
                                  (8'h9d) : reg1954) : $unsigned(forvar2111))));
                      reg2170 <= (-$signed((8'ha9)));
                      reg2171 <= forvar2084[(3'h6):(2'h2)];
                    end
                end
              if (($signed(forvar2028[(2'h3):(1'h1)]) ?
                  reg2188 : $unsigned(reg2035)))
                begin
                  for (forvar2172 = (1'h0); (forvar2172 < (1'h1)); forvar2172 = (forvar2172 + (1'h1)))
                    begin
                      reg2173 <= (reg1969 & $unsigned({{reg2160}}));
                      reg2174 <= (reg2010[(2'h3):(2'h2)] ?
                          (-reg2059[(1'h0):(1'h0)]) : $unsigned($signed($signed(forvar2173))));
                    end
                end
              else
                begin
                  for (forvar2172 = (1'h0); (forvar2172 < (2'h3)); forvar2172 = (forvar2172 + (1'h1)))
                    begin
                      reg2173 <= (|reg2109);
                      reg2174 <= $unsigned(forvar2065);
                    end
                end
            end
          else
            begin
              if (((~|{reg2216[(4'h8):(1'h0)]}) ?
                  (^$signed((8'hb8))) : ($unsigned((reg2063 ?
                      reg2086 : reg1929)) ^~ {{reg2059}})))
                begin
                  reg2163 <= $unsigned((&((forvar1963 ?
                      forvar2208 : reg2171) && (reg2164 ^ reg1980))));
                  for (forvar2164 = (1'h0); (forvar2164 < (2'h2)); forvar2164 = (forvar2164 + (1'h1)))
                    begin
                      reg2165 <= (reg2044 ?
                          reg1944[(2'h2):(2'h2)] : $signed((~|$signed(forvar2162))));
                      reg2166 <= $signed((^forvar2028));
                    end
                end
              else
                begin
                  for (forvar2163 = (1'h0); (forvar2163 < (1'h1)); forvar2163 = (forvar2163 + (1'h1)))
                    begin
                      reg2164 <= reg2201;
                      reg2165 <= $unsigned((8'ha6));
                      reg2166 <= reg2011[(3'h7):(2'h2)];
                      reg2167 <= reg2150;
                    end
                  if ($unsigned((~&(~^forvar1939))))
                    begin
                      reg2168 <= forvar2022[(3'h6):(3'h6)];
                      reg2169 <= reg2057;
                      reg2170 <= ($unsigned(forvar2173[(2'h3):(1'h1)]) ?
                          (~$signed(((8'had) <<< (8'hae)))) : ((^(reg2152 ^~ reg2110)) >> reg2002[(4'h8):(2'h2)]));
                      reg2171 <= reg2165[(3'h6):(3'h4)];
                    end
                  else
                    begin
                      reg2168 <= reg1972;
                      reg2169 <= $signed($signed(((|forvar2103) ?
                          reg2198 : (reg2005 <= reg2058))));
                      reg2170 <= (($unsigned(wire1924[(1'h1):(1'h0)]) ?
                              {(^reg2086)} : ($signed(reg2118) != (~|forvar1948))) ?
                          (~|forvar2132) : reg2164);
                    end
                  for (forvar2172 = (1'h0); (forvar2172 < (1'h0)); forvar2172 = (forvar2172 + (1'h1)))
                    begin
                      reg2173 <= (reg2207[(2'h2):(2'h2)] ?
                          {$signed($unsigned(reg2047))} : forvar2103[(2'h3):(2'h3)]);
                    end
                end
              for (forvar2174 = (1'h0); (forvar2174 < (2'h3)); forvar2174 = (forvar2174 + (1'h1)))
                begin
                  reg2175 <= reg1988[(1'h0):(1'h0)];
                  reg2176 <= forvar2102;
                end
            end
        end
      if (((((forvar2020 ?
              forvar2022 : (8'hab)) >>> forvar2174[(2'h2):(1'h0)]) || reg2074[(1'h1):(1'h1)]) ?
          (($unsigned(reg1979) >>> (&reg1972)) >= ({forvar1939} > forvar2179)) : (8'ha5)))
        begin
          for (forvar2228 = (1'h0); (forvar2228 < (1'h0)); forvar2228 = (forvar2228 + (1'h1)))
            begin
              for (forvar2229 = (1'h0); (forvar2229 < (1'h1)); forvar2229 = (forvar2229 + (1'h1)))
                begin
                  if (reg1950)
                    begin
                      reg2230 <= reg1991;
                      reg2231 <= forvar2213[(2'h3):(1'h1)];
                      reg2232 <= (reg2050 + ((^~reg1949[(1'h1):(1'h1)]) > $signed((|reg2010))));
                    end
                  else
                    begin
                      reg2230 <= ($unsigned(reg1954[(4'h8):(3'h4)]) >> $unsigned(((-reg2146) & reg2172)));
                    end
                  if ($unsigned(($unsigned((forvar2086 && reg1977)) ~^ ((!forvar2047) ?
                      (reg1966 && (8'haf)) : $signed(reg2211)))))
                    begin
                      reg2233 <= $signed(reg2151);
                      reg2234 <= (((~^$signed(forvar2041)) && ({reg2079} ?
                          (^forvar2083) : {reg2080})) ^~ (~&$signed({reg2093})));
                    end
                  else
                    begin
                      reg2233 <= (~&$unsigned(({reg1954} ~^ $unsigned((8'hb7)))));
                      reg2234 <= $signed({$unsigned(reg1965)});
                    end
                  if ($signed({$signed(reg1957[(4'hd):(4'h9)])}))
                    begin
                      reg2235 <= forvar2212[(1'h1):(1'h0)];
                      reg2236 <= $signed((reg2161 ^~ $signed((forvar2091 ?
                          wire1924 : reg2221))));
                    end
                  else
                    begin
                      reg2235 <= reg2177;
                      reg2236 <= ((8'haa) != ((reg1957 * (reg1962 ?
                          forvar2028 : (8'ha9))) >= (reg2119[(2'h2):(1'h1)] ?
                          reg2219 : (~^(8'haa)))));
                      reg2237 <= reg1976;
                    end
                  for (forvar2238 = (1'h0); (forvar2238 < (1'h1)); forvar2238 = (forvar2238 + (1'h1)))
                    begin
                      reg2239 <= {(reg2093 ?
                              ((forvar2212 > (8'hb7)) <= (reg2197 ?
                                  reg2204 : reg2184)) : $signed((reg2006 ?
                                  forvar1930 : reg1938)))};
                      reg2240 <= ($signed(({reg2207} ?
                              (reg2102 ?
                                  reg2074 : forvar2106) : reg2052[(2'h2):(1'h0)])) ?
                          reg1996 : $signed($unsigned(((8'hb4) || reg2094))));
                      reg2241 <= forvar2035[(3'h4):(3'h4)];
                      reg2242 <= ((forvar2187 < $unsigned(forvar1959[(4'ha):(2'h3)])) - reg1939);
                    end
                end
              for (forvar2243 = (1'h0); (forvar2243 < (2'h3)); forvar2243 = (forvar2243 + (1'h1)))
                begin
                  if ({{$signed(reg2091[(1'h1):(1'h1)])}})
                    begin
                      reg2244 <= ({({forvar2052} * reg1940)} ?
                          forvar1941[(1'h0):(1'h0)] : reg2240[(3'h7):(1'h1)]);
                      reg2245 <= ((!reg2079) >= $signed((((8'hb1) ?
                              (8'h9d) : reg2192) ?
                          reg2242 : ((8'hb4) & reg1948))));
                    end
                  else
                    begin
                      reg2244 <= reg1935;
                      reg2245 <= reg2090[(3'h4):(3'h4)];
                      reg2246 <= ($signed(reg2146[(3'h4):(2'h3)]) ?
                          $signed($unsigned($signed(reg2114))) : (&forvar2201[(1'h0):(1'h0)]));
                    end
                end
            end
          for (forvar2247 = (1'h0); (forvar2247 < (2'h3)); forvar2247 = (forvar2247 + (1'h1)))
            begin
              for (forvar2248 = (1'h0); (forvar2248 < (2'h3)); forvar2248 = (forvar2248 + (1'h1)))
                begin
                  reg2249 <= ($signed((8'ha4)) ^~ reg1979[(2'h2):(1'h0)]);
                  for (forvar2250 = (1'h0); (forvar2250 < (1'h1)); forvar2250 = (forvar2250 + (1'h1)))
                    begin
                      reg2251 <= $signed((~&reg1967));
                      reg2252 <= reg1955;
                      reg2253 <= $signed($unsigned($signed((reg2131 ?
                          (8'ha7) : reg2051))));
                      reg2254 <= reg1973[(2'h2):(1'h1)];
                    end
                  for (forvar2255 = (1'h0); (forvar2255 < (1'h1)); forvar2255 = (forvar2255 + (1'h1)))
                    begin
                      reg2256 <= $signed((reg2000 != reg1938[(4'h8):(3'h7)]));
                      reg2257 <= ((reg2029[(4'h8):(1'h0)] + forvar2065[(2'h3):(2'h3)]) ?
                          {(^~$unsigned(reg2090))} : (-(reg2043 ?
                              $signed((8'hb2)) : reg2008[(1'h1):(1'h0)])));
                      reg2258 <= forvar1943[(2'h2):(1'h0)];
                    end
                  if ((($signed(forvar1943[(2'h2):(1'h0)]) ?
                      $signed({forvar2174}) : reg2171[(3'h7):(3'h7)]) - $unsigned($unsigned($signed(wire1925)))))
                    begin
                      reg2259 <= {($signed((reg2088 ? reg2039 : reg2024)) ?
                              (~$unsigned(forvar2103)) : reg1947[(1'h0):(1'h0)])};
                      reg2260 <= forvar1999[(2'h3):(2'h2)];
                      reg2261 <= (wire1925[(3'h5):(3'h5)] && $unsigned((!$unsigned(reg2064))));
                      reg2262 <= $signed($unsigned(reg2071));
                    end
                  else
                    begin
                      reg2259 <= $signed($unsigned((reg2003[(1'h0):(1'h0)] ?
                          (reg2259 > forvar1970) : (|reg2170))));
                      reg2260 <= (&(~(~^reg2182)));
                      reg2261 <= (reg1980 - $unsigned($unsigned({reg2109})));
                    end
                end
            end
          if (reg1991[(4'h8):(3'h5)])
            begin
              for (forvar2263 = (1'h0); (forvar2263 < (2'h3)); forvar2263 = (forvar2263 + (1'h1)))
                begin
                  for (forvar2264 = (1'h0); (forvar2264 < (1'h0)); forvar2264 = (forvar2264 + (1'h1)))
                    begin
                      reg2265 <= $signed($signed(((~^forvar2049) ?
                          reg2112[(3'h4):(2'h2)] : {reg1935})));
                      reg2266 <= ($unsigned(reg1949) + $unsigned(reg2222));
                      reg2267 <= (8'hb7);
                      reg2268 <= (reg2037[(1'h0):(1'h0)] >= $signed(($unsigned(reg1995) >= {(8'hb9)})));
                    end
                  reg2269 <= $unsigned($unsigned(($signed(forvar2040) ?
                      $signed(reg2138) : {(8'hac)})));
                end
            end
          else
            begin
              for (forvar2263 = (1'h0); (forvar2263 < (1'h0)); forvar2263 = (forvar2263 + (1'h1)))
                begin
                  for (forvar2264 = (1'h0); (forvar2264 < (2'h3)); forvar2264 = (forvar2264 + (1'h1)))
                    begin
                      reg2265 <= ((~|(forvar2030 || forvar2040)) << (((reg2089 ?
                                  wire1924 : reg1982) ?
                              {wire1928} : {(8'hae)}) ?
                          {(reg2102 >>> reg2009)} : {{reg2024}}));
                      reg2266 <= ($unsigned((reg2010 <= $unsigned(reg2261))) || $unsigned(reg2090));
                      reg2267 <= reg2230;
                      reg2268 <= (reg2039 + reg1941[(1'h1):(1'h1)]);
                    end
                end
              if ((8'hba))
                begin
                  for (forvar2269 = (1'h0); (forvar2269 < (2'h2)); forvar2269 = (forvar2269 + (1'h1)))
                    begin
                      reg2270 <= (^{{(!reg1992)}});
                    end
                  reg2271 <= $unsigned((-reg2121));
                  reg2272 <= (reg2016 ?
                      ((reg1994 ?
                          reg2195[(4'h8):(3'h4)] : reg2036[(1'h1):(1'h0)]) ^ $unsigned($signed(reg2020))) : reg1957[(4'h8):(2'h2)]);
                end
              else
                begin
                  reg2269 <= ((^reg2204) != ({$signed(forvar2263)} ^ reg2268));
                  for (forvar2270 = (1'h0); (forvar2270 < (2'h2)); forvar2270 = (forvar2270 + (1'h1)))
                    begin
                      reg2271 <= (reg1994 ?
                          ($signed((forvar2115 <<< forvar2220)) ?
                              (reg2202 ?
                                  reg2002 : $signed(reg1936)) : ((reg1938 ?
                                  reg2204 : reg1985) - (forvar1936 > forvar2023))) : reg2085[(3'h7):(3'h7)]);
                      reg2272 <= ((((forvar2023 ? forvar2106 : reg2237) ?
                                  reg2225[(1'h1):(1'h0)] : (~^reg2114)) ?
                              $signed((~^reg1955)) : ((forvar2179 == reg2135) >>> (reg1992 ?
                                  reg1962 : reg2053))) ?
                          reg2125 : ((8'hb7) == $unsigned($unsigned(forvar2020))));
                      reg2273 <= reg2226;
                      reg2274 <= (^~reg2107);
                    end
                end
            end
        end
      else
        begin
          for (forvar2228 = (1'h0); (forvar2228 < (1'h1)); forvar2228 = (forvar2228 + (1'h1)))
            begin
              for (forvar2229 = (1'h0); (forvar2229 < (2'h3)); forvar2229 = (forvar2229 + (1'h1)))
                begin
                  reg2230 <= (!reg2265[(3'h7):(3'h7)]);
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg2147[(4'hb):(3'h4)])
        begin
          reg2275 <= (reg2186 ?
              reg1984[(1'h0):(1'h0)] : ($signed((~reg2035)) ?
                  ((forvar2182 | forvar2264) ?
                      ((8'hb0) ?
                          reg2253 : forvar1934) : forvar2022[(3'h4):(2'h3)]) : $signed((~&reg2088))));
          for (forvar2276 = (1'h0); (forvar2276 < (2'h2)); forvar2276 = (forvar2276 + (1'h1)))
            begin
              reg2277 <= ((&({forvar2050} ?
                      $signed(forvar1962) : (~forvar1931))) ?
                  $signed((~|$signed(forvar2028))) : $unsigned(reg2271[(3'h5):(2'h3)]));
              reg2278 <= ((8'hba) >> $unsigned((^~(!reg2185))));
            end
          for (forvar2279 = (1'h0); (forvar2279 < (2'h2)); forvar2279 = (forvar2279 + (1'h1)))
            begin
              for (forvar2280 = (1'h0); (forvar2280 < (1'h0)); forvar2280 = (forvar2280 + (1'h1)))
                begin
                  for (forvar2281 = (1'h0); (forvar2281 < (2'h3)); forvar2281 = (forvar2281 + (1'h1)))
                    begin
                      reg2282 <= forvar2243[(3'h5):(1'h1)];
                      reg2283 <= reg2211[(4'h8):(2'h3)];
                    end
                  reg2284 <= (reg1973[(3'h4):(3'h4)] && reg1934);
                  for (forvar2285 = (1'h0); (forvar2285 < (2'h2)); forvar2285 = (forvar2285 + (1'h1)))
                    begin
                      reg2286 <= {forvar1998};
                      reg2287 <= forvar2208[(4'h8):(3'h6)];
                      reg2288 <= (reg1994[(1'h0):(1'h0)] ?
                          $unsigned($signed(reg2186)) : (~&(reg1957 & $unsigned(reg2172))));
                      reg2289 <= forvar2022[(2'h3):(2'h2)];
                    end
                end
              if ((($signed((reg2186 * reg2258)) >>> $signed(forvar2172)) & $unsigned(forvar2106[(1'h0):(1'h0)])))
                begin
                  for (forvar2290 = (1'h0); (forvar2290 < (1'h1)); forvar2290 = (forvar2290 + (1'h1)))
                    begin
                      reg2291 <= {$signed($signed(((8'ha1) ^~ forvar2075)))};
                      reg2292 <= $unsigned($unsigned(((&reg2036) ?
                          (forvar2164 ? reg2166 : (8'hb4)) : forvar2290)));
                    end
                  if ($signed(((forvar2264 <<< (^reg2118)) ^ {reg2067[(1'h1):(1'h0)]})))
                    begin
                      reg2293 <= {($unsigned((^reg2283)) + reg2232)};
                      reg2294 <= reg1929[(4'hb):(3'h5)];
                    end
                  else
                    begin
                      reg2293 <= ($unsigned(reg2009[(4'h9):(3'h5)]) ?
                          (~{(reg2091 - reg1993)}) : reg1967);
                      reg2294 <= reg1987[(4'h9):(2'h3)];
                    end
                  for (forvar2295 = (1'h0); (forvar2295 < (1'h1)); forvar2295 = (forvar2295 + (1'h1)))
                    begin
                      reg2296 <= (reg2006[(3'h6):(2'h3)] ?
                          $signed($unsigned($unsigned(forvar2065))) : ($signed((8'ha8)) ?
                              reg2190 : forvar2279));
                      reg2297 <= $signed(((8'hb1) <<< (-reg2139[(4'he):(3'h7)])));
                      reg2298 <= reg2123[(2'h2):(2'h2)];
                    end
                  if ($signed(forvar2075[(4'hd):(3'h4)]))
                    begin
                      reg2299 <= (8'hb2);
                      reg2300 <= ((~(~^(forvar2264 ?
                              forvar2013 : forvar1933))) ?
                          $signed((~^reg2141)) : (&forvar2033));
                      reg2301 <= $signed({reg1989[(1'h1):(1'h0)]});
                    end
                  else
                    begin
                      reg2299 <= $signed({reg2253[(3'h7):(3'h4)]});
                    end
                end
              else
                begin
                  if (({({reg2016} ?
                          {reg2038} : $signed(reg2036))} << forvar2065))
                    begin
                      reg2290 <= (-((&$signed(forvar2015)) >>> (~forvar2172)));
                      reg2291 <= (8'hb6);
                    end
                  else
                    begin
                      reg2290 <= $signed($unsigned({$unsigned((8'ha6))}));
                      reg2291 <= ($unsigned({reg2151}) ?
                          $signed(reg2232[(1'h1):(1'h1)]) : $unsigned(forvar1948[(2'h2):(2'h2)]));
                      reg2292 <= ((((reg2089 ?
                              reg1968 : (8'hb8)) >= $unsigned(reg2059)) * reg2284[(2'h2):(1'h0)]) ?
                          reg1986[(3'h4):(2'h3)] : ((((8'ha1) ?
                                      reg2244 : reg2156) ?
                                  (^reg1965) : $unsigned(reg1958)) ?
                              (reg2267 >= reg2180) : forvar2082));
                      reg2293 <= (^(8'h9d));
                    end
                  reg2294 <= reg2209[(2'h2):(1'h0)];
                  if ($signed($signed(reg2044)))
                    begin
                      reg2295 <= $signed((^(^reg2036)));
                      reg2296 <= (^$unsigned(($unsigned(reg2139) <= $unsigned(reg2180))));
                    end
                  else
                    begin
                      reg2295 <= (8'h9e);
                      reg2296 <= (~^$unsigned(forvar2132[(4'hc):(2'h3)]));
                      reg2297 <= $unsigned(reg2282);
                    end
                  for (forvar2298 = (1'h0); (forvar2298 < (1'h1)); forvar2298 = (forvar2298 + (1'h1)))
                    begin
                      reg2299 <= (!((~&(reg2251 && (8'h9c))) < ($signed(reg2119) == reg1976)));
                      reg2300 <= ((+($signed(reg2025) >>> (reg2086 != forvar2143))) ?
                          ($unsigned({reg2128}) * $signed(reg2172[(2'h2):(1'h0)])) : (~|reg2221));
                      reg2301 <= (reg2110 | $signed((&reg2251[(2'h3):(2'h3)])));
                      reg2302 <= $unsigned(reg1941[(2'h3):(2'h3)]);
                    end
                end
            end
        end
      else
        begin
          if ($signed(forvar2168))
            begin
              for (forvar2275 = (1'h0); (forvar2275 < (1'h0)); forvar2275 = (forvar2275 + (1'h1)))
                begin
                  for (forvar2276 = (1'h0); (forvar2276 < (2'h2)); forvar2276 = (forvar2276 + (1'h1)))
                    begin
                      reg2277 <= $unsigned($signed($signed((forvar2247 | forvar2128))));
                    end
                  if ((^~reg2146))
                    begin
                      reg2278 <= $signed({$signed($signed(reg1941))});
                      reg2279 <= forvar1934;
                    end
                  else
                    begin
                      reg2278 <= $signed(reg2279);
                    end
                end
              reg2280 <= forvar2205[(2'h3):(2'h3)];
              for (forvar2281 = (1'h0); (forvar2281 < (2'h3)); forvar2281 = (forvar2281 + (1'h1)))
                begin
                  for (forvar2282 = (1'h0); (forvar2282 < (2'h3)); forvar2282 = (forvar2282 + (1'h1)))
                    begin
                      reg2283 <= reg2252[(3'h5):(3'h4)];
                      reg2284 <= (|((~^(reg2101 >>> reg2072)) ?
                          $signed({(8'hb1)}) : (reg1939 ?
                              (|(8'hac)) : $unsigned(reg1958))));
                      reg2285 <= $signed((forvar2047[(5'h10):(4'he)] ?
                          $unsigned({reg1951}) : {(~&reg1951)}));
                      reg2286 <= (+(+$signed((&reg1971))));
                    end
                  for (forvar2287 = (1'h0); (forvar2287 < (2'h2)); forvar2287 = (forvar2287 + (1'h1)))
                    begin
                      reg2288 <= reg2256;
                    end
                end
              for (forvar2289 = (1'h0); (forvar2289 < (1'h1)); forvar2289 = (forvar2289 + (1'h1)))
                begin
                  for (forvar2290 = (1'h0); (forvar2290 < (1'h1)); forvar2290 = (forvar2290 + (1'h1)))
                    begin
                      reg2291 <= (($signed((reg2299 | (8'hb6))) ^ ((reg2171 || reg2161) || $unsigned(reg2201))) == (^~(8'hab)));
                      reg2292 <= (8'haf);
                    end
                  for (forvar2293 = (1'h0); (forvar2293 < (2'h2)); forvar2293 = (forvar2293 + (1'h1)))
                    begin
                      reg2294 <= $unsigned(($unsigned((8'hb7)) > (~|reg2084)));
                      reg2295 <= (reg1969[(3'h5):(2'h3)] > $unsigned((~|forvar2290)));
                    end
                  for (forvar2296 = (1'h0); (forvar2296 < (1'h0)); forvar2296 = (forvar2296 + (1'h1)))
                    begin
                      reg2297 <= reg1981;
                      reg2298 <= $unsigned($signed((+$unsigned(forvar2250))));
                      reg2299 <= (~^$signed((8'had)));
                      reg2300 <= (~&reg2025[(3'h7):(3'h6)]);
                    end
                end
            end
          else
            begin
              for (forvar2275 = (1'h0); (forvar2275 < (2'h2)); forvar2275 = (forvar2275 + (1'h1)))
                begin
                  reg2276 <= {$signed((reg2125 <= reg2077))};
                  if ((~|$signed(((+reg1994) ?
                      (reg2113 ? reg1949 : reg2173) : $signed((8'haf))))))
                    begin
                      reg2277 <= (reg2041[(3'h4):(2'h3)] ?
                          {forvar2213} : $signed({$unsigned(forvar2028)}));
                    end
                  else
                    begin
                      reg2277 <= {(reg2067 ?
                              {(forvar2295 * reg2044)} : (reg2290[(4'ha):(3'h5)] && (+forvar2030)))};
                    end
                  reg2278 <= $unsigned($unsigned(reg2280));
                  reg2279 <= (!reg1975);
                end
              reg2280 <= {reg1950};
              for (forvar2281 = (1'h0); (forvar2281 < (1'h1)); forvar2281 = (forvar2281 + (1'h1)))
                begin
                  if ($signed((&(~|$signed(reg1938)))))
                    begin
                      reg2282 <= $signed($signed((!$unsigned(forvar2275))));
                    end
                  else
                    begin
                      reg2282 <= (((!(~&reg1985)) ?
                              (~&(reg1934 ? reg2042 : reg1931)) : {{reg2126}}) ?
                          (8'hba) : forvar2145[(3'h5):(1'h1)]);
                    end
                  for (forvar2283 = (1'h0); (forvar2283 < (2'h2)); forvar2283 = (forvar2283 + (1'h1)))
                    begin
                      reg2284 <= {(~^reg2244[(1'h0):(1'h0)])};
                    end
                end
              if ($unsigned((^forvar1933[(4'h8):(3'h7)])))
                begin
                  if ((~^$signed($signed(((8'ha1) ? reg2039 : reg1937)))))
                    begin
                      reg2285 <= ({$unsigned(reg2038)} ?
                          (~^(&(8'ha2))) : $signed((reg1950 ?
                              $signed(forvar2228) : (reg1976 ?
                                  (8'hba) : forvar2023))));
                      reg2286 <= $unsigned(reg2167[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2285 <= reg1941;
                      reg2286 <= ($signed({(8'ha3)}) ?
                          {((reg2137 ? reg2063 : reg2301) ?
                                  $unsigned(forvar2269) : (reg2225 - reg2171))} : ($signed(reg2105[(2'h3):(2'h3)]) ?
                              (reg2276[(3'h7):(3'h5)] > (forvar1963 * reg2081)) : reg2268));
                    end
                end
              else
                begin
                  if (reg2183[(3'h5):(2'h2)])
                    begin
                      reg2285 <= ({((^~(8'ha7)) ?
                                  $signed(reg2128) : {reg2181})} ?
                          {(-$signed(forvar2084))} : (forvar2132 ?
                              $unsigned({reg2069}) : $signed(((8'hb3) ?
                                  forvar1999 : reg2271))));
                      reg2286 <= {($unsigned($signed(reg2094)) != $signed({reg2254}))};
                    end
                  else
                    begin
                      reg2285 <= $signed((($signed((8'ha5)) ?
                              ((8'ha9) > reg1962) : (~^(8'hba))) ?
                          reg2284 : reg2141));
                      reg2286 <= forvar2015[(4'h8):(3'h6)];
                      reg2287 <= (|(^(^$unsigned((8'ha6)))));
                      reg2288 <= reg2020;
                    end
                  for (forvar2289 = (1'h0); (forvar2289 < (2'h2)); forvar2289 = (forvar2289 + (1'h1)))
                    begin
                      reg2290 <= (-$unsigned({(reg2173 | forvar1948)}));
                      reg2291 <= {($signed(reg2138) ?
                              reg2276[(1'h0):(1'h0)] : ($signed(reg2045) << forvar2004[(2'h2):(2'h2)]))};
                      reg2292 <= {$unsigned(wire1928[(3'h5):(2'h3)])};
                    end
                  if ($unsigned($unsigned(reg1937[(3'h5):(1'h1)])))
                    begin
                      reg2293 <= (8'ha2);
                    end
                  else
                    begin
                      reg2293 <= (^reg2002[(3'h7):(2'h2)]);
                      reg2294 <= $unsigned(({(reg2071 >> forvar2100)} ?
                          $unsigned((reg1975 ?
                              forvar2035 : reg2175)) : (-$unsigned(forvar2145))));
                      reg2295 <= reg2279[(3'h4):(3'h4)];
                      reg2296 <= $unsigned({$unsigned(reg2120)});
                    end
                  reg2297 <= ($signed(forvar2293) ? forvar2173 : (8'had));
                end
            end
          for (forvar2301 = (1'h0); (forvar2301 < (2'h2)); forvar2301 = (forvar2301 + (1'h1)))
            begin
              reg2302 <= (~(reg2117[(3'h4):(1'h0)] > forvar2084));
              for (forvar2303 = (1'h0); (forvar2303 < (2'h2)); forvar2303 = (forvar2303 + (1'h1)))
                begin
                  if ($unsigned($unsigned($signed($unsigned(reg2054)))))
                    begin
                      reg2304 <= forvar2023;
                      reg2305 <= forvar2133;
                    end
                  else
                    begin
                      reg2304 <= reg2191[(2'h3):(1'h0)];
                      reg2305 <= $signed(reg2305);
                      reg2306 <= ((!$unsigned($signed(reg1970))) ?
                          $unsigned(($unsigned(reg2268) < {reg2121})) : ((|reg2180) ?
                              reg1986[(3'h6):(1'h0)] : ((~reg2147) ?
                                  $unsigned(reg2108) : (reg1957 - reg2021))));
                    end
                  if (reg2191[(3'h4):(2'h3)])
                    begin
                      reg2307 <= (reg1977[(3'h5):(1'h0)] && ((8'hb5) * {reg2084}));
                      reg2308 <= $signed($unsigned($signed({reg2104})));
                      reg2309 <= reg2146[(4'hf):(2'h2)];
                    end
                  else
                    begin
                      reg2307 <= reg2056[(1'h0):(1'h0)];
                      reg2308 <= ($signed((&(forvar2264 ^~ (8'ha8)))) ?
                          (reg2273[(3'h6):(2'h2)] & reg2035) : (~|forvar1931));
                      reg2309 <= (&($unsigned((reg2174 > forvar2028)) ^~ forvar2001));
                      reg2310 <= (~forvar2065);
                    end
                end
              for (forvar2311 = (1'h0); (forvar2311 < (1'h0)); forvar2311 = (forvar2311 + (1'h1)))
                begin
                  reg2312 <= ((({forvar1970} + $unsigned(reg2267)) ?
                      reg2306[(2'h2):(1'h1)] : ({reg2197} ?
                          (reg2183 | reg2155) : reg1996)) * (^~$signed($signed((8'hb8)))));
                  for (forvar2313 = (1'h0); (forvar2313 < (2'h2)); forvar2313 = (forvar2313 + (1'h1)))
                    begin
                      reg2314 <= ($signed({{wire1928}}) ?
                          forvar2004[(3'h4):(3'h4)] : $signed((-(~^reg2084))));
                      reg2315 <= $signed({forvar1980[(2'h3):(1'h0)]});
                    end
                  for (forvar2316 = (1'h0); (forvar2316 < (2'h3)); forvar2316 = (forvar2316 + (1'h1)))
                    begin
                      reg2317 <= reg1935;
                    end
                  if ($unsigned($signed((!$unsigned(reg2162)))))
                    begin
                      reg2318 <= reg2061;
                      reg2319 <= {{({reg2226} >= reg2227[(3'h6):(3'h6)])}};
                      reg2320 <= $unsigned((-($unsigned((8'ha0)) ?
                          $unsigned(reg2235) : $unsigned(reg2092))));
                    end
                  else
                    begin
                      reg2318 <= ((((reg2251 ?
                                  forvar1983 : (8'hb9)) ^ reg2220) ?
                              ((~|(8'hab)) ?
                                  $unsigned(forvar2287) : $unsigned(forvar2293)) : reg2008) ?
                          ((~&reg2190) ?
                              reg2025[(3'h5):(3'h5)] : (reg2015 ^ reg2184)) : (((8'hb9) ?
                              ((8'ha7) ?
                                  forvar2095 : forvar2162) : {forvar2128}) >= forvar2179[(2'h2):(2'h2)]));
                      reg2319 <= ({reg2283} ?
                          (^~$unsigned($signed((8'ha2)))) : ((^(&reg2270)) << forvar1943[(1'h1):(1'h1)]));
                      reg2320 <= $signed((^$unsigned((forvar2030 >> reg2156))));
                    end
                end
            end
          for (forvar2321 = (1'h0); (forvar2321 < (1'h0)); forvar2321 = (forvar2321 + (1'h1)))
            begin
              for (forvar2322 = (1'h0); (forvar2322 < (1'h1)); forvar2322 = (forvar2322 + (1'h1)))
                begin
                  for (forvar2323 = (1'h0); (forvar2323 < (1'h0)); forvar2323 = (forvar2323 + (1'h1)))
                    begin
                      reg2324 <= reg2016;
                    end
                  for (forvar2325 = (1'h0); (forvar2325 < (2'h3)); forvar2325 = (forvar2325 + (1'h1)))
                    begin
                      reg2326 <= ((reg2175 ^~ reg2201) == {reg2189});
                      reg2327 <= forvar1956[(3'h5):(1'h0)];
                      reg2328 <= $unsigned((($signed(reg2203) ?
                              (reg1975 ? forvar2321 : (8'hb1)) : reg2251) ?
                          reg2059 : (reg2277[(1'h1):(1'h1)] ~^ reg2269)));
                      reg2329 <= $unsigned($signed(($signed(reg2163) | (-reg2125))));
                    end
                  for (forvar2330 = (1'h0); (forvar2330 < (1'h1)); forvar2330 = (forvar2330 + (1'h1)))
                    begin
                      reg2331 <= reg2047;
                      reg2332 <= reg2183[(1'h0):(1'h0)];
                      reg2333 <= forvar2220[(3'h5):(2'h3)];
                    end
                  reg2334 <= $signed((!reg2029[(4'h9):(2'h2)]));
                end
              if ((8'hb9))
                begin
                  if ((~forvar2187))
                    begin
                      reg2335 <= $unsigned((reg2037[(1'h1):(1'h0)] ~^ {$signed(reg2285)}));
                      reg2336 <= forvar2091;
                      reg2337 <= reg2012[(2'h3):(1'h0)];
                      reg2338 <= ((($unsigned(reg2186) && $unsigned(reg2172)) & $unsigned(reg1997[(4'hb):(3'h5)])) >= {(~&(reg2283 >= reg2107))});
                    end
                  else
                    begin
                      reg2335 <= (-(reg2215 ?
                          ((wire1924 ?
                              forvar1931 : reg2207) >> (~&reg2108)) : $unsigned(reg2318)));
                      reg2336 <= forvar2095;
                      reg2337 <= (~|{(^((8'h9d) ? reg1963 : reg2010))});
                    end
                  for (forvar2339 = (1'h0); (forvar2339 < (1'h0)); forvar2339 = (forvar2339 + (1'h1)))
                    begin
                      reg2340 <= $signed((reg2003 >= reg2234[(2'h2):(1'h0)]));
                      reg2341 <= ($unsigned($unsigned((reg2068 ?
                              (8'h9e) : (8'ha1)))) ?
                          reg2123 : reg2214[(3'h5):(1'h0)]);
                      reg2342 <= forvar2106;
                    end
                end
              else
                begin
                  for (forvar2335 = (1'h0); (forvar2335 < (1'h1)); forvar2335 = (forvar2335 + (1'h1)))
                    begin
                      reg2336 <= {{(~^forvar2058)}};
                      reg2337 <= (forvar2275 < reg2058[(4'ha):(2'h3)]);
                      reg2338 <= (((~$signed(reg2314)) != $signed((forvar2051 ?
                              reg1950 : (8'hac)))) ?
                          (~&(reg2016[(3'h4):(2'h3)] * $signed(forvar2091))) : ($signed((reg2182 <<< forvar2091)) >>> (~|reg1929[(2'h3):(1'h1)])));
                      reg2339 <= (~&(~|$unsigned((forvar2323 ?
                          forvar2075 : reg2149))));
                    end
                  reg2340 <= ((reg2314 > reg2037[(3'h5):(3'h4)]) < $unsigned((-reg2140[(1'h1):(1'h0)])));
                  if (forvar2126[(2'h2):(2'h2)])
                    begin
                      reg2341 <= (reg2109[(4'h9):(1'h1)] ?
                          (|((reg2054 ? forvar1956 : reg2289) ?
                              $unsigned(forvar2167) : (+reg2097))) : reg2148);
                      reg2342 <= (($signed($unsigned(forvar1956)) ?
                          $signed({forvar2208}) : $unsigned((~^reg2080))) > (~^((reg1948 ^~ reg2052) != forvar2264[(2'h3):(2'h2)])));
                      reg2343 <= reg2020[(2'h2):(1'h0)];
                      reg2344 <= $signed($unsigned(forvar2145));
                    end
                  else
                    begin
                      reg2341 <= reg2184[(3'h7):(1'h0)];
                      reg2342 <= $unsigned(forvar2078);
                      reg2343 <= {$signed($signed((forvar1970 > reg1991)))};
                      reg2344 <= forvar2050[(4'he):(2'h3)];
                    end
                  reg2345 <= reg2187[(1'h1):(1'h0)];
                end
            end
          if ({($unsigned((reg2181 ? reg2222 : reg2257)) - $signed({reg2117}))})
            begin
              for (forvar2346 = (1'h0); (forvar2346 < (1'h0)); forvar2346 = (forvar2346 + (1'h1)))
                begin
                  reg2347 <= ($unsigned((reg2332 ?
                      $signed(reg2074) : forvar2124)) >> (($unsigned((8'hac)) ?
                          (forvar1956 | reg2235) : (reg2262 ?
                              reg1968 : forvar2033)) ?
                      ((reg1947 ?
                          (8'haf) : (8'ha1)) || $signed((8'ha0))) : forvar1967));
                end
              if ({forvar1947})
                begin
                  reg2348 <= forvar2283[(1'h1):(1'h1)];
                end
              else
                begin
                  reg2348 <= reg2251[(2'h3):(1'h0)];
                  if ($signed(reg2257[(3'h4):(1'h1)]))
                    begin
                      reg2349 <= (!reg1938);
                      reg2350 <= forvar2095;
                      reg2351 <= $signed($unsigned($unsigned($unsigned(forvar2011))));
                    end
                  else
                    begin
                      reg2349 <= $signed((!$unsigned(forvar2164[(3'h6):(3'h5)])));
                      reg2350 <= (&$unsigned((~forvar2086[(4'hb):(4'ha)])));
                      reg2351 <= ($signed($unsigned({(8'hb4)})) - reg2081[(2'h2):(1'h0)]);
                      reg2352 <= {(^$unsigned((~^reg2217)))};
                    end
                  reg2353 <= (~&($unsigned($unsigned(reg1954)) && ((&reg2334) ?
                      $unsigned(forvar2096) : ((8'hb3) ?
                          forvar2053 : reg2155))));
                end
              if (reg2224[(1'h1):(1'h0)])
                begin
                  for (forvar2354 = (1'h0); (forvar2354 < (2'h3)); forvar2354 = (forvar2354 + (1'h1)))
                    begin
                      reg2355 <= reg2147;
                      reg2356 <= reg2256;
                    end
                  if ((&((forvar2323 ?
                          reg2024[(4'ha):(4'h9)] : reg2298[(4'h9):(3'h5)]) ?
                      ($signed(reg2227) ?
                          {reg2270} : (forvar2179 ?
                              reg2335 : reg2307)) : (+$signed(reg2317)))))
                    begin
                      reg2357 <= ((-(~|forvar2011[(2'h3):(2'h2)])) == reg2215);
                      reg2358 <= ($signed((&$signed(reg2230))) ?
                          ({$unsigned(reg2279)} > {$unsigned((8'h9e))}) : (-reg1986));
                      reg2359 <= (^~(+((reg2197 ?
                          forvar2143 : forvar2172) <= $signed(reg2320))));
                      reg2360 <= $unsigned($unsigned($signed(((8'hb6) | forvar2143))));
                    end
                  else
                    begin
                      reg2357 <= ((($signed(reg2296) ?
                              $unsigned(forvar2083) : $unsigned((8'hb8))) ?
                          $signed($signed(reg2018)) : ($signed(reg2174) ?
                              (reg1951 ?
                                  reg2242 : reg2057) : reg2120[(2'h3):(1'h0)])) ^ $signed({$signed((8'hb7))}));
                      reg2358 <= ((forvar2279[(2'h3):(1'h1)] != forvar1999) ?
                          $signed({$signed(forvar2023)}) : reg2051);
                    end
                end
              else
                begin
                  if (forvar1933)
                    begin
                      reg2354 <= $unsigned(reg2021);
                    end
                  else
                    begin
                      reg2354 <= wire1927;
                    end
                  for (forvar2355 = (1'h0); (forvar2355 < (1'h0)); forvar2355 = (forvar2355 + (1'h1)))
                    begin
                      reg2356 <= (+{($signed(forvar2083) < $unsigned(reg2091))});
                    end
                  for (forvar2357 = (1'h0); (forvar2357 < (2'h2)); forvar2357 = (forvar2357 + (1'h1)))
                    begin
                      reg2358 <= (8'ha3);
                    end
                  for (forvar2359 = (1'h0); (forvar2359 < (2'h2)); forvar2359 = (forvar2359 + (1'h1)))
                    begin
                      reg2360 <= $unsigned((reg2173 ~^ reg2131[(1'h0):(1'h0)]));
                    end
                end
            end
          else
            begin
              reg2346 <= $signed($unsigned(((^~wire1925) ?
                  reg2135[(2'h3):(1'h0)] : (reg2266 <<< reg2357))));
              reg2347 <= $signed((~((+(8'hb6)) >= reg1957[(3'h5):(2'h3)])));
              for (forvar2348 = (1'h0); (forvar2348 < (1'h1)); forvar2348 = (forvar2348 + (1'h1)))
                begin
                  for (forvar2349 = (1'h0); (forvar2349 < (2'h2)); forvar2349 = (forvar2349 + (1'h1)))
                    begin
                      reg2350 <= $signed(reg2059);
                    end
                end
              for (forvar2351 = (1'h0); (forvar2351 < (1'h1)); forvar2351 = (forvar2351 + (1'h1)))
                begin
                  for (forvar2352 = (1'h0); (forvar2352 < (2'h2)); forvar2352 = (forvar2352 + (1'h1)))
                    begin
                      reg2353 <= $signed(reg2253);
                    end
                  reg2354 <= $unsigned(reg2338[(4'hc):(3'h6)]);
                  reg2355 <= ((~&reg2138[(3'h4):(3'h4)]) ?
                      ($signed({forvar2269}) == ($unsigned(forvar2163) && ((8'hac) > (8'ha8)))) : $signed(($unsigned(reg2239) ?
                          {(8'had)} : forvar2210[(2'h2):(1'h1)])));
                  if ($signed(reg2230))
                    begin
                      reg2356 <= ((^~reg2130[(1'h1):(1'h0)]) == forvar2168[(3'h6):(1'h1)]);
                    end
                  else
                    begin
                      reg2356 <= ((((reg2173 <<< reg2203) ?
                                  forvar2212[(4'hb):(4'h8)] : (~&(8'hb5))) ?
                              {(forvar2058 ? reg1955 : forvar2316)} : reg1987) ?
                          $unsigned((|{reg2085})) : $signed({reg2191[(3'h5):(2'h2)]}));
                      reg2357 <= (8'hae);
                    end
                end
            end
        end
      for (forvar2361 = (1'h0); (forvar2361 < (2'h3)); forvar2361 = (forvar2361 + (1'h1)))
        begin
          for (forvar2362 = (1'h0); (forvar2362 < (1'h0)); forvar2362 = (forvar2362 + (1'h1)))
            begin
              for (forvar2363 = (1'h0); (forvar2363 < (1'h1)); forvar2363 = (forvar2363 + (1'h1)))
                begin
                  for (forvar2364 = (1'h0); (forvar2364 < (2'h3)); forvar2364 = (forvar2364 + (1'h1)))
                    begin
                      reg2365 <= $signed({$unsigned((~&reg2089))});
                      reg2366 <= $unsigned(reg2282[(2'h3):(2'h3)]);
                      reg2367 <= (reg1957[(3'h4):(3'h4)] ?
                          reg1993[(1'h1):(1'h1)] : $unsigned($unsigned((forvar2041 ?
                              forvar2023 : reg2090))));
                    end
                  for (forvar2368 = (1'h0); (forvar2368 < (2'h3)); forvar2368 = (forvar2368 + (1'h1)))
                    begin
                      reg2369 <= $signed((!(-{(8'h9c)})));
                    end
                end
            end
          if (($unsigned($unsigned((forvar2349 ? forvar2346 : reg2302))) ?
              $signed(reg2260[(2'h2):(1'h1)]) : $unsigned($signed($signed(forvar2339)))))
            begin
              if ($signed({(+$unsigned(reg2044))}))
                begin
                  if ($signed(forvar2022[(3'h6):(2'h2)]))
                    begin
                      reg2370 <= {$unsigned({(reg2181 ? reg2300 : reg2304)})};
                      reg2371 <= $unsigned(((^(~|reg1986)) && (((8'hb7) ~^ (8'hac)) > ((8'ha8) ?
                          (8'hb7) : reg1931))));
                      reg2372 <= $unsigned(($signed(reg2134[(4'hb):(3'h7)]) ?
                          $signed((^~reg2193)) : ($signed(reg2119) ?
                              {reg2052} : $signed(reg2341))));
                    end
                  else
                    begin
                      reg2370 <= (^~$unsigned($signed((8'hb8))));
                    end
                  for (forvar2373 = (1'h0); (forvar2373 < (1'h0)); forvar2373 = (forvar2373 + (1'h1)))
                    begin
                      reg2374 <= (+reg2183);
                      reg2375 <= ({{reg2081[(3'h7):(2'h2)]}} <= $signed(forvar2362[(3'h5):(1'h1)]));
                      reg2376 <= {$unsigned(reg1980)};
                    end
                  if (forvar2095[(2'h3):(2'h2)])
                    begin
                      reg2377 <= (8'ha3);
                    end
                  else
                    begin
                      reg2377 <= reg1945[(4'hb):(3'h7)];
                      reg2378 <= ((({(8'hb4)} ?
                          (reg2182 ? (8'hb7) : (8'hb2)) : (reg2357 ?
                              (8'ha8) : reg2258)) || ($unsigned((8'hb2)) ?
                          (8'hb2) : {reg2051})) == (forvar1963[(3'h5):(2'h2)] * (reg2271 >> $unsigned(forvar2301))));
                    end
                end
              else
                begin
                  for (forvar2370 = (1'h0); (forvar2370 < (2'h2)); forvar2370 = (forvar2370 + (1'h1)))
                    begin
                      reg2371 <= (~(+reg2089));
                    end
                  reg2372 <= $unsigned((~|$signed($signed(reg2224))));
                end
              for (forvar2379 = (1'h0); (forvar2379 < (1'h1)); forvar2379 = (forvar2379 + (1'h1)))
                begin
                  reg2380 <= {reg2108};
                  reg2381 <= $unsigned($unsigned((reg2349[(3'h4):(1'h1)] ?
                      (forvar2164 || reg1935) : (forvar1959 + reg2012))));
                end
            end
          else
            begin
              for (forvar2370 = (1'h0); (forvar2370 < (1'h1)); forvar2370 = (forvar2370 + (1'h1)))
                begin
                  for (forvar2371 = (1'h0); (forvar2371 < (1'h1)); forvar2371 = (forvar2371 + (1'h1)))
                    begin
                      reg2372 <= ((((&forvar2287) ?
                          (reg2063 ^ forvar2283) : reg2102[(1'h0):(1'h0)]) - {$signed(reg2134)}) | reg2319[(2'h2):(1'h1)]);
                      reg2373 <= $unsigned((8'h9c));
                      reg2374 <= $signed((forvar2335 >= $signed(reg2051)));
                    end
                  reg2375 <= (~^reg2067);
                  if ((($signed((&reg2312)) * (8'h9e)) ?
                      ($signed({reg2113}) > ((8'ha7) ?
                          $signed(reg2256) : (^~(8'hb3)))) : (forvar2177[(3'h7):(3'h5)] - reg2312)))
                    begin
                      reg2376 <= (reg2279 ?
                          (((reg2118 ? reg2257 : forvar2167) ?
                                  $signed(reg2338) : reg1978) ?
                              reg2193[(3'h7):(3'h6)] : (wire1928 != (forvar2321 ?
                                  (8'hb8) : reg2340))) : reg1981[(2'h3):(1'h0)]);
                      reg2377 <= $signed((^~(|$signed(reg2274))));
                      reg2378 <= $unsigned(({(reg2081 >= forvar2095)} ?
                          (~|(~(8'hb7))) : $unsigned(forvar1938)));
                    end
                  else
                    begin
                      reg2376 <= (forvar2279[(2'h3):(2'h3)] ?
                          $unsigned(({forvar1976} ?
                              forvar2028 : reg2012)) : (-$unsigned($unsigned((8'had)))));
                    end
                end
            end
        end
      if ((-$signed(((-forvar2363) ?
          ((8'hb9) ? reg2161 : reg2226) : (reg1929 ? forvar2339 : reg2290)))))
        begin
          for (forvar2382 = (1'h0); (forvar2382 < (1'h1)); forvar2382 = (forvar2382 + (1'h1)))
            begin
              for (forvar2383 = (1'h0); (forvar2383 < (1'h0)); forvar2383 = (forvar2383 + (1'h1)))
                begin
                  reg2384 <= reg1932;
                end
              reg2385 <= {reg1954};
              for (forvar2386 = (1'h0); (forvar2386 < (1'h0)); forvar2386 = (forvar2386 + (1'h1)))
                begin
                  for (forvar2387 = (1'h0); (forvar2387 < (2'h2)); forvar2387 = (forvar2387 + (1'h1)))
                    begin
                      reg2388 <= reg2261[(1'h1):(1'h0)];
                      reg2389 <= forvar2187[(4'h8):(3'h4)];
                      reg2390 <= reg2014[(3'h5):(3'h4)];
                      reg2391 <= forvar2285;
                    end
                  for (forvar2392 = (1'h0); (forvar2392 < (1'h1)); forvar2392 = (forvar2392 + (1'h1)))
                    begin
                      reg2393 <= (!$unsigned($unsigned((reg2147 ?
                          reg1952 : forvar2368))));
                    end
                end
              for (forvar2394 = (1'h0); (forvar2394 < (1'h0)); forvar2394 = (forvar2394 + (1'h1)))
                begin
                  for (forvar2395 = (1'h0); (forvar2395 < (2'h2)); forvar2395 = (forvar2395 + (1'h1)))
                    begin
                      reg2396 <= $signed(reg2198);
                    end
                  reg2397 <= forvar1971[(3'h5):(2'h2)];
                  reg2398 <= {reg2258[(1'h0):(1'h0)]};
                  for (forvar2399 = (1'h0); (forvar2399 < (2'h3)); forvar2399 = (forvar2399 + (1'h1)))
                    begin
                      reg2400 <= (8'ha3);
                      reg2401 <= forvar2132[(4'ha):(3'h4)];
                      reg2402 <= $unsigned(reg2050[(1'h1):(1'h1)]);
                    end
                end
            end
          reg2403 <= $unsigned((({reg2000} ?
              $signed(forvar2091) : (forvar2395 >= (8'haf))) ^ $unsigned($signed(reg2152))));
          if (((({reg2275} ? $signed(forvar2084) : $unsigned((8'ha6))) ?
              ($unsigned(reg2291) ^~ $signed(reg2079)) : {reg2014}) << $unsigned((reg1980 ^ (reg2315 >>> reg2339)))))
            begin
              if ((reg2179 <= {(~$unsigned(forvar2357))}))
                begin
                  reg2404 <= reg2225;
                  if (((|reg2242[(2'h2):(1'h1)]) ?
                      ((reg2164 < reg2236[(1'h0):(1'h0)]) << $signed((|(8'haa)))) : {reg1946}))
                    begin
                      reg2405 <= {$signed(forvar1948)};
                      reg2406 <= ({reg2045[(1'h0):(1'h0)]} ?
                          ($unsigned($signed((8'h9e))) | {(reg2233 + forvar1970)}) : $signed(reg2112));
                      reg2407 <= ((~&$signed($unsigned(reg2396))) ?
                          (-($signed(reg1932) ^ reg2206[(1'h0):(1'h0)])) : (~|((reg2016 >> (8'ha7)) ?
                              $unsigned(reg2355) : (+forvar2128))));
                      reg2408 <= (((~^reg2109) > forvar2373[(4'h9):(3'h6)]) ?
                          (((reg2171 << forvar2349) + (reg2165 | forvar2383)) >>> ($unsigned(forvar2269) ?
                              (reg2274 * reg2123) : $unsigned(forvar2371))) : ((-(reg2158 ?
                              forvar2049 : (8'hac))) >>> reg2179));
                    end
                  else
                    begin
                      reg2405 <= forvar2035[(3'h5):(3'h5)];
                      reg2406 <= $signed($signed(((reg2038 ?
                              reg1938 : reg2032) ?
                          forvar2001[(4'hb):(4'hb)] : $signed(forvar2052))));
                    end
                  reg2409 <= (8'h9c);
                  if ({(((&reg2275) ? reg1929 : (~^reg2089)) & wire1926)})
                    begin
                      reg2410 <= ($signed((^~$unsigned(reg1951))) ?
                          (~|reg2373) : (!$unsigned(reg2089[(2'h2):(2'h2)])));
                      reg2411 <= ($unsigned($unsigned(forvar2157[(4'hb):(2'h3)])) > forvar2280);
                      reg2412 <= ({reg2320[(1'h1):(1'h1)]} ?
                          (^forvar2325[(4'hb):(4'hb)]) : (~&(~&{(8'ha9)})));
                    end
                  else
                    begin
                      reg2410 <= reg2178[(4'hb):(4'hb)];
                      reg2411 <= $unsigned((reg2168[(2'h3):(2'h3)] ?
                          (~&$signed(forvar1936)) : (+(reg1929 ?
                              (8'ha0) : reg1951))));
                      reg2412 <= reg2164[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar2404 = (1'h0); (forvar2404 < (1'h0)); forvar2404 = (forvar2404 + (1'h1)))
                    begin
                      reg2405 <= ((~^((reg2140 ?
                          reg2347 : reg2335) ~^ $signed(forvar2280))) >>> reg2179);
                      reg2406 <= (~^$signed((reg2118[(1'h1):(1'h1)] ?
                          (reg2272 ?
                              forvar2382 : forvar2096) : (reg2215 ^ reg2051))));
                      reg2407 <= {reg1929[(5'h10):(4'hc)]};
                      reg2408 <= $unsigned(reg2138[(1'h0):(1'h0)]);
                    end
                  for (forvar2409 = (1'h0); (forvar2409 < (2'h2)); forvar2409 = (forvar2409 + (1'h1)))
                    begin
                      reg2410 <= (8'ha2);
                      reg2411 <= reg2175[(1'h0):(1'h0)];
                      reg2412 <= (8'haf);
                    end
                  for (forvar2413 = (1'h0); (forvar2413 < (1'h0)); forvar2413 = (forvar2413 + (1'h1)))
                    begin
                      reg2414 <= (reg2276[(1'h1):(1'h0)] >> reg2081[(4'hd):(3'h4)]);
                      reg2415 <= $unsigned((~^(&reg2149)));
                    end
                end
              if ({$unsigned({reg2061[(4'hb):(2'h3)]})})
                begin
                  for (forvar2416 = (1'h0); (forvar2416 < (2'h3)); forvar2416 = (forvar2416 + (1'h1)))
                    begin
                      reg2417 <= (forvar2362 ?
                          (+reg2188) : $unsigned($unsigned($unsigned(reg2142))));
                    end
                  for (forvar2418 = (1'h0); (forvar2418 < (2'h2)); forvar2418 = (forvar2418 + (1'h1)))
                    begin
                      reg2419 <= (~^$signed({forvar2201[(4'ha):(3'h6)]}));
                      reg2420 <= ($signed(forvar2136[(2'h3):(2'h3)]) ?
                          $signed(reg2211[(2'h3):(2'h2)]) : $signed((((8'h9e) ?
                              (8'hba) : reg1953) ^ $signed(reg1970))));
                      reg2421 <= forvar1962;
                    end
                  for (forvar2422 = (1'h0); (forvar2422 < (2'h2)); forvar2422 = (forvar2422 + (1'h1)))
                    begin
                      reg2423 <= {forvar2363[(1'h1):(1'h0)]};
                      reg2424 <= $unsigned(reg2254);
                    end
                end
              else
                begin
                  if ((($unsigned($unsigned((8'ha6))) ?
                          $signed((~^reg2183)) : forvar2187) ?
                      reg2293[(4'hc):(4'ha)] : {($signed((8'ha5)) ?
                              ((8'haf) == reg2180) : (8'hb8))}))
                    begin
                      reg2416 <= (^($unsigned(forvar2349) << ($signed(reg2189) ?
                          (reg2086 || reg2258) : reg2107)));
                    end
                  else
                    begin
                      reg2416 <= ($signed(reg2027) ?
                          {$signed(reg2416)} : {$signed(reg2396[(4'h9):(4'h8)])});
                      reg2417 <= reg2155;
                      reg2418 <= reg2126[(1'h1):(1'h0)];
                      reg2419 <= ((($signed(reg1947) & (~reg2270)) >> reg2417[(4'hc):(4'ha)]) & ((+reg2166[(4'hb):(4'h8)]) ?
                          forvar2082 : (reg2003 && (8'hb6))));
                    end
                  for (forvar2420 = (1'h0); (forvar2420 < (1'h0)); forvar2420 = (forvar2420 + (1'h1)))
                    begin
                      reg2421 <= reg1929;
                      reg2422 <= reg2328[(3'h4):(1'h0)];
                      reg2423 <= reg2008;
                    end
                  if ((&(&reg2293)))
                    begin
                      reg2424 <= {reg1961[(3'h4):(2'h2)]};
                      reg2425 <= {reg1932[(3'h4):(1'h1)]};
                      reg2426 <= reg1969[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg2424 <= reg2223;
                      reg2425 <= ($unsigned($unsigned(((8'h9f) ?
                              reg2353 : forvar2321))) ?
                          forvar2395 : reg2152);
                      reg2426 <= reg2181[(3'h6):(2'h2)];
                    end
                  if ($unsigned($signed((8'hab))))
                    begin
                      reg2427 <= ($signed({$signed(wire1925)}) <= $unsigned(reg2221[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg2427 <= (!((forvar2220[(2'h3):(1'h1)] ?
                              (+reg1993) : (-forvar1998)) ?
                          (&forvar2196) : forvar2020[(3'h5):(1'h1)]));
                    end
                end
              if (($unsigned(forvar2047[(4'hf):(3'h4)]) != $unsigned(reg2202[(4'ha):(3'h6)])))
                begin
                  if ((~&$unsigned({$unsigned(reg2314)})))
                    begin
                      reg2428 <= (reg2001 >> reg2348);
                      reg2429 <= (reg2375[(1'h0):(1'h0)] ^~ reg2426[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg2428 <= $unsigned((((reg2184 ? forvar2177 : (8'hb2)) ?
                              $unsigned(reg2424) : (!forvar2287)) ?
                          (-(forvar2285 - (8'ha9))) : $unsigned({forvar1941})));
                      reg2429 <= $signed($unsigned(reg2371[(2'h3):(1'h1)]));
                    end
                  for (forvar2430 = (1'h0); (forvar2430 < (1'h1)); forvar2430 = (forvar2430 + (1'h1)))
                    begin
                      reg2431 <= $signed($unsigned(reg2376[(2'h2):(1'h1)]));
                      reg2432 <= $unsigned(((reg2201 ?
                              $unsigned((8'had)) : $signed((8'h9e))) ?
                          forvar2133 : (^~(^~reg1987))));
                      reg2433 <= reg2409;
                      reg2434 <= reg2200;
                    end
                  reg2435 <= (forvar2373[(3'h4):(2'h3)] <= (8'hb1));
                  for (forvar2436 = (1'h0); (forvar2436 < (1'h0)); forvar2436 = (forvar2436 + (1'h1)))
                    begin
                      reg2437 <= reg2046;
                    end
                end
              else
                begin
                  for (forvar2428 = (1'h0); (forvar2428 < (1'h1)); forvar2428 = (forvar2428 + (1'h1)))
                    begin
                      reg2429 <= reg2046;
                    end
                end
            end
          else
            begin
              for (forvar2404 = (1'h0); (forvar2404 < (2'h2)); forvar2404 = (forvar2404 + (1'h1)))
                begin
                  if ($unsigned(forvar1959))
                    begin
                      reg2405 <= $signed((((reg2221 < (8'haf)) > $unsigned((8'ha7))) || reg2355[(2'h2):(1'h1)]));
                      reg2406 <= reg2053[(4'ha):(3'h6)];
                    end
                  else
                    begin
                      reg2405 <= (+reg2103);
                      reg2406 <= (((8'hae) ?
                              $signed((reg2345 ?
                                  reg2216 : reg2188)) : (reg2225[(3'h5):(1'h1)] ?
                                  reg2283 : $unsigned(reg2431))) ?
                          {$signed($unsigned(reg2279))} : ((~^(reg2069 ?
                              reg2000 : reg2226)) ^ $unsigned((reg2134 >= forvar2082))));
                      reg2407 <= {(&((8'haa) * {reg2140}))};
                      reg2408 <= (~(forvar2177 ?
                          reg2029[(2'h2):(1'h1)] : (^$signed(reg2042))));
                    end
                end
              for (forvar2409 = (1'h0); (forvar2409 < (2'h3)); forvar2409 = (forvar2409 + (1'h1)))
                begin
                  if (((((forvar2128 ? reg2037 : reg2240) && (^forvar2281)) ?
                          {wire1924[(1'h0):(1'h0)]} : $unsigned($signed(forvar2196))) ?
                      $signed({(^~reg1964)}) : $unsigned(reg2410[(1'h0):(1'h0)])))
                    begin
                      reg2410 <= $unsigned($signed(reg2266[(3'h4):(3'h4)]));
                      reg2411 <= $signed((8'ha9));
                      reg2412 <= ($unsigned((^~reg1967[(1'h1):(1'h0)])) <= $signed({(reg2393 && forvar2095)}));
                    end
                  else
                    begin
                      reg2410 <= $unsigned({{$signed(forvar2162)}});
                      reg2411 <= ($unsigned(reg2165[(1'h1):(1'h0)]) < ((~^(-reg1977)) >= $signed($unsigned(reg2203))));
                      reg2412 <= reg2335[(4'hc):(3'h6)];
                    end
                end
              for (forvar2413 = (1'h0); (forvar2413 < (1'h0)); forvar2413 = (forvar2413 + (1'h1)))
                begin
                  for (forvar2414 = (1'h0); (forvar2414 < (1'h1)); forvar2414 = (forvar2414 + (1'h1)))
                    begin
                      reg2415 <= forvar2290;
                      reg2416 <= ({$signed(reg2055[(3'h5):(3'h4)])} ^~ reg2254);
                      reg2417 <= (reg1946[(3'h6):(3'h6)] ?
                          (((reg2276 ? reg2053 : (8'ha7)) ^~ reg2389) ?
                              reg2337[(1'h1):(1'h0)] : $signed(reg2401)) : (~$unsigned((forvar1963 || reg2289))));
                      reg2418 <= $unsigned({((forvar2053 ^ reg2114) < $unsigned(reg2044))});
                    end
                end
            end
          reg2438 <= ((({reg2314} <= (|reg2219)) ^ {(reg1993 << forvar2196)}) ?
              $signed((forvar2083[(3'h7):(3'h5)] ?
                  forvar2023 : (forvar2041 > reg2088))) : (forvar2359 <<< {$unsigned(reg2079)}));
        end
      else
        begin
          for (forvar2382 = (1'h0); (forvar2382 < (1'h1)); forvar2382 = (forvar2382 + (1'h1)))
            begin
              if (reg2283[(3'h5):(1'h1)])
                begin
                  if (($signed($unsigned(((8'ha3) <= reg2426))) <= (((reg1947 << reg2227) ?
                          reg2245 : $unsigned(reg2205)) ?
                      forvar2285[(1'h1):(1'h1)] : (^(wire1925 ^ reg2433)))))
                    begin
                      reg2383 <= $unsigned((((reg2054 ?
                              reg2286 : reg2244) ~^ (|reg2334)) ?
                          forvar2174[(3'h7):(3'h4)] : reg2207));
                    end
                  else
                    begin
                      reg2383 <= (|{$signed((~|reg2035))});
                    end
                end
              else
                begin
                  for (forvar2383 = (1'h0); (forvar2383 < (1'h1)); forvar2383 = (forvar2383 + (1'h1)))
                    begin
                      reg2384 <= (reg2326[(3'h7):(1'h1)] <<< $unsigned(((!reg2268) + reg2094[(2'h2):(1'h1)])));
                    end
                  reg2385 <= reg2306[(2'h3):(2'h3)];
                  for (forvar2386 = (1'h0); (forvar2386 < (1'h1)); forvar2386 = (forvar2386 + (1'h1)))
                    begin
                      reg2387 <= ($signed({{forvar2298}}) ?
                          ((reg2333 * $unsigned(reg2354)) + reg2155[(3'h5):(1'h1)]) : reg2317[(4'h9):(3'h4)]);
                      reg2388 <= $unsigned(reg2005[(4'hc):(3'h7)]);
                      reg2389 <= ($signed($unsigned($unsigned(reg2037))) ?
                          reg2118[(1'h0):(1'h0)] : forvar2048);
                      reg2390 <= $signed((!(&((8'ha8) ?
                          forvar2053 : reg2219))));
                    end
                  if (($signed($unsigned(((8'h9d) ? (8'hb4) : reg1979))) ?
                      $signed((~|{forvar2212})) : {(^~$unsigned(reg2026))}))
                    begin
                      reg2391 <= (&(8'h9e));
                      reg2392 <= reg2052;
                      reg2393 <= $signed($unsigned($unsigned(forvar2177[(4'hb):(1'h1)])));
                      reg2394 <= (((~&(+(8'ha1))) ?
                              reg2400 : $signed($unsigned(forvar2103))) ?
                          ((-reg2318[(2'h2):(2'h2)]) ?
                              ($unsigned((8'ha1)) ^~ (reg2137 ?
                                  reg2424 : reg2268)) : forvar2349[(3'h6):(1'h1)]) : $signed(reg2400));
                    end
                  else
                    begin
                      reg2391 <= $unsigned(($unsigned($signed(reg2398)) > $unsigned($unsigned((8'haa)))));
                    end
                end
              if ($signed($signed({(8'hb4)})))
                begin
                  for (forvar2395 = (1'h0); (forvar2395 < (2'h2)); forvar2395 = (forvar2395 + (1'h1)))
                    begin
                      reg2396 <= ((~^$signed(reg2434[(1'h0):(1'h0)])) ^~ (&$unsigned($signed(reg2069))));
                    end
                  if ($signed(forvar2270))
                    begin
                      reg2397 <= forvar1974;
                      reg2398 <= ((((~reg1994) | (reg2335 & forvar2050)) >>> forvar2004[(2'h2):(2'h2)]) >= (reg2183 >= $signed(reg2046[(3'h4):(1'h1)])));
                      reg2399 <= ((~^(reg2002[(3'h6):(2'h3)] ?
                          (^reg2187) : reg1985[(1'h0):(1'h0)])) >>> reg2301[(4'h9):(2'h2)]);
                      reg2400 <= reg2158[(4'h8):(2'h3)];
                    end
                  else
                    begin
                      reg2397 <= $unsigned(($unsigned(reg1934[(3'h6):(1'h1)]) >>> $unsigned((forvar1998 ?
                          reg2179 : reg2270))));
                      reg2398 <= forvar2172;
                    end
                  reg2401 <= $signed((~&{(^(8'ha0))}));
                  for (forvar2402 = (1'h0); (forvar2402 < (1'h0)); forvar2402 = (forvar2402 + (1'h1)))
                    begin
                      reg2403 <= $signed($signed(reg2280));
                      reg2404 <= (-($unsigned(((8'ha4) & reg1934)) >>> $signed((reg2275 | (8'ha2)))));
                      reg2405 <= reg2012[(3'h5):(3'h4)];
                    end
                end
              else
                begin
                  reg2395 <= $unsigned(({reg2351} ?
                      $unsigned($unsigned(reg2105)) : $signed(forvar2048)));
                end
              reg2406 <= reg2094[(1'h0):(1'h0)];
            end
          for (forvar2407 = (1'h0); (forvar2407 < (2'h2)); forvar2407 = (forvar2407 + (1'h1)))
            begin
              reg2408 <= (~^reg2290[(4'he):(4'hc)]);
              reg2409 <= $signed({(!$unsigned(reg2287))});
            end
          if ({{(reg2278[(2'h3):(1'h0)] ? reg1957[(4'h8):(2'h2)] : (8'haf))}})
            begin
              for (forvar2410 = (1'h0); (forvar2410 < (2'h2)); forvar2410 = (forvar2410 + (1'h1)))
                begin
                  reg2411 <= ((reg2373 ?
                      {forvar2162[(4'hc):(4'h8)]} : ((reg2027 ?
                          forvar2392 : (8'haf)) != $unsigned((8'ha8)))) ^ $signed(($unsigned((8'ha4)) ?
                      $unsigned(forvar2229) : forvar2282)));
                  if ($unsigned($signed(forvar2111[(1'h1):(1'h0)])))
                    begin
                      reg2412 <= (reg2178 <= reg2306[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2412 <= $unsigned(($signed((~&(8'hac))) ?
                          (-forvar2322) : ((|forvar2275) == $unsigned(reg2087))));
                      reg2413 <= reg1970;
                    end
                end
              if ((^~((~&(8'h9f)) ?
                  ((^reg2312) && (reg2169 * forvar2136)) : forvar2418[(4'hd):(2'h2)])))
                begin
                  if ($signed($signed((~$unsigned(reg2241)))))
                    begin
                      reg2414 <= forvar2213;
                      reg2415 <= reg1991[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2414 <= reg2127;
                      reg2415 <= (~&reg2419);
                      reg2416 <= ((^$unsigned($unsigned(forvar2132))) || (((forvar1967 ?
                          reg2091 : forvar2168) - (reg1951 - reg1962)) >>> ($unsigned(reg2223) >> $signed((8'ha0)))));
                      reg2417 <= forvar2296;
                    end
                  if (($signed({(forvar1980 ?
                          reg2215 : reg2336)}) ^~ {reg1985[(1'h1):(1'h0)]}))
                    begin
                      reg2418 <= (((~|reg2192) ?
                          $signed((forvar2287 ?
                              reg2312 : reg1992)) : $signed((^reg2156))) <= ($signed((reg2018 ?
                          forvar1930 : forvar2351)) * reg2347));
                      reg2419 <= reg2015[(3'h4):(2'h2)];
                      reg2420 <= {(forvar2373[(4'h9):(3'h5)] ?
                              $unsigned($unsigned(forvar2330)) : ((reg1950 ?
                                      (8'ha6) : reg2310) ?
                                  forvar1931 : $signed(forvar2311)))};
                      reg2421 <= {reg2294};
                    end
                  else
                    begin
                      reg2418 <= forvar2078;
                      reg2419 <= (reg2271 ?
                          $unsigned(reg2061[(4'hb):(4'h9)]) : (reg2377 ?
                              ((reg2433 ?
                                  reg2001 : reg2348) - {reg2005}) : reg2385));
                      reg2420 <= reg2206[(4'he):(4'h9)];
                    end
                  if ($unsigned({$signed(forvar1948)}))
                    begin
                      reg2422 <= reg2431;
                      reg2423 <= ($unsigned({reg2413[(1'h1):(1'h1)]}) >> forvar2167[(4'h8):(3'h4)]);
                    end
                  else
                    begin
                      reg2422 <= ({reg2025[(3'h7):(1'h1)]} ^~ reg2270[(3'h4):(2'h3)]);
                      reg2423 <= $unsigned({((8'ha0) ?
                              (-reg2089) : forvar2173[(3'h7):(3'h7)])});
                      reg2424 <= ((&((|forvar2316) + reg2301)) ^ $signed(((reg2108 ?
                              reg2138 : forvar2386) ?
                          reg2130[(1'h0):(1'h0)] : ((8'hb8) * reg2135))));
                    end
                end
              else
                begin
                  for (forvar2414 = (1'h0); (forvar2414 < (1'h0)); forvar2414 = (forvar2414 + (1'h1)))
                    begin
                      reg2415 <= ($signed(forvar2413) ?
                          $signed(forvar2106) : reg2416[(1'h1):(1'h0)]);
                      reg2416 <= $signed({reg2355});
                      reg2417 <= $unsigned((~^reg2403));
                      reg2418 <= (($signed(reg2293) ?
                          reg2245 : $signed((&(8'haa)))) ~^ reg2365[(3'h4):(1'h0)]);
                    end
                end
              for (forvar2425 = (1'h0); (forvar2425 < (1'h1)); forvar2425 = (forvar2425 + (1'h1)))
                begin
                  for (forvar2426 = (1'h0); (forvar2426 < (1'h1)); forvar2426 = (forvar2426 + (1'h1)))
                    begin
                      reg2427 <= $signed($unsigned({(|reg2127)}));
                      reg2428 <= ($unsigned(($signed(reg1955) < forvar2285)) ?
                          (-(8'ha0)) : (~$unsigned((reg2415 > reg2428))));
                    end
                  if ((($unsigned((reg2231 & (8'ha3))) >>> ((reg2112 << (8'hab)) ?
                      (reg2120 << reg2072) : forvar2210[(1'h0):(1'h0)])) >= (-(~^{forvar1998}))))
                    begin
                      reg2429 <= $signed($unsigned($unsigned((reg2315 << reg2295))));
                      reg2430 <= reg2162[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2429 <= {$signed(reg2224)};
                      reg2430 <= (({$unsigned(reg2167)} ?
                              forvar2075 : reg2064) ?
                          (reg2110[(2'h2):(1'h1)] > forvar2066[(3'h4):(3'h4)]) : reg2119);
                    end
                end
              for (forvar2431 = (1'h0); (forvar2431 < (1'h1)); forvar2431 = (forvar2431 + (1'h1)))
                begin
                  for (forvar2432 = (1'h0); (forvar2432 < (1'h0)); forvar2432 = (forvar2432 + (1'h1)))
                    begin
                      reg2433 <= ((forvar2364[(3'h4):(3'h4)] || $unsigned(((8'hb5) ?
                              (8'h9c) : reg2168))) ?
                          reg2090[(2'h3):(2'h2)] : $signed($unsigned((~&(8'haf)))));
                    end
                  for (forvar2434 = (1'h0); (forvar2434 < (1'h0)); forvar2434 = (forvar2434 + (1'h1)))
                    begin
                      reg2435 <= $unsigned(reg1970);
                      reg2436 <= ($unsigned(($signed(reg2198) ?
                              (+reg2146) : (^reg2126))) ?
                          $signed((reg2349 ^ $signed((8'haf)))) : $unsigned((reg2415 ?
                              reg2181[(3'h5):(3'h5)] : (|(8'ha5)))));
                      reg2437 <= (({(forvar2213 < forvar2168)} ?
                          (!reg2047[(4'he):(4'ha)]) : reg2422[(4'h8):(3'h7)]) > $signed($signed((+reg1945))));
                      reg2438 <= (~forvar2228);
                    end
                  reg2439 <= forvar2157[(3'h4):(1'h0)];
                end
            end
          else
            begin
              reg2410 <= forvar1939;
            end
          if ($signed(({$unsigned(forvar2407)} >= reg2384)))
            begin
              reg2440 <= $signed($signed($signed(forvar2322)));
              if (($unsigned(($unsigned(reg2118) >>> (forvar2023 * reg2370))) ?
                  $signed(((reg2070 != (8'ha5)) ?
                      (-forvar1941) : $unsigned(forvar2157))) : ($signed($unsigned(forvar2124)) ?
                      (|$unsigned(reg1938)) : ($signed(reg2424) > (8'hb0)))))
                begin
                  if ((^~forvar2040[(3'h4):(1'h0)]))
                    begin
                      reg2441 <= (forvar2255 <= $unsigned(($signed(reg2318) ^~ reg2347[(1'h0):(1'h0)])));
                      reg2442 <= ($unsigned(reg2162) ?
                          reg2164[(4'h8):(3'h7)] : reg2176);
                      reg2443 <= reg2327[(1'h0):(1'h0)];
                      reg2444 <= (reg2202 ?
                          (~(!(reg2352 ^~ reg1929))) : (~^(reg2423 <= (reg2417 ?
                              forvar2290 : (8'h9f)))));
                    end
                  else
                    begin
                      reg2441 <= forvar2263;
                      reg2442 <= reg2044;
                    end
                  if ((($unsigned((&forvar2228)) << (+$unsigned(reg2260))) + {$unsigned((forvar2164 ?
                          (8'hb0) : forvar1934))}))
                    begin
                      reg2445 <= ((((forvar2124 >> forvar2247) ?
                              $unsigned(reg2286) : (!reg2258)) ?
                          reg2192[(2'h3):(2'h2)] : {$signed(reg2401)}) <= $signed((~&(forvar2420 <<< reg2431))));
                      reg2446 <= ($signed((~(forvar2316 ?
                              (8'hac) : forvar2111))) ?
                          $unsigned(reg2268) : reg1942[(3'h6):(3'h5)]);
                      reg2447 <= {reg2129};
                      reg2448 <= (reg2431[(2'h2):(1'h1)] ?
                          $unsigned({reg2152[(3'h5):(1'h0)]}) : reg2239);
                    end
                  else
                    begin
                      reg2445 <= $signed(reg2267);
                      reg2446 <= (|(~^(reg2306 * (~&reg2410))));
                      reg2447 <= $unsigned(reg2430[(1'h1):(1'h1)]);
                      reg2448 <= $signed(forvar2276);
                    end
                  if ($unsigned({$signed((reg1977 ? reg2089 : reg2201))}))
                    begin
                      reg2449 <= (~&((8'hb5) + (~{forvar2035})));
                      reg2450 <= reg2093;
                      reg2451 <= (~^reg2307);
                      reg2452 <= (($signed((8'hb3)) == reg2101[(1'h0):(1'h0)]) ?
                          ($unsigned(((8'hba) ?
                              (8'ha6) : reg2227)) < $signed(forvar1983[(1'h0):(1'h0)])) : (~|reg1975));
                    end
                  else
                    begin
                      reg2449 <= reg2052;
                      reg2450 <= ((^reg2406[(4'ha):(2'h2)]) ?
                          ((reg2351[(1'h1):(1'h1)] ?
                              $signed(reg2405) : ((8'ha0) <<< reg2340)) < $unsigned((8'ha3))) : (reg2200 ?
                              forvar2359[(4'hf):(2'h2)] : (^~$signed(forvar2128))));
                      reg2451 <= $unsigned($signed($signed((reg1944 ?
                          forvar2418 : reg2014))));
                      reg2452 <= $signed((($signed(reg2441) ?
                              $unsigned(forvar2126) : ((8'haf) <= reg2194)) ?
                          $unsigned($signed(reg2020)) : reg2103));
                    end
                  if (forvar2322)
                    begin
                      reg2453 <= forvar2122[(1'h0):(1'h0)];
                      reg2454 <= ((($unsigned(forvar1999) ?
                          forvar2410[(3'h4):(3'h4)] : (~^forvar2143)) - $signed(reg2269[(3'h5):(3'h4)])) << reg2054[(2'h2):(1'h0)]);
                      reg2455 <= {(((reg2237 >> (8'hb4)) ?
                                  (reg2440 & forvar2011) : (reg2398 ?
                                      reg2449 : reg2284)) ?
                              forvar2283[(4'h8):(3'h7)] : $signed(reg2110[(1'h0):(1'h0)]))};
                      reg2456 <= reg2219[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg2453 <= (&($signed((reg2113 ? reg2056 : reg2092)) ?
                          (reg2043 >> (-reg2349)) : ({(8'ha9)} * forvar2316)));
                      reg2454 <= reg2450[(4'h8):(1'h0)];
                      reg2455 <= (((reg2165[(1'h0):(1'h0)] ^ $signed(forvar1983)) == $signed($unsigned(reg2150))) + (8'haa));
                    end
                end
              else
                begin
                  for (forvar2441 = (1'h0); (forvar2441 < (2'h3)); forvar2441 = (forvar2441 + (1'h1)))
                    begin
                      reg2442 <= (8'hb6);
                      reg2443 <= {reg1945[(3'h6):(3'h4)]};
                      reg2444 <= $unsigned(($signed($signed((8'h9f))) ?
                          reg2334[(2'h3):(1'h1)] : reg2403[(1'h0):(1'h0)]));
                      reg2445 <= $signed(((-reg2080) < $signed($signed(forvar2162))));
                    end
                  if ($unsigned($unsigned((8'hb8))))
                    begin
                      reg2446 <= ((reg2401 ?
                              $unsigned((reg2207 << reg2258)) : (reg2050[(3'h7):(2'h2)] ?
                                  {(8'hb7)} : $unsigned((8'ha6)))) ?
                          (~reg2309) : $signed($unsigned(((8'ha6) ?
                              wire1924 : (8'had)))));
                      reg2447 <= $signed((reg1937 & (reg2186[(1'h1):(1'h1)] ?
                          (~(8'hb9)) : $signed((8'ha2)))));
                      reg2448 <= reg2003;
                      reg2449 <= $unsigned((-(+$unsigned(reg2010))));
                    end
                  else
                    begin
                      reg2446 <= ($signed($signed(forvar1936[(1'h1):(1'h0)])) ?
                          forvar2434[(1'h1):(1'h1)] : $unsigned($unsigned((~|reg2064))));
                    end
                  for (forvar2450 = (1'h0); (forvar2450 < (1'h1)); forvar2450 = (forvar2450 + (1'h1)))
                    begin
                      reg2451 <= $unsigned($signed($signed($signed(reg2239))));
                      reg2452 <= ((~&forvar2392) << {$unsigned((reg2354 ?
                              (8'ha8) : reg2109))});
                      reg2453 <= ((reg2099 ?
                              (~(reg1936 ? (8'haf) : reg2310)) : forvar1967) ?
                          ($unsigned($signed(reg2374)) >>> ({(8'h9c)} ?
                              reg2150[(4'h9):(1'h0)] : $signed(reg1990))) : reg2237);
                    end
                  reg2454 <= {reg1958};
                end
            end
          else
            begin
              for (forvar2440 = (1'h0); (forvar2440 < (2'h2)); forvar2440 = (forvar2440 + (1'h1)))
                begin
                  for (forvar2441 = (1'h0); (forvar2441 < (1'h0)); forvar2441 = (forvar2441 + (1'h1)))
                    begin
                      reg2442 <= forvar2212[(4'h9):(3'h5)];
                      reg2443 <= (~|forvar2086);
                      reg2444 <= $unsigned({$unsigned($signed(reg2052))});
                      reg2445 <= {(|forvar2281)};
                    end
                  for (forvar2446 = (1'h0); (forvar2446 < (2'h2)); forvar2446 = (forvar2446 + (1'h1)))
                    begin
                      reg2447 <= reg2191[(4'h8):(3'h4)];
                    end
                  for (forvar2448 = (1'h0); (forvar2448 < (1'h0)); forvar2448 = (forvar2448 + (1'h1)))
                    begin
                      reg2449 <= reg2158;
                      reg2450 <= forvar2115[(3'h6):(1'h0)];
                    end
                  for (forvar2451 = (1'h0); (forvar2451 < (2'h3)); forvar2451 = (forvar2451 + (1'h1)))
                    begin
                      reg2452 <= (8'ha9);
                      reg2453 <= (~reg1996);
                      reg2454 <= reg2434[(3'h7):(3'h7)];
                      reg2455 <= ($unsigned(reg1975) ?
                          (|$unsigned($unsigned(reg2042))) : {($unsigned((8'hb5)) ?
                                  (forvar2168 ? (8'ha8) : reg2098) : reg2224)});
                    end
                end
              if (reg2215)
                begin
                  for (forvar2456 = (1'h0); (forvar2456 < (2'h2)); forvar2456 = (forvar2456 + (1'h1)))
                    begin
                      reg2457 <= (($signed($signed(reg2331)) <= (-$signed(reg2262))) & (~forvar1948[(3'h6):(2'h3)]));
                      reg2458 <= ((|forvar2362[(4'ha):(1'h0)]) >= (reg2254[(1'h1):(1'h0)] ?
                          {$unsigned(forvar2228)} : $signed((reg2344 ?
                              reg2365 : reg2397))));
                      reg2459 <= forvar2351[(4'h9):(2'h2)];
                      reg2460 <= reg2375;
                    end
                  for (forvar2461 = (1'h0); (forvar2461 < (2'h2)); forvar2461 = (forvar2461 + (1'h1)))
                    begin
                      reg2462 <= (~|(+((reg2155 <<< (8'hb7)) ?
                          $signed((8'had)) : (reg2347 == (8'ha1)))));
                      reg2463 <= (+(8'hba));
                    end
                  if (($signed($unsigned((!forvar2270))) * $signed($signed((forvar2431 ?
                      reg2416 : (8'hb9))))))
                    begin
                      reg2464 <= reg2396;
                    end
                  else
                    begin
                      reg2464 <= $signed(reg2326[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar2456 = (1'h0); (forvar2456 < (2'h2)); forvar2456 = (forvar2456 + (1'h1)))
                    begin
                      reg2457 <= ((reg1995[(1'h1):(1'h0)] <= ($signed(reg1991) ?
                              reg2459[(3'h6):(1'h1)] : {(8'ha8)})) ?
                          forvar2187 : forvar2325[(4'hb):(4'h9)]);
                    end
                end
            end
        end
    end
  assign wire2465 = $signed($unsigned(forvar1974[(4'hb):(4'h8)]));
  always
    @(posedge clk) begin
      for (forvar2466 = (1'h0); (forvar2466 < (1'h0)); forvar2466 = (forvar2466 + (1'h1)))
        begin
          if ($unsigned({($signed(reg2074) ? {reg2280} : reg2090)}))
            begin
              for (forvar2467 = (1'h0); (forvar2467 < (1'h0)); forvar2467 = (forvar2467 + (1'h1)))
                begin
                  if ($unsigned({forvar2162}))
                    begin
                      reg2468 <= (reg2346[(2'h2):(1'h1)] - $unsigned((^~reg2304[(3'h4):(1'h1)])));
                      reg2469 <= forvar2395;
                      reg2470 <= forvar2023;
                      reg2471 <= ((-reg2186) <<< reg2123);
                    end
                  else
                    begin
                      reg2468 <= $unsigned(($signed((^reg2236)) ?
                          reg2094[(1'h1):(1'h0)] : $unsigned({forvar2410})));
                    end
                  for (forvar2472 = (1'h0); (forvar2472 < (1'h1)); forvar2472 = (forvar2472 + (1'h1)))
                    begin
                      reg2473 <= $unsigned(((|reg2453[(4'h9):(1'h0)]) > $unsigned($signed(reg2374))));
                    end
                  reg2474 <= ($unsigned(((forvar2001 ?
                          reg2221 : forvar2352) < (^~reg1983))) ?
                      $signed($unsigned(reg2412)) : (8'h9d));
                end
              for (forvar2475 = (1'h0); (forvar2475 < (2'h2)); forvar2475 = (forvar2475 + (1'h1)))
                begin
                  for (forvar2476 = (1'h0); (forvar2476 < (2'h3)); forvar2476 = (forvar2476 + (1'h1)))
                    begin
                      reg2477 <= reg2302[(3'h4):(2'h3)];
                      reg2478 <= (reg2107[(3'h4):(1'h0)] ?
                          $signed(reg2266) : reg2119[(1'h1):(1'h0)]);
                    end
                  for (forvar2479 = (1'h0); (forvar2479 < (2'h2)); forvar2479 = (forvar2479 + (1'h1)))
                    begin
                      reg2480 <= (^~forvar2162[(3'h5):(2'h3)]);
                      reg2481 <= (^~$signed(reg2092[(2'h3):(1'h1)]));
                    end
                  for (forvar2482 = (1'h0); (forvar2482 < (1'h0)); forvar2482 = (forvar2482 + (1'h1)))
                    begin
                      reg2483 <= ($signed((forvar2354[(1'h0):(1'h0)] + (!forvar2028))) & ((-(forvar2311 ?
                              reg2009 : reg2182)) ?
                          reg2404 : (8'hb5)));
                    end
                  for (forvar2484 = (1'h0); (forvar2484 < (1'h1)); forvar2484 = (forvar2484 + (1'h1)))
                    begin
                      reg2485 <= reg2180;
                      reg2486 <= (reg2319[(1'h0):(1'h0)] ?
                          reg2112[(1'h1):(1'h1)] : forvar2355[(3'h4):(1'h0)]);
                    end
                end
              if (reg1974)
                begin
                  for (forvar2487 = (1'h0); (forvar2487 < (1'h0)); forvar2487 = (forvar2487 + (1'h1)))
                    begin
                      reg2488 <= forvar2007[(1'h1):(1'h0)];
                      reg2489 <= (~&reg2092[(1'h1):(1'h1)]);
                    end
                  reg2490 <= $unsigned({(reg2378[(1'h1):(1'h0)] || (reg2314 > reg2291))});
                end
              else
                begin
                  if (reg1983)
                    begin
                      reg2487 <= reg1978[(4'h9):(3'h6)];
                      reg2488 <= reg2418;
                    end
                  else
                    begin
                      reg2487 <= $unsigned($unsigned((~^(reg2261 ?
                          forvar2382 : (8'ha7)))));
                      reg2488 <= $signed((forvar2322[(1'h0):(1'h0)] ?
                          ((^reg2346) | (~^forvar2015)) : ({forvar2436} ?
                              (+forvar1962) : forvar2290[(2'h2):(1'h0)])));
                    end
                  for (forvar2489 = (1'h0); (forvar2489 < (1'h1)); forvar2489 = (forvar2489 + (1'h1)))
                    begin
                      reg2490 <= (!(($unsigned(reg2188) ?
                          reg1932 : forvar2370[(3'h4):(1'h1)]) >= (forvar2410 & (^(8'hb4)))));
                      reg2491 <= $unsigned((((reg2016 ? (8'hb0) : reg2404) ?
                              reg2413[(3'h4):(1'h0)] : $signed((8'hb8))) ?
                          $unsigned((8'ha4)) : {(reg2331 ?
                                  reg2446 : (8'ha4))}));
                      reg2492 <= $unsigned({$signed(forvar2243)});
                      reg2493 <= (!{(~(&reg1993))});
                    end
                  if ((({(reg2148 ? (8'ha0) : forvar2383)} ?
                      reg2427 : reg2088[(3'h4):(1'h1)]) >= (~{$signed(forvar2484)})))
                    begin
                      reg2494 <= reg2165;
                    end
                  else
                    begin
                      reg2494 <= $unsigned((8'hb0));
                      reg2495 <= $unsigned(reg2053);
                    end
                end
              for (forvar2496 = (1'h0); (forvar2496 < (2'h2)); forvar2496 = (forvar2496 + (1'h1)))
                begin
                  for (forvar2497 = (1'h0); (forvar2497 < (2'h3)); forvar2497 = (forvar2497 + (1'h1)))
                    begin
                      reg2498 <= reg2205[(3'h4):(2'h3)];
                      reg2499 <= reg2200;
                      reg2500 <= (~&reg2407);
                    end
                  for (forvar2501 = (1'h0); (forvar2501 < (1'h0)); forvar2501 = (forvar2501 + (1'h1)))
                    begin
                      reg2502 <= ($signed(((reg1942 ~^ forvar2201) > (~reg2449))) ?
                          reg2329 : (-forvar1939[(3'h4):(1'h0)]));
                      reg2503 <= $signed((reg1964 >> (~&forvar2354)));
                      reg2504 <= ((reg2314 ~^ reg1986[(3'h6):(3'h4)]) > $unsigned(reg2306[(2'h2):(1'h1)]));
                      reg2505 <= (($signed(reg2017) ?
                              (reg2443 ?
                                  reg2080 : $signed(reg2357)) : reg2460) ?
                          reg2431 : (~&forvar2487));
                    end
                  for (forvar2506 = (1'h0); (forvar2506 < (2'h2)); forvar2506 = (forvar2506 + (1'h1)))
                    begin
                      reg2507 <= {$unsigned((+reg2412))};
                      reg2508 <= $unsigned((~$signed(forvar1933)));
                      reg2509 <= (8'had);
                    end
                  for (forvar2510 = (1'h0); (forvar2510 < (1'h1)); forvar2510 = (forvar2510 + (1'h1)))
                    begin
                      reg2511 <= $unsigned(($unsigned((wire1927 ?
                          (8'hae) : reg2039)) < forvar2387));
                    end
                end
            end
          else
            begin
              if ((^~reg2326[(3'h7):(3'h5)]))
                begin
                  for (forvar2467 = (1'h0); (forvar2467 < (2'h3)); forvar2467 = (forvar2467 + (1'h1)))
                    begin
                      reg2468 <= ($signed($unsigned({reg2105})) > $unsigned($unsigned((^~forvar1948))));
                    end
                  reg2469 <= (&($signed((~&reg2413)) < $unsigned($signed(reg2252))));
                end
              else
                begin
                  if ($signed($unsigned({reg1996[(4'hb):(3'h7)]})))
                    begin
                      reg2467 <= (reg2276 != reg1947);
                      reg2468 <= (|forvar2357);
                      reg2469 <= $unsigned($signed(($unsigned((8'hb4)) ?
                          $signed(forvar2311) : $unsigned((8'ha2)))));
                    end
                  else
                    begin
                      reg2467 <= (reg2014 >= $signed(reg2148[(4'h9):(2'h2)]));
                      reg2468 <= ((!reg2284) ?
                          forvar2028[(1'h0):(1'h0)] : $unsigned(forvar2348[(1'h0):(1'h0)]));
                      reg2469 <= ((((~&forvar2166) ?
                              {reg2102} : (~&reg2216)) < (&(reg2425 ?
                              forvar2255 : reg2312))) ?
                          (~|((!reg2424) ?
                              reg1958 : $unsigned(reg2418))) : reg2371[(3'h5):(1'h1)]);
                    end
                  reg2470 <= forvar2062[(1'h0):(1'h0)];
                  for (forvar2471 = (1'h0); (forvar2471 < (2'h3)); forvar2471 = (forvar2471 + (1'h1)))
                    begin
                      reg2472 <= $unsigned($unsigned((forvar2028[(2'h3):(2'h3)] ?
                          reg1996 : {(8'ha9)})));
                    end
                end
              if (forvar2348)
                begin
                  reg2473 <= $unsigned($unsigned({forvar2162}));
                  if (($unsigned((reg2072[(1'h1):(1'h1)] ~^ {reg2188})) <<< $signed(reg2061[(4'h8):(1'h1)])))
                    begin
                      reg2474 <= forvar2325[(4'ha):(3'h4)];
                      reg2475 <= (~&reg2486);
                      reg2476 <= $unsigned(($signed((reg2305 ?
                              reg2341 : (8'hb5))) ?
                          $signed((reg2123 ^ reg2204)) : (reg2002 <= {forvar2011})));
                    end
                  else
                    begin
                      reg2474 <= (+((forvar2414 <<< (~|reg2092)) ?
                          $unsigned($unsigned(forvar2053)) : $signed((~(8'hb7)))));
                      reg2475 <= reg2462[(1'h0):(1'h0)];
                      reg2476 <= $signed({(^~(forvar2436 ?
                              reg2398 : forvar2323))});
                      reg2477 <= reg2352[(4'ha):(1'h1)];
                    end
                end
              else
                begin
                  if (($unsigned(((reg2032 ? reg2260 : (8'hb8)) <= reg2107)) ?
                      $signed((forvar2280 * reg2342[(4'h8):(2'h2)])) : $signed((forvar2001 > ((8'ha7) * reg1957)))))
                    begin
                      reg2473 <= (8'hb0);
                      reg2474 <= $signed(((|((8'hae) >>> reg2492)) ?
                          $signed((forvar2418 ?
                              reg2077 : forvar2040)) : $unsigned(reg2261)));
                    end
                  else
                    begin
                      reg2473 <= {(!($signed((8'h9f)) ~^ (reg2385 != (8'had))))};
                    end
                  for (forvar2475 = (1'h0); (forvar2475 < (2'h2)); forvar2475 = (forvar2475 + (1'h1)))
                    begin
                      reg2476 <= $unsigned($unsigned(reg2344[(1'h1):(1'h0)]));
                    end
                end
            end
          reg2512 <= ($unsigned(forvar2116[(3'h5):(3'h5)]) ?
              (-((reg2347 > (8'hba)) != forvar2313[(2'h2):(2'h2)])) : {$signed(reg2056)});
          for (forvar2513 = (1'h0); (forvar2513 < (2'h3)); forvar2513 = (forvar2513 + (1'h1)))
            begin
              if (((&reg2031) <<< (+(~&wire1926[(3'h5):(2'h2)]))))
                begin
                  for (forvar2514 = (1'h0); (forvar2514 < (1'h0)); forvar2514 = (forvar2514 + (1'h1)))
                    begin
                      reg2515 <= (($signed({(8'ha1)}) ?
                              (8'ha5) : {$unsigned(reg2003)}) ?
                          $unsigned(($signed(forvar2124) <= $unsigned(reg2071))) : reg2236);
                      reg2516 <= (+(8'hb1));
                      reg2517 <= $signed($unsigned(({reg2200} ?
                          (+reg2059) : (+(8'hb5)))));
                    end
                  for (forvar2518 = (1'h0); (forvar2518 < (2'h3)); forvar2518 = (forvar2518 + (1'h1)))
                    begin
                      reg2519 <= reg1983[(2'h3):(2'h2)];
                      reg2520 <= $signed(forvar1956);
                      reg2521 <= reg2314;
                    end
                  if ((8'hae))
                    begin
                      reg2522 <= $unsigned($signed((reg2107 < $unsigned(reg2350))));
                    end
                  else
                    begin
                      reg2522 <= forvar2020;
                    end
                  for (forvar2523 = (1'h0); (forvar2523 < (1'h1)); forvar2523 = (forvar2523 + (1'h1)))
                    begin
                      reg2524 <= (forvar2111[(1'h1):(1'h1)] == forvar2205[(3'h4):(2'h3)]);
                      reg2525 <= reg2317[(3'h5):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar2514 = (1'h0); (forvar2514 < (2'h2)); forvar2514 = (forvar2514 + (1'h1)))
                    begin
                      reg2515 <= reg1979;
                      reg2516 <= ({$unsigned(reg2072)} ?
                          (8'hac) : $unsigned(($unsigned(reg2097) && forvar2162[(4'ha):(4'h9)])));
                      reg2517 <= $unsigned(forvar2399[(1'h0):(1'h0)]);
                    end
                  reg2518 <= reg1963;
                  for (forvar2519 = (1'h0); (forvar2519 < (1'h1)); forvar2519 = (forvar2519 + (1'h1)))
                    begin
                      reg2520 <= reg2258;
                      reg2521 <= (!{$signed($unsigned(reg1944))});
                    end
                  if (reg1936)
                    begin
                      reg2522 <= (~^$unsigned(reg2254[(2'h2):(2'h2)]));
                      reg2523 <= $unsigned((|reg2273[(2'h2):(2'h2)]));
                      reg2524 <= $unsigned(($signed(reg1954[(2'h2):(1'h1)]) | $unsigned((reg1978 >>> forvar2301))));
                    end
                  else
                    begin
                      reg2522 <= ((({forvar2467} >= (forvar2102 >> reg2067)) ^~ reg2152) || (+(|{reg1938})));
                      reg2523 <= $signed($signed(reg2376));
                      reg2524 <= (^forvar2301);
                    end
                end
            end
          for (forvar2526 = (1'h0); (forvar2526 < (2'h3)); forvar2526 = (forvar2526 + (1'h1)))
            begin
              if ((($unsigned($signed(forvar2028)) ?
                      ($unsigned(reg2367) <<< reg2038) : ($signed(forvar2210) + reg2489[(2'h3):(1'h0)])) ?
                  {reg2222[(3'h5):(2'h3)]} : $unsigned((reg2070 ^~ reg2200))))
                begin
                  reg2527 <= (8'h9f);
                  for (forvar2528 = (1'h0); (forvar2528 < (1'h1)); forvar2528 = (forvar2528 + (1'h1)))
                    begin
                      reg2529 <= reg2056;
                      reg2530 <= reg1994;
                    end
                  for (forvar2531 = (1'h0); (forvar2531 < (2'h2)); forvar2531 = (forvar2531 + (1'h1)))
                    begin
                      reg2532 <= (+((+(forvar2298 ?
                          (8'ha1) : forvar2349)) >= (forvar1962 > (reg2471 ?
                          forvar2392 : forvar2420))));
                    end
                  if ({(((forvar2167 ? reg2192 : wire1927) && (forvar2040 ?
                          reg2245 : forvar2279)) && ((reg2507 ?
                          forvar2399 : reg2408) || (reg2192 ^ reg2109)))})
                    begin
                      reg2533 <= reg2098;
                      reg2534 <= ({{(reg1985 == reg2489)}} ?
                          reg2221 : $signed(reg2284));
                      reg2535 <= reg2226[(1'h1):(1'h0)];
                      reg2536 <= $signed($unsigned(($unsigned(reg2486) ?
                          $signed(reg2252) : (reg2020 ? reg2234 : reg2388))));
                    end
                  else
                    begin
                      reg2533 <= $unsigned($unsigned($signed($unsigned(forvar2287))));
                    end
                end
              else
                begin
                  for (forvar2527 = (1'h0); (forvar2527 < (1'h1)); forvar2527 = (forvar2527 + (1'h1)))
                    begin
                      reg2528 <= (~&(|(|reg2242)));
                      reg2529 <= forvar2409;
                      reg2530 <= $unsigned({reg1990[(1'h1):(1'h1)]});
                      reg2531 <= $signed($unsigned(reg2071));
                    end
                  if (reg1970[(3'h5):(2'h3)])
                    begin
                      reg2532 <= reg2242;
                    end
                  else
                    begin
                      reg2532 <= (~(reg2450 ?
                          $unsigned(forvar2451[(1'h1):(1'h1)]) : $signed($unsigned((8'had)))));
                      reg2533 <= ($signed(forvar2434) ?
                          reg2458[(2'h2):(1'h1)] : (reg2312[(2'h2):(1'h1)] != ($signed(forvar2519) ~^ {reg2431})));
                      reg2534 <= reg2487[(2'h3):(2'h2)];
                      reg2535 <= (8'ha1);
                    end
                  for (forvar2536 = (1'h0); (forvar2536 < (1'h1)); forvar2536 = (forvar2536 + (1'h1)))
                    begin
                      reg2537 <= {(~^{$unsigned(reg2160)})};
                      reg2538 <= reg2488;
                    end
                end
              if (($unsigned((reg1937 ?
                      forvar2373[(1'h0):(1'h0)] : $signed(reg2060))) ?
                  (~&$unsigned(reg2272[(1'h1):(1'h1)])) : reg2152))
                begin
                  if ((~^($signed($signed(reg1990)) >> reg2258)))
                    begin
                      reg2539 <= (^~(~|$signed($signed(forvar2434))));
                      reg2540 <= $signed({((reg2164 ^~ forvar2179) >> $signed(forvar2220))});
                      reg2541 <= $signed({(^~reg1979)});
                    end
                  else
                    begin
                      reg2539 <= (8'h9c);
                      reg2540 <= $signed($unsigned(((forvar1936 ~^ (8'hb1)) >>> (+reg2091))));
                      reg2541 <= reg2140[(3'h5):(1'h0)];
                      reg2542 <= {(reg1931 ?
                              $unsigned((reg2104 != (8'hb5))) : $unsigned(reg2232[(1'h0):(1'h0)]))};
                    end
                  for (forvar2543 = (1'h0); (forvar2543 < (1'h1)); forvar2543 = (forvar2543 + (1'h1)))
                    begin
                      reg2544 <= (^({$unsigned((8'hb1))} > reg1993[(2'h2):(1'h0)]));
                      reg2545 <= reg2088[(4'h8):(1'h1)];
                      reg2546 <= reg2079;
                      reg2547 <= reg2384[(1'h1):(1'h1)];
                    end
                  if (($signed(reg2098[(3'h7):(2'h3)]) ?
                      $unsigned($unsigned(reg2034[(2'h3):(1'h0)])) : $signed($unsigned({reg2445}))))
                    begin
                      reg2548 <= {reg2523[(4'ha):(3'h7)]};
                    end
                  else
                    begin
                      reg2548 <= $signed($signed($unsigned((forvar2285 && (8'hba)))));
                      reg2549 <= ($signed(({reg2320} ?
                              $signed(reg2087) : reg1982)) ?
                          forvar2426 : $unsigned(forvar1963));
                    end
                end
              else
                begin
                  for (forvar2539 = (1'h0); (forvar2539 < (1'h1)); forvar2539 = (forvar2539 + (1'h1)))
                    begin
                      reg2540 <= reg2050[(4'h9):(3'h7)];
                      reg2541 <= ({reg2442} ? reg2271[(1'h0):(1'h0)] : reg2025);
                      reg2542 <= ((&((forvar2062 >> reg2380) <<< $signed(reg2037))) ?
                          reg2518 : ({(+reg2021)} ?
                              forvar2451 : ((^reg2327) <= (reg2128 || reg2198))));
                    end
                end
              for (forvar2550 = (1'h0); (forvar2550 < (2'h2)); forvar2550 = (forvar2550 + (1'h1)))
                begin
                  for (forvar2551 = (1'h0); (forvar2551 < (1'h0)); forvar2551 = (forvar2551 + (1'h1)))
                    begin
                      reg2552 <= ({$unsigned((&reg2417))} <<< (reg2373 ?
                          (&(forvar2475 ?
                              (8'hb0) : forvar2536)) : $signed(reg2256)));
                      reg2553 <= (+$unsigned(($signed(reg2324) ?
                          $signed(forvar2229) : reg2357[(3'h6):(1'h1)])));
                      reg2554 <= (^($signed($unsigned(reg2446)) ?
                          reg1938 : ((!reg2423) ?
                              (forvar2475 ? reg2390 : reg2552) : (&(8'hb9)))));
                      reg2555 <= $signed((forvar1970[(3'h6):(2'h3)] ?
                          (8'hb7) : (~^reg2493[(3'h4):(3'h4)])));
                    end
                  for (forvar2556 = (1'h0); (forvar2556 < (1'h1)); forvar2556 = (forvar2556 + (1'h1)))
                    begin
                      reg2557 <= reg2480;
                      reg2558 <= ($unsigned($unsigned((-forvar2466))) ?
                          ((8'ha0) >= $signed((forvar2392 + reg2172))) : $signed({$signed(forvar2330)}));
                      reg2559 <= $signed(reg2140);
                      reg2560 <= {reg2161[(3'h5):(1'h0)]};
                    end
                  reg2561 <= $unsigned($unsigned((reg2318 <= (reg2442 << reg2256))));
                end
              for (forvar2562 = (1'h0); (forvar2562 < (2'h3)); forvar2562 = (forvar2562 + (1'h1)))
                begin
                  if ((^($unsigned(reg2013[(3'h4):(1'h1)]) ?
                      (reg2101 >>> (forvar2102 >= forvar2475)) : reg2103)))
                    begin
                      reg2563 <= (&(~^reg2355));
                      reg2564 <= reg2449;
                    end
                  else
                    begin
                      reg2563 <= (forvar2348 ?
                          $signed({$signed(reg2394)}) : ((~$unsigned(reg2046)) ^ {((8'had) & reg2369)}));
                      reg2564 <= (8'haf);
                      reg2565 <= (({{(8'hba)}} ?
                              (!(reg2546 & forvar2162)) : (&(reg2135 > reg2279))) ?
                          $signed($signed({reg2152})) : reg2401[(2'h2):(1'h1)]);
                      reg2566 <= ($unsigned(reg2539[(2'h3):(1'h0)]) ?
                          $signed(forvar2187[(2'h3):(2'h3)]) : $signed($signed(reg2193[(3'h7):(3'h7)])));
                    end
                  if ((~|$unsigned((|(reg2525 << reg2324)))))
                    begin
                      reg2567 <= $signed((forvar2052 ?
                          $unsigned((|forvar2279)) : (^~{reg2314})));
                    end
                  else
                    begin
                      reg2567 <= (^~{(&$unsigned(forvar2539))});
                      reg2568 <= reg1981;
                      reg2569 <= (forvar2164[(4'h8):(1'h0)] & (($signed((8'ha0)) ?
                              reg1978 : reg2538[(1'h0):(1'h0)]) ?
                          forvar2382 : $unsigned((reg2294 ?
                              reg2104 : forvar2153))));
                      reg2570 <= (~^$signed((reg2411[(3'h7):(1'h0)] ?
                          reg2186 : (+forvar2015))));
                    end
                  if ($signed($signed($unsigned((reg2357 ?
                      reg2416 : (8'ha5))))))
                    begin
                      reg2571 <= ({$unsigned((reg2377 || forvar2539))} == {((-(8'hb3)) ?
                              (~^reg2195) : reg2163)});
                    end
                  else
                    begin
                      reg2571 <= {$unsigned(reg2442[(4'he):(2'h3)])};
                      reg2572 <= ({$signed((reg2384 ?
                              reg2375 : forvar2351))} <= (forvar2075 >> $signed(reg2182)));
                      reg2573 <= reg2291;
                      reg2574 <= {((-reg2467) ?
                              reg2265[(4'ha):(2'h2)] : {$signed(wire1927)})};
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(forvar2293[(4'h8):(3'h7)])))
        begin
          for (forvar2575 = (1'h0); (forvar2575 < (1'h0)); forvar2575 = (forvar2575 + (1'h1)))
            begin
              if ($unsigned(reg2119[(3'h7):(3'h7)]))
                begin
                  for (forvar2576 = (1'h0); (forvar2576 < (1'h0)); forvar2576 = (forvar2576 + (1'h1)))
                    begin
                      reg2577 <= (8'haf);
                      reg2578 <= reg2367[(1'h0):(1'h0)];
                      reg2579 <= reg2154[(2'h2):(1'h0)];
                      reg2580 <= (^$unsigned(forvar2373[(4'h9):(4'h8)]));
                    end
                  for (forvar2581 = (1'h0); (forvar2581 < (2'h2)); forvar2581 = (forvar2581 + (1'h1)))
                    begin
                      reg2582 <= forvar2096;
                    end
                  reg2583 <= reg2003;
                end
              else
                begin
                  reg2576 <= reg2211;
                  for (forvar2577 = (1'h0); (forvar2577 < (1'h1)); forvar2577 = (forvar2577 + (1'h1)))
                    begin
                      reg2578 <= ((reg2319 ^ ((~&(8'hb8)) <<< $signed(reg2504))) * ((-forvar2392[(1'h1):(1'h0)]) < $signed((reg2003 < (8'ha8)))));
                      reg2579 <= (&((((8'h9e) ?
                              reg1969 : (8'ha0)) ^~ (!forvar2075)) ?
                          ((^(8'ha6)) <= (+(8'h9d))) : $signed(reg2296[(3'h5):(1'h0)])));
                      reg2580 <= $unsigned($signed(reg2473[(3'h4):(3'h4)]));
                      reg2581 <= $signed($signed(reg2101));
                    end
                  if ((^~(-(reg2565 ?
                      (reg2419 <= reg2110) : forvar2420[(4'ha):(3'h7)]))))
                    begin
                      reg2582 <= (~^(reg2268[(1'h1):(1'h1)] ?
                          $signed($unsigned((8'hb2))) : {$unsigned(forvar2526)}));
                      reg2583 <= {(-(~^(~|reg2544)))};
                      reg2584 <= $unsigned(reg1981);
                      reg2585 <= $signed($unsigned({(reg2121 ?
                              (8'ha4) : forvar1943)}));
                    end
                  else
                    begin
                      reg2582 <= forvar2581[(1'h1):(1'h0)];
                      reg2583 <= reg2103[(1'h1):(1'h0)];
                    end
                  for (forvar2586 = (1'h0); (forvar2586 < (1'h0)); forvar2586 = (forvar2586 + (1'h1)))
                    begin
                      reg2587 <= ($signed((8'h9d)) ~^ $unsigned(((reg2284 && (8'h9d)) <<< $unsigned(reg1990))));
                      reg2588 <= $signed({reg2308[(4'ha):(2'h2)]});
                      reg2589 <= ({$signed($unsigned(reg2162))} == reg2015[(3'h5):(1'h0)]);
                      reg2590 <= ((((reg2189 < (8'ha3)) ?
                          (reg2572 ?
                              reg2227 : reg2275) : reg2343) || ($signed(forvar2432) || {reg2428})) - ((((8'hb2) ?
                                  reg2503 : forvar2451) ?
                              $signed(forvar2263) : (forvar2373 ?
                                  forvar2506 : reg2487)) ?
                          (forvar2243[(1'h1):(1'h0)] ?
                              reg2155 : (reg2419 ^~ reg2503)) : $unsigned({(8'haa)})));
                    end
                end
            end
        end
      else
        begin
          reg2575 <= reg2395;
          for (forvar2576 = (1'h0); (forvar2576 < (2'h2)); forvar2576 = (forvar2576 + (1'h1)))
            begin
              reg2577 <= (((~&(reg2205 ? forvar2440 : reg2507)) ?
                      $signed(reg2225[(2'h3):(2'h2)]) : ($signed(forvar2163) >>> forvar2487)) ?
                  reg2036[(1'h1):(1'h0)] : {(^(+forvar2100))});
              for (forvar2578 = (1'h0); (forvar2578 < (1'h1)); forvar2578 = (forvar2578 + (1'h1)))
                begin
                  if ({forvar1971[(3'h7):(3'h4)]})
                    begin
                      reg2579 <= (((^reg2326) ?
                          $signed((^reg1984)) : $unsigned(reg2232)) >>> $unsigned($signed($signed(reg2318))));
                      reg2580 <= forvar2100[(2'h2):(1'h0)];
                      reg2581 <= $unsigned($signed(reg2029));
                      reg2582 <= (~&$unsigned({(&reg2201)}));
                    end
                  else
                    begin
                      reg2579 <= reg2219;
                      reg2580 <= (forvar2166 <= (reg2319[(3'h4):(2'h2)] ?
                          (!$unsigned(forvar2082)) : reg2306));
                    end
                end
            end
          for (forvar2583 = (1'h0); (forvar2583 < (1'h1)); forvar2583 = (forvar2583 + (1'h1)))
            begin
              for (forvar2584 = (1'h0); (forvar2584 < (1'h1)); forvar2584 = (forvar2584 + (1'h1)))
                begin
                  for (forvar2585 = (1'h0); (forvar2585 < (2'h2)); forvar2585 = (forvar2585 + (1'h1)))
                    begin
                      reg2586 <= ((^~forvar2434) >= {{(~|(8'ha3))}});
                    end
                end
              for (forvar2587 = (1'h0); (forvar2587 < (2'h3)); forvar2587 = (forvar2587 + (1'h1)))
                begin
                  reg2588 <= (|reg2535);
                  for (forvar2589 = (1'h0); (forvar2589 < (1'h1)); forvar2589 = (forvar2589 + (1'h1)))
                    begin
                      reg2590 <= (&reg2452[(1'h0):(1'h0)]);
                      reg2591 <= $signed($unsigned(reg2138[(1'h1):(1'h0)]));
                      reg2592 <= reg2343;
                      reg2593 <= (forvar2096 || reg2191);
                    end
                  for (forvar2594 = (1'h0); (forvar2594 < (1'h0)); forvar2594 = (forvar2594 + (1'h1)))
                    begin
                      reg2595 <= (($signed($unsigned(reg1991)) & reg2579) ?
                          $unsigned((8'haf)) : (forvar2475[(2'h2):(2'h2)] < $signed((^reg1963))));
                      reg2596 <= reg2536[(2'h2):(1'h0)];
                      reg2597 <= reg2230[(2'h3):(1'h1)];
                      reg2598 <= (~&(($unsigned(reg2047) ?
                              (reg2242 * reg2318) : {forvar2325}) ?
                          $signed($unsigned(reg2571)) : $unsigned((reg1936 ?
                              forvar1963 : forvar2228))));
                    end
                  if (((&$unsigned(reg2519[(1'h0):(1'h0)])) * (8'haa)))
                    begin
                      reg2599 <= (~|reg2166[(2'h3):(1'h0)]);
                      reg2600 <= reg2067;
                      reg2601 <= (($signed($signed(reg2422)) ^~ (-(forvar2335 << forvar2379))) ?
                          reg2286 : {(^~(~^reg2319))});
                      reg2602 <= $signed($signed((8'hac)));
                    end
                  else
                    begin
                      reg2599 <= reg2450[(3'h5):(2'h3)];
                      reg2600 <= (|(+((reg2582 * reg2293) > {(8'hb7)})));
                    end
                end
            end
        end
      for (forvar2603 = (1'h0); (forvar2603 < (2'h3)); forvar2603 = (forvar2603 + (1'h1)))
        begin
          for (forvar2604 = (1'h0); (forvar2604 < (1'h0)); forvar2604 = (forvar2604 + (1'h1)))
            begin
              for (forvar2605 = (1'h0); (forvar2605 < (2'h2)); forvar2605 = (forvar2605 + (1'h1)))
                begin
                  for (forvar2606 = (1'h0); (forvar2606 < (1'h1)); forvar2606 = (forvar2606 + (1'h1)))
                    begin
                      reg2607 <= (forvar2298 + (8'haa));
                      reg2608 <= forvar2355;
                      reg2609 <= (~^($unsigned(reg2236[(1'h1):(1'h1)]) ?
                          (&(reg2140 ?
                              reg2017 : reg2569)) : (&$signed(reg2230))));
                    end
                  reg2610 <= reg2427[(3'h5):(2'h2)];
                end
            end
          reg2611 <= reg2344;
          for (forvar2612 = (1'h0); (forvar2612 < (2'h3)); forvar2612 = (forvar2612 + (1'h1)))
            begin
              if (forvar2086[(4'ha):(4'h8)])
                begin
                  for (forvar2613 = (1'h0); (forvar2613 < (1'h1)); forvar2613 = (forvar2613 + (1'h1)))
                    begin
                      reg2614 <= reg2369[(4'h8):(4'h8)];
                    end
                  reg2615 <= $unsigned($unsigned(($unsigned(reg2300) + (&reg2277))));
                end
              else
                begin
                  if ((~&(($unsigned((8'hb2)) ? {(8'hb5)} : $signed((8'hb3))) ?
                      ((|forvar2577) ?
                          (^~reg2602) : {forvar2182}) : ((~&reg2495) | forvar2095[(2'h3):(1'h1)]))))
                    begin
                      reg2613 <= ((^reg2535[(1'h1):(1'h1)]) ?
                          reg2532[(4'ha):(1'h0)] : $unsigned(((8'h9e) || (forvar2428 ?
                              reg2129 : reg2218))));
                      reg2614 <= reg2252[(3'h5):(1'h1)];
                      reg2615 <= reg2103;
                      reg2616 <= reg2200;
                    end
                  else
                    begin
                      reg2613 <= forvar2613[(2'h3):(2'h3)];
                      reg2614 <= $unsigned($unsigned(($unsigned(forvar2528) != reg2279[(1'h0):(1'h0)])));
                    end
                end
              if (reg2054[(1'h1):(1'h0)])
                begin
                  if ($signed((({reg2460} ?
                          ((8'ha0) ?
                              (8'ha6) : reg2488) : reg2044[(2'h2):(1'h0)]) ?
                      reg2337 : $unsigned((&reg2596)))))
                    begin
                      reg2617 <= $unsigned(($unsigned(reg2232) ?
                          (reg2425 ?
                              reg2371 : (forvar2510 != reg2370)) : (&$unsigned(forvar2604))));
                    end
                  else
                    begin
                      reg2617 <= $signed($signed((-reg2428[(2'h3):(2'h2)])));
                      reg2618 <= (^$signed(reg2200));
                      reg2619 <= (8'h9f);
                    end
                end
              else
                begin
                  reg2617 <= {(reg2318 >> $signed($signed(reg1993)))};
                  for (forvar2618 = (1'h0); (forvar2618 < (1'h0)); forvar2618 = (forvar2618 + (1'h1)))
                    begin
                      reg2619 <= {$unsigned(forvar2187)};
                      reg2620 <= $signed((8'ha2));
                      reg2621 <= ($signed((+$signed(reg1951))) ?
                          reg2554[(1'h0):(1'h0)] : $unsigned(($unsigned(reg1946) ?
                              (forvar1936 ? reg1977 : (8'hb3)) : (-reg2113))));
                    end
                  if ($signed(((~^{forvar2410}) ?
                      reg2025 : forvar2612[(4'hc):(3'h7)])))
                    begin
                      reg2622 <= reg1948;
                      reg2623 <= (reg2413[(2'h3):(2'h3)] - reg2142[(4'ha):(2'h3)]);
                    end
                  else
                    begin
                      reg2622 <= (|$signed($signed($signed(reg1965))));
                    end
                  for (forvar2624 = (1'h0); (forvar2624 < (1'h0)); forvar2624 = (forvar2624 + (1'h1)))
                    begin
                      reg2625 <= {($unsigned((8'hb1)) * $signed($unsigned(reg2074)))};
                      reg2626 <= reg2058;
                      reg2627 <= forvar1936;
                    end
                end
              if ((8'hac))
                begin
                  for (forvar2628 = (1'h0); (forvar2628 < (1'h1)); forvar2628 = (forvar2628 + (1'h1)))
                    begin
                      reg2629 <= $unsigned((((reg2306 && (8'hba)) ?
                              ((8'hb8) << forvar2618) : (&reg1993)) ?
                          (8'hb6) : $signed(((8'haa) * reg2061))));
                    end
                  for (forvar2630 = (1'h0); (forvar2630 < (1'h0)); forvar2630 = (forvar2630 + (1'h1)))
                    begin
                      reg2631 <= (!$unsigned((~$unsigned(forvar2167))));
                      reg2632 <= reg2503;
                    end
                  if ((8'ha8))
                    begin
                      reg2633 <= forvar2577;
                      reg2634 <= (|reg2393);
                      reg2635 <= $signed($unsigned(((forvar2461 ^ reg2528) ?
                          $unsigned(reg2591) : (forvar2143 ?
                              forvar1939 : forvar2428))));
                      reg2636 <= reg2302;
                    end
                  else
                    begin
                      reg2633 <= reg2591[(4'h8):(3'h5)];
                      reg2634 <= reg2189;
                      reg2635 <= reg2231[(3'h6):(2'h2)];
                    end
                  reg2637 <= ({(reg2220 ? $signed(reg2481) : reg2402)} ?
                      {$signed((^~reg2352))} : forvar2023[(2'h2):(1'h0)]);
                end
              else
                begin
                  for (forvar2628 = (1'h0); (forvar2628 < (1'h1)); forvar2628 = (forvar2628 + (1'h1)))
                    begin
                      reg2629 <= {(~|reg2359)};
                    end
                  if ({(!(reg2434 <= (reg2046 ? reg2627 : forvar2311)))})
                    begin
                      reg2630 <= reg1933[(3'h6):(3'h5)];
                      reg2631 <= reg2424;
                    end
                  else
                    begin
                      reg2630 <= reg2394[(3'h4):(2'h3)];
                      reg2631 <= $signed($unsigned(reg2554[(2'h3):(2'h3)]));
                    end
                end
            end
          for (forvar2638 = (1'h0); (forvar2638 < (2'h3)); forvar2638 = (forvar2638 + (1'h1)))
            begin
              if ($unsigned((&(!$signed(reg2487)))))
                begin
                  for (forvar2639 = (1'h0); (forvar2639 < (2'h3)); forvar2639 = (forvar2639 + (1'h1)))
                    begin
                      reg2640 <= ($unsigned((~^reg2273[(2'h2):(1'h1)])) & ((forvar2311[(2'h2):(1'h1)] ?
                              (&forvar2583) : (reg2352 == (8'hb3))) ?
                          $signed(reg2595) : reg2312));
                      reg2641 <= (forvar2173[(4'hb):(2'h2)] << $unsigned($unsigned((forvar2450 << (8'hb9)))));
                      reg2642 <= ((8'ha8) || ($unsigned(reg2359[(4'hd):(3'h5)]) ?
                          reg2244[(2'h3):(2'h2)] : $signed({forvar2414})));
                      reg2643 <= ((reg2305 < $unsigned((~forvar2436))) ?
                          (~^((reg2129 - (8'hac)) ?
                              reg1985[(2'h3):(1'h0)] : (8'ha1))) : reg2457[(4'he):(3'h7)]);
                    end
                  reg2644 <= $unsigned((^(|$signed(forvar2349))));
                  reg2645 <= (&wire1926);
                  for (forvar2646 = (1'h0); (forvar2646 < (2'h2)); forvar2646 = (forvar2646 + (1'h1)))
                    begin
                      reg2647 <= ((($unsigned(reg2067) >= (8'h9c)) ?
                          reg2421[(4'hb):(4'h9)] : (8'haa)) * (&$signed(reg2365[(1'h0):(1'h0)])));
                      reg2648 <= {{$signed((~|reg2121))}};
                      reg2649 <= ({reg2564} <<< {(^~$unsigned((8'hb8)))});
                      reg2650 <= ({reg2128[(4'h9):(2'h2)]} || reg1957);
                    end
                end
              else
                begin
                  reg2639 <= ((~reg2191) ?
                      $unsigned($signed($unsigned(reg2430))) : ((^~reg2447) ?
                          $unsigned(reg2630) : $signed(reg2309[(3'h7):(1'h0)])));
                end
              for (forvar2651 = (1'h0); (forvar2651 < (1'h0)); forvar2651 = (forvar2651 + (1'h1)))
                begin
                  if (reg2622)
                    begin
                      reg2652 <= $signed((!$signed($signed(reg2156))));
                      reg2653 <= ($unsigned(((8'hb4) || $unsigned(reg2380))) <= ($signed((reg2161 ?
                              (8'hac) : (8'hb5))) ?
                          ($signed((8'hab)) ?
                              {(8'h9d)} : reg2265) : $signed((reg2006 - reg2249))));
                    end
                  else
                    begin
                      reg2652 <= $unsigned($signed({reg2545[(3'h5):(2'h2)]}));
                    end
                  for (forvar2654 = (1'h0); (forvar2654 < (2'h3)); forvar2654 = (forvar2654 + (1'h1)))
                    begin
                      reg2655 <= forvar1936[(1'h0):(1'h0)];
                      reg2656 <= reg1986;
                      reg2657 <= (-$signed(($signed(reg2165) && (forvar2179 ?
                          reg2107 : reg2131))));
                    end
                  for (forvar2658 = (1'h0); (forvar2658 < (1'h1)); forvar2658 = (forvar2658 + (1'h1)))
                    begin
                      reg2659 <= {$unsigned(((reg2128 <<< reg2585) ?
                              (reg2003 ? forvar2208 : reg2272) : (^~reg2584)))};
                    end
                end
            end
        end
    end
  assign wire2660 = ($unsigned($unsigned(forvar2078)) >>> reg2310);
  assign wire2661 = ((&($signed(reg2246) || reg2345)) || (((8'ha1) >> reg2163) ^~ $unsigned(reg2537[(2'h2):(1'h1)])));
  assign wire2662 = reg2591;
  assign wire2663 = (reg2342[(5'h10):(3'h7)] ?
                        reg2477[(1'h0):(1'h0)] : $unsigned(reg2613));
  assign wire2664 = reg2205;
  assign wire2665 = $unsigned(({(~&(8'hae))} && reg2038));
  assign wire2666 = (~|(reg2038 ~^ $signed((reg2223 | forvar2414))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1509
#(parameter param1734 = (!(~|({(8'hb6)} ? (~^(8'h9d)) : (!(8'h9d))))))
(y, clk, wire1510, wire1511, wire1512, wire1513);
  output wire [(32'h33a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire1510;
  input wire [(4'hf):(1'h0)] wire1511;
  input wire [(4'he):(1'h0)] wire1512;
  input wire signed [(4'hb):(1'h0)] wire1513;
  wire signed [(2'h3):(1'h0)] wire1733;
  reg [(4'h8):(1'h0)] reg1732 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1731 = (1'h0);
  reg [(4'hd):(1'h0)] reg1730 = (1'h0);
  reg [(3'h4):(1'h0)] reg1729 = (1'h0);
  reg [(3'h4):(1'h0)] reg1728 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1727 = (1'h0);
  reg [(2'h3):(1'h0)] reg1726 = (1'h0);
  reg [(4'h8):(1'h0)] reg1725 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1724 = (1'h0);
  reg [(4'h8):(1'h0)] reg1723 = (1'h0);
  reg [(3'h4):(1'h0)] reg1722 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1721 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1720 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1719 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1718 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1717 = (1'h0);
  reg [(2'h3):(1'h0)] reg1716 = (1'h0);
  reg [(2'h3):(1'h0)] reg1715 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1714 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1713 = (1'h0);
  reg [(4'h9):(1'h0)] reg1712 = (1'h0);
  reg [(4'ha):(1'h0)] reg1711 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1710 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1709 = (1'h0);
  reg [(4'h9):(1'h0)] reg1708 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1707 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1705 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1701 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1706 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1705 = (1'h0);
  reg [(5'h10):(1'h0)] reg1704 = (1'h0);
  reg [(5'h10):(1'h0)] reg1703 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1702 = (1'h0);
  reg [(4'hf):(1'h0)] reg1701 = (1'h0);
  reg [(4'hb):(1'h0)] reg1700 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1699 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1698 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1697 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1694 = (1'h0);
  reg [(3'h6):(1'h0)] reg1696 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1695 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1694 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1693 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1692 = (1'h0);
  reg [(3'h7):(1'h0)] reg1691 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1690 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1689 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1688 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1687 = (1'h0);
  reg [(2'h3):(1'h0)] reg1686 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1685 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1684 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1683 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1682 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1675 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1666 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1662 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1674 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1672 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1670 = (1'h0);
  reg [(2'h2):(1'h0)] reg1668 = (1'h0);
  reg [(4'h8):(1'h0)] reg1678 = (1'h0);
  reg [(3'h6):(1'h0)] reg1676 = (1'h0);
  reg [(2'h2):(1'h0)] reg1681 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1680 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1679 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1678 = (1'h0);
  reg [(5'h10):(1'h0)] reg1677 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1676 = (1'h0);
  reg [(3'h7):(1'h0)] reg1675 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1674 = (1'h0);
  reg [(4'hf):(1'h0)] reg1673 = (1'h0);
  reg [(4'h8):(1'h0)] reg1672 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1671 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1670 = (1'h0);
  reg [(2'h3):(1'h0)] reg1669 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1667 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1666 = (1'h0);
  reg [(3'h4):(1'h0)] reg1664 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1663 = (1'h0);
  reg [(2'h2):(1'h0)] reg1665 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1664 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1663 = (1'h0);
  reg [(4'he):(1'h0)] forvar1662 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1661 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1660 = (1'h0);
  reg [(3'h5):(1'h0)] reg1659 = (1'h0);
  reg [(4'ha):(1'h0)] reg1658 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1657 = (1'h0);
  reg [(2'h2):(1'h0)] reg1656 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1655 = (1'h0);
  reg [(3'h5):(1'h0)] reg1654 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1653 = (1'h0);
  reg [(2'h2):(1'h0)] reg1652 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1651 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1650 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1649 = (1'h0);
  wire [(3'h5):(1'h0)] wire1514;
  wire signed [(5'h10):(1'h0)] wire1647;
  assign y = {wire1733,
                 reg1732,
                 reg1731,
                 reg1730,
                 reg1729,
                 reg1728,
                 reg1727,
                 reg1726,
                 reg1725,
                 forvar1724,
                 reg1723,
                 reg1722,
                 reg1721,
                 reg1720,
                 reg1719,
                 forvar1718,
                 reg1717,
                 reg1716,
                 reg1715,
                 forvar1714,
                 forvar1713,
                 reg1712,
                 reg1711,
                 forvar1710,
                 reg1709,
                 reg1708,
                 reg1707,
                 forvar1705,
                 forvar1701,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1703,
                 reg1702,
                 reg1701,
                 reg1700,
                 reg1699,
                 forvar1698,
                 reg1697,
                 forvar1694,
                 reg1696,
                 reg1695,
                 reg1694,
                 forvar1693,
                 reg1692,
                 reg1691,
                 forvar1690,
                 reg1689,
                 reg1688,
                 reg1687,
                 reg1686,
                 forvar1685,
                 reg1684,
                 forvar1683,
                 reg1682,
                 forvar1675,
                 forvar1666,
                 reg1662,
                 reg1674,
                 forvar1672,
                 reg1670,
                 reg1668,
                 reg1678,
                 reg1676,
                 reg1681,
                 reg1680,
                 reg1679,
                 forvar1678,
                 reg1677,
                 forvar1676,
                 reg1675,
                 forvar1674,
                 reg1673,
                 reg1672,
                 reg1671,
                 forvar1670,
                 reg1669,
                 forvar1668,
                 reg1667,
                 reg1666,
                 reg1664,
                 forvar1663,
                 reg1665,
                 forvar1664,
                 reg1663,
                 forvar1662,
                 reg1661,
                 reg1660,
                 reg1659,
                 reg1658,
                 reg1657,
                 reg1656,
                 reg1655,
                 reg1654,
                 reg1653,
                 reg1652,
                 forvar1651,
                 forvar1650,
                 forvar1649,
                 wire1514,
                 wire1647,
                 (1'h0)};
  assign wire1514 = ((((~|(8'hb2)) | {(8'h9e)}) ?
                            (wire1512 >= (wire1511 ?
                                wire1511 : (8'hb7))) : wire1511[(4'hc):(4'ha)]) ?
                        (~^wire1513) : ($unsigned(wire1510[(4'h9):(1'h1)]) ^~ $unsigned(wire1511)));
  module1515 modinst1648 (.clk(clk), .y(wire1647), .wire1517(wire1510), .wire1516(wire1511), .wire1520(wire1512), .wire1519(wire1513), .wire1518(wire1514));
  always
    @(posedge clk) begin
      for (forvar1649 = (1'h0); (forvar1649 < (2'h2)); forvar1649 = (forvar1649 + (1'h1)))
        begin
          for (forvar1650 = (1'h0); (forvar1650 < (1'h1)); forvar1650 = (forvar1650 + (1'h1)))
            begin
              if ((~|wire1511))
                begin
                  for (forvar1651 = (1'h0); (forvar1651 < (2'h2)); forvar1651 = (forvar1651 + (1'h1)))
                    begin
                      reg1652 <= {$unsigned(((forvar1651 >>> forvar1649) << forvar1650))};
                      reg1653 <= ($unsigned(($signed(wire1510) ?
                          (~(8'haa)) : $signed(forvar1650))) >> (((forvar1651 >>> wire1510) >> wire1647[(3'h6):(2'h3)]) ^ $signed(forvar1649)));
                      reg1654 <= $signed({wire1511[(4'h9):(2'h2)]});
                    end
                  if ((forvar1649 | (({reg1652} < (8'ha3)) << (&$unsigned(wire1514)))))
                    begin
                      reg1655 <= $unsigned(($signed(wire1513) ?
                          wire1647[(4'h8):(3'h7)] : ((reg1654 || reg1652) >> (wire1510 ?
                              forvar1650 : wire1513))));
                      reg1656 <= {{forvar1649}};
                      reg1657 <= $signed(forvar1651);
                    end
                  else
                    begin
                      reg1655 <= (!$unsigned((|(forvar1650 ?
                          forvar1651 : reg1656))));
                      reg1656 <= $unsigned(reg1653[(1'h0):(1'h0)]);
                      reg1657 <= wire1513;
                    end
                  if ({($unsigned($signed(wire1511)) != reg1655[(2'h2):(1'h0)])})
                    begin
                      reg1658 <= (($unsigned((8'hb6)) ?
                          forvar1651[(1'h1):(1'h0)] : wire1510[(3'h6):(2'h3)]) + (wire1510 ?
                          $unsigned(forvar1649) : (8'h9c)));
                      reg1659 <= $unsigned(wire1513[(4'h8):(1'h0)]);
                    end
                  else
                    begin
                      reg1658 <= ({{reg1655}} <<< ($signed((forvar1650 ?
                              wire1510 : reg1656)) ?
                          wire1511 : wire1513[(2'h3):(2'h3)]));
                      reg1659 <= ($signed((8'ha5)) ?
                          (^~reg1658[(2'h2):(2'h2)]) : {(|reg1652[(1'h0):(1'h0)])});
                      reg1660 <= reg1656[(2'h2):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar1651 = (1'h0); (forvar1651 < (1'h0)); forvar1651 = (forvar1651 + (1'h1)))
                    begin
                      reg1652 <= (8'hba);
                      reg1653 <= ($unsigned(wire1513[(4'ha):(3'h4)]) ?
                          $signed(($unsigned(reg1654) ?
                              $signed(reg1659) : {wire1510})) : $signed(((reg1657 * wire1511) ?
                              wire1514 : (&(8'hb3)))));
                      reg1654 <= $unsigned((&{$signed(forvar1651)}));
                      reg1655 <= reg1657[(3'h5):(2'h3)];
                    end
                end
              reg1661 <= (reg1657[(1'h1):(1'h1)] <= wire1510[(4'he):(4'hd)]);
            end
        end
      if ((^~(((8'h9d) ?
          $signed(wire1514) : forvar1650) < reg1657[(2'h2):(2'h2)])))
        begin
          if ((8'hab))
            begin
              for (forvar1662 = (1'h0); (forvar1662 < (1'h0)); forvar1662 = (forvar1662 + (1'h1)))
                begin
                  reg1663 <= forvar1651[(1'h1):(1'h1)];
                  for (forvar1664 = (1'h0); (forvar1664 < (1'h1)); forvar1664 = (forvar1664 + (1'h1)))
                    begin
                      reg1665 <= ((wire1511 << (^{wire1513})) - {$unsigned((|forvar1649))});
                    end
                end
            end
          else
            begin
              for (forvar1662 = (1'h0); (forvar1662 < (1'h0)); forvar1662 = (forvar1662 + (1'h1)))
                begin
                  for (forvar1663 = (1'h0); (forvar1663 < (1'h1)); forvar1663 = (forvar1663 + (1'h1)))
                    begin
                      reg1664 <= $unsigned(((~&$signed(reg1653)) ?
                          (reg1659 < {reg1659}) : $signed(reg1661[(1'h1):(1'h0)])));
                      reg1665 <= $unsigned(reg1658[(2'h3):(1'h1)]);
                      reg1666 <= $unsigned((|$signed(reg1660[(4'ha):(3'h4)])));
                      reg1667 <= $signed(wire1513);
                    end
                  for (forvar1668 = (1'h0); (forvar1668 < (2'h3)); forvar1668 = (forvar1668 + (1'h1)))
                    begin
                      reg1669 <= $signed($signed({forvar1663[(4'ha):(2'h3)]}));
                    end
                end
              if (wire1647[(4'ha):(4'ha)])
                begin
                  for (forvar1670 = (1'h0); (forvar1670 < (1'h0)); forvar1670 = (forvar1670 + (1'h1)))
                    begin
                      reg1671 <= $unsigned(reg1653[(2'h3):(1'h0)]);
                      reg1672 <= $unsigned((((forvar1664 <= (8'hb0)) ?
                              (!reg1661) : {wire1512}) ?
                          $unsigned((reg1655 ^ reg1653)) : ((reg1667 ?
                              (8'ha1) : reg1661) >> (reg1656 ?
                              wire1514 : (8'h9d)))));
                      reg1673 <= {forvar1663[(3'h4):(1'h1)]};
                    end
                  for (forvar1674 = (1'h0); (forvar1674 < (1'h1)); forvar1674 = (forvar1674 + (1'h1)))
                    begin
                      reg1675 <= reg1666;
                    end
                  for (forvar1676 = (1'h0); (forvar1676 < (2'h2)); forvar1676 = (forvar1676 + (1'h1)))
                    begin
                      reg1677 <= $unsigned(reg1655[(1'h1):(1'h1)]);
                    end
                  for (forvar1678 = (1'h0); (forvar1678 < (1'h1)); forvar1678 = (forvar1678 + (1'h1)))
                    begin
                      reg1679 <= (forvar1649[(4'ha):(1'h1)] >= ($unsigned($signed(reg1671)) ?
                          (reg1663 ?
                              $unsigned((8'ha2)) : {forvar1651}) : forvar1678));
                      reg1680 <= (^~($signed(reg1672[(1'h1):(1'h1)]) ?
                          wire1647[(4'hc):(3'h6)] : ((~|wire1514) ?
                              (reg1679 + wire1510) : $signed((8'ha6)))));
                      reg1681 <= forvar1674;
                    end
                end
              else
                begin
                  for (forvar1670 = (1'h0); (forvar1670 < (1'h0)); forvar1670 = (forvar1670 + (1'h1)))
                    begin
                      reg1671 <= $signed($unsigned($signed($unsigned(reg1667))));
                      reg1672 <= $signed((+(~|(8'hac))));
                      reg1673 <= forvar1678;
                    end
                  for (forvar1674 = (1'h0); (forvar1674 < (2'h2)); forvar1674 = (forvar1674 + (1'h1)))
                    begin
                      reg1675 <= $signed(reg1666);
                      reg1676 <= {reg1657};
                      reg1677 <= reg1673[(1'h0):(1'h0)];
                      reg1678 <= reg1657;
                    end
                end
            end
        end
      else
        begin
          if (reg1677[(3'h6):(3'h6)])
            begin
              if (reg1666[(3'h4):(2'h2)])
                begin
                  for (forvar1662 = (1'h0); (forvar1662 < (1'h1)); forvar1662 = (forvar1662 + (1'h1)))
                    begin
                      reg1663 <= $signed(($unsigned((reg1675 ^ forvar1676)) ~^ reg1659[(3'h5):(1'h1)]));
                      reg1664 <= reg1680;
                    end
                  if (((+(!$unsigned(reg1652))) | $unsigned(wire1510[(4'ha):(2'h2)])))
                    begin
                      reg1665 <= wire1511[(4'ha):(2'h3)];
                      reg1666 <= (((8'haa) ?
                              $unsigned({reg1672}) : ((~&wire1514) ?
                                  wire1510[(1'h1):(1'h1)] : reg1672[(1'h0):(1'h0)])) ?
                          (($signed((8'ha1)) ?
                              reg1680 : $signed((8'hb5))) < reg1656[(1'h0):(1'h0)]) : (-(~&$signed((8'had)))));
                      reg1667 <= {((&(8'ha4)) ?
                              $signed({wire1647}) : forvar1650[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg1665 <= reg1663[(4'h8):(1'h0)];
                      reg1666 <= (+$signed($unsigned((reg1664 * (8'h9e)))));
                      reg1667 <= $unsigned((reg1677[(4'h8):(3'h6)] != $signed({reg1658})));
                      reg1668 <= reg1673[(4'he):(3'h7)];
                    end
                  if ((&$unsigned((((8'haf) >> forvar1663) ?
                      wire1513[(1'h1):(1'h0)] : $unsigned(reg1653)))))
                    begin
                      reg1669 <= forvar1674[(1'h0):(1'h0)];
                      reg1670 <= $signed((($signed(forvar1678) ?
                          ((8'hb9) ?
                              reg1659 : forvar1663) : reg1669[(1'h1):(1'h0)]) ^~ reg1658));
                      reg1671 <= reg1655[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1669 <= reg1659;
                      reg1670 <= $signed((((^~reg1666) ~^ (reg1677 ?
                              reg1657 : (8'had))) ?
                          (reg1659 ?
                              (reg1655 + (8'ha8)) : $unsigned(forvar1674)) : forvar1664[(1'h1):(1'h1)]));
                      reg1671 <= $unsigned(reg1680[(2'h2):(2'h2)]);
                    end
                  for (forvar1672 = (1'h0); (forvar1672 < (1'h1)); forvar1672 = (forvar1672 + (1'h1)))
                    begin
                      reg1673 <= ({((-reg1655) ?
                              reg1658 : (wire1510 << forvar1650))} + (reg1665[(1'h0):(1'h0)] ?
                          reg1653 : ($unsigned(reg1665) ?
                              (reg1663 > forvar1649) : {reg1679})));
                      reg1674 <= reg1672;
                      reg1675 <= $unsigned({{wire1647[(4'hc):(4'hc)]}});
                      reg1676 <= reg1656[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if (($unsigned((~$unsigned(reg1672))) ^ $signed(($signed(reg1679) ?
                      ((8'hab) ^~ forvar1676) : $signed(reg1677)))))
                    begin
                      reg1662 <= (({(forvar1651 ?
                              forvar1664 : reg1653)} ^ (+{(8'ha5)})) * (^((forvar1676 >> reg1681) > reg1670)));
                      reg1663 <= (^$unsigned($unsigned(wire1647)));
                    end
                  else
                    begin
                      reg1662 <= $unsigned(reg1656[(2'h2):(2'h2)]);
                    end
                end
            end
          else
            begin
              for (forvar1662 = (1'h0); (forvar1662 < (1'h1)); forvar1662 = (forvar1662 + (1'h1)))
                begin
                  if ({$signed(((reg1666 ~^ (8'ha6)) ?
                          (~reg1674) : forvar1674[(1'h1):(1'h0)]))})
                    begin
                      reg1663 <= (+(((forvar1676 ? reg1658 : forvar1676) ?
                              ((8'ha0) ?
                                  reg1657 : (8'haa)) : forvar1678[(3'h6):(1'h0)]) ?
                          ((forvar1663 >= reg1666) ^ reg1660) : (forvar1672 << $signed(reg1656))));
                    end
                  else
                    begin
                      reg1663 <= $unsigned($unsigned($unsigned((~|reg1681))));
                      reg1664 <= forvar1674[(3'h5):(1'h1)];
                    end
                  reg1665 <= reg1668[(1'h0):(1'h0)];
                  for (forvar1666 = (1'h0); (forvar1666 < (2'h2)); forvar1666 = (forvar1666 + (1'h1)))
                    begin
                      reg1667 <= (^(!((reg1676 ? forvar1668 : wire1514) ?
                          (reg1679 && (8'hb5)) : (~|(8'hb9)))));
                      reg1668 <= (8'hac);
                      reg1669 <= ($signed(reg1654) ?
                          ((forvar1649 ?
                                  $unsigned(wire1647) : $signed(reg1655)) ?
                              (-(~(8'h9f))) : $unsigned($unsigned((8'hb7)))) : (forvar1678 - $signed((reg1680 >> forvar1672))));
                      reg1670 <= ($unsigned($unsigned(reg1671)) >= $signed(((forvar1662 & reg1673) ?
                          $unsigned((8'h9f)) : (!reg1678))));
                    end
                end
              if ((($signed($unsigned(reg1672)) << $signed({forvar1663})) - (8'hba)))
                begin
                  if ($unsigned($signed($signed((reg1666 * forvar1670)))))
                    begin
                      reg1671 <= $unsigned($unsigned({$unsigned(reg1678)}));
                    end
                  else
                    begin
                      reg1671 <= (~^(($unsigned(reg1672) >= {(8'hab)}) ?
                          (reg1661[(1'h0):(1'h0)] ?
                              (-reg1672) : reg1676) : (8'ha3)));
                      reg1672 <= $signed(((reg1655 >= wire1647) - (((8'hae) == forvar1651) ?
                          $unsigned(reg1679) : forvar1678)));
                    end
                  if (forvar1650[(1'h1):(1'h1)])
                    begin
                      reg1673 <= (&$signed($unsigned(forvar1649)));
                      reg1674 <= $unsigned(reg1666);
                      reg1675 <= forvar1651[(2'h2):(1'h0)];
                      reg1676 <= (((^~wire1511[(3'h6):(1'h0)]) ?
                          (^reg1672) : {(wire1513 >> (8'hb3))}) <= ((~&{(8'hb6)}) ^ ((8'h9f) >> $signed(reg1658))));
                    end
                  else
                    begin
                      reg1673 <= reg1676[(3'h5):(2'h2)];
                    end
                  if (((&{$unsigned(forvar1666)}) ?
                      (forvar1649[(3'h5):(3'h5)] ^ ((forvar1664 ?
                          (8'hb3) : reg1675) ^~ (forvar1664 & reg1670))) : (^((reg1673 == reg1671) && $unsigned(reg1667)))))
                    begin
                      reg1677 <= ($signed(((^~wire1514) < $unsigned((8'hb4)))) >> (~reg1658[(2'h2):(1'h0)]));
                      reg1678 <= forvar1664;
                    end
                  else
                    begin
                      reg1677 <= {forvar1676};
                      reg1678 <= (~(~^({reg1658} ?
                          $signed(reg1660) : $unsigned(reg1652))));
                      reg1679 <= $signed(forvar1666[(3'h6):(3'h6)]);
                    end
                  reg1680 <= reg1669;
                end
              else
                begin
                  if (((reg1669 ?
                          forvar1670 : ($unsigned(forvar1668) >>> (&forvar1664))) ?
                      forvar1650[(3'h4):(1'h0)] : (({reg1661} ?
                          reg1654[(2'h3):(2'h2)] : forvar1651) * (~reg1663))))
                    begin
                      reg1671 <= $unsigned(({(reg1653 ?
                              wire1510 : (8'hb6))} >> reg1671));
                      reg1672 <= ($signed($signed((reg1670 ?
                          reg1671 : (8'hb8)))) <= $unsigned(reg1668));
                      reg1673 <= {$unsigned((((8'had) ^~ reg1677) - reg1664[(1'h1):(1'h0)]))};
                    end
                  else
                    begin
                      reg1671 <= (~|($unsigned((wire1514 | reg1676)) ?
                          reg1663 : {(&reg1670)}));
                      reg1672 <= $signed($signed((8'hb4)));
                      reg1673 <= ((8'ha2) ?
                          (forvar1678[(2'h3):(2'h3)] ?
                              {(reg1652 || reg1653)} : forvar1649[(2'h3):(1'h1)]) : (((|reg1669) ?
                                  forvar1668[(4'hb):(1'h1)] : $unsigned(forvar1672)) ?
                              (|(&reg1679)) : (&((8'ha3) ?
                                  reg1654 : reg1681))));
                      reg1674 <= (8'h9f);
                    end
                  for (forvar1675 = (1'h0); (forvar1675 < (1'h1)); forvar1675 = (forvar1675 + (1'h1)))
                    begin
                      reg1676 <= (&$signed(reg1669));
                      reg1677 <= (-forvar1649);
                      reg1678 <= forvar1672;
                    end
                  if (reg1681)
                    begin
                      reg1679 <= ({$signed(((8'h9c) ? forvar1670 : reg1664))} ?
                          {wire1511[(4'h8):(1'h1)]} : {(~$unsigned(reg1656))});
                      reg1680 <= $unsigned(reg1676);
                    end
                  else
                    begin
                      reg1679 <= forvar1651[(2'h2):(1'h1)];
                      reg1680 <= forvar1662;
                      reg1681 <= (|$signed((&(wire1514 ? reg1676 : reg1667))));
                      reg1682 <= reg1653;
                    end
                end
              for (forvar1683 = (1'h0); (forvar1683 < (1'h0)); forvar1683 = (forvar1683 + (1'h1)))
                begin
                  reg1684 <= ((wire1512[(4'ha):(2'h2)] & {{reg1653}}) || (forvar1676[(1'h1):(1'h1)] >>> (^~reg1671[(1'h1):(1'h1)])));
                  for (forvar1685 = (1'h0); (forvar1685 < (1'h0)); forvar1685 = (forvar1685 + (1'h1)))
                    begin
                      reg1686 <= (!forvar1662[(4'he):(1'h1)]);
                      reg1687 <= (^wire1513[(1'h1):(1'h1)]);
                      reg1688 <= ((reg1673[(1'h0):(1'h0)] ?
                              (^(reg1654 ^~ forvar1664)) : reg1669[(1'h1):(1'h1)]) ?
                          {$signed($unsigned(reg1656))} : (($signed(reg1669) ?
                              forvar1663 : $signed(reg1654)) >> {$unsigned(reg1658)}));
                      reg1689 <= {(($signed(forvar1670) << $unsigned((8'ha1))) <<< ((forvar1672 ?
                              reg1654 : forvar1685) && reg1668))};
                    end
                  for (forvar1690 = (1'h0); (forvar1690 < (1'h1)); forvar1690 = (forvar1690 + (1'h1)))
                    begin
                      reg1691 <= ($signed(((8'hb3) && $unsigned(forvar1650))) ^~ (&forvar1670));
                      reg1692 <= (+{(~|(reg1661 >> reg1674))});
                    end
                end
            end
          for (forvar1693 = (1'h0); (forvar1693 < (1'h0)); forvar1693 = (forvar1693 + (1'h1)))
            begin
              if (wire1513)
                begin
                  if ((-{forvar1650}))
                    begin
                      reg1694 <= {reg1678};
                      reg1695 <= {(forvar1678[(4'h8):(4'h8)] ?
                              reg1660 : reg1686)};
                    end
                  else
                    begin
                      reg1694 <= ((^reg1674[(1'h0):(1'h0)]) ?
                          forvar1690[(1'h1):(1'h1)] : (reg1687[(3'h6):(3'h6)] + {wire1510[(1'h1):(1'h0)]}));
                      reg1695 <= (reg1688[(4'h8):(3'h6)] ?
                          (((+forvar1666) ^ $signed(reg1657)) ?
                              {forvar1693[(3'h4):(1'h1)]} : (8'ha9)) : wire1512[(4'hd):(1'h0)]);
                      reg1696 <= (~&$unsigned($signed(forvar1676)));
                    end
                end
              else
                begin
                  for (forvar1694 = (1'h0); (forvar1694 < (2'h2)); forvar1694 = (forvar1694 + (1'h1)))
                    begin
                      reg1695 <= forvar1650;
                      reg1696 <= (!(~|forvar1670));
                      reg1697 <= reg1672;
                    end
                  for (forvar1698 = (1'h0); (forvar1698 < (1'h1)); forvar1698 = (forvar1698 + (1'h1)))
                    begin
                      reg1699 <= $unsigned($unsigned($signed((8'hb8))));
                      reg1700 <= (wire1511 ^ $signed((^~(~^reg1686))));
                    end
                end
              if ($unsigned($signed($unsigned((~&reg1675)))))
                begin
                  reg1701 <= (~&($unsigned({reg1664}) ?
                      {forvar1698} : $unsigned((forvar1675 ?
                          reg1664 : (8'h9c)))));
                  if ({$signed((reg1677[(3'h7):(3'h7)] * (forvar1683 < forvar1694)))})
                    begin
                      reg1702 <= ((^forvar1651[(1'h1):(1'h0)]) < ($unsigned($signed(reg1687)) | (8'hba)));
                      reg1703 <= forvar1662[(4'hb):(3'h7)];
                      reg1704 <= $signed((^~reg1697));
                    end
                  else
                    begin
                      reg1702 <= (!forvar1674);
                      reg1703 <= {(~&{forvar1664})};
                    end
                  if (($signed($signed((forvar1649 ^ (8'ha6)))) ?
                      (reg1700[(4'h9):(3'h7)] ?
                          reg1671 : reg1664) : $unsigned(((forvar1693 ~^ forvar1683) ?
                          wire1511[(3'h6):(2'h2)] : $unsigned(forvar1675)))))
                    begin
                      reg1705 <= ({$signed(reg1684[(3'h6):(3'h6)])} == reg1703);
                    end
                  else
                    begin
                      reg1705 <= $signed(((reg1684[(3'h6):(3'h6)] ~^ reg1703) & (reg1680 ?
                          reg1664[(2'h2):(1'h0)] : $unsigned(reg1692))));
                    end
                  reg1706 <= ($unsigned(((reg1657 ?
                      reg1692 : reg1659) || $unsigned(reg1694))) || $unsigned((+$unsigned(reg1679))));
                end
              else
                begin
                  for (forvar1701 = (1'h0); (forvar1701 < (2'h3)); forvar1701 = (forvar1701 + (1'h1)))
                    begin
                      reg1702 <= (reg1660[(4'hc):(3'h5)] ^ {(-(forvar1685 ?
                              reg1662 : reg1661))});
                      reg1703 <= reg1697[(2'h2):(2'h2)];
                      reg1704 <= forvar1678[(3'h4):(1'h0)];
                    end
                  for (forvar1705 = (1'h0); (forvar1705 < (2'h2)); forvar1705 = (forvar1705 + (1'h1)))
                    begin
                      reg1706 <= ({reg1682} ?
                          (8'hb8) : $signed(($unsigned(reg1663) >>> (reg1702 | reg1663))));
                      reg1707 <= ((&(^(&reg1681))) ?
                          $signed($unsigned((+forvar1662))) : $unsigned((!reg1703[(3'h5):(1'h1)])));
                      reg1708 <= (~&$signed({reg1652[(1'h0):(1'h0)]}));
                      reg1709 <= $unsigned((!(reg1663 ?
                          (8'hb7) : (reg1655 == reg1703))));
                    end
                  for (forvar1710 = (1'h0); (forvar1710 < (2'h2)); forvar1710 = (forvar1710 + (1'h1)))
                    begin
                      reg1711 <= $unsigned($unsigned(($unsigned(reg1691) != (~|reg1704))));
                      reg1712 <= ($signed(wire1514) ?
                          $signed(wire1512) : (~|(~(8'ha2))));
                    end
                end
              for (forvar1713 = (1'h0); (forvar1713 < (1'h1)); forvar1713 = (forvar1713 + (1'h1)))
                begin
                  for (forvar1714 = (1'h0); (forvar1714 < (2'h3)); forvar1714 = (forvar1714 + (1'h1)))
                    begin
                      reg1715 <= $unsigned((~&reg1687[(3'h7):(3'h5)]));
                    end
                  if ($unsigned({$unsigned($signed(reg1668))}))
                    begin
                      reg1716 <= wire1514;
                    end
                  else
                    begin
                      reg1716 <= reg1700;
                      reg1717 <= ($unsigned($unsigned($signed(forvar1685))) ?
                          $unsigned({(~^forvar1675)}) : ((reg1668 >= forvar1672[(2'h3):(2'h3)]) ?
                              reg1667[(1'h1):(1'h1)] : reg1686[(2'h3):(1'h1)]));
                    end
                  for (forvar1718 = (1'h0); (forvar1718 < (1'h1)); forvar1718 = (forvar1718 + (1'h1)))
                    begin
                      reg1719 <= (8'hb1);
                    end
                end
              if ((reg1659[(2'h3):(2'h2)] ?
                  $signed(forvar1664[(3'h4):(1'h1)]) : $unsigned(reg1711)))
                begin
                  if ($unsigned({$signed((|reg1708))}))
                    begin
                      reg1720 <= reg1719;
                      reg1721 <= (~|(-reg1697[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1720 <= reg1679[(1'h1):(1'h1)];
                      reg1721 <= $unsigned($signed({(reg1682 ?
                              forvar1714 : reg1706)}));
                    end
                  reg1722 <= $unsigned(reg1656);
                end
              else
                begin
                  if ($unsigned((~$signed(forvar1678[(2'h3):(2'h3)]))))
                    begin
                      reg1720 <= $signed(reg1670);
                      reg1721 <= $unsigned((~^$unsigned(reg1673)));
                      reg1722 <= {{forvar1713}};
                      reg1723 <= $signed(($signed($unsigned(reg1684)) ?
                          (~reg1659[(3'h4):(2'h3)]) : reg1657[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg1720 <= {($unsigned((~^reg1670)) && forvar1663[(4'ha):(3'h6)])};
                      reg1721 <= (reg1686 ?
                          {$signed((forvar1701 ?
                                  (8'hb4) : reg1665))} : ((^~(~&reg1692)) ~^ reg1681));
                      reg1722 <= reg1665;
                      reg1723 <= reg1668[(1'h0):(1'h0)];
                    end
                  for (forvar1724 = (1'h0); (forvar1724 < (2'h3)); forvar1724 = (forvar1724 + (1'h1)))
                    begin
                      reg1725 <= wire1647[(2'h3):(2'h3)];
                      reg1726 <= (((^~$unsigned((8'h9e))) * (~|$unsigned(reg1673))) ?
                          reg1676 : ({(+(8'ha5))} - forvar1668[(2'h3):(1'h1)]));
                      reg1727 <= $signed($unsigned((~^reg1676)));
                    end
                  reg1728 <= (-$signed((~&$signed((8'h9d)))));
                  if (reg1672[(4'h8):(1'h0)])
                    begin
                      reg1729 <= wire1510;
                      reg1730 <= wire1512;
                      reg1731 <= $unsigned((forvar1672 ?
                          reg1694[(3'h5):(2'h2)] : reg1709));
                      reg1732 <= reg1672;
                    end
                  else
                    begin
                      reg1729 <= reg1677[(4'h9):(2'h2)];
                    end
                end
            end
        end
    end
  assign wire1733 = {reg1703[(4'h9):(4'h9)]};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module591  (y, clk, wire596, wire595, wire594, wire593, wire592);
  output wire [(32'h1023):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire596;
  input wire [(4'hc):(1'h0)] wire595;
  input wire [(4'hb):(1'h0)] wire594;
  input wire signed [(3'h4):(1'h0)] wire593;
  input wire [(5'h10):(1'h0)] wire592;
  wire [(4'h8):(1'h0)] wire1144;
  wire [(2'h3):(1'h0)] wire1143;
  wire [(2'h3):(1'h0)] wire1142;
  reg [(3'h6):(1'h0)] reg1130 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1128 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1126 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1121 = (1'h0);
  reg [(3'h5):(1'h0)] reg1119 = (1'h0);
  reg [(4'ha):(1'h0)] reg1114 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1111 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1141 = (1'h0);
  reg [(4'h8):(1'h0)] reg1140 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1139 = (1'h0);
  reg [(2'h2):(1'h0)] reg1138 = (1'h0);
  reg [(3'h7):(1'h0)] reg1137 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1136 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1135 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1134 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1133 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1132 = (1'h0);
  reg [(4'hb):(1'h0)] reg1131 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1130 = (1'h0);
  reg [(4'he):(1'h0)] reg1129 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1128 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1127 = (1'h0);
  reg [(4'hf):(1'h0)] reg1126 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1125 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1124 = (1'h0);
  reg [(3'h6):(1'h0)] reg1123 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1122 = (1'h0);
  reg [(4'ha):(1'h0)] reg1121 = (1'h0);
  reg [(4'hd):(1'h0)] reg1120 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1119 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1118 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1117 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1116 = (1'h0);
  reg [(3'h6):(1'h0)] reg1115 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1114 = (1'h0);
  reg [(3'h6):(1'h0)] reg1108 = (1'h0);
  reg [(5'h10):(1'h0)] reg1113 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1112 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1111 = (1'h0);
  reg [(3'h4):(1'h0)] reg1110 = (1'h0);
  reg [(3'h6):(1'h0)] reg1109 = (1'h0);
  reg [(4'he):(1'h0)] forvar1108 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1107 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1087 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1081 = (1'h0);
  reg [(4'hb):(1'h0)] reg1083 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1082 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1079 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1072 = (1'h0);
  reg [(5'h10):(1'h0)] reg1093 = (1'h0);
  reg [(4'h8):(1'h0)] reg1106 = (1'h0);
  reg [(3'h6):(1'h0)] reg1105 = (1'h0);
  reg [(4'hd):(1'h0)] reg1104 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1103 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1102 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1101 = (1'h0);
  reg [(4'h8):(1'h0)] reg1100 = (1'h0);
  reg [(3'h4):(1'h0)] reg1099 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1098 = (1'h0);
  reg [(4'hd):(1'h0)] reg1097 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1096 = (1'h0);
  reg [(2'h3):(1'h0)] reg1095 = (1'h0);
  reg [(4'hf):(1'h0)] reg1094 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1093 = (1'h0);
  reg [(3'h7):(1'h0)] reg1092 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1091 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1090 = (1'h0);
  reg [(2'h2):(1'h0)] reg1089 = (1'h0);
  reg [(3'h4):(1'h0)] reg1088 = (1'h0);
  reg [(3'h6):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1086 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1085 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1083 = (1'h0);
  reg [(4'ha):(1'h0)] reg1082 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1081 = (1'h0);
  reg [(4'h9):(1'h0)] reg1080 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1079 = (1'h0);
  reg [(4'h9):(1'h0)] reg1078 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1077 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1076 = (1'h0);
  reg [(4'hb):(1'h0)] reg1075 = (1'h0);
  reg [(4'hb):(1'h0)] reg1074 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1073 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1072 = (1'h0);
  reg [(4'h8):(1'h0)] reg1071 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1064 = (1'h0);
  reg [(4'h8):(1'h0)] reg1070 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1069 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1068 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1055 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1065 = (1'h0);
  reg [(4'h9):(1'h0)] reg1067 = (1'h0);
  reg [(2'h2):(1'h0)] reg1062 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1060 = (1'h0);
  reg [(2'h2):(1'h0)] reg1066 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1065 = (1'h0);
  reg [(5'h10):(1'h0)] reg1064 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1063 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1062 = (1'h0);
  reg [(4'h9):(1'h0)] reg1061 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1060 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1059 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1058 = (1'h0);
  reg [(3'h4):(1'h0)] reg1057 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1056 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1055 = (1'h0);
  reg [(2'h2):(1'h0)] reg1054 = (1'h0);
  reg [(4'he):(1'h0)] reg1053 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1052 = (1'h0);
  reg [(4'hf):(1'h0)] reg1051 = (1'h0);
  reg [(4'ha):(1'h0)] reg1050 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1049 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1048 = (1'h0);
  reg [(3'h4):(1'h0)] reg1041 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1038 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1036 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1047 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1046 = (1'h0);
  reg [(3'h6):(1'h0)] reg1045 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1044 = (1'h0);
  reg [(5'h10):(1'h0)] reg1043 = (1'h0);
  reg [(4'hf):(1'h0)] reg1042 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1041 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1040 = (1'h0);
  reg [(4'hd):(1'h0)] reg1039 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1038 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1037 = (1'h0);
  reg [(3'h5):(1'h0)] reg1036 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1035 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1034 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1033 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1032 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1031 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1030 = (1'h0);
  reg [(4'he):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1028 = (1'h0);
  reg [(3'h7):(1'h0)] reg1027 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1026 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1025 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1024 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1023 = (1'h0);
  reg [(2'h2):(1'h0)] reg1022 = (1'h0);
  reg [(5'h10):(1'h0)] reg1021 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1020 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1019 = (1'h0);
  reg [(3'h5):(1'h0)] reg1018 = (1'h0);
  reg [(4'hd):(1'h0)] reg1017 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1016 = (1'h0);
  reg [(2'h3):(1'h0)] reg1015 = (1'h0);
  reg [(4'hf):(1'h0)] reg1014 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1013 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1012 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1011 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1010 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1009 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1008 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1007 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1003 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1002 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1006 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1005 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1004 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1003 = (1'h0);
  reg [(4'h9):(1'h0)] reg1002 = (1'h0);
  reg [(4'h9):(1'h0)] reg1001 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1000 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar999 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg998 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg999 = (1'h0);
  reg [(4'he):(1'h0)] forvar998 = (1'h0);
  reg [(4'h8):(1'h0)] forvar997 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg946 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg945 = (1'h0);
  reg [(4'h8):(1'h0)] forvar944 = (1'h0);
  reg [(2'h3):(1'h0)] reg941 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar940 = (1'h0);
  reg [(5'h10):(1'h0)] forvar934 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg992 = (1'h0);
  reg [(5'h10):(1'h0)] forvar985 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg996 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg995 = (1'h0);
  reg [(3'h6):(1'h0)] reg994 = (1'h0);
  reg [(4'hd):(1'h0)] reg993 = (1'h0);
  reg [(3'h6):(1'h0)] forvar992 = (1'h0);
  reg [(4'hf):(1'h0)] reg991 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg990 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar989 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg988 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg987 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg986 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg985 = (1'h0);
  reg [(3'h5):(1'h0)] reg984 = (1'h0);
  reg [(4'ha):(1'h0)] reg983 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg982 = (1'h0);
  reg [(4'he):(1'h0)] reg981 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg980 = (1'h0);
  reg [(5'h10):(1'h0)] reg979 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg978 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar977 = (1'h0);
  reg [(4'he):(1'h0)] reg976 = (1'h0);
  reg [(3'h7):(1'h0)] forvar975 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg974 = (1'h0);
  reg [(4'hf):(1'h0)] reg973 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg972 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar970 = (1'h0);
  reg [(4'hd):(1'h0)] reg971 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg970 = (1'h0);
  reg [(4'hb):(1'h0)] forvar969 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar930 = (1'h0);
  reg [(4'ha):(1'h0)] reg968 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg967 = (1'h0);
  reg [(3'h7):(1'h0)] reg966 = (1'h0);
  reg [(2'h3):(1'h0)] forvar965 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg964 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg963 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg962 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg961 = (1'h0);
  reg [(4'hc):(1'h0)] forvar960 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar959 = (1'h0);
  reg [(5'h10):(1'h0)] reg958 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg957 = (1'h0);
  reg [(3'h6):(1'h0)] reg956 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg955 = (1'h0);
  reg [(5'h10):(1'h0)] reg954 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg953 = (1'h0);
  reg [(4'hb):(1'h0)] reg952 = (1'h0);
  reg [(4'ha):(1'h0)] forvar951 = (1'h0);
  reg [(3'h7):(1'h0)] reg950 = (1'h0);
  reg [(4'h8):(1'h0)] reg949 = (1'h0);
  reg [(4'hb):(1'h0)] reg948 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg947 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar946 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar945 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg944 = (1'h0);
  reg [(4'ha):(1'h0)] reg943 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg942 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar941 = (1'h0);
  reg [(3'h6):(1'h0)] reg940 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar939 = (1'h0);
  reg [(2'h2):(1'h0)] forvar935 = (1'h0);
  reg [(5'h10):(1'h0)] reg933 = (1'h0);
  reg [(4'h9):(1'h0)] reg931 = (1'h0);
  reg [(3'h6):(1'h0)] reg939 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg938 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg937 = (1'h0);
  reg [(5'h10):(1'h0)] reg936 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg935 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg934 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar933 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg932 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar931 = (1'h0);
  reg [(3'h5):(1'h0)] reg930 = (1'h0);
  reg [(4'hd):(1'h0)] reg929 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg928 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg927 = (1'h0);
  reg [(3'h6):(1'h0)] reg926 = (1'h0);
  reg [(3'h4):(1'h0)] reg925 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar921 = (1'h0);
  reg [(4'hd):(1'h0)] forvar916 = (1'h0);
  reg [(3'h6):(1'h0)] reg913 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar911 = (1'h0);
  reg [(4'ha):(1'h0)] forvar908 = (1'h0);
  reg [(4'h9):(1'h0)] forvar904 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg902 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar907 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar903 = (1'h0);
  reg [(4'hc):(1'h0)] reg901 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar899 = (1'h0);
  reg [(5'h10):(1'h0)] forvar889 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg885 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar896 = (1'h0);
  reg [(4'hb):(1'h0)] reg894 = (1'h0);
  reg [(4'hf):(1'h0)] forvar892 = (1'h0);
  reg signed [(4'he):(1'h0)] reg891 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar888 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg887 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg886 = (1'h0);
  reg [(4'ha):(1'h0)] forvar914 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg924 = (1'h0);
  reg [(2'h3):(1'h0)] reg923 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg915 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg922 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg921 = (1'h0);
  reg [(3'h4):(1'h0)] reg920 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg919 = (1'h0);
  reg [(4'he):(1'h0)] reg918 = (1'h0);
  reg [(4'he):(1'h0)] reg917 = (1'h0);
  reg [(4'ha):(1'h0)] reg916 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar915 = (1'h0);
  reg [(5'h10):(1'h0)] reg914 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar913 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg912 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg911 = (1'h0);
  reg signed [(4'he):(1'h0)] reg910 = (1'h0);
  reg [(4'hf):(1'h0)] reg909 = (1'h0);
  reg signed [(4'he):(1'h0)] reg908 = (1'h0);
  reg [(4'ha):(1'h0)] reg907 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg906 = (1'h0);
  reg [(2'h2):(1'h0)] reg905 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg904 = (1'h0);
  reg [(3'h6):(1'h0)] reg903 = (1'h0);
  reg [(2'h2):(1'h0)] forvar902 = (1'h0);
  reg [(4'h9):(1'h0)] forvar901 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg899 = (1'h0);
  reg [(4'he):(1'h0)] reg898 = (1'h0);
  reg [(3'h4):(1'h0)] reg897 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg896 = (1'h0);
  reg [(5'h10):(1'h0)] reg895 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar894 = (1'h0);
  reg [(4'hf):(1'h0)] reg893 = (1'h0);
  reg [(4'h8):(1'h0)] reg892 = (1'h0);
  reg [(2'h2):(1'h0)] forvar891 = (1'h0);
  reg [(4'h8):(1'h0)] reg890 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg889 = (1'h0);
  reg [(3'h5):(1'h0)] reg888 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar887 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar886 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar885 = (1'h0);
  reg [(4'he):(1'h0)] forvar837 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar836 = (1'h0);
  reg [(3'h5):(1'h0)] reg834 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar831 = (1'h0);
  reg [(3'h7):(1'h0)] forvar827 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg826 = (1'h0);
  reg [(4'hb):(1'h0)] forvar825 = (1'h0);
  reg [(2'h3):(1'h0)] reg822 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar820 = (1'h0);
  reg [(4'hb):(1'h0)] forvar818 = (1'h0);
  reg [(3'h5):(1'h0)] reg813 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg807 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar806 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg804 = (1'h0);
  reg [(4'he):(1'h0)] forvar802 = (1'h0);
  reg [(4'h8):(1'h0)] forvar801 = (1'h0);
  reg [(3'h6):(1'h0)] reg800 = (1'h0);
  reg [(3'h7):(1'h0)] forvar799 = (1'h0);
  reg [(4'he):(1'h0)] reg796 = (1'h0);
  reg [(4'h8):(1'h0)] forvar795 = (1'h0);
  reg [(4'h9):(1'h0)] reg794 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar792 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar791 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg884 = (1'h0);
  reg [(3'h5):(1'h0)] forvar883 = (1'h0);
  reg [(2'h2):(1'h0)] reg882 = (1'h0);
  reg [(4'hf):(1'h0)] forvar881 = (1'h0);
  reg [(3'h4):(1'h0)] forvar880 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar879 = (1'h0);
  reg [(4'hb):(1'h0)] forvar868 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg866 = (1'h0);
  reg [(4'hd):(1'h0)] reg878 = (1'h0);
  reg [(4'hc):(1'h0)] reg877 = (1'h0);
  reg [(4'hc):(1'h0)] forvar876 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg875 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar874 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg872 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg874 = (1'h0);
  reg [(3'h4):(1'h0)] reg873 = (1'h0);
  reg [(4'h9):(1'h0)] forvar872 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg871 = (1'h0);
  reg [(4'h8):(1'h0)] reg870 = (1'h0);
  reg [(4'h8):(1'h0)] reg869 = (1'h0);
  reg signed [(4'he):(1'h0)] reg868 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg867 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar866 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg865 = (1'h0);
  reg [(3'h4):(1'h0)] forvar864 = (1'h0);
  reg [(5'h10):(1'h0)] forvar863 = (1'h0);
  reg [(4'hc):(1'h0)] reg862 = (1'h0);
  reg [(4'hb):(1'h0)] reg861 = (1'h0);
  reg [(4'hb):(1'h0)] forvar860 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg859 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg858 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar857 = (1'h0);
  reg [(4'h9):(1'h0)] reg856 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg855 = (1'h0);
  reg [(4'hc):(1'h0)] forvar854 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg853 = (1'h0);
  reg [(3'h6):(1'h0)] reg852 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg851 = (1'h0);
  reg [(4'he):(1'h0)] reg850 = (1'h0);
  reg [(4'hd):(1'h0)] reg849 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg848 = (1'h0);
  reg [(3'h4):(1'h0)] reg847 = (1'h0);
  reg [(3'h4):(1'h0)] reg846 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg845 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg843 = (1'h0);
  reg [(4'hb):(1'h0)] reg842 = (1'h0);
  reg signed [(4'he):(1'h0)] reg841 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg840 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg839 = (1'h0);
  reg [(4'hc):(1'h0)] reg838 = (1'h0);
  reg [(3'h7):(1'h0)] reg837 = (1'h0);
  reg [(4'he):(1'h0)] reg836 = (1'h0);
  reg [(4'he):(1'h0)] reg835 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar834 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg833 = (1'h0);
  reg [(2'h2):(1'h0)] reg832 = (1'h0);
  reg [(3'h4):(1'h0)] reg831 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg830 = (1'h0);
  reg [(3'h6):(1'h0)] reg829 = (1'h0);
  reg [(2'h3):(1'h0)] reg828 = (1'h0);
  reg signed [(4'he):(1'h0)] reg827 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar826 = (1'h0);
  reg [(4'hb):(1'h0)] forvar814 = (1'h0);
  reg [(4'hd):(1'h0)] reg825 = (1'h0);
  reg [(3'h6):(1'h0)] reg824 = (1'h0);
  reg signed [(4'he):(1'h0)] reg823 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar822 = (1'h0);
  reg [(4'hd):(1'h0)] reg821 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg820 = (1'h0);
  reg [(4'hf):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg818 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg817 = (1'h0);
  reg [(3'h7):(1'h0)] reg816 = (1'h0);
  reg [(4'hb):(1'h0)] reg815 = (1'h0);
  reg [(2'h2):(1'h0)] reg814 = (1'h0);
  reg [(4'h8):(1'h0)] forvar813 = (1'h0);
  reg [(3'h6):(1'h0)] reg812 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar811 = (1'h0);
  reg [(4'ha):(1'h0)] reg810 = (1'h0);
  reg signed [(4'he):(1'h0)] reg809 = (1'h0);
  reg [(4'hb):(1'h0)] reg808 = (1'h0);
  reg [(4'hd):(1'h0)] forvar807 = (1'h0);
  reg [(4'h8):(1'h0)] reg806 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg805 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar804 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg803 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg802 = (1'h0);
  reg [(4'hb):(1'h0)] reg801 = (1'h0);
  reg [(4'he):(1'h0)] forvar800 = (1'h0);
  reg [(3'h4):(1'h0)] reg799 = (1'h0);
  reg [(2'h3):(1'h0)] reg798 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg797 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar796 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg795 = (1'h0);
  reg [(5'h10):(1'h0)] forvar794 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg793 = (1'h0);
  reg signed [(4'he):(1'h0)] reg792 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg791 = (1'h0);
  reg signed [(4'he):(1'h0)] reg790 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg789 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg788 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar787 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar786 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar785 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire783;
  wire signed [(4'h8):(1'h0)] wire599;
  wire [(3'h5):(1'h0)] wire598;
  wire [(5'h10):(1'h0)] wire597;
  assign y = {wire1144,
                 wire1143,
                 wire1142,
                 reg1130,
                 forvar1128,
                 forvar1126,
                 forvar1121,
                 reg1119,
                 reg1114,
                 forvar1111,
                 reg1141,
                 reg1140,
                 forvar1139,
                 reg1138,
                 reg1137,
                 reg1136,
                 forvar1135,
                 reg1134,
                 reg1133,
                 reg1132,
                 reg1131,
                 forvar1130,
                 reg1129,
                 reg1128,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1123,
                 reg1122,
                 reg1121,
                 reg1120,
                 forvar1119,
                 reg1118,
                 reg1117,
                 reg1116,
                 reg1115,
                 forvar1114,
                 reg1108,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1110,
                 reg1109,
                 forvar1108,
                 forvar1107,
                 forvar1087,
                 forvar1081,
                 reg1083,
                 forvar1082,
                 forvar1079,
                 reg1072,
                 reg1093,
                 reg1106,
                 reg1105,
                 reg1104,
                 forvar1103,
                 reg1102,
                 reg1101,
                 reg1100,
                 reg1099,
                 forvar1098,
                 reg1097,
                 reg1096,
                 reg1095,
                 reg1094,
                 forvar1093,
                 reg1092,
                 reg1091,
                 reg1090,
                 reg1089,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 reg1084,
                 forvar1083,
                 reg1082,
                 reg1081,
                 reg1080,
                 reg1079,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1075,
                 reg1074,
                 reg1073,
                 forvar1072,
                 reg1071,
                 forvar1064,
                 reg1070,
                 reg1069,
                 reg1068,
                 reg1055,
                 forvar1065,
                 reg1067,
                 reg1062,
                 forvar1060,
                 reg1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 forvar1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1057,
                 forvar1056,
                 forvar1055,
                 reg1054,
                 reg1053,
                 reg1052,
                 reg1051,
                 reg1050,
                 forvar1049,
                 forvar1048,
                 reg1041,
                 reg1038,
                 forvar1036,
                 reg1047,
                 reg1046,
                 reg1045,
                 forvar1044,
                 reg1043,
                 reg1042,
                 forvar1041,
                 reg1040,
                 reg1039,
                 forvar1038,
                 forvar1037,
                 reg1036,
                 reg1035,
                 forvar1034,
                 reg1033,
                 reg1032,
                 forvar1031,
                 reg1030,
                 reg1029,
                 reg1028,
                 reg1027,
                 forvar1026,
                 forvar1025,
                 forvar1024,
                 forvar1023,
                 reg1022,
                 reg1021,
                 reg1020,
                 reg1019,
                 reg1018,
                 reg1017,
                 forvar1016,
                 reg1015,
                 reg1014,
                 reg1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1008,
                 forvar1007,
                 reg1003,
                 forvar1002,
                 reg1006,
                 reg1005,
                 reg1004,
                 forvar1003,
                 reg1002,
                 reg1001,
                 reg1000,
                 forvar999,
                 reg998,
                 reg999,
                 forvar998,
                 forvar997,
                 reg946,
                 reg945,
                 forvar944,
                 reg941,
                 forvar940,
                 forvar934,
                 reg992,
                 forvar985,
                 reg996,
                 reg995,
                 reg994,
                 reg993,
                 forvar992,
                 reg991,
                 reg990,
                 forvar989,
                 reg988,
                 reg987,
                 reg986,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg981,
                 reg980,
                 reg979,
                 reg978,
                 forvar977,
                 reg976,
                 forvar975,
                 reg974,
                 reg973,
                 reg972,
                 forvar970,
                 reg971,
                 reg970,
                 forvar969,
                 forvar930,
                 reg968,
                 reg967,
                 reg966,
                 forvar965,
                 reg964,
                 reg963,
                 reg962,
                 reg961,
                 forvar960,
                 forvar959,
                 reg958,
                 reg957,
                 reg956,
                 reg955,
                 reg954,
                 reg953,
                 reg952,
                 forvar951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 forvar946,
                 forvar945,
                 reg944,
                 reg943,
                 reg942,
                 forvar941,
                 reg940,
                 forvar939,
                 forvar935,
                 reg933,
                 reg931,
                 reg939,
                 reg938,
                 reg937,
                 reg936,
                 reg935,
                 reg934,
                 forvar933,
                 reg932,
                 forvar931,
                 reg930,
                 reg929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 forvar921,
                 forvar916,
                 reg913,
                 forvar911,
                 forvar908,
                 forvar904,
                 reg902,
                 forvar907,
                 forvar903,
                 reg901,
                 forvar899,
                 forvar889,
                 reg885,
                 forvar896,
                 reg894,
                 forvar892,
                 reg891,
                 forvar888,
                 reg887,
                 reg886,
                 forvar914,
                 reg924,
                 reg923,
                 reg915,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 forvar915,
                 reg914,
                 forvar913,
                 reg912,
                 reg911,
                 reg910,
                 reg909,
                 reg908,
                 reg907,
                 reg906,
                 reg905,
                 reg904,
                 reg903,
                 forvar902,
                 forvar901,
                 reg900,
                 reg899,
                 reg898,
                 reg897,
                 reg896,
                 reg895,
                 forvar894,
                 reg893,
                 reg892,
                 forvar891,
                 reg890,
                 reg889,
                 reg888,
                 forvar887,
                 forvar886,
                 forvar885,
                 forvar837,
                 forvar836,
                 reg834,
                 forvar831,
                 forvar827,
                 reg826,
                 forvar825,
                 reg822,
                 forvar820,
                 forvar818,
                 reg813,
                 reg807,
                 forvar806,
                 reg804,
                 forvar802,
                 forvar801,
                 reg800,
                 forvar799,
                 reg796,
                 forvar795,
                 reg794,
                 forvar792,
                 forvar791,
                 reg884,
                 forvar883,
                 reg882,
                 forvar881,
                 forvar880,
                 forvar879,
                 forvar868,
                 reg866,
                 reg878,
                 reg877,
                 forvar876,
                 reg875,
                 forvar874,
                 reg872,
                 reg874,
                 reg873,
                 forvar872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 reg867,
                 forvar866,
                 reg865,
                 forvar864,
                 forvar863,
                 reg862,
                 reg861,
                 forvar860,
                 reg859,
                 reg858,
                 forvar857,
                 reg856,
                 reg855,
                 forvar854,
                 reg853,
                 reg852,
                 reg851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 reg845,
                 reg844,
                 reg843,
                 reg842,
                 reg841,
                 reg840,
                 reg839,
                 reg838,
                 reg837,
                 reg836,
                 reg835,
                 forvar834,
                 reg833,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 reg827,
                 forvar826,
                 forvar814,
                 reg825,
                 reg824,
                 reg823,
                 forvar822,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 forvar813,
                 reg812,
                 forvar811,
                 reg810,
                 reg809,
                 reg808,
                 forvar807,
                 reg806,
                 reg805,
                 forvar804,
                 reg803,
                 reg802,
                 reg801,
                 forvar800,
                 reg799,
                 reg798,
                 reg797,
                 forvar796,
                 reg795,
                 forvar794,
                 reg793,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 reg788,
                 forvar787,
                 forvar786,
                 forvar785,
                 wire783,
                 wire599,
                 wire598,
                 wire597,
                 (1'h0)};
  assign wire597 = (($unsigned({wire595}) ?
                           $unsigned($signed(wire594)) : wire595[(1'h1):(1'h1)]) ?
                       wire594[(4'hb):(4'hb)] : (^$unsigned((+wire595))));
  assign wire598 = (($unsigned($signed(wire592)) ^~ {(wire595 || wire594)}) ?
                       wire593[(3'h4):(2'h2)] : wire592);
  assign wire599 = ($signed($signed(wire593[(2'h3):(2'h3)])) || (($unsigned(wire595) ?
                       $unsigned(wire595) : (&(8'hab))) ^~ {wire594[(4'hb):(3'h5)]}));
  module600 modinst784 (.wire603(wire595), .wire601(wire599), .wire602(wire597), .y(wire783), .clk(clk), .wire604(wire592));
  always
    @(posedge clk) begin
      if ((((^~(wire595 && (8'ha6))) ? wire593 : wire592) ?
          $unsigned(($unsigned(wire597) ~^ (wire593 ~^ wire598))) : ($unsigned($unsigned(wire598)) ?
              ($unsigned(wire599) ?
                  (wire593 | wire598) : $signed(wire595)) : $unsigned((wire597 >> wire597)))))
        begin
          for (forvar785 = (1'h0); (forvar785 < (2'h3)); forvar785 = (forvar785 + (1'h1)))
            begin
              for (forvar786 = (1'h0); (forvar786 < (2'h2)); forvar786 = (forvar786 + (1'h1)))
                begin
                  for (forvar787 = (1'h0); (forvar787 < (1'h1)); forvar787 = (forvar787 + (1'h1)))
                    begin
                      reg788 <= ((wire598 ?
                          (~|(wire592 <<< (8'hb7))) : wire597[(3'h5):(1'h1)]) ^ ({(wire593 != wire593)} != $unsigned(wire597)));
                      reg789 <= {wire595};
                      reg790 <= $unsigned(wire599);
                    end
                  if ((^$signed(wire783[(1'h0):(1'h0)])))
                    begin
                      reg791 <= wire597[(3'h7):(1'h0)];
                      reg792 <= wire599[(3'h7):(3'h5)];
                      reg793 <= (((wire594[(1'h1):(1'h0)] > wire596[(4'h9):(1'h0)]) ?
                          (+wire598) : $unsigned((~&(8'hac)))) | reg791);
                    end
                  else
                    begin
                      reg791 <= $unsigned(({((8'ha2) | forvar787)} ?
                          ($unsigned(wire592) ?
                              reg792 : ((8'ha4) ?
                                  wire592 : forvar785)) : $unsigned(reg790[(4'h8):(3'h5)])));
                      reg792 <= reg792[(1'h0):(1'h0)];
                    end
                  for (forvar794 = (1'h0); (forvar794 < (1'h1)); forvar794 = (forvar794 + (1'h1)))
                    begin
                      reg795 <= $unsigned(reg789[(2'h2):(1'h1)]);
                    end
                end
              for (forvar796 = (1'h0); (forvar796 < (1'h1)); forvar796 = (forvar796 + (1'h1)))
                begin
                  if (wire599[(3'h4):(3'h4)])
                    begin
                      reg797 <= ((reg795[(3'h7):(3'h4)] && wire599) & (~&$signed((wire595 * forvar796))));
                      reg798 <= (-{(~{wire783})});
                      reg799 <= reg789;
                    end
                  else
                    begin
                      reg797 <= (({$signed(reg791)} ?
                              $unsigned((reg789 ?
                                  wire599 : reg792)) : $signed($unsigned((8'hac)))) ?
                          (reg792 ?
                              wire593[(1'h1):(1'h1)] : ((reg793 ^~ wire597) >> (~|reg789))) : (^forvar785));
                      reg798 <= wire596[(4'h9):(4'h9)];
                      reg799 <= (|wire597);
                    end
                  for (forvar800 = (1'h0); (forvar800 < (2'h2)); forvar800 = (forvar800 + (1'h1)))
                    begin
                      reg801 <= ((8'hba) == (wire597 ?
                          (|{(8'hb2)}) : reg795[(2'h2):(1'h1)]));
                      reg802 <= (-(((|reg797) - reg790) ?
                          $signed((forvar787 ?
                              forvar794 : reg797)) : (&(^reg789))));
                      reg803 <= ((wire593 <= $unsigned(reg790)) != $signed(((+reg801) - forvar794)));
                    end
                  for (forvar804 = (1'h0); (forvar804 < (1'h1)); forvar804 = (forvar804 + (1'h1)))
                    begin
                      reg805 <= $unsigned((~&wire594[(1'h1):(1'h0)]));
                      reg806 <= (^(^($unsigned(forvar800) >= (~&wire596))));
                    end
                end
              for (forvar807 = (1'h0); (forvar807 < (1'h0)); forvar807 = (forvar807 + (1'h1)))
                begin
                  reg808 <= wire596;
                  if ($signed((((&wire597) ?
                          (wire598 ? wire599 : wire594) : {reg792}) ?
                      wire596[(4'h9):(1'h1)] : $signed(wire597))))
                    begin
                      reg809 <= wire594[(1'h0):(1'h0)];
                      reg810 <= (^~(8'ha1));
                    end
                  else
                    begin
                      reg809 <= (~&(+{{forvar800}}));
                      reg810 <= (wire598[(3'h5):(3'h5)] && (reg788 || $signed(wire592[(3'h4):(2'h2)])));
                    end
                  for (forvar811 = (1'h0); (forvar811 < (2'h2)); forvar811 = (forvar811 + (1'h1)))
                    begin
                      reg812 <= (^~forvar786);
                    end
                end
            end
          for (forvar813 = (1'h0); (forvar813 < (1'h0)); forvar813 = (forvar813 + (1'h1)))
            begin
              if ((~^$unsigned((8'h9c))))
                begin
                  if (reg812[(1'h1):(1'h0)])
                    begin
                      reg814 <= $signed((($unsigned(reg798) ?
                          forvar794 : (forvar796 ?
                              forvar796 : forvar811)) & ((^~reg791) != $signed((8'h9e)))));
                    end
                  else
                    begin
                      reg814 <= forvar811;
                      reg815 <= forvar786;
                      reg816 <= $signed((reg795[(3'h6):(3'h6)] != ((|reg814) << {reg802})));
                      reg817 <= reg812[(3'h5):(3'h4)];
                    end
                  if (reg810[(4'h8):(3'h5)])
                    begin
                      reg818 <= {(8'hb9)};
                    end
                  else
                    begin
                      reg818 <= reg797;
                      reg819 <= $unsigned(((reg810 ?
                          wire783[(1'h1):(1'h1)] : {reg798}) ~^ $signed({reg795})));
                      reg820 <= reg799;
                    end
                  reg821 <= ((reg788[(4'h8):(3'h7)] >> {{wire594}}) ?
                      reg801[(1'h1):(1'h1)] : $unsigned(wire783));
                  for (forvar822 = (1'h0); (forvar822 < (2'h2)); forvar822 = (forvar822 + (1'h1)))
                    begin
                      reg823 <= $signed((&$unsigned((reg792 ^~ (8'hb3)))));
                      reg824 <= $unsigned($unsigned($unsigned($signed((8'hb8)))));
                      reg825 <= $signed(($unsigned(reg820[(2'h2):(2'h2)]) >> (~&$signed((8'h9f)))));
                    end
                end
              else
                begin
                  for (forvar814 = (1'h0); (forvar814 < (1'h0)); forvar814 = (forvar814 + (1'h1)))
                    begin
                      reg815 <= (!wire599);
                      reg816 <= $signed(wire596);
                      reg817 <= reg814[(1'h0):(1'h0)];
                      reg818 <= $unsigned((-$unsigned(reg802)));
                    end
                  reg819 <= $unsigned(forvar800);
                end
              for (forvar826 = (1'h0); (forvar826 < (2'h2)); forvar826 = (forvar826 + (1'h1)))
                begin
                  if (((~&reg792[(3'h4):(3'h4)]) ?
                      ($signed($signed(forvar796)) ?
                          reg803 : forvar822) : (wire596[(1'h1):(1'h1)] ?
                          ($unsigned(reg803) ?
                              reg814[(1'h1):(1'h0)] : (reg805 - forvar813)) : $signed($signed(reg799)))))
                    begin
                      reg827 <= forvar796[(3'h5):(2'h3)];
                      reg828 <= forvar794;
                      reg829 <= (+$signed(((reg808 + wire595) ?
                          reg815[(1'h1):(1'h0)] : $unsigned(forvar826))));
                    end
                  else
                    begin
                      reg827 <= (({(reg820 == reg824)} ?
                          ($signed(forvar796) * (-reg810)) : (&forvar794[(4'hf):(2'h3)])) && forvar787);
                    end
                  if (({(|$unsigned((8'ha5)))} ?
                      $unsigned(wire596) : ($unsigned(reg808[(1'h1):(1'h0)]) ?
                          reg788[(3'h7):(1'h0)] : forvar796)))
                    begin
                      reg830 <= (~^((~forvar804) ?
                          wire597[(1'h0):(1'h0)] : forvar796));
                      reg831 <= (wire593[(2'h3):(2'h3)] >= ({reg827[(2'h3):(2'h2)]} ?
                          ({wire599} ?
                              $signed(wire594) : (^~reg803)) : $unsigned($signed(reg814))));
                      reg832 <= reg821[(3'h7):(2'h3)];
                      reg833 <= {reg788};
                    end
                  else
                    begin
                      reg830 <= ((!$unsigned($unsigned((8'hb2)))) ^~ reg829);
                    end
                  for (forvar834 = (1'h0); (forvar834 < (1'h1)); forvar834 = (forvar834 + (1'h1)))
                    begin
                      reg835 <= ($signed((!$unsigned(reg793))) >= ($signed((^(8'hb6))) && $unsigned((reg806 ?
                          reg820 : wire598))));
                      reg836 <= $unsigned((reg802[(1'h1):(1'h0)] ?
                          (8'hac) : (~&(forvar834 ? (8'ha7) : reg809))));
                      reg837 <= reg824[(1'h0):(1'h0)];
                      reg838 <= (reg790[(2'h2):(1'h1)] ?
                          $signed($signed(reg808)) : reg791);
                    end
                  if ($signed({reg830[(2'h3):(2'h3)]}))
                    begin
                      reg839 <= $unsigned({(+(~|wire599))});
                      reg840 <= ((forvar800[(4'ha):(2'h3)] ?
                          (8'hb0) : {reg832[(1'h0):(1'h0)]}) + $unsigned($unsigned((reg805 == forvar822))));
                      reg841 <= ($unsigned($signed($unsigned(reg820))) | (+{(wire593 - (8'hb9))}));
                    end
                  else
                    begin
                      reg839 <= $signed(reg814);
                    end
                end
              if ($unsigned((|(forvar813[(1'h0):(1'h0)] >> (~reg839)))))
                begin
                  reg842 <= $signed($signed((reg797[(1'h0):(1'h0)] ?
                      (^reg803) : reg814[(1'h1):(1'h1)])));
                end
              else
                begin
                  if ($signed({($signed((8'ha6)) ?
                          forvar786[(3'h4):(3'h4)] : $unsigned(wire597))}))
                    begin
                      reg842 <= forvar811;
                      reg843 <= $signed((~^(~$signed(reg809))));
                      reg844 <= (reg802 ?
                          {(^~(forvar804 ?
                                  (8'hac) : reg806))} : reg809[(4'he):(2'h2)]);
                      reg845 <= reg829;
                    end
                  else
                    begin
                      reg842 <= (((~|(-reg789)) ?
                              ((~^reg830) ?
                                  (reg788 * (8'ha1)) : reg798[(2'h3):(1'h1)]) : ((reg797 >>> reg830) <<< forvar826)) ?
                          {(!{(8'ha9)})} : (($signed(reg842) ?
                                  ((8'ha6) ?
                                      (8'ha7) : reg795) : (~|forvar811)) ?
                              $signed((^forvar814)) : $signed(forvar811[(3'h5):(1'h1)])));
                      reg843 <= $signed((8'h9d));
                      reg844 <= reg820;
                    end
                  if ($unsigned($signed((reg819[(3'h4):(1'h0)] << forvar813))))
                    begin
                      reg846 <= {((~^(forvar813 < (8'ha6))) ?
                              $unsigned($unsigned(reg836)) : (^~((8'haa) ?
                                  reg802 : forvar822)))};
                    end
                  else
                    begin
                      reg846 <= reg841[(4'h9):(2'h3)];
                      reg847 <= (((~|forvar814[(2'h2):(1'h1)]) || reg795[(1'h0):(1'h0)]) ?
                          {$unsigned($signed(reg832))} : reg802[(1'h0):(1'h0)]);
                      reg848 <= ((|$signed((-reg802))) >> ((8'hae) + (forvar804[(2'h2):(2'h2)] ?
                          (&reg827) : reg827[(4'h8):(1'h1)])));
                      reg849 <= {(!reg839[(1'h1):(1'h1)])};
                    end
                  if ((wire597 ?
                      ($unsigned((forvar811 ?
                          reg842 : (8'hba))) ^~ reg789[(3'h4):(1'h0)]) : (reg806[(2'h3):(1'h0)] ?
                          (~&forvar834) : (reg829[(3'h6):(2'h3)] ?
                              wire598 : (wire593 == forvar794)))))
                    begin
                      reg850 <= $signed(((!forvar813) || reg795));
                      reg851 <= (wire783 <= $signed($unsigned($unsigned((8'hb9)))));
                      reg852 <= wire598;
                      reg853 <= $unsigned((($unsigned(reg812) ?
                              (&reg837) : (reg849 ~^ reg820)) ?
                          (~|(^reg820)) : {(reg793 >= forvar811)}));
                    end
                  else
                    begin
                      reg850 <= ((forvar796 ? forvar800 : forvar807) ?
                          forvar826 : $signed(reg844));
                    end
                end
              for (forvar854 = (1'h0); (forvar854 < (2'h2)); forvar854 = (forvar854 + (1'h1)))
                begin
                  if ((({(&wire783)} >> $signed($signed(reg842))) ?
                      reg790 : reg828[(2'h3):(1'h0)]))
                    begin
                      reg855 <= wire594;
                      reg856 <= ((reg814 - ($unsigned(reg832) != ((8'ha8) + reg827))) ?
                          (reg851 ^~ reg805[(1'h1):(1'h0)]) : (reg846 ^~ forvar796[(3'h6):(3'h6)]));
                    end
                  else
                    begin
                      reg855 <= {$unsigned($unsigned(((8'hb2) ?
                              wire592 : reg820)))};
                    end
                  for (forvar857 = (1'h0); (forvar857 < (1'h0)); forvar857 = (forvar857 + (1'h1)))
                    begin
                      reg858 <= (|$signed((~&$signed(reg846))));
                    end
                  reg859 <= $signed(($signed($unsigned(reg810)) + ((~^reg853) - reg792)));
                  for (forvar860 = (1'h0); (forvar860 < (2'h2)); forvar860 = (forvar860 + (1'h1)))
                    begin
                      reg861 <= ({((^~wire592) & (!reg845))} ?
                          reg815 : ({(^~forvar811)} ?
                              ({reg827} == (+reg821)) : reg850[(4'h9):(2'h3)]));
                      reg862 <= (~^($signed(reg846) ?
                          wire594[(4'hb):(2'h3)] : (8'hb4)));
                    end
                end
            end
          if (((^(+(~^forvar813))) ?
              $signed(forvar826) : {$signed((forvar796 ^~ forvar796))}))
            begin
              for (forvar863 = (1'h0); (forvar863 < (2'h3)); forvar863 = (forvar863 + (1'h1)))
                begin
                  for (forvar864 = (1'h0); (forvar864 < (1'h0)); forvar864 = (forvar864 + (1'h1)))
                    begin
                      reg865 <= (reg851[(2'h2):(1'h1)] ^~ reg853[(3'h7):(2'h3)]);
                    end
                  for (forvar866 = (1'h0); (forvar866 < (2'h3)); forvar866 = (forvar866 + (1'h1)))
                    begin
                      reg867 <= ((~^(((8'ha8) ? reg845 : (8'hb7)) * (8'hb6))) ?
                          (&reg835) : (!({(8'ha6)} || forvar814)));
                      reg868 <= $signed((reg853 ?
                          $signed((reg803 >>> reg808)) : reg818));
                      reg869 <= ({$unsigned(forvar813)} << (-$unsigned($signed(reg815))));
                      reg870 <= reg848;
                    end
                end
              if ((forvar826 + (+{reg819[(2'h3):(2'h2)]})))
                begin
                  reg871 <= ($unsigned($unsigned((forvar863 != reg839))) ?
                      $unsigned($signed($signed(reg859))) : reg815[(3'h5):(1'h1)]);
                  for (forvar872 = (1'h0); (forvar872 < (2'h3)); forvar872 = (forvar872 + (1'h1)))
                    begin
                      reg873 <= reg815[(2'h2):(2'h2)];
                    end
                  reg874 <= reg829;
                end
              else
                begin
                  if (($signed((~&reg816)) ^~ $signed((reg844[(3'h4):(1'h1)] ?
                      $signed(reg799) : forvar822[(4'hb):(4'h8)]))))
                    begin
                      reg871 <= reg795[(4'h8):(2'h3)];
                      reg872 <= reg874[(1'h1):(1'h1)];
                      reg873 <= (!((reg792[(4'h8):(3'h7)] ?
                              (&forvar800) : (reg795 ? reg798 : forvar794)) ?
                          $signed((8'ha0)) : (!wire595[(4'h9):(4'h9)])));
                    end
                  else
                    begin
                      reg871 <= reg827;
                      reg872 <= ((8'ha7) >= $unsigned($unsigned((~|reg791))));
                    end
                  for (forvar874 = (1'h0); (forvar874 < (1'h0)); forvar874 = (forvar874 + (1'h1)))
                    begin
                      reg875 <= $unsigned($signed((~&(|reg852))));
                    end
                end
              for (forvar876 = (1'h0); (forvar876 < (2'h2)); forvar876 = (forvar876 + (1'h1)))
                begin
                  if (({reg836[(4'hb):(4'h8)]} ?
                      ((reg868[(3'h4):(1'h0)] ?
                          reg840 : $signed((8'ha1))) * ((^wire595) ?
                          $unsigned(reg798) : {reg808})) : {($unsigned((8'hb9)) >> ((8'ha5) | reg825))}))
                    begin
                      reg877 <= $unsigned(({$signed(reg832)} ?
                          $signed(wire597[(4'hb):(4'hb)]) : ($unsigned((8'ha8)) << (&reg828))));
                      reg878 <= ((~|((&forvar787) ?
                              ((8'hb8) ?
                                  reg855 : forvar785) : reg842[(3'h6):(2'h3)])) ?
                          $unsigned($unsigned((reg842 * reg835))) : {(8'hb5)});
                    end
                  else
                    begin
                      reg877 <= {$signed((8'hb6))};
                    end
                end
            end
          else
            begin
              for (forvar863 = (1'h0); (forvar863 < (1'h0)); forvar863 = (forvar863 + (1'h1)))
                begin
                  for (forvar864 = (1'h0); (forvar864 < (2'h2)); forvar864 = (forvar864 + (1'h1)))
                    begin
                      reg865 <= $signed((8'haf));
                      reg866 <= (reg821 ?
                          $signed(forvar863[(2'h3):(1'h0)]) : $unsigned(reg848));
                      reg867 <= (!((((8'hb9) ^ reg870) ?
                              forvar786 : $signed(forvar874)) ?
                          (+$signed(reg792)) : (^~(forvar872 || (8'ha6)))));
                    end
                  for (forvar868 = (1'h0); (forvar868 < (2'h3)); forvar868 = (forvar868 + (1'h1)))
                    begin
                      reg869 <= reg842;
                      reg870 <= reg846[(3'h4):(3'h4)];
                      reg871 <= ((reg865 ^ (8'h9e)) & ((|{reg840}) ?
                          forvar876 : reg852[(3'h5):(2'h2)]));
                    end
                  reg872 <= $signed($unsigned(({reg824} ?
                      ((8'hb8) ? reg799 : reg873) : forvar813)));
                  reg873 <= (reg812[(3'h6):(2'h2)] - (8'had));
                end
            end
          for (forvar879 = (1'h0); (forvar879 < (2'h2)); forvar879 = (forvar879 + (1'h1)))
            begin
              for (forvar880 = (1'h0); (forvar880 < (1'h1)); forvar880 = (forvar880 + (1'h1)))
                begin
                  for (forvar881 = (1'h0); (forvar881 < (2'h2)); forvar881 = (forvar881 + (1'h1)))
                    begin
                      reg882 <= (&(forvar804 < $signed($unsigned(reg847))));
                    end
                  for (forvar883 = (1'h0); (forvar883 < (2'h3)); forvar883 = (forvar883 + (1'h1)))
                    begin
                      reg884 <= {(reg836 ? forvar883 : (!wire599))};
                    end
                end
            end
        end
      else
        begin
          for (forvar785 = (1'h0); (forvar785 < (2'h3)); forvar785 = (forvar785 + (1'h1)))
            begin
              for (forvar786 = (1'h0); (forvar786 < (2'h2)); forvar786 = (forvar786 + (1'h1)))
                begin
                  for (forvar787 = (1'h0); (forvar787 < (2'h3)); forvar787 = (forvar787 + (1'h1)))
                    begin
                      reg788 <= {reg797};
                      reg789 <= reg846[(2'h3):(1'h0)];
                      reg790 <= (~wire596);
                    end
                end
              for (forvar791 = (1'h0); (forvar791 < (1'h1)); forvar791 = (forvar791 + (1'h1)))
                begin
                  for (forvar792 = (1'h0); (forvar792 < (2'h2)); forvar792 = (forvar792 + (1'h1)))
                    begin
                      reg793 <= $signed(reg790);
                      reg794 <= $unsigned((reg846[(2'h3):(1'h1)] - (|reg830[(1'h0):(1'h0)])));
                    end
                  for (forvar795 = (1'h0); (forvar795 < (1'h1)); forvar795 = (forvar795 + (1'h1)))
                    begin
                      reg796 <= (~&$signed((reg871 | (forvar864 ?
                          (8'hac) : reg869))));
                      reg797 <= (-$signed(forvar813[(1'h0):(1'h0)]));
                      reg798 <= (~^(~($signed(reg839) > reg844[(3'h5):(2'h2)])));
                    end
                  for (forvar799 = (1'h0); (forvar799 < (2'h3)); forvar799 = (forvar799 + (1'h1)))
                    begin
                      reg800 <= forvar868;
                    end
                end
            end
          if (reg877[(1'h0):(1'h0)])
            begin
              for (forvar801 = (1'h0); (forvar801 < (2'h3)); forvar801 = (forvar801 + (1'h1)))
                begin
                  for (forvar802 = (1'h0); (forvar802 < (2'h3)); forvar802 = (forvar802 + (1'h1)))
                    begin
                      reg803 <= reg831[(2'h3):(2'h2)];
                      reg804 <= $unsigned($unsigned((~|$signed((8'hae)))));
                    end
                  reg805 <= ((-((reg841 ? forvar872 : forvar794) ?
                      $unsigned(reg823) : $unsigned(reg825))) ^ $signed(forvar879));
                  for (forvar806 = (1'h0); (forvar806 < (1'h1)); forvar806 = (forvar806 + (1'h1)))
                    begin
                      reg807 <= reg844;
                      reg808 <= $signed((-($unsigned(reg796) ?
                          $signed(reg850) : reg871[(2'h2):(2'h2)])));
                      reg809 <= {(~$unsigned((reg853 ? (8'ha6) : forvar864)))};
                      reg810 <= (forvar826 ^~ reg817);
                    end
                  for (forvar811 = (1'h0); (forvar811 < (2'h3)); forvar811 = (forvar811 + (1'h1)))
                    begin
                      reg812 <= $unsigned($signed(forvar876[(3'h7):(2'h3)]));
                      reg813 <= forvar807[(3'h7):(3'h7)];
                    end
                end
              for (forvar814 = (1'h0); (forvar814 < (1'h0)); forvar814 = (forvar814 + (1'h1)))
                begin
                  if ((reg805 | $signed(((&forvar864) == (reg873 ?
                      reg804 : reg865)))))
                    begin
                      reg815 <= {{$unsigned((forvar864 - forvar866))}};
                      reg816 <= $unsigned(forvar881);
                      reg817 <= $signed((^{reg858}));
                    end
                  else
                    begin
                      reg815 <= (($unsigned((-(8'ha9))) ?
                              (reg804[(1'h1):(1'h1)] ?
                                  (8'hab) : $signed((8'hae))) : wire597) ?
                          forvar786[(3'h4):(2'h2)] : $signed({reg808}));
                      reg816 <= $signed((reg851[(2'h2):(1'h0)] ?
                          (8'hb6) : forvar857[(2'h2):(1'h0)]));
                      reg817 <= reg882;
                    end
                  for (forvar818 = (1'h0); (forvar818 < (2'h3)); forvar818 = (forvar818 + (1'h1)))
                    begin
                      reg819 <= (~&(^~{reg882}));
                    end
                  for (forvar820 = (1'h0); (forvar820 < (1'h0)); forvar820 = (forvar820 + (1'h1)))
                    begin
                      reg821 <= ($signed(($signed(reg856) ^~ reg839[(1'h0):(1'h0)])) ?
                          forvar785[(1'h1):(1'h0)] : forvar799);
                      reg822 <= (^{(~&(reg866 ~^ reg866))});
                      reg823 <= ($signed(((forvar883 ? (8'ha5) : forvar881) ?
                              reg843[(4'hf):(3'h7)] : forvar826)) ?
                          forvar822[(4'ha):(1'h1)] : $signed($unsigned(reg840[(2'h3):(1'h0)])));
                      reg824 <= $signed(reg815[(4'h9):(1'h1)]);
                    end
                end
            end
          else
            begin
              for (forvar801 = (1'h0); (forvar801 < (1'h0)); forvar801 = (forvar801 + (1'h1)))
                begin
                  for (forvar802 = (1'h0); (forvar802 < (2'h3)); forvar802 = (forvar802 + (1'h1)))
                    begin
                      reg803 <= (($signed((~^reg792)) ?
                          reg809[(4'hc):(3'h7)] : (^$signed(reg859))) != ($unsigned($unsigned(reg839)) >= reg821));
                    end
                  for (forvar804 = (1'h0); (forvar804 < (2'h3)); forvar804 = (forvar804 + (1'h1)))
                    begin
                      reg805 <= $unsigned(reg835);
                      reg806 <= (forvar795 != (&forvar806));
                    end
                end
            end
          for (forvar825 = (1'h0); (forvar825 < (1'h1)); forvar825 = (forvar825 + (1'h1)))
            begin
              reg826 <= (&(^(~|$signed(forvar796))));
              if (((~{{forvar822}}) ?
                  $unsigned($signed(reg841)) : (reg867 ?
                      $unsigned((&forvar866)) : $signed(reg810))))
                begin
                  for (forvar827 = (1'h0); (forvar827 < (1'h1)); forvar827 = (forvar827 + (1'h1)))
                    begin
                      reg828 <= $unsigned($unsigned(((reg810 ?
                          (8'h9e) : reg828) ^~ reg839)));
                      reg829 <= forvar792[(3'h7):(3'h4)];
                      reg830 <= forvar883[(3'h5):(1'h0)];
                    end
                  for (forvar831 = (1'h0); (forvar831 < (1'h1)); forvar831 = (forvar831 + (1'h1)))
                    begin
                      reg832 <= wire593[(1'h0):(1'h0)];
                      reg833 <= wire593;
                      reg834 <= $signed($unsigned($unsigned(((8'hac) ?
                          reg815 : reg848))));
                      reg835 <= $unsigned((forvar831 ?
                          ((wire595 ~^ (8'ha2)) + $signed(reg867)) : $signed((reg861 >= (8'ha6)))));
                    end
                end
              else
                begin
                  reg827 <= $signed($signed(reg798));
                  if ({$unsigned($unsigned({forvar814}))})
                    begin
                      reg828 <= $unsigned($unsigned(((reg844 ?
                              forvar820 : reg819) ?
                          (reg819 ? reg798 : reg872) : $signed(reg858))));
                      reg829 <= ({($unsigned((8'hb1)) ?
                                  $signed(wire592) : reg827)} ?
                          {{(forvar831 <<< reg799)}} : $signed($unsigned(forvar831[(4'ha):(2'h2)])));
                    end
                  else
                    begin
                      reg828 <= forvar834[(3'h7):(2'h3)];
                      reg829 <= ($signed((((8'hb5) ? reg841 : wire597) ?
                              (reg841 & reg795) : (wire596 <<< reg804))) ?
                          reg789 : $signed(reg812));
                    end
                end
            end
          for (forvar836 = (1'h0); (forvar836 < (2'h2)); forvar836 = (forvar836 + (1'h1)))
            begin
              if ($signed(forvar881[(1'h1):(1'h0)]))
                begin
                  reg837 <= (^($unsigned(reg806[(1'h1):(1'h1)]) > forvar868[(3'h7):(2'h2)]));
                  reg838 <= {$signed(({(8'hb4)} ?
                          $unsigned(reg818) : {reg882}))};
                end
              else
                begin
                  for (forvar837 = (1'h0); (forvar837 < (1'h0)); forvar837 = (forvar837 + (1'h1)))
                    begin
                      reg838 <= $unsigned($signed(((forvar792 ?
                              reg867 : forvar866) ?
                          reg812[(3'h5):(3'h5)] : $signed((8'hba)))));
                      reg839 <= reg869;
                      reg840 <= $unsigned(($signed($signed(wire596)) > reg796));
                      reg841 <= ({(^~(forvar806 ? forvar827 : reg848))} ?
                          $unsigned(reg856) : reg804);
                    end
                end
            end
        end
      if ($unsigned((+forvar864)))
        begin
          for (forvar885 = (1'h0); (forvar885 < (2'h3)); forvar885 = (forvar885 + (1'h1)))
            begin
              for (forvar886 = (1'h0); (forvar886 < (1'h1)); forvar886 = (forvar886 + (1'h1)))
                begin
                  for (forvar887 = (1'h0); (forvar887 < (1'h0)); forvar887 = (forvar887 + (1'h1)))
                    begin
                      reg888 <= reg875[(2'h2):(1'h0)];
                      reg889 <= reg873[(1'h0):(1'h0)];
                      reg890 <= ((-$unsigned(forvar814)) ?
                          wire598[(1'h0):(1'h0)] : reg826[(3'h4):(3'h4)]);
                    end
                  for (forvar891 = (1'h0); (forvar891 < (1'h1)); forvar891 = (forvar891 + (1'h1)))
                    begin
                      reg892 <= {($unsigned((forvar879 ? reg851 : reg828)) ?
                              forvar794 : {(forvar836 ? (8'ha5) : reg794)})};
                    end
                  reg893 <= $unsigned($unsigned(((forvar806 * (8'ha0)) << (~|forvar857))));
                end
              if (reg791[(3'h6):(2'h2)])
                begin
                  for (forvar894 = (1'h0); (forvar894 < (2'h3)); forvar894 = (forvar894 + (1'h1)))
                    begin
                      reg895 <= $unsigned($unsigned((reg812[(1'h1):(1'h0)] ?
                          (wire593 <<< reg790) : $signed(reg838))));
                      reg896 <= ((-(forvar883 ?
                          forvar795 : (wire783 <= reg874))) == forvar799[(2'h3):(1'h0)]);
                    end
                  reg897 <= (((~(reg890 && reg888)) ?
                      ((8'hb2) <<< reg865) : $unsigned((reg870 ?
                          wire595 : reg851))) ^~ $signed(forvar891[(1'h1):(1'h0)]));
                end
              else
                begin
                  for (forvar894 = (1'h0); (forvar894 < (2'h3)); forvar894 = (forvar894 + (1'h1)))
                    begin
                      reg895 <= (forvar801 ?
                          (forvar887[(1'h0):(1'h0)] ?
                              $signed((8'ha9)) : (+reg797)) : (~|$signed((reg798 ?
                              reg801 : reg801))));
                      reg896 <= $signed((~&((reg789 && reg796) <= ((8'ha1) ?
                          reg812 : (8'ha5)))));
                      reg897 <= {$signed(({reg893} ~^ reg844))};
                    end
                  if ((8'hb8))
                    begin
                      reg898 <= ($signed((!$unsigned(reg809))) ?
                          (&reg835[(1'h1):(1'h0)]) : {$unsigned((forvar887 ?
                                  (8'ha7) : (8'hb7)))});
                      reg899 <= (^~($unsigned($signed(reg867)) >>> ($unsigned((8'haa)) | (reg796 ?
                          (8'hae) : forvar872))));
                    end
                  else
                    begin
                      reg898 <= (reg809[(2'h2):(2'h2)] ?
                          $signed((+reg893)) : ((8'ha7) ?
                              ((forvar854 ? reg874 : reg827) ?
                                  (reg888 ? reg843 : reg831) : (reg795 ?
                                      reg819 : (8'hb5))) : reg833[(3'h6):(1'h0)]));
                      reg899 <= wire593;
                      reg900 <= (($unsigned((wire592 == forvar792)) ^~ $unsigned($signed(forvar799))) | $signed(forvar820));
                    end
                end
              for (forvar901 = (1'h0); (forvar901 < (1'h0)); forvar901 = (forvar901 + (1'h1)))
                begin
                  for (forvar902 = (1'h0); (forvar902 < (1'h1)); forvar902 = (forvar902 + (1'h1)))
                    begin
                      reg903 <= $unsigned($signed((8'h9f)));
                      reg904 <= reg836[(2'h2):(1'h1)];
                      reg905 <= reg789;
                      reg906 <= (8'ha4);
                    end
                  if ($unsigned(wire592))
                    begin
                      reg907 <= (8'hb3);
                    end
                  else
                    begin
                      reg907 <= (forvar834[(4'h9):(1'h0)] ?
                          (+($signed(wire598) ^~ reg853[(4'h9):(3'h4)])) : $signed(($signed(forvar786) ?
                              (!reg812) : $unsigned(forvar831))));
                      reg908 <= $unsigned($unsigned(reg906[(3'h7):(3'h7)]));
                      reg909 <= $unsigned($unsigned(forvar872[(2'h3):(1'h1)]));
                      reg910 <= $unsigned(({forvar874} ?
                          $signed({forvar864}) : $signed($signed(reg815))));
                    end
                end
              reg911 <= forvar881[(4'h9):(3'h4)];
            end
          reg912 <= $signed(reg870);
          if (($signed($signed((reg833 + reg868))) ?
              (($signed(forvar881) ?
                      ((8'ha4) > reg823) : (reg798 ? (8'h9d) : reg796)) ?
                  (reg895 & (+reg821)) : reg818[(4'hd):(3'h5)]) : (!(!$unsigned(reg802)))))
            begin
              if ((~|(^$signed(reg823))))
                begin
                  for (forvar913 = (1'h0); (forvar913 < (1'h1)); forvar913 = (forvar913 + (1'h1)))
                    begin
                      reg914 <= (reg850[(4'ha):(3'h6)] && (~^$unsigned(reg849)));
                    end
                  for (forvar915 = (1'h0); (forvar915 < (1'h1)); forvar915 = (forvar915 + (1'h1)))
                    begin
                      reg916 <= (^reg853[(4'hc):(3'h6)]);
                      reg917 <= {$unsigned(((wire598 - forvar836) > (~^reg888)))};
                      reg918 <= ($unsigned((~&{(8'hae)})) <<< $unsigned(((~&reg791) ?
                          (~forvar786) : (reg878 * (8'hab)))));
                      reg919 <= (^~(forvar880 == ((&forvar792) ?
                          $signed((8'hb8)) : {reg793})));
                    end
                  if (reg890[(2'h2):(2'h2)])
                    begin
                      reg920 <= $unsigned((!((reg851 >> forvar800) >> reg897)));
                      reg921 <= (({$signed(reg910)} ?
                              (((8'hab) ? reg918 : forvar887) & (forvar887 ?
                                  reg844 : (8'hba))) : (forvar800 < $unsigned(forvar786))) ?
                          (-{(|reg877)}) : $unsigned(((forvar864 ^~ reg847) ?
                              (~reg844) : reg793)));
                      reg922 <= reg799[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg920 <= $signed((~|(^~(&reg873))));
                      reg921 <= forvar826;
                      reg922 <= (-{$signed((forvar799 ? reg877 : (8'h9c)))});
                    end
                end
              else
                begin
                  for (forvar913 = (1'h0); (forvar913 < (1'h0)); forvar913 = (forvar913 + (1'h1)))
                    begin
                      reg914 <= $signed((!(~&(reg820 < forvar854))));
                      reg915 <= ((reg838[(4'h8):(2'h3)] | $signed($signed(reg874))) ?
                          $unsigned(($unsigned(forvar825) && $unsigned(reg803))) : ((reg800 & forvar820) ?
                              $signed((forvar880 ^~ forvar806)) : ((&forvar887) ^ $unsigned((8'had)))));
                    end
                end
              reg923 <= $unsigned({$signed(((8'ha2) == (8'had)))});
              reg924 <= (reg851 ^ $signed((((8'ha0) ? reg809 : reg899) ?
                  forvar826 : (reg845 ? forvar818 : reg911))));
            end
          else
            begin
              for (forvar913 = (1'h0); (forvar913 < (1'h0)); forvar913 = (forvar913 + (1'h1)))
                begin
                  for (forvar914 = (1'h0); (forvar914 < (1'h1)); forvar914 = (forvar914 + (1'h1)))
                    begin
                      reg915 <= $signed(reg866[(4'h8):(1'h1)]);
                      reg916 <= $signed($signed((~|((8'hb0) * reg815))));
                      reg917 <= $signed(forvar881);
                      reg918 <= (forvar836 ? (~reg908) : (~|$signed(reg803)));
                    end
                  reg919 <= {(reg840[(4'h9):(3'h7)] ?
                          $signed($unsigned(reg813)) : {(forvar879 || reg908)})};
                end
            end
        end
      else
        begin
          if ((^(((reg832 ? forvar887 : reg918) ?
                  (reg841 ? forvar837 : reg893) : (8'ha4)) ?
              (-(!forvar807)) : forvar914)))
            begin
              for (forvar885 = (1'h0); (forvar885 < (2'h2)); forvar885 = (forvar885 + (1'h1)))
                begin
                  reg886 <= $signed(((~&reg824[(2'h3):(2'h3)]) ~^ reg888[(1'h0):(1'h0)]));
                end
              if ((|(8'hab)))
                begin
                  reg887 <= $signed($signed((^~(&forvar883))));
                  for (forvar888 = (1'h0); (forvar888 < (1'h0)); forvar888 = (forvar888 + (1'h1)))
                    begin
                      reg889 <= ((~|((wire783 ?
                              reg803 : (8'hab)) != $signed((8'ha6)))) ?
                          forvar834 : $signed($unsigned({forvar802})));
                      reg890 <= forvar914[(4'h8):(2'h2)];
                      reg891 <= {reg912[(1'h1):(1'h1)]};
                    end
                  for (forvar892 = (1'h0); (forvar892 < (1'h0)); forvar892 = (forvar892 + (1'h1)))
                    begin
                      reg893 <= {(~^((+reg847) ?
                              reg796 : ((8'hb1) ? reg874 : forvar874)))};
                      reg894 <= (|($signed({forvar857}) & $unsigned(reg790[(3'h5):(1'h1)])));
                    end
                end
              else
                begin
                  if ($unsigned(({$signed((8'hb9))} ^~ forvar827)))
                    begin
                      reg887 <= reg850;
                    end
                  else
                    begin
                      reg887 <= {{(forvar872 + $unsigned(reg791))}};
                      reg888 <= $signed((-wire783[(2'h2):(1'h1)]));
                      reg889 <= {$unsigned(($signed(forvar796) < (forvar887 | forvar818)))};
                      reg890 <= $signed($unsigned(((+(8'hb3)) >> reg814[(1'h0):(1'h0)])));
                    end
                  for (forvar891 = (1'h0); (forvar891 < (2'h2)); forvar891 = (forvar891 + (1'h1)))
                    begin
                      reg892 <= ((reg910 != ((reg915 && reg827) ?
                          {reg900} : {reg850})) ~^ (^~($signed((8'h9e)) ?
                          (8'ha1) : (forvar795 ? forvar880 : (8'ha0)))));
                    end
                  if ({(^~reg903[(3'h5):(2'h3)])})
                    begin
                      reg893 <= $signed($unsigned(reg836));
                      reg894 <= (~($unsigned((|reg830)) ?
                          ((forvar796 > (8'hb0)) ^ $unsigned(reg893)) : (reg835[(1'h1):(1'h1)] | (reg868 == reg849))));
                      reg895 <= reg812;
                    end
                  else
                    begin
                      reg893 <= reg903[(3'h6):(3'h6)];
                      reg894 <= ($signed((+forvar902)) << {(-(&reg882))});
                      reg895 <= {$signed({forvar820})};
                    end
                  for (forvar896 = (1'h0); (forvar896 < (2'h2)); forvar896 = (forvar896 + (1'h1)))
                    begin
                      reg897 <= reg900;
                      reg898 <= reg873;
                    end
                end
              reg899 <= $signed(reg804[(2'h2):(2'h2)]);
              reg900 <= $signed((8'h9e));
            end
          else
            begin
              reg885 <= (&(($unsigned(forvar863) ?
                  (forvar787 ?
                      reg856 : (8'ha1)) : (8'hac)) ~^ $signed((~&reg873))));
              if ((|forvar820))
                begin
                  reg886 <= {(8'h9c)};
                  if (wire596)
                    begin
                      reg887 <= $signed(forvar792);
                    end
                  else
                    begin
                      reg887 <= (^~(forvar876 ?
                          reg829 : (forvar795[(3'h5):(2'h2)] ?
                              $unsigned(reg795) : (|reg919))));
                      reg888 <= (^reg887[(1'h1):(1'h1)]);
                      reg889 <= forvar888;
                      reg890 <= (~|($unsigned((reg906 ? reg912 : (8'hb1))) ?
                          reg917 : ($signed(reg819) ?
                              (8'haf) : (forvar837 ? (8'hb1) : reg912))));
                    end
                  reg891 <= (^~(reg817[(2'h3):(1'h1)] ^ reg809));
                  for (forvar892 = (1'h0); (forvar892 < (1'h0)); forvar892 = (forvar892 + (1'h1)))
                    begin
                      reg893 <= ($signed($unsigned(((8'ha2) ^ wire593))) ?
                          forvar801[(3'h7):(1'h1)] : {{forvar885[(3'h4):(2'h3)]}});
                      reg894 <= (reg850[(3'h4):(2'h3)] <<< $unsigned((reg834[(2'h3):(2'h3)] ?
                          wire592 : reg798[(2'h2):(1'h1)])));
                      reg895 <= ((~|(~&$signed((8'hb2)))) || ({{reg812}} >= reg789));
                    end
                end
              else
                begin
                  for (forvar886 = (1'h0); (forvar886 < (1'h1)); forvar886 = (forvar886 + (1'h1)))
                    begin
                      reg887 <= reg835[(2'h3):(2'h2)];
                      reg888 <= (reg865 - forvar872[(4'h8):(3'h4)]);
                    end
                  for (forvar889 = (1'h0); (forvar889 < (1'h1)); forvar889 = (forvar889 + (1'h1)))
                    begin
                      reg890 <= (|$signed((reg827[(4'hc):(2'h2)] ?
                          (reg829 ?
                              forvar785 : reg861) : reg820[(4'he):(3'h4)])));
                      reg891 <= $unsigned(wire598[(2'h2):(2'h2)]);
                      reg892 <= {(forvar881 ?
                              reg812 : ({forvar787} && $signed(forvar785)))};
                      reg893 <= $unsigned((&forvar837));
                    end
                  for (forvar894 = (1'h0); (forvar894 < (2'h3)); forvar894 = (forvar894 + (1'h1)))
                    begin
                      reg895 <= (+$signed(reg829));
                      reg896 <= $signed(reg861[(2'h2):(1'h0)]);
                      reg897 <= $unsigned(($signed(forvar801) ?
                          $unsigned($unsigned((8'hab))) : ((forvar864 ?
                              reg830 : forvar864) != (reg831 == reg819))));
                      reg898 <= (((~(forvar915 ? wire598 : reg911)) <= reg800) ?
                          reg794 : $signed({(reg832 == reg845)}));
                    end
                  for (forvar899 = (1'h0); (forvar899 < (2'h2)); forvar899 = (forvar899 + (1'h1)))
                    begin
                      reg900 <= $unsigned(forvar795[(3'h5):(2'h3)]);
                      reg901 <= (&(reg866 ? reg891 : reg921));
                    end
                end
            end
          if ({((reg801[(3'h4):(1'h0)] ? reg813 : {reg844}) ?
                  {$unsigned(reg834)} : reg841[(2'h3):(1'h1)])})
            begin
              for (forvar902 = (1'h0); (forvar902 < (2'h3)); forvar902 = (forvar902 + (1'h1)))
                begin
                  for (forvar903 = (1'h0); (forvar903 < (1'h1)); forvar903 = (forvar903 + (1'h1)))
                    begin
                      reg904 <= (+$unsigned(reg915));
                      reg905 <= reg843;
                      reg906 <= forvar822[(3'h6):(2'h2)];
                    end
                  for (forvar907 = (1'h0); (forvar907 < (1'h1)); forvar907 = (forvar907 + (1'h1)))
                    begin
                      reg908 <= reg816[(3'h5):(2'h3)];
                    end
                  reg909 <= reg868;
                  if ((forvar800[(4'ha):(1'h1)] ^~ (reg799 ~^ (|$signed(forvar857)))))
                    begin
                      reg910 <= reg856;
                      reg911 <= forvar885[(2'h2):(1'h0)];
                      reg912 <= {(((forvar799 ?
                                  reg869 : (8'hb9)) ^ ((8'h9c) >> reg865)) ?
                              {reg845} : $signed($unsigned(reg822)))};
                    end
                  else
                    begin
                      reg910 <= {$unsigned({$unsigned(reg924)})};
                      reg911 <= (reg867[(3'h7):(3'h6)] ?
                          (-((~&(8'ha6)) ~^ {reg866})) : (reg874[(4'h8):(2'h3)] * reg831[(1'h1):(1'h1)]));
                      reg912 <= $signed({$unsigned((reg871 ?
                              (8'ha2) : forvar806))});
                    end
                end
              for (forvar913 = (1'h0); (forvar913 < (2'h3)); forvar913 = (forvar913 + (1'h1)))
                begin
                  for (forvar914 = (1'h0); (forvar914 < (1'h1)); forvar914 = (forvar914 + (1'h1)))
                    begin
                      reg915 <= (8'hb8);
                      reg916 <= ($signed(reg882) ?
                          $signed(forvar894) : {forvar807});
                      reg917 <= {(forvar902 ?
                              reg797 : $signed($signed(reg911)))};
                      reg918 <= (~^forvar881[(3'h7):(3'h5)]);
                    end
                  if (($unsigned($unsigned($unsigned(reg801))) <<< $unsigned($unsigned(forvar802[(4'hc):(4'h9)]))))
                    begin
                      reg919 <= forvar801[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg919 <= {(reg803 <<< ({reg806} ?
                              $signed(reg837) : $unsigned((8'hb6))))};
                    end
                  reg920 <= (8'h9c);
                end
              reg921 <= $signed(((!reg872) ?
                  ($signed(reg909) ?
                      $signed(reg795) : $unsigned(reg847)) : (reg799[(2'h2):(2'h2)] == reg914[(4'he):(2'h3)])));
            end
          else
            begin
              reg902 <= (~&(reg899 ?
                  ((~&reg873) ?
                      ((8'ha4) ?
                          (8'haf) : reg859) : $unsigned(forvar902)) : ($signed(forvar868) << (reg886 ?
                      (8'hb5) : reg789))));
              for (forvar903 = (1'h0); (forvar903 < (1'h0)); forvar903 = (forvar903 + (1'h1)))
                begin
                  for (forvar904 = (1'h0); (forvar904 < (1'h0)); forvar904 = (forvar904 + (1'h1)))
                    begin
                      reg905 <= forvar863;
                    end
                  if ({((forvar804 < $signed(reg790)) ?
                          $signed((reg871 ?
                              (8'ha9) : wire593)) : forvar795[(3'h6):(3'h6)])})
                    begin
                      reg906 <= (({$signed(forvar818)} <<< $signed(forvar826)) ~^ reg852[(3'h4):(1'h0)]);
                      reg907 <= ($signed(forvar913) ?
                          (reg907[(3'h6):(1'h0)] ?
                              $signed((+reg835)) : $unsigned($unsigned(forvar787))) : ({$unsigned(forvar836)} | reg915));
                    end
                  else
                    begin
                      reg906 <= $signed(reg852[(3'h5):(1'h0)]);
                      reg907 <= ($signed($signed($signed(forvar901))) ?
                          reg895[(3'h7):(2'h2)] : reg820);
                    end
                  for (forvar908 = (1'h0); (forvar908 < (2'h3)); forvar908 = (forvar908 + (1'h1)))
                    begin
                      reg909 <= ($unsigned($unsigned(reg845[(3'h7):(3'h7)])) >= (~&$signed(reg878[(4'hb):(4'ha)])));
                      reg910 <= (^reg902[(2'h2):(2'h2)]);
                    end
                end
              if ($unsigned($signed($signed((8'hab)))))
                begin
                  for (forvar911 = (1'h0); (forvar911 < (1'h1)); forvar911 = (forvar911 + (1'h1)))
                    begin
                      reg912 <= $unsigned((forvar903[(1'h1):(1'h0)] ?
                          {(reg904 ^~ reg841)} : {$unsigned(reg830)}));
                      reg913 <= reg793[(1'h0):(1'h0)];
                      reg914 <= $unsigned($unsigned(reg842[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  if ($signed({((reg838 ?
                          reg888 : reg815) - (reg866 >= forvar831))}))
                    begin
                      reg911 <= forvar881;
                      reg912 <= reg919;
                      reg913 <= (8'hab);
                    end
                  else
                    begin
                      reg911 <= (forvar913[(1'h1):(1'h1)] ?
                          (forvar792 <= reg849[(4'hd):(3'h4)]) : (reg856[(4'h8):(3'h4)] <= (reg873[(1'h1):(1'h0)] ?
                              $signed((8'hb3)) : (forvar908 < reg922))));
                      reg912 <= (-$signed(forvar891));
                    end
                end
              for (forvar915 = (1'h0); (forvar915 < (2'h2)); forvar915 = (forvar915 + (1'h1)))
                begin
                  for (forvar916 = (1'h0); (forvar916 < (1'h1)); forvar916 = (forvar916 + (1'h1)))
                    begin
                      reg917 <= $signed(((~(8'hab)) << reg872));
                      reg918 <= {$unsigned((~|(forvar887 ?
                              forvar894 : (8'ha6))))};
                      reg919 <= ($unsigned($signed(reg893[(1'h1):(1'h0)])) == reg865[(1'h1):(1'h1)]);
                      reg920 <= $signed((^reg885));
                    end
                  for (forvar921 = (1'h0); (forvar921 < (1'h1)); forvar921 = (forvar921 + (1'h1)))
                    begin
                      reg922 <= $signed($signed($signed($signed(forvar791))));
                      reg923 <= ($signed(($unsigned(reg923) ?
                          ((8'ha1) >>> reg836) : (forvar801 >>> forvar802))) || {(reg807[(1'h1):(1'h0)] ?
                              (8'hab) : (forvar795 * forvar907))});
                    end
                  if (($signed(forvar822) - reg793[(2'h2):(1'h1)]))
                    begin
                      reg924 <= (^$signed(reg817[(4'h8):(2'h2)]));
                      reg925 <= $unsigned($signed(($signed(reg835) <<< $unsigned((8'ha9)))));
                    end
                  else
                    begin
                      reg924 <= reg873;
                      reg925 <= forvar807[(2'h2):(1'h1)];
                      reg926 <= (|reg827[(4'ha):(3'h6)]);
                    end
                  if ((($signed(((8'h9e) | reg829)) ?
                          ((reg790 ? reg924 : forvar907) ?
                              {reg805} : (^~forvar860)) : {(!forvar866)}) ?
                      $unsigned($signed($signed((8'hac)))) : forvar896[(2'h2):(1'h0)]))
                    begin
                      reg927 <= $signed($signed(((reg798 >> wire596) == (!(8'ha1)))));
                      reg928 <= (!(~|(8'hba)));
                    end
                  else
                    begin
                      reg927 <= ({forvar802[(2'h2):(1'h0)]} != $signed((~|(forvar814 * forvar907))));
                      reg928 <= (&$unsigned((reg891 ?
                          (reg888 ? reg867 : reg882) : reg902)));
                      reg929 <= reg911;
                    end
                end
            end
        end
      if (forvar792)
        begin
          if ($unsigned({{{reg829}}}))
            begin
              reg930 <= ((forvar863[(4'he):(2'h3)] ?
                  ({reg817} ?
                      $unsigned(forvar894) : (reg871 ?
                          wire595 : reg850)) : (~$signed(reg910))) || (((wire597 ?
                          reg805 : reg825) ?
                      (reg804 ? forvar864 : reg912) : $unsigned((8'h9f))) ?
                  reg796[(3'h5):(2'h3)] : $unsigned(reg869)));
              if (($signed((forvar886 ~^ $signed((8'hb1)))) ^~ $unsigned(reg824)))
                begin
                  for (forvar931 = (1'h0); (forvar931 < (1'h0)); forvar931 = (forvar931 + (1'h1)))
                    begin
                      reg932 <= reg884[(1'h1):(1'h1)];
                    end
                  for (forvar933 = (1'h0); (forvar933 < (2'h2)); forvar933 = (forvar933 + (1'h1)))
                    begin
                      reg934 <= ($unsigned((forvar785 ?
                          (reg835 ? reg816 : reg821) : (reg821 ?
                              reg858 : (8'ha1)))) << ($unsigned(reg797[(1'h0):(1'h0)]) ?
                          {$unsigned(reg800)} : $signed({forvar872})));
                      reg935 <= {$signed(reg790[(1'h1):(1'h0)])};
                    end
                  if (reg798)
                    begin
                      reg936 <= $signed(($signed($unsigned(wire783)) ?
                          ((reg810 == reg912) ?
                              (^~reg897) : (^~reg894)) : (reg894 < $signed(reg920))));
                      reg937 <= $signed($unsigned($unsigned($unsigned(reg884))));
                      reg938 <= $signed($unsigned(((forvar787 << (8'hb4)) <= (forvar885 ?
                          wire783 : reg925))));
                      reg939 <= (reg845 < (reg805[(1'h1):(1'h1)] & $signed(forvar826[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg936 <= forvar904;
                      reg937 <= ($unsigned(forvar795) > (-($unsigned((8'hb9)) >= $signed(reg918))));
                      reg938 <= $unsigned(($signed(((8'ha1) <<< reg878)) > {reg888[(2'h3):(2'h3)]}));
                      reg939 <= {forvar894[(3'h5):(1'h0)]};
                    end
                end
              else
                begin
                  if ((!$signed((!reg789[(1'h1):(1'h1)]))))
                    begin
                      reg931 <= reg923;
                      reg932 <= $unsigned((8'h9c));
                      reg933 <= $unsigned($signed($unsigned(reg832[(1'h1):(1'h1)])));
                      reg934 <= ((-(+(reg877 >= reg809))) << ($signed(reg917) ?
                          (-(-forvar894)) : (((8'hac) * reg853) ?
                              $unsigned(reg839) : (reg827 != reg907))));
                    end
                  else
                    begin
                      reg931 <= $signed(($signed(reg902) <= $signed($unsigned(reg819))));
                      reg932 <= $signed(((+$unsigned(reg833)) == {(forvar864 <= reg795)}));
                      reg933 <= (+(8'ha5));
                    end
                  for (forvar935 = (1'h0); (forvar935 < (1'h0)); forvar935 = (forvar935 + (1'h1)))
                    begin
                      reg936 <= $unsigned(reg809[(3'h5):(2'h3)]);
                      reg937 <= ((((reg793 ? forvar911 : reg826) ?
                              ((8'ha3) == reg922) : (~&reg917)) ?
                          {(&reg833)} : (reg888 ?
                              {reg805} : $signed(reg848))) << $signed((^(+(8'hac)))));
                      reg938 <= ($unsigned($unsigned((|reg902))) ?
                          (((^forvar786) ?
                              {reg825} : $signed(reg837)) - (forvar794[(4'he):(4'h8)] != reg797[(1'h0):(1'h0)])) : (~(-$signed(reg861))));
                    end
                  for (forvar939 = (1'h0); (forvar939 < (2'h3)); forvar939 = (forvar939 + (1'h1)))
                    begin
                      reg940 <= {(((~&forvar916) ?
                              $unsigned(reg923) : forvar911[(3'h4):(2'h3)]) - ((forvar935 <= reg910) ?
                              reg930[(1'h0):(1'h0)] : (+(8'ha6))))};
                    end
                  for (forvar941 = (1'h0); (forvar941 < (1'h0)); forvar941 = (forvar941 + (1'h1)))
                    begin
                      reg942 <= {{$signed(reg830[(2'h3):(1'h0)])}};
                      reg943 <= $unsigned(($signed($unsigned(forvar854)) >>> {$signed(reg925)}));
                      reg944 <= (reg890 ?
                          $unsigned((~&reg858[(3'h5):(3'h5)])) : (({reg831} ?
                              (+forvar921) : reg882[(1'h1):(1'h0)]) ~^ (+$signed(reg790))));
                    end
                end
              for (forvar945 = (1'h0); (forvar945 < (2'h3)); forvar945 = (forvar945 + (1'h1)))
                begin
                  for (forvar946 = (1'h0); (forvar946 < (1'h1)); forvar946 = (forvar946 + (1'h1)))
                    begin
                      reg947 <= ({(8'hac)} != $unsigned(reg802[(2'h3):(2'h2)]));
                      reg948 <= (reg894[(2'h3):(1'h1)] ?
                          $unsigned(((!reg882) ?
                              (reg872 << reg884) : ((8'hb8) ?
                                  forvar911 : (8'hb4)))) : $unsigned(reg913[(3'h5):(2'h2)]));
                      reg949 <= $signed(forvar796);
                      reg950 <= reg795[(3'h6):(1'h0)];
                    end
                  for (forvar951 = (1'h0); (forvar951 < (1'h0)); forvar951 = (forvar951 + (1'h1)))
                    begin
                      reg952 <= wire783;
                      reg953 <= (~^($signed(reg926[(3'h5):(2'h3)]) < $unsigned((reg821 - forvar802))));
                      reg954 <= $unsigned((8'hab));
                      reg955 <= {(8'hb8)};
                    end
                  if ({reg849[(4'h9):(2'h2)]})
                    begin
                      reg956 <= reg833;
                      reg957 <= reg852;
                    end
                  else
                    begin
                      reg956 <= reg931[(1'h1):(1'h0)];
                    end
                  reg958 <= $unsigned({forvar907[(3'h5):(2'h2)]});
                end
              for (forvar959 = (1'h0); (forvar959 < (2'h3)); forvar959 = (forvar959 + (1'h1)))
                begin
                  for (forvar960 = (1'h0); (forvar960 < (2'h2)); forvar960 = (forvar960 + (1'h1)))
                    begin
                      reg961 <= (8'hb7);
                      reg962 <= reg929;
                      reg963 <= {reg861[(4'hb):(3'h6)]};
                      reg964 <= ($signed((reg834[(2'h2):(1'h1)] ?
                              reg830[(3'h7):(3'h6)] : {forvar811})) ?
                          {forvar864} : (^$signed((&reg849))));
                    end
                  for (forvar965 = (1'h0); (forvar965 < (2'h3)); forvar965 = (forvar965 + (1'h1)))
                    begin
                      reg966 <= forvar915;
                      reg967 <= (((8'h9d) & reg892) == $unsigned(reg886));
                    end
                  reg968 <= (!($signed(forvar807) * ({reg842} ?
                      (reg796 ? reg922 : forvar939) : $signed(forvar941))));
                end
            end
          else
            begin
              for (forvar930 = (1'h0); (forvar930 < (2'h3)); forvar930 = (forvar930 + (1'h1)))
                begin
                  if (((!$unsigned(reg947)) ?
                      ((^~$signed(forvar864)) >= ((reg823 << reg855) ?
                          (reg850 > reg829) : (8'h9d))) : reg916))
                    begin
                      reg931 <= (($unsigned((+forvar827)) ^~ $unsigned(reg805[(3'h4):(2'h2)])) ?
                          reg803 : (reg907 | forvar916[(3'h6):(3'h4)]));
                      reg932 <= $unsigned((({reg917} ?
                              (reg832 ?
                                  forvar801 : reg875) : $unsigned(reg884)) ?
                          $signed(forvar887[(3'h5):(1'h0)]) : ((8'ha0) ^~ $signed(forvar791))));
                      reg933 <= {(reg809[(3'h5):(2'h2)] ?
                              ($signed(reg851) ?
                                  ((8'hb4) ?
                                      (8'had) : reg890) : forvar800) : reg805[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg931 <= reg835;
                      reg932 <= $signed(($signed(reg858) ?
                          (~^(reg831 ?
                              reg871 : forvar814)) : reg815[(3'h4):(3'h4)]));
                    end
                end
            end
          for (forvar969 = (1'h0); (forvar969 < (2'h2)); forvar969 = (forvar969 + (1'h1)))
            begin
              if (wire595[(3'h7):(3'h5)])
                begin
                  reg970 <= (reg874[(3'h6):(3'h6)] ?
                      $signed($signed(((8'ha4) >>> forvar837))) : reg821[(4'hd):(3'h6)]);
                  reg971 <= reg802[(1'h1):(1'h1)];
                end
              else
                begin
                  for (forvar970 = (1'h0); (forvar970 < (1'h1)); forvar970 = (forvar970 + (1'h1)))
                    begin
                      reg971 <= (($unsigned(reg901) ?
                          forvar901[(3'h7):(2'h2)] : (8'ha3)) - reg939);
                    end
                  if ((((~^((8'hb0) < reg858)) ?
                          reg915[(3'h5):(3'h4)] : reg897[(3'h4):(3'h4)]) ?
                      $signed($signed((&forvar868))) : ($signed((reg934 ?
                          reg889 : reg906)) ^ ((reg861 ? (8'h9c) : reg967) ?
                          ((8'hb4) ? forvar820 : reg920) : (+forvar914)))))
                    begin
                      reg972 <= reg820;
                      reg973 <= reg821[(2'h2):(2'h2)];
                      reg974 <= ($unsigned(forvar913[(3'h4):(3'h4)]) ?
                          $unsigned($signed($unsigned(reg810))) : {reg866});
                    end
                  else
                    begin
                      reg972 <= $unsigned({((forvar894 ?
                              forvar811 : reg807) < (reg974 ?
                              forvar960 : reg961))});
                      reg973 <= (|forvar904);
                      reg974 <= ((($unsigned(forvar935) ?
                          (reg837 & forvar914) : {forvar874}) ^ $unsigned((8'ha0))) < ((~^$unsigned(reg806)) & $signed(reg884[(2'h2):(1'h1)])));
                    end
                  for (forvar975 = (1'h0); (forvar975 < (1'h1)); forvar975 = (forvar975 + (1'h1)))
                    begin
                      reg976 <= forvar921[(3'h6):(3'h4)];
                    end
                end
            end
          for (forvar977 = (1'h0); (forvar977 < (2'h2)); forvar977 = (forvar977 + (1'h1)))
            begin
              reg978 <= (!(|$signed(forvar896[(3'h5):(1'h0)])));
              if ((($signed($unsigned(reg833)) ?
                  (-$unsigned(reg958)) : reg915) >> $unsigned(reg833)))
                begin
                  reg979 <= forvar863;
                  if ({reg888})
                    begin
                      reg980 <= $signed(((^~reg845[(1'h0):(1'h0)]) == (~|$signed(reg797))));
                      reg981 <= $unsigned(reg942[(3'h4):(1'h1)]);
                      reg982 <= (~&(^~forvar965));
                      reg983 <= (~$signed(reg943[(3'h4):(1'h0)]));
                    end
                  else
                    begin
                      reg980 <= reg940;
                    end
                  reg984 <= ($signed(forvar887) ?
                      (($signed(reg862) ?
                          (forvar866 >> reg866) : reg943[(4'ha):(1'h1)]) + reg833[(3'h7):(1'h1)]) : {$unsigned(((8'hb9) ?
                              reg943 : reg809))});
                end
              else
                begin
                  if ($unsigned($unsigned(reg798[(2'h3):(2'h2)])))
                    begin
                      reg979 <= (($signed((8'ha6)) ?
                              $signed((reg944 ?
                                  (8'hab) : reg915)) : ($unsigned(forvar787) ?
                                  (forvar894 > wire783) : (forvar911 | reg823))) ?
                          $unsigned(forvar941[(2'h2):(2'h2)]) : $signed($unsigned({forvar785})));
                    end
                  else
                    begin
                      reg979 <= $signed((reg928 ? forvar876 : reg976));
                      reg980 <= $unsigned((({reg823} ?
                          reg912 : (reg828 ^ reg903)) >> reg897));
                    end
                  if ((^$unsigned(reg819[(2'h3):(2'h3)])))
                    begin
                      reg981 <= $unsigned($signed(((reg982 ?
                          forvar813 : forvar806) <<< $signed(reg902))));
                      reg982 <= $signed($signed(({reg924} - $signed(reg906))));
                      reg983 <= reg798[(1'h0):(1'h0)];
                      reg984 <= forvar876[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg981 <= $unsigned({$signed((reg830 != reg842))});
                      reg982 <= $signed((-reg819));
                      reg983 <= reg927;
                    end
                end
              if (forvar886[(4'h8):(2'h3)])
                begin
                  if ((8'ha9))
                    begin
                      reg985 <= reg922;
                      reg986 <= {$unsigned({(8'ha6)})};
                      reg987 <= $unsigned(reg986);
                      reg988 <= $unsigned($signed(forvar883));
                    end
                  else
                    begin
                      reg985 <= forvar904;
                      reg986 <= $signed(($signed($signed(reg793)) ^ $unsigned(reg948)));
                      reg987 <= forvar903;
                      reg988 <= {$signed({$signed((8'hae))})};
                    end
                  for (forvar989 = (1'h0); (forvar989 < (2'h2)); forvar989 = (forvar989 + (1'h1)))
                    begin
                      reg990 <= $signed(((reg861[(3'h6):(3'h5)] && (forvar892 != reg979)) ?
                          (((8'had) ^ forvar975) <= (^reg809)) : $unsigned((reg962 ?
                              reg902 : forvar970))));
                    end
                  reg991 <= $unsigned($unsigned((~|(&(8'hb0)))));
                  for (forvar992 = (1'h0); (forvar992 < (2'h2)); forvar992 = (forvar992 + (1'h1)))
                    begin
                      reg993 <= reg801;
                      reg994 <= forvar903[(2'h2):(1'h0)];
                      reg995 <= $unsigned({reg929});
                      reg996 <= $signed($unsigned(($signed((8'hb8)) ?
                          ((8'ha0) >> reg892) : $unsigned(reg801))));
                    end
                end
              else
                begin
                  for (forvar985 = (1'h0); (forvar985 < (1'h1)); forvar985 = (forvar985 + (1'h1)))
                    begin
                      reg986 <= reg830[(4'ha):(3'h7)];
                    end
                  reg987 <= reg856;
                  reg988 <= reg859;
                  for (forvar989 = (1'h0); (forvar989 < (2'h2)); forvar989 = (forvar989 + (1'h1)))
                    begin
                      reg990 <= {((~&(reg957 ~^ forvar787)) >> {reg943[(3'h7):(3'h7)]})};
                      reg991 <= $signed($signed(($unsigned(reg830) ?
                          $signed(forvar804) : (reg950 | (8'h9d)))));
                      reg992 <= ((reg922[(2'h3):(1'h0)] ?
                          ((reg944 ?
                              forvar827 : (8'hb0)) ^ (forvar807 >>> reg841)) : $signed((reg966 ?
                              reg852 : (8'h9f)))) == $signed(forvar834));
                      reg993 <= ($unsigned($signed($signed(forvar946))) & reg986[(4'ha):(3'h4)]);
                    end
                end
            end
        end
      else
        begin
          reg930 <= $unsigned($signed(reg942[(3'h4):(1'h1)]));
          for (forvar931 = (1'h0); (forvar931 < (2'h2)); forvar931 = (forvar931 + (1'h1)))
            begin
              reg932 <= wire597[(4'ha):(3'h5)];
              for (forvar933 = (1'h0); (forvar933 < (2'h3)); forvar933 = (forvar933 + (1'h1)))
                begin
                  for (forvar934 = (1'h0); (forvar934 < (2'h3)); forvar934 = (forvar934 + (1'h1)))
                    begin
                      reg935 <= $unsigned($unsigned($signed((forvar804 < forvar827))));
                      reg936 <= (8'ha6);
                      reg937 <= $signed($unsigned({$unsigned(forvar951)}));
                      reg938 <= (reg894[(2'h3):(1'h1)] ?
                          (~&$unsigned($signed(reg897))) : {(!reg849)});
                    end
                end
              reg939 <= forvar985;
              for (forvar940 = (1'h0); (forvar940 < (2'h3)); forvar940 = (forvar940 + (1'h1)))
                begin
                  if (($signed(($signed(reg845) ?
                      reg898 : (+forvar902))) != (-{reg874[(2'h2):(2'h2)]})))
                    begin
                      reg941 <= {(reg943 > (&forvar989))};
                      reg942 <= reg826[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg941 <= reg832;
                      reg942 <= (^~($signed((reg872 ? forvar880 : (8'hb1))) ?
                          $unsigned($unsigned(reg917)) : (~|$unsigned(reg831))));
                      reg943 <= (+({reg906} ?
                          (forvar892[(4'ha):(3'h7)] * (reg895 ?
                              reg808 : reg970)) : $signed({reg937})));
                    end
                  for (forvar944 = (1'h0); (forvar944 < (2'h2)); forvar944 = (forvar944 + (1'h1)))
                    begin
                      reg945 <= forvar874[(4'ha):(4'h8)];
                      reg946 <= ($unsigned(((|(8'ha5)) >>> $unsigned(wire592))) ?
                          ({$unsigned(reg916)} != {(+(8'ha1))}) : reg848[(3'h6):(2'h3)]);
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar997 = (1'h0); (forvar997 < (1'h0)); forvar997 = (forvar997 + (1'h1)))
        begin
          if ($signed($unsigned($signed($unsigned(reg822)))))
            begin
              for (forvar998 = (1'h0); (forvar998 < (1'h0)); forvar998 = (forvar998 + (1'h1)))
                begin
                  reg999 <= ($signed((~&{(8'h9c)})) == $unsigned($unsigned($unsigned(reg920))));
                end
            end
          else
            begin
              if (reg987)
                begin
                  reg998 <= ((($signed(reg893) ?
                      (wire595 ? reg921 : reg922) : forvar836) && (~&(reg985 ?
                      (8'had) : reg862))) == $unsigned($unsigned((!reg862))));
                  for (forvar999 = (1'h0); (forvar999 < (2'h2)); forvar999 = (forvar999 + (1'h1)))
                    begin
                      reg1000 <= ($signed(reg998[(3'h7):(1'h1)]) ?
                          ({{forvar946}} ? reg833 : (^forvar822)) : forvar931);
                      reg1001 <= reg878[(3'h6):(2'h3)];
                      reg1002 <= $unsigned(($unsigned(wire592[(2'h3):(1'h0)]) < (forvar874 > (^~reg920))));
                    end
                  for (forvar1003 = (1'h0); (forvar1003 < (2'h2)); forvar1003 = (forvar1003 + (1'h1)))
                    begin
                      reg1004 <= (&reg941);
                      reg1005 <= (reg822 ?
                          $unsigned({$unsigned(reg889)}) : ({(reg941 <= (8'ha1))} ?
                              $unsigned((reg906 ?
                                  reg984 : reg820)) : $unsigned(reg810[(2'h2):(2'h2)])));
                      reg1006 <= forvar826[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  if ($signed((|{$unsigned(reg946)})))
                    begin
                      reg998 <= (~reg841);
                      reg999 <= (|(($signed(forvar904) == reg1005) < reg912));
                      reg1000 <= ($unsigned(($signed(reg889) ^~ (forvar921 <<< reg926))) >>> (reg953 - $unsigned((reg802 ?
                          reg796 : reg982))));
                      reg1001 <= reg887;
                    end
                  else
                    begin
                      reg998 <= reg820;
                      reg999 <= ((!(+(wire595 + forvar944))) ?
                          reg842[(3'h6):(2'h3)] : (~|(reg916 ?
                              $signed(reg884) : forvar969[(3'h6):(2'h2)])));
                    end
                  for (forvar1002 = (1'h0); (forvar1002 < (1'h1)); forvar1002 = (forvar1002 + (1'h1)))
                    begin
                      reg1003 <= $unsigned(($signed((~^reg907)) ?
                          $unsigned(reg885) : $signed(reg816[(3'h7):(3'h5)])));
                      reg1004 <= forvar883;
                    end
                end
              for (forvar1007 = (1'h0); (forvar1007 < (1'h1)); forvar1007 = (forvar1007 + (1'h1)))
                begin
                  if ($unsigned({{$signed(reg824)}}))
                    begin
                      reg1008 <= (8'ha6);
                      reg1009 <= reg994[(3'h4):(2'h3)];
                      reg1010 <= ((!(forvar892[(4'hb):(3'h6)] ?
                              (reg987 ~^ reg850) : (|reg849))) ?
                          (+$unsigned(reg916)) : (reg861 == $unsigned((reg938 ^~ reg929))));
                      reg1011 <= ($signed($unsigned({(8'hac)})) - (~^$unsigned(reg821[(3'h6):(1'h1)])));
                    end
                  else
                    begin
                      reg1008 <= reg861[(2'h2):(1'h0)];
                      reg1009 <= reg932;
                      reg1010 <= $unsigned({(~^forvar880[(1'h1):(1'h1)])});
                    end
                  if ($signed($unsigned(((forvar896 ?
                      forvar1003 : forvar791) ^ (^(8'hb0))))))
                    begin
                      reg1012 <= $unsigned((^(reg944 ?
                          (8'had) : $unsigned(reg840))));
                      reg1013 <= $unsigned((~|reg979[(4'hc):(4'h9)]));
                      reg1014 <= $unsigned($signed(((reg878 >= forvar970) ?
                          forvar892 : (reg928 ? reg859 : reg1003))));
                    end
                  else
                    begin
                      reg1012 <= $signed(((~^(reg916 ? reg856 : reg919)) ?
                          $signed(reg804) : $signed((reg902 ?
                              reg828 : reg867))));
                      reg1013 <= reg988[(1'h1):(1'h1)];
                      reg1014 <= $unsigned(($signed((reg887 >= reg963)) && $unsigned(forvar881[(3'h6):(1'h1)])));
                      reg1015 <= $signed($unsigned($unsigned($signed(forvar904))));
                    end
                  for (forvar1016 = (1'h0); (forvar1016 < (1'h0)); forvar1016 = (forvar1016 + (1'h1)))
                    begin
                      reg1017 <= ((($unsigned(reg868) ~^ $signed(reg869)) ?
                          $unsigned((^reg941)) : ($unsigned((8'hb7)) ?
                              forvar796[(3'h4):(1'h1)] : (8'haa))) >>> $unsigned($signed(reg835)));
                      reg1018 <= (reg1004 ?
                          reg884 : (((8'hb0) >= {reg837}) ^~ (+(reg867 ?
                              forvar876 : reg976))));
                      reg1019 <= (wire599 ?
                          (~($unsigned(reg877) ?
                              forvar787[(2'h2):(1'h1)] : {(8'hab)})) : (~|((&reg925) != reg804[(1'h1):(1'h0)])));
                      reg1020 <= $unsigned((8'h9f));
                    end
                end
            end
          reg1021 <= $unsigned(forvar901);
          reg1022 <= {(((reg924 ?
                  forvar801 : reg802) << (~forvar881)) || (((8'ha4) ?
                      forvar883 : reg870) ?
                  ((8'hba) - reg919) : $signed(forvar818)))};
        end
      for (forvar1023 = (1'h0); (forvar1023 < (1'h0)); forvar1023 = (forvar1023 + (1'h1)))
        begin
          for (forvar1024 = (1'h0); (forvar1024 < (1'h0)); forvar1024 = (forvar1024 + (1'h1)))
            begin
              for (forvar1025 = (1'h0); (forvar1025 < (2'h2)); forvar1025 = (forvar1025 + (1'h1)))
                begin
                  for (forvar1026 = (1'h0); (forvar1026 < (1'h1)); forvar1026 = (forvar1026 + (1'h1)))
                    begin
                      reg1027 <= {(^~(((8'h9f) ? reg800 : forvar933) ?
                              (reg930 && wire595) : forvar916))};
                      reg1028 <= $signed(reg832);
                      reg1029 <= (reg967[(2'h3):(2'h2)] ?
                          reg911[(1'h0):(1'h0)] : {(^~(+wire598))});
                    end
                  reg1030 <= ((~^reg886[(4'ha):(4'ha)]) * reg831);
                  for (forvar1031 = (1'h0); (forvar1031 < (1'h1)); forvar1031 = (forvar1031 + (1'h1)))
                    begin
                      reg1032 <= (8'ha5);
                      reg1033 <= $unsigned((~&forvar827[(1'h0):(1'h0)]));
                    end
                  for (forvar1034 = (1'h0); (forvar1034 < (2'h2)); forvar1034 = (forvar1034 + (1'h1)))
                    begin
                      reg1035 <= (reg894[(4'hb):(3'h6)] ?
                          (!($signed((8'ha2)) ?
                              reg941[(2'h2):(1'h1)] : (~|forvar879))) : (~^(((8'ha2) ?
                              (8'ha9) : reg983) ^~ (reg930 ^ (8'ha8)))));
                    end
                end
            end
          if ($unsigned(forvar831))
            begin
              reg1036 <= reg868[(3'h7):(2'h3)];
              for (forvar1037 = (1'h0); (forvar1037 < (1'h0)); forvar1037 = (forvar1037 + (1'h1)))
                begin
                  for (forvar1038 = (1'h0); (forvar1038 < (1'h0)); forvar1038 = (forvar1038 + (1'h1)))
                    begin
                      reg1039 <= (($signed(reg852) ?
                          $signed(forvar814) : $signed({reg830})) == (((8'hb4) ?
                          reg866[(4'hd):(4'h8)] : reg1020) | (~$signed(reg836))));
                      reg1040 <= $unsigned(forvar827[(2'h3):(2'h2)]);
                    end
                  for (forvar1041 = (1'h0); (forvar1041 < (2'h2)); forvar1041 = (forvar1041 + (1'h1)))
                    begin
                      reg1042 <= forvar814;
                      reg1043 <= (((^$unsigned(reg963)) ~^ (8'hb7)) ?
                          ((+(reg793 + forvar837)) & $signed({(8'ha2)})) : {{$signed((8'hb1))}});
                    end
                  for (forvar1044 = (1'h0); (forvar1044 < (2'h2)); forvar1044 = (forvar1044 + (1'h1)))
                    begin
                      reg1045 <= $signed($signed((^(reg822 > reg825))));
                      reg1046 <= $unsigned((8'hb8));
                      reg1047 <= (reg846[(2'h3):(1'h0)] & reg895[(2'h2):(1'h0)]);
                    end
                end
            end
          else
            begin
              for (forvar1036 = (1'h0); (forvar1036 < (1'h0)); forvar1036 = (forvar1036 + (1'h1)))
                begin
                  for (forvar1037 = (1'h0); (forvar1037 < (2'h3)); forvar1037 = (forvar1037 + (1'h1)))
                    begin
                      reg1038 <= ((+(&$signed(reg967))) & forvar826[(2'h2):(2'h2)]);
                      reg1039 <= $signed($unsigned(forvar1024[(2'h3):(1'h1)]));
                      reg1040 <= forvar960[(4'ha):(3'h7)];
                      reg1041 <= reg806[(1'h1):(1'h0)];
                    end
                  if ($unsigned(({forvar889} < reg925)))
                    begin
                      reg1042 <= $signed($unsigned(forvar913));
                      reg1043 <= {(+(~|((8'ha7) ? reg964 : forvar935)))};
                    end
                  else
                    begin
                      reg1042 <= ((($unsigned(forvar960) ^ (reg819 ?
                              reg885 : reg791)) | (!$unsigned(forvar811))) ?
                          $signed(($signed(reg1046) <= (^~forvar826))) : {$unsigned((reg1005 ?
                                  (8'hb6) : (8'h9c)))});
                      reg1043 <= reg833;
                    end
                end
            end
          for (forvar1048 = (1'h0); (forvar1048 < (1'h1)); forvar1048 = (forvar1048 + (1'h1)))
            begin
              for (forvar1049 = (1'h0); (forvar1049 < (1'h0)); forvar1049 = (forvar1049 + (1'h1)))
                begin
                  if (reg953[(1'h1):(1'h0)])
                    begin
                      reg1050 <= forvar1031[(1'h0):(1'h0)];
                      reg1051 <= $unsigned(reg967[(2'h3):(2'h2)]);
                      reg1052 <= (($unsigned(reg866[(4'hc):(3'h5)]) ?
                              forvar940[(1'h0):(1'h0)] : (-(reg986 < reg952))) ?
                          $unsigned($unsigned($unsigned(reg871))) : (($signed((8'h9d)) ?
                                  $unsigned(reg832) : $signed(reg927)) ?
                              $unsigned((forvar880 ?
                                  (8'h9f) : reg973)) : $unsigned((&reg829))));
                    end
                  else
                    begin
                      reg1050 <= $unsigned((reg1003 ?
                          (+reg1029[(1'h1):(1'h0)]) : forvar831[(1'h1):(1'h1)]));
                    end
                end
              reg1053 <= {(8'h9d)};
              reg1054 <= (+{$unsigned(reg918)});
            end
        end
      if (($unsigned($signed(reg1039)) >>> (8'h9e)))
        begin
          if ($signed(reg1032[(1'h0):(1'h0)]))
            begin
              for (forvar1055 = (1'h0); (forvar1055 < (2'h3)); forvar1055 = (forvar1055 + (1'h1)))
                begin
                  for (forvar1056 = (1'h0); (forvar1056 < (2'h2)); forvar1056 = (forvar1056 + (1'h1)))
                    begin
                      reg1057 <= ($signed({{reg912}}) ?
                          reg825[(2'h3):(2'h3)] : (~^{forvar860[(4'ha):(3'h4)]}));
                    end
                  reg1058 <= $unsigned(({(8'ha1)} ?
                      ($signed(forvar825) ?
                          (forvar911 == reg985) : (8'ha3)) : reg1021));
                  if ({$unsigned(((reg873 ?
                          forvar896 : reg916) || $unsigned(forvar916)))})
                    begin
                      reg1059 <= ($signed(reg813) ?
                          $unsigned((forvar813 || (8'hae))) : reg901[(3'h5):(2'h2)]);
                      reg1060 <= {$signed(((~|(8'haf)) + (forvar930 ~^ reg1000)))};
                      reg1061 <= $unsigned($signed({reg816[(3'h4):(1'h1)]}));
                    end
                  else
                    begin
                      reg1059 <= ((reg896[(1'h0):(1'h0)] <= (((8'h9e) ?
                                  forvar881 : (8'h9d)) ?
                              $unsigned(forvar951) : $signed((8'h9d)))) ?
                          reg1008 : (^$unsigned(reg910[(4'hc):(4'h8)])));
                      reg1060 <= (~^(~&({forvar1007} ?
                          $signed(reg794) : ((8'ha8) ? (8'h9d) : forvar891))));
                    end
                  for (forvar1062 = (1'h0); (forvar1062 < (1'h1)); forvar1062 = (forvar1062 + (1'h1)))
                    begin
                      reg1063 <= forvar820[(3'h5):(2'h2)];
                      reg1064 <= ((reg918[(4'hd):(4'h9)] ~^ $signed($unsigned((8'hb8)))) ?
                          (8'ha4) : reg1008[(5'h10):(1'h0)]);
                      reg1065 <= $unsigned((({reg982} ?
                              $signed(reg1051) : $unsigned(reg1043)) ?
                          wire783[(1'h0):(1'h0)] : (+reg847[(1'h0):(1'h0)])));
                      reg1066 <= ((reg1045[(3'h4):(3'h4)] | $signed((forvar880 ?
                          wire596 : forvar885))) && (reg935[(2'h3):(2'h3)] + (^(^forvar800))));
                    end
                end
            end
          else
            begin
              for (forvar1055 = (1'h0); (forvar1055 < (2'h2)); forvar1055 = (forvar1055 + (1'h1)))
                begin
                  for (forvar1056 = (1'h0); (forvar1056 < (2'h3)); forvar1056 = (forvar1056 + (1'h1)))
                    begin
                      reg1057 <= ((~|reg1053) ?
                          (~(~&$unsigned(forvar887))) : (reg936 ?
                              (((8'hb0) ?
                                  forvar885 : forvar791) && $signed(reg870)) : $unsigned((-(8'hb5)))));
                      reg1058 <= ($signed($signed(reg986[(4'hb):(4'hb)])) >>> ($unsigned({reg827}) & forvar1002));
                    end
                  reg1059 <= $unsigned({$signed(forvar796[(3'h5):(2'h2)])});
                end
              if ({forvar945[(3'h5):(1'h1)]})
                begin
                  for (forvar1060 = (1'h0); (forvar1060 < (2'h3)); forvar1060 = (forvar1060 + (1'h1)))
                    begin
                      reg1061 <= $signed($unsigned(({forvar989} ?
                          (~reg1020) : $unsigned(reg816))));
                    end
                  if ({($unsigned((|reg849)) ?
                          $signed($unsigned(forvar889)) : $signed((wire597 ?
                              reg1027 : (8'had))))})
                    begin
                      reg1062 <= (reg795[(3'h7):(1'h0)] || (forvar834 ~^ reg967));
                    end
                  else
                    begin
                      reg1062 <= (forvar799 ?
                          (((reg801 > (8'hb7)) ?
                              (~reg910) : (+reg869)) <= {(reg1035 ?
                                  forvar822 : reg937)}) : (!(8'ha3)));
                      reg1063 <= (8'h9e);
                    end
                  if (reg801)
                    begin
                      reg1064 <= ((|(8'haf)) + ((reg887 ?
                              $unsigned(forvar941) : $unsigned(reg788)) ?
                          forvar997 : $signed($signed(forvar885))));
                      reg1065 <= (~&(reg998 ? $signed(reg943) : (|{reg839})));
                    end
                  else
                    begin
                      reg1064 <= ({reg888} ?
                          $unsigned(reg865[(1'h1):(1'h1)]) : reg927);
                      reg1065 <= reg829[(1'h0):(1'h0)];
                    end
                  if ((|reg944[(3'h6):(1'h0)]))
                    begin
                      reg1066 <= reg994[(2'h2):(2'h2)];
                      reg1067 <= reg1038;
                    end
                  else
                    begin
                      reg1066 <= (reg852 ?
                          ((&reg825[(2'h3):(2'h3)]) ?
                              $signed(reg939[(1'h0):(1'h0)]) : ((forvar876 ~^ reg818) ~^ $unsigned(reg1014))) : forvar837[(2'h2):(2'h2)]);
                      reg1067 <= (8'hb0);
                    end
                end
              else
                begin
                  for (forvar1060 = (1'h0); (forvar1060 < (1'h1)); forvar1060 = (forvar1060 + (1'h1)))
                    begin
                      reg1061 <= ($signed((~|reg918[(3'h7):(1'h0)])) * $signed((reg871[(3'h4):(1'h1)] ?
                          (~|forvar894) : (forvar876 ? reg835 : forvar1055))));
                    end
                  if ($signed({forvar940}))
                    begin
                      reg1062 <= $unsigned((reg1054 ?
                          ((reg868 ?
                              reg912 : reg794) > (8'h9f)) : $signed($unsigned(reg937))));
                      reg1063 <= (~|reg923[(2'h3):(1'h1)]);
                      reg1064 <= {$unsigned(((forvar997 ~^ forvar891) ^~ reg985))};
                    end
                  else
                    begin
                      reg1062 <= ($signed((((8'ha1) >= (8'ha2)) + reg916[(1'h1):(1'h1)])) & (~&({(8'h9e)} ?
                          forvar1037[(1'h0):(1'h0)] : {reg1040})));
                      reg1063 <= $unsigned((8'ha6));
                      reg1064 <= reg986[(4'hd):(4'h9)];
                    end
                  for (forvar1065 = (1'h0); (forvar1065 < (1'h1)); forvar1065 = (forvar1065 + (1'h1)))
                    begin
                      reg1066 <= forvar804;
                    end
                end
            end
        end
      else
        begin
          if ((^reg869[(4'h8):(3'h5)]))
            begin
              reg1055 <= ((8'hba) > forvar915[(3'h6):(2'h3)]);
            end
          else
            begin
              reg1055 <= reg911[(2'h2):(2'h2)];
              for (forvar1056 = (1'h0); (forvar1056 < (1'h1)); forvar1056 = (forvar1056 + (1'h1)))
                begin
                  reg1057 <= ({$signed((forvar785 * reg796))} ?
                      reg933 : ((~|(reg927 ? (8'ha2) : forvar1024)) ?
                          forvar998[(2'h2):(2'h2)] : (reg871[(3'h7):(1'h0)] * (|forvar1056))));
                  if (forvar899)
                    begin
                      reg1058 <= $signed({(+(&forvar876))});
                    end
                  else
                    begin
                      reg1058 <= forvar1044[(3'h4):(1'h0)];
                    end
                  reg1059 <= ((forvar1062 ?
                      $signed((reg954 & reg869)) : ((reg899 && reg994) ?
                          reg809[(4'ha):(1'h0)] : $signed((8'hb0)))) && ($signed({reg1065}) ?
                      $unsigned(reg836) : (!(&reg872))));
                end
              if ((~&$signed((((8'haa) && (8'hab)) ?
                  reg832[(1'h0):(1'h0)] : reg1039))))
                begin
                  for (forvar1060 = (1'h0); (forvar1060 < (2'h2)); forvar1060 = (forvar1060 + (1'h1)))
                    begin
                      reg1061 <= $unsigned($unsigned(((-(8'hb8)) ^ (reg931 ?
                          forvar1034 : (8'hb3)))));
                      reg1062 <= reg822;
                      reg1063 <= ({(~&reg849)} * {reg940[(3'h6):(3'h4)]});
                      reg1064 <= $unsigned({forvar1016});
                    end
                  for (forvar1065 = (1'h0); (forvar1065 < (2'h3)); forvar1065 = (forvar1065 + (1'h1)))
                    begin
                      reg1066 <= forvar960[(4'h8):(4'h8)];
                    end
                  if (reg797[(1'h0):(1'h0)])
                    begin
                      reg1067 <= ((~^reg919) * $unsigned($signed((reg905 > (8'hb5)))));
                      reg1068 <= ((8'h9c) ?
                          (!((reg841 ? wire594 : reg1057) ?
                              forvar939[(2'h3):(2'h2)] : (reg953 ?
                                  reg808 : forvar1036))) : (({reg931} << forvar785[(3'h6):(1'h1)]) ?
                              ($signed(reg825) >> reg855) : $signed(reg1041[(2'h3):(2'h3)])));
                    end
                  else
                    begin
                      reg1067 <= reg830;
                      reg1068 <= forvar837;
                      reg1069 <= (+$signed(((reg1042 != forvar799) ?
                          reg835[(4'hc):(4'h8)] : forvar1041[(3'h7):(3'h7)])));
                      reg1070 <= {({forvar1049} == (((8'hba) <<< reg992) ?
                              $unsigned(reg837) : forvar908[(2'h2):(1'h0)]))};
                    end
                end
              else
                begin
                  for (forvar1060 = (1'h0); (forvar1060 < (2'h3)); forvar1060 = (forvar1060 + (1'h1)))
                    begin
                      reg1061 <= reg1040;
                      reg1062 <= (|$signed({$signed(wire597)}));
                      reg1063 <= $unsigned(((~&(forvar806 ?
                              (8'ha4) : (8'hb4))) ?
                          forvar827[(3'h6):(3'h6)] : ({forvar1060} > (reg885 ?
                              forvar1048 : forvar891))));
                    end
                  for (forvar1064 = (1'h0); (forvar1064 < (1'h0)); forvar1064 = (forvar1064 + (1'h1)))
                    begin
                      reg1065 <= reg923[(1'h1):(1'h0)];
                      reg1066 <= wire596[(1'h0):(1'h0)];
                      reg1067 <= (reg931 ?
                          wire783[(2'h3):(2'h3)] : reg1045[(1'h1):(1'h1)]);
                    end
                end
              reg1071 <= (^~reg928);
            end
          if (reg796[(2'h3):(2'h2)])
            begin
              if (reg912)
                begin
                  for (forvar1072 = (1'h0); (forvar1072 < (1'h1)); forvar1072 = (forvar1072 + (1'h1)))
                    begin
                      reg1073 <= reg793[(2'h2):(1'h1)];
                      reg1074 <= $unsigned(forvar818[(4'h8):(2'h2)]);
                      reg1075 <= ($unsigned((reg795[(3'h4):(2'h3)] ?
                              forvar1049[(2'h3):(1'h0)] : (-reg788))) ?
                          reg869[(3'h4):(1'h0)] : (($unsigned(reg819) && (reg861 + reg1066)) ?
                              ((8'hb6) ?
                                  $unsigned(forvar794) : reg1015) : $signed((reg964 == reg835))));
                      reg1076 <= $signed(reg983);
                    end
                end
              else
                begin
                  for (forvar1072 = (1'h0); (forvar1072 < (1'h0)); forvar1072 = (forvar1072 + (1'h1)))
                    begin
                      reg1073 <= $signed({$unsigned(reg1038[(4'h9):(1'h1)])});
                      reg1074 <= ({$unsigned((reg874 ?
                              (8'h9f) : reg866))} << {{(wire596 & (8'hae))}});
                      reg1075 <= reg1073[(1'h0):(1'h0)];
                      reg1076 <= ($unsigned({forvar879}) ?
                          forvar975[(3'h5):(1'h0)] : (reg927[(2'h3):(1'h1)] && $unsigned((~^reg912))));
                    end
                  if ((|forvar934[(4'ha):(2'h3)]))
                    begin
                      reg1077 <= (&$signed(forvar801[(1'h0):(1'h0)]));
                      reg1078 <= ($signed({reg884}) >= (!$signed((~reg1074))));
                    end
                  else
                    begin
                      reg1077 <= (^~$signed({reg979[(4'hc):(1'h0)]}));
                    end
                  if (forvar1049[(2'h3):(2'h2)])
                    begin
                      reg1079 <= reg888;
                    end
                  else
                    begin
                      reg1079 <= reg1057[(3'h4):(1'h0)];
                      reg1080 <= (^$unsigned({(wire595 ?
                              forvar891 : (8'ha0))}));
                      reg1081 <= ((~&(reg933[(4'hc):(3'h6)] ?
                          (reg1047 ?
                              reg872 : reg853) : reg957)) + ((forvar959[(3'h5):(1'h1)] + (+reg911)) > reg943));
                      reg1082 <= forvar879;
                    end
                end
              for (forvar1083 = (1'h0); (forvar1083 < (2'h3)); forvar1083 = (forvar1083 + (1'h1)))
                begin
                  if (forvar864[(1'h0):(1'h0)])
                    begin
                      reg1084 <= (8'had);
                    end
                  else
                    begin
                      reg1084 <= (~^forvar945[(2'h3):(2'h3)]);
                      reg1085 <= $unsigned(($unsigned(((8'ha8) ?
                              reg894 : forvar1055)) ?
                          ($signed(reg1076) ?
                              (reg1036 ?
                                  reg939 : forvar864) : $signed(reg1063)) : $unsigned((8'hb1))));
                      reg1086 <= reg911[(1'h1):(1'h0)];
                      reg1087 <= forvar857[(2'h3):(2'h3)];
                    end
                  if ({((reg893 ?
                          (forvar1037 ?
                              reg1058 : (8'hac)) : reg987[(3'h4):(2'h2)]) << reg1027[(1'h1):(1'h1)])})
                    begin
                      reg1088 <= $signed((~^reg810[(4'h9):(2'h2)]));
                      reg1089 <= reg1052;
                      reg1090 <= (($unsigned(forvar1041) >= $unsigned((reg914 ^~ reg862))) <<< reg794);
                      reg1091 <= (((-$signed(forvar1007)) >= {$signed((8'h9e))}) ?
                          $unsigned({(forvar901 ?
                                  reg949 : forvar997)}) : reg848[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg1088 <= reg884[(1'h1):(1'h1)];
                      reg1089 <= (~&$signed(forvar868[(1'h1):(1'h1)]));
                      reg1090 <= (reg1047 ?
                          forvar800[(2'h3):(2'h2)] : (~reg821));
                    end
                end
              reg1092 <= reg1063;
              if (reg866[(4'ha):(1'h0)])
                begin
                  for (forvar1093 = (1'h0); (forvar1093 < (1'h0)); forvar1093 = (forvar1093 + (1'h1)))
                    begin
                      reg1094 <= $unsigned(forvar935[(1'h1):(1'h1)]);
                      reg1095 <= (&$unsigned($signed((~(8'hb3)))));
                      reg1096 <= ((8'hb5) >>> {wire599});
                      reg1097 <= (~^(reg979[(3'h7):(1'h1)] || (^(reg948 <<< forvar977))));
                    end
                  for (forvar1098 = (1'h0); (forvar1098 < (1'h0)); forvar1098 = (forvar1098 + (1'h1)))
                    begin
                      reg1099 <= $signed((~|{reg906}));
                      reg1100 <= (^$signed((reg846 << (^~reg1077))));
                      reg1101 <= ($unsigned(forvar887[(2'h3):(1'h1)]) ?
                          $unsigned(forvar800[(3'h4):(2'h2)]) : ($signed(reg1059[(4'h8):(1'h0)]) * reg1027[(3'h5):(1'h0)]));
                      reg1102 <= $unsigned((-({reg941} ?
                          (forvar886 | forvar915) : (reg1076 - reg819))));
                    end
                  for (forvar1103 = (1'h0); (forvar1103 < (2'h3)); forvar1103 = (forvar1103 + (1'h1)))
                    begin
                      reg1104 <= $unsigned((~|{(reg963 ?
                              reg956 : forvar1056)}));
                    end
                  if (reg1014)
                    begin
                      reg1105 <= $unsigned((&$unsigned({forvar1034})));
                    end
                  else
                    begin
                      reg1105 <= ($signed((8'ha9)) ~^ $unsigned(($unsigned(reg825) <= (reg885 && reg877))));
                      reg1106 <= {$signed((reg931[(1'h1):(1'h0)] ~^ (forvar904 >> forvar1026)))};
                    end
                end
              else
                begin
                  if ((+{(8'haa)}))
                    begin
                      reg1093 <= (reg1046[(3'h6):(2'h3)] < {((reg798 ?
                                  forvar1048 : reg931) ?
                              (&forvar887) : (forvar872 ? reg894 : reg798))});
                      reg1094 <= {(!(forvar951 ^ (reg1005 ~^ reg1061)))};
                      reg1095 <= (|$unsigned(reg792[(3'h4):(2'h2)]));
                      reg1096 <= $signed($unsigned($signed((reg1074 ?
                          reg996 : forvar965))));
                    end
                  else
                    begin
                      reg1093 <= $signed($unsigned(($unsigned(reg1039) + (^~reg866))));
                    end
                end
            end
          else
            begin
              if (($signed((~&(^~reg829))) ?
                  (reg890[(3'h4):(3'h4)] ?
                      forvar977 : (reg998[(1'h1):(1'h1)] ?
                          $signed(forvar791) : (wire596 ?
                              reg914 : (8'hb4)))) : (^~{reg1009[(1'h0):(1'h0)]})))
                begin
                  if (((wire599[(2'h3):(2'h2)] ?
                          forvar901 : ((~|(8'haa)) | forvar860[(3'h7):(3'h7)])) ?
                      forvar891[(1'h1):(1'h1)] : (forvar977[(1'h0):(1'h0)] << $unsigned(reg958))))
                    begin
                      reg1072 <= {((forvar903 ~^ reg1005[(1'h0):(1'h0)]) ?
                              reg1089[(1'h1):(1'h0)] : (forvar985 ?
                                  (reg797 != reg1069) : (~|forvar951)))};
                      reg1073 <= reg944;
                    end
                  else
                    begin
                      reg1072 <= $unsigned((reg950 << $signed((~|reg954))));
                      reg1073 <= $unsigned(($unsigned(((8'hb9) ?
                              (8'hb3) : forvar874)) ?
                          $signed(reg1065) : reg824));
                      reg1074 <= (-({(reg967 == forvar921)} | $unsigned($signed(reg801))));
                    end
                  if ($unsigned(reg798[(1'h1):(1'h0)]))
                    begin
                      reg1075 <= ($signed($unsigned((forvar921 + reg865))) ?
                          $signed($unsigned((~^forvar903))) : reg799[(2'h3):(2'h3)]);
                      reg1076 <= (reg928[(3'h4):(3'h4)] ?
                          reg800 : forvar887[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg1075 <= (^$unsigned(forvar1025));
                      reg1076 <= (-($unsigned(reg796) <= reg923));
                    end
                  if ($signed(reg899))
                    begin
                      reg1077 <= (reg809 >= $signed(reg1090));
                      reg1078 <= forvar977;
                    end
                  else
                    begin
                      reg1077 <= forvar1031[(1'h1):(1'h1)];
                    end
                  for (forvar1079 = (1'h0); (forvar1079 < (1'h0)); forvar1079 = (forvar1079 + (1'h1)))
                    begin
                      reg1080 <= $signed($unsigned(((forvar1079 || reg1019) ^~ (forvar868 ?
                          forvar872 : reg1010))));
                    end
                end
              else
                begin
                  if ($unsigned(forvar939))
                    begin
                      reg1072 <= ({$signed(reg836[(3'h7):(3'h4)])} ?
                          (+reg875[(1'h0):(1'h0)]) : ($unsigned($signed(reg1004)) ?
                              ((reg892 ? reg889 : forvar885) ?
                                  $signed(forvar876) : {reg1004}) : forvar945[(1'h0):(1'h0)]));
                      reg1073 <= $unsigned($unsigned((|forvar872[(3'h4):(3'h4)])));
                      reg1074 <= (forvar1093 ?
                          $unsigned((|reg900)) : reg1054[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1072 <= (^$unsigned($unsigned($signed(forvar863))));
                      reg1073 <= reg833[(3'h7):(3'h7)];
                      reg1074 <= reg924;
                    end
                end
              if ((&reg926[(2'h3):(2'h2)]))
                begin
                  reg1081 <= (~&reg833[(4'ha):(4'h9)]);
                  for (forvar1082 = (1'h0); (forvar1082 < (1'h0)); forvar1082 = (forvar1082 + (1'h1)))
                    begin
                      reg1083 <= (((~|$signed(forvar826)) >= ((^~reg889) ?
                              (reg1000 ? (8'haa) : reg835) : reg920)) ?
                          reg1022 : {($signed(reg919) ?
                                  (^reg829) : ((8'hae) ? (8'hb3) : reg1086))});
                      reg1084 <= (~^(reg1094[(3'h5):(3'h4)] ^~ $signed((reg837 >>> reg802))));
                      reg1085 <= (($unsigned(reg1010) >> $signed((~^(8'hb2)))) & forvar998);
                    end
                end
              else
                begin
                  for (forvar1081 = (1'h0); (forvar1081 < (1'h1)); forvar1081 = (forvar1081 + (1'h1)))
                    begin
                      reg1082 <= ($signed($unsigned((^forvar1065))) > (forvar792 ?
                          ((reg1076 ?
                              forvar886 : reg954) * $unsigned(reg986)) : ((forvar1079 ?
                              reg1081 : forvar857) ^ (~&reg962))));
                      reg1083 <= $unsigned(((|reg1004) | (&(~&reg1069))));
                      reg1084 <= (+$signed(reg1008));
                    end
                  reg1085 <= {(+(+$unsigned(reg1104)))};
                  reg1086 <= ((|(~((8'hb8) ?
                      reg852 : reg809))) * $unsigned(forvar914[(4'h9):(3'h7)]));
                end
              if (reg884[(1'h1):(1'h1)])
                begin
                  for (forvar1087 = (1'h0); (forvar1087 < (1'h1)); forvar1087 = (forvar1087 + (1'h1)))
                    begin
                      reg1088 <= forvar796[(1'h1):(1'h0)];
                      reg1089 <= (~(((&forvar868) >>> forvar1060[(1'h0):(1'h0)]) ?
                          forvar945[(4'he):(1'h1)] : (~|wire593[(1'h0):(1'h0)])));
                      reg1090 <= reg816;
                    end
                end
              else
                begin
                  for (forvar1087 = (1'h0); (forvar1087 < (2'h3)); forvar1087 = (forvar1087 + (1'h1)))
                    begin
                      reg1088 <= {reg1039};
                      reg1089 <= ($signed($unsigned((-reg812))) == ((forvar887[(1'h0):(1'h0)] >= reg974) ?
                          $signed((reg918 ?
                              reg821 : (8'hb3))) : $unsigned((forvar794 * forvar944))));
                      reg1090 <= $unsigned(((!(~&reg979)) ?
                          ((~|reg994) ?
                              (!forvar1065) : ((8'h9f) >> reg1069)) : $unsigned(reg1018)));
                      reg1091 <= (+{(|(&forvar836))});
                    end
                  reg1092 <= $unsigned(forvar960[(4'h8):(3'h4)]);
                  if ($signed((forvar1065 ?
                      reg853[(3'h6):(1'h1)] : ((~^forvar1023) < (~|forvar916)))))
                    begin
                      reg1093 <= {reg899[(4'hc):(4'h8)]};
                    end
                  else
                    begin
                      reg1093 <= $unsigned(($unsigned(forvar992) ?
                          {forvar1036[(2'h3):(2'h3)]} : {(~reg1018)}));
                      reg1094 <= $unsigned(reg877[(3'h5):(2'h3)]);
                      reg1095 <= {$unsigned($unsigned($signed(forvar791)))};
                    end
                end
            end
        end
      for (forvar1107 = (1'h0); (forvar1107 < (1'h0)); forvar1107 = (forvar1107 + (1'h1)))
        begin
          if ((((~reg1011) < ((reg884 ? forvar885 : reg835) ?
              {(8'ha8)} : (^~reg915))) >>> (($unsigned(reg1078) << reg983) ?
              (!$unsigned(reg1065)) : forvar985[(2'h3):(2'h2)])))
            begin
              if (forvar1107[(4'hd):(4'hd)])
                begin
                  for (forvar1108 = (1'h0); (forvar1108 < (2'h2)); forvar1108 = (forvar1108 + (1'h1)))
                    begin
                      reg1109 <= $signed(($unsigned($unsigned(forvar876)) <<< $unsigned($signed(reg955))));
                      reg1110 <= reg1071;
                    end
                  if ($signed(((((8'had) ? reg1068 : reg948) ?
                      reg911 : {(8'hac)}) >= forvar1007[(1'h0):(1'h0)])))
                    begin
                      reg1111 <= (~$unsigned((+(reg821 ? reg1000 : wire592))));
                      reg1112 <= {reg843[(4'h8):(1'h0)]};
                    end
                  else
                    begin
                      reg1111 <= ({$unsigned({reg823})} >>> reg905[(1'h1):(1'h0)]);
                      reg1112 <= $signed($unsigned(($unsigned(reg914) ?
                          {(8'hb6)} : reg967[(1'h0):(1'h0)])));
                      reg1113 <= reg906[(2'h3):(1'h0)];
                    end
                end
              else
                begin
                  reg1108 <= ($signed(((-forvar1025) && forvar826[(2'h2):(1'h1)])) ?
                      $signed($unsigned((^reg829))) : ({(8'h9f)} || reg898));
                end
              for (forvar1114 = (1'h0); (forvar1114 < (1'h0)); forvar1114 = (forvar1114 + (1'h1)))
                begin
                  if (($signed($signed((~&forvar965))) ?
                      $signed(($unsigned(reg948) ?
                          {reg1102} : (reg926 ?
                              forvar939 : reg921))) : $unsigned(forvar814[(1'h0):(1'h0)])))
                    begin
                      reg1115 <= forvar934[(3'h4):(3'h4)];
                      reg1116 <= forvar1025;
                      reg1117 <= $unsigned(reg828[(2'h2):(1'h0)]);
                      reg1118 <= ((forvar1079[(1'h0):(1'h0)] != (reg923[(2'h3):(1'h1)] ?
                          reg992 : reg877[(3'h7):(3'h4)])) - (forvar902[(2'h2):(2'h2)] ?
                          (reg939 && forvar787) : ((^~forvar891) ?
                              $unsigned(reg1110) : $unsigned(reg1084))));
                    end
                  else
                    begin
                      reg1115 <= (!reg817[(4'h8):(2'h3)]);
                      reg1116 <= $signed((8'hba));
                    end
                  for (forvar1119 = (1'h0); (forvar1119 < (1'h1)); forvar1119 = (forvar1119 + (1'h1)))
                    begin
                      reg1120 <= $signed(({$signed(forvar1065)} && $unsigned($unsigned(reg851))));
                    end
                  if (forvar1083)
                    begin
                      reg1121 <= ($unsigned((reg862 >= forvar794[(2'h3):(1'h0)])) ?
                          reg1012[(4'he):(4'h9)] : $unsigned(({forvar913} ?
                              $signed(reg885) : $unsigned(reg847))));
                      reg1122 <= reg966;
                      reg1123 <= (~forvar1060);
                      reg1124 <= forvar854[(4'hc):(3'h5)];
                    end
                  else
                    begin
                      reg1121 <= (reg922[(3'h4):(3'h4)] * reg984);
                      reg1122 <= (((~^{reg972}) ?
                              $unsigned((reg948 != forvar1083)) : (8'ha8)) ?
                          $signed(reg816) : reg988);
                      reg1123 <= reg1097[(3'h6):(1'h1)];
                    end
                  if (({$unsigned((|forvar899))} ?
                      $unsigned($unsigned(forvar892[(4'hd):(3'h4)])) : (&(forvar899 ?
                          $unsigned(forvar836) : reg1009))))
                    begin
                      reg1125 <= reg968[(3'h6):(1'h0)];
                    end
                  else
                    begin
                      reg1125 <= (8'h9f);
                      reg1126 <= $unsigned(forvar1055[(1'h1):(1'h0)]);
                      reg1127 <= (forvar818[(1'h1):(1'h0)] ?
                          reg1101 : $signed(reg827[(1'h1):(1'h1)]));
                      reg1128 <= $signed(reg928);
                    end
                end
              reg1129 <= (~&$signed({$unsigned(reg930)}));
              for (forvar1130 = (1'h0); (forvar1130 < (2'h2)); forvar1130 = (forvar1130 + (1'h1)))
                begin
                  if (reg994[(2'h2):(1'h1)])
                    begin
                      reg1131 <= (($unsigned($signed(reg909)) << reg1002[(1'h0):(1'h0)]) || $unsigned($signed(((8'ha0) ?
                          reg896 : forvar901))));
                      reg1132 <= (&(8'hb3));
                      reg1133 <= (~&(forvar1049[(2'h2):(1'h1)] ?
                          reg1036 : (+reg1013)));
                      reg1134 <= $unsigned($unsigned($unsigned((8'ha1))));
                    end
                  else
                    begin
                      reg1131 <= (~reg1074[(3'h5):(1'h1)]);
                    end
                  for (forvar1135 = (1'h0); (forvar1135 < (2'h3)); forvar1135 = (forvar1135 + (1'h1)))
                    begin
                      reg1136 <= reg903[(3'h6):(1'h0)];
                      reg1137 <= $unsigned(forvar902);
                      reg1138 <= reg814;
                    end
                  for (forvar1139 = (1'h0); (forvar1139 < (2'h2)); forvar1139 = (forvar1139 + (1'h1)))
                    begin
                      reg1140 <= $signed($unsigned((^(~(8'hb5)))));
                      reg1141 <= {wire598};
                    end
                end
            end
          else
            begin
              for (forvar1108 = (1'h0); (forvar1108 < (1'h1)); forvar1108 = (forvar1108 + (1'h1)))
                begin
                  if ({$unsigned($unsigned($signed(reg1138)))})
                    begin
                      reg1109 <= forvar915[(3'h5):(2'h2)];
                      reg1110 <= (forvar827[(1'h0):(1'h0)] ?
                          $signed(reg910[(3'h7):(1'h1)]) : $unsigned(($unsigned(reg910) ?
                              (^~reg817) : forvar946)));
                    end
                  else
                    begin
                      reg1109 <= $signed(((((8'haa) ~^ reg1077) ?
                              ((8'hb1) ? reg801 : reg1008) : ((8'haf) ?
                                  reg1066 : reg1039)) ?
                          $unsigned(forvar997[(3'h4):(2'h2)]) : $unsigned($unsigned((8'haa)))));
                    end
                  for (forvar1111 = (1'h0); (forvar1111 < (1'h0)); forvar1111 = (forvar1111 + (1'h1)))
                    begin
                      reg1112 <= ((reg1039[(3'h4):(2'h2)] < ((&wire593) >>> $signed((8'hb8)))) ?
                          $signed($signed((forvar913 ?
                              wire594 : reg1077))) : ((|{reg898}) ?
                              reg874 : reg1015[(1'h0):(1'h0)]));
                      reg1113 <= (!forvar888[(3'h7):(2'h3)]);
                      reg1114 <= forvar791;
                    end
                  if (reg895)
                    begin
                      reg1115 <= $signed($unsigned(((!reg1131) >> forvar822[(4'ha):(3'h6)])));
                    end
                  else
                    begin
                      reg1115 <= reg1128[(3'h4):(1'h1)];
                      reg1116 <= ($signed(((forvar934 == reg868) ?
                          (~&reg1105) : reg1089)) == ({forvar879[(3'h4):(2'h3)]} || (forvar885[(1'h0):(1'h0)] == ((8'haf) ?
                          reg1029 : reg853))));
                      reg1117 <= ($signed($signed(forvar868[(2'h2):(2'h2)])) ?
                          forvar959 : {forvar806});
                      reg1118 <= (~reg1127[(3'h6):(3'h4)]);
                    end
                  if ($unsigned($signed(($unsigned(reg1038) < $unsigned(reg900)))))
                    begin
                      reg1119 <= reg1129;
                      reg1120 <= (~^((reg935 & reg976[(1'h0):(1'h0)]) >> ((forvar880 ?
                          reg1134 : reg1101) >> $unsigned(reg1076))));
                    end
                  else
                    begin
                      reg1119 <= {(reg885[(4'h9):(4'h8)] ?
                              {(|forvar1098)} : reg800[(3'h4):(1'h0)])};
                    end
                end
              if ((8'haa))
                begin
                  if (reg1038[(4'h8):(1'h0)])
                    begin
                      reg1121 <= reg1125[(3'h6):(3'h4)];
                      reg1122 <= reg1041[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1121 <= $signed(reg1059);
                      reg1122 <= reg981;
                    end
                  if ((forvar1049 - ($unsigned((forvar1055 ^~ reg943)) - $unsigned((reg834 + (8'ha8))))))
                    begin
                      reg1123 <= reg1050[(3'h4):(2'h3)];
                      reg1124 <= (~(reg855 > forvar834[(4'h9):(1'h1)]));
                    end
                  else
                    begin
                      reg1123 <= $signed($unsigned($signed((reg803 ?
                          reg971 : reg1050))));
                      reg1124 <= (|(($signed(reg1133) || (wire596 ?
                          forvar1044 : (8'h9f))) ^~ (^~(wire592 ?
                          reg1030 : wire596))));
                      reg1125 <= (reg1126 + (reg862 ?
                          $unsigned(reg1087[(3'h5):(2'h2)]) : $signed($signed(reg901))));
                    end
                  if (((reg973 >= {(~reg918)}) ?
                      reg1087[(1'h1):(1'h0)] : $unsigned($unsigned((forvar904 < reg882)))))
                    begin
                      reg1126 <= (((|(!(8'ha5))) << reg924) <<< (8'ha7));
                      reg1127 <= $signed((+((reg948 ? reg995 : (8'ha0)) ?
                          reg908 : (8'hae))));
                      reg1128 <= $unsigned(reg1006);
                    end
                  else
                    begin
                      reg1126 <= (!($unsigned((forvar799 ?
                          forvar914 : reg992)) ^ $signed(reg1070)));
                      reg1127 <= reg940;
                    end
                end
              else
                begin
                  for (forvar1121 = (1'h0); (forvar1121 < (2'h2)); forvar1121 = (forvar1121 + (1'h1)))
                    begin
                      reg1122 <= reg1127[(1'h1):(1'h0)];
                      reg1123 <= $signed((((reg1102 ? reg875 : (8'hb4)) ?
                          (8'hb5) : $signed(reg984)) ^ (~reg803)));
                      reg1124 <= $signed($unsigned(({reg818} && $signed((8'hb3)))));
                      reg1125 <= reg855[(3'h7):(3'h5)];
                    end
                  for (forvar1126 = (1'h0); (forvar1126 < (2'h3)); forvar1126 = (forvar1126 + (1'h1)))
                    begin
                      reg1127 <= forvar818;
                    end
                  for (forvar1128 = (1'h0); (forvar1128 < (1'h0)); forvar1128 = (forvar1128 + (1'h1)))
                    begin
                      reg1129 <= ((8'hb4) >>> $unsigned({forvar1038[(1'h1):(1'h0)]}));
                      reg1130 <= (reg983 ?
                          $signed(((!forvar975) ?
                              (reg1081 ?
                                  reg869 : reg1060) : (+reg796))) : {(^~{reg1117})});
                      reg1131 <= (~|(({(8'haf)} >>> reg852[(3'h4):(1'h1)]) <<< ({reg855} ?
                          $unsigned(reg948) : (reg903 ? reg1002 : forvar866))));
                      reg1132 <= ($unsigned($unsigned(reg875[(3'h6):(3'h4)])) ?
                          ((+$unsigned(reg1004)) ?
                              (reg920[(3'h4):(1'h1)] && (&reg1093)) : ((reg972 ?
                                  (8'ha5) : reg805) - (+reg806))) : (-$signed({(8'ha5)})));
                    end
                end
              reg1133 <= {((8'hb5) || $signed($unsigned(forvar1007)))};
            end
        end
    end
  assign wire1142 = reg872;
  assign wire1143 = $signed({($unsigned((8'hac)) ?
                            ((8'haf) && forvar892) : (forvar913 ?
                                reg887 : reg847))});
  assign wire1144 = $signed(forvar1139);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module600  (y, clk, wire604, wire603, wire602, wire601);
  output wire [(32'h7e1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire604;
  input wire signed [(3'h4):(1'h0)] wire603;
  input wire [(5'h10):(1'h0)] wire602;
  input wire signed [(4'h8):(1'h0)] wire601;
  wire signed [(3'h5):(1'h0)] wire782;
  wire signed [(3'h6):(1'h0)] wire781;
  wire [(4'hf):(1'h0)] wire780;
  wire signed [(4'he):(1'h0)] wire779;
  reg [(4'ha):(1'h0)] reg778 = (1'h0);
  reg [(3'h4):(1'h0)] forvar770 = (1'h0);
  reg [(3'h5):(1'h0)] reg769 = (1'h0);
  reg [(4'he):(1'h0)] reg777 = (1'h0);
  reg [(2'h2):(1'h0)] reg776 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg775 = (1'h0);
  reg [(2'h2):(1'h0)] reg774 = (1'h0);
  reg [(2'h2):(1'h0)] reg773 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg772 = (1'h0);
  reg [(4'hd):(1'h0)] reg771 = (1'h0);
  reg [(3'h7):(1'h0)] reg770 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar769 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg765 = (1'h0);
  reg [(4'h8):(1'h0)] reg768 = (1'h0);
  reg [(2'h2):(1'h0)] reg767 = (1'h0);
  reg [(5'h10):(1'h0)] reg766 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar765 = (1'h0);
  reg signed [(4'he):(1'h0)] reg764 = (1'h0);
  reg [(3'h6):(1'h0)] reg763 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar762 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg761 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg760 = (1'h0);
  reg [(3'h4):(1'h0)] reg759 = (1'h0);
  reg [(4'he):(1'h0)] reg758 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar757 = (1'h0);
  reg [(4'ha):(1'h0)] reg756 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg755 = (1'h0);
  reg [(3'h6):(1'h0)] reg754 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg753 = (1'h0);
  reg [(3'h7):(1'h0)] reg752 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg751 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar750 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg749 = (1'h0);
  reg [(4'h9):(1'h0)] reg748 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg747 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg746 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg745 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar741 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar736 = (1'h0);
  reg [(2'h3):(1'h0)] reg744 = (1'h0);
  reg [(4'he):(1'h0)] reg743 = (1'h0);
  reg [(4'h8):(1'h0)] reg742 = (1'h0);
  reg [(3'h6):(1'h0)] reg741 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg740 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg739 = (1'h0);
  reg [(3'h7):(1'h0)] reg738 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg737 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg736 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg735 = (1'h0);
  reg [(4'he):(1'h0)] reg734 = (1'h0);
  reg [(3'h5):(1'h0)] reg733 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg732 = (1'h0);
  reg [(4'hb):(1'h0)] reg731 = (1'h0);
  reg [(4'hf):(1'h0)] reg730 = (1'h0);
  reg [(4'h8):(1'h0)] reg729 = (1'h0);
  reg [(4'hb):(1'h0)] forvar728 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg727 = (1'h0);
  reg [(3'h4):(1'h0)] reg726 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg725 = (1'h0);
  reg [(4'hb):(1'h0)] reg724 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar723 = (1'h0);
  reg [(4'hf):(1'h0)] forvar722 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg721 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg720 = (1'h0);
  reg [(4'h9):(1'h0)] reg719 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg718 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg717 = (1'h0);
  reg [(4'he):(1'h0)] reg716 = (1'h0);
  reg [(4'hb):(1'h0)] reg715 = (1'h0);
  reg [(3'h6):(1'h0)] reg714 = (1'h0);
  reg [(3'h7):(1'h0)] forvar713 = (1'h0);
  reg [(4'h8):(1'h0)] reg712 = (1'h0);
  reg [(3'h5):(1'h0)] reg711 = (1'h0);
  reg [(4'hd):(1'h0)] reg710 = (1'h0);
  reg [(3'h5):(1'h0)] reg709 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg708 = (1'h0);
  reg [(4'hf):(1'h0)] forvar707 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg706 = (1'h0);
  reg [(4'he):(1'h0)] forvar705 = (1'h0);
  reg [(5'h10):(1'h0)] reg704 = (1'h0);
  reg signed [(4'he):(1'h0)] reg703 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg702 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg701 = (1'h0);
  reg [(4'hd):(1'h0)] reg700 = (1'h0);
  reg [(3'h5):(1'h0)] forvar699 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg698 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg697 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar696 = (1'h0);
  reg [(2'h3):(1'h0)] forvar695 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar694 = (1'h0);
  reg [(4'hb):(1'h0)] reg693 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg692 = (1'h0);
  reg [(2'h2):(1'h0)] reg691 = (1'h0);
  reg [(3'h7):(1'h0)] forvar690 = (1'h0);
  reg [(2'h3):(1'h0)] reg689 = (1'h0);
  reg [(4'h9):(1'h0)] reg688 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar687 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar686 = (1'h0);
  reg [(3'h5):(1'h0)] reg681 = (1'h0);
  reg [(3'h5):(1'h0)] reg685 = (1'h0);
  reg [(4'hd):(1'h0)] reg684 = (1'h0);
  reg signed [(4'he):(1'h0)] reg683 = (1'h0);
  reg [(2'h2):(1'h0)] reg682 = (1'h0);
  reg [(3'h6):(1'h0)] forvar681 = (1'h0);
  reg [(4'hb):(1'h0)] reg680 = (1'h0);
  reg [(4'h9):(1'h0)] reg679 = (1'h0);
  reg [(4'h9):(1'h0)] reg678 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg677 = (1'h0);
  reg [(4'hb):(1'h0)] forvar676 = (1'h0);
  reg [(4'he):(1'h0)] forvar670 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar659 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar653 = (1'h0);
  reg [(4'he):(1'h0)] forvar645 = (1'h0);
  reg [(2'h3):(1'h0)] forvar648 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar654 = (1'h0);
  reg [(3'h7):(1'h0)] forvar652 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg650 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg649 = (1'h0);
  reg [(2'h2):(1'h0)] forvar641 = (1'h0);
  reg [(3'h6):(1'h0)] forvar639 = (1'h0);
  reg [(4'h9):(1'h0)] forvar631 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg629 = (1'h0);
  reg [(4'hc):(1'h0)] reg628 = (1'h0);
  reg [(4'hd):(1'h0)] forvar627 = (1'h0);
  reg [(4'he):(1'h0)] reg623 = (1'h0);
  reg [(4'ha):(1'h0)] reg622 = (1'h0);
  reg [(3'h7):(1'h0)] forvar620 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar617 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg618 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar615 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar612 = (1'h0);
  reg [(4'hc):(1'h0)] forvar607 = (1'h0);
  reg [(4'hc):(1'h0)] forvar606 = (1'h0);
  reg [(4'ha):(1'h0)] forvar673 = (1'h0);
  reg [(3'h7):(1'h0)] forvar669 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar665 = (1'h0);
  reg [(2'h2):(1'h0)] reg664 = (1'h0);
  reg [(5'h10):(1'h0)] forvar660 = (1'h0);
  reg [(3'h6):(1'h0)] reg672 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar671 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg666 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg675 = (1'h0);
  reg [(2'h3):(1'h0)] reg674 = (1'h0);
  reg [(4'ha):(1'h0)] reg673 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar672 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg671 = (1'h0);
  reg [(4'hb):(1'h0)] reg670 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg669 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg668 = (1'h0);
  reg [(4'hf):(1'h0)] reg667 = (1'h0);
  reg [(4'h8):(1'h0)] forvar666 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg665 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar664 = (1'h0);
  reg [(2'h3):(1'h0)] reg663 = (1'h0);
  reg [(4'hf):(1'h0)] reg662 = (1'h0);
  reg [(3'h5):(1'h0)] forvar661 = (1'h0);
  reg [(3'h6):(1'h0)] reg660 = (1'h0);
  reg signed [(4'he):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg658 = (1'h0);
  reg [(2'h2):(1'h0)] reg657 = (1'h0);
  reg [(4'h8):(1'h0)] reg656 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg655 = (1'h0);
  reg [(4'hb):(1'h0)] reg654 = (1'h0);
  reg [(4'h9):(1'h0)] reg653 = (1'h0);
  reg [(2'h2):(1'h0)] reg652 = (1'h0);
  reg [(2'h2):(1'h0)] reg651 = (1'h0);
  reg [(5'h10):(1'h0)] forvar650 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar649 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg648 = (1'h0);
  reg [(4'hb):(1'h0)] reg647 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar644 = (1'h0);
  reg [(4'he):(1'h0)] forvar642 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg638 = (1'h0);
  reg [(4'hf):(1'h0)] reg637 = (1'h0);
  reg [(4'hc):(1'h0)] reg646 = (1'h0);
  reg [(5'h10):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg644 = (1'h0);
  reg [(4'ha):(1'h0)] reg643 = (1'h0);
  reg [(5'h10):(1'h0)] reg642 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg641 = (1'h0);
  reg [(4'h8):(1'h0)] reg640 = (1'h0);
  reg [(3'h6):(1'h0)] reg639 = (1'h0);
  reg [(4'hc):(1'h0)] forvar638 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar637 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg635 = (1'h0);
  reg [(2'h2):(1'h0)] reg634 = (1'h0);
  reg [(5'h10):(1'h0)] reg633 = (1'h0);
  reg [(3'h5):(1'h0)] reg632 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg631 = (1'h0);
  reg [(2'h2):(1'h0)] reg630 = (1'h0);
  reg [(4'ha):(1'h0)] forvar629 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar628 = (1'h0);
  reg [(3'h5):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg626 = (1'h0);
  reg [(4'hf):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg624 = (1'h0);
  reg [(4'hc):(1'h0)] forvar623 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar622 = (1'h0);
  reg [(3'h7):(1'h0)] reg621 = (1'h0);
  reg [(4'hc):(1'h0)] reg620 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg619 = (1'h0);
  reg [(5'h10):(1'h0)] forvar618 = (1'h0);
  reg [(4'hf):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg616 = (1'h0);
  reg [(3'h5):(1'h0)] reg615 = (1'h0);
  reg [(5'h10):(1'h0)] reg614 = (1'h0);
  reg [(4'he):(1'h0)] reg613 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg612 = (1'h0);
  reg [(3'h6):(1'h0)] forvar611 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar610 = (1'h0);
  reg [(2'h2):(1'h0)] reg611 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar608 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg610 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg609 = (1'h0);
  reg [(4'hc):(1'h0)] reg608 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg607 = (1'h0);
  reg [(3'h4):(1'h0)] reg606 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire605;
  assign y = {wire782,
                 wire781,
                 wire780,
                 wire779,
                 reg778,
                 forvar770,
                 reg769,
                 reg777,
                 reg776,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 forvar769,
                 reg765,
                 reg768,
                 reg767,
                 reg766,
                 forvar765,
                 reg764,
                 reg763,
                 forvar762,
                 reg761,
                 reg760,
                 reg759,
                 reg758,
                 forvar757,
                 reg756,
                 reg755,
                 reg754,
                 reg753,
                 reg752,
                 reg751,
                 forvar750,
                 reg749,
                 reg748,
                 reg747,
                 reg746,
                 reg745,
                 forvar741,
                 forvar736,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 reg740,
                 reg739,
                 reg738,
                 reg737,
                 reg736,
                 reg735,
                 reg734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 reg729,
                 forvar728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 forvar723,
                 forvar722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 forvar713,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 reg708,
                 forvar707,
                 reg706,
                 forvar705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg700,
                 forvar699,
                 reg698,
                 reg697,
                 forvar696,
                 forvar695,
                 forvar694,
                 reg693,
                 reg692,
                 reg691,
                 forvar690,
                 reg689,
                 reg688,
                 forvar687,
                 forvar686,
                 reg681,
                 reg685,
                 reg684,
                 reg683,
                 reg682,
                 forvar681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 forvar676,
                 forvar670,
                 forvar659,
                 forvar653,
                 forvar645,
                 forvar648,
                 forvar654,
                 forvar652,
                 reg650,
                 reg649,
                 forvar641,
                 forvar639,
                 forvar631,
                 reg629,
                 reg628,
                 forvar627,
                 reg623,
                 reg622,
                 forvar620,
                 forvar617,
                 reg618,
                 forvar615,
                 forvar612,
                 forvar607,
                 forvar606,
                 forvar673,
                 forvar669,
                 forvar665,
                 reg664,
                 forvar660,
                 reg672,
                 forvar671,
                 reg666,
                 reg675,
                 reg674,
                 reg673,
                 forvar672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 reg667,
                 forvar666,
                 reg665,
                 forvar664,
                 reg663,
                 reg662,
                 forvar661,
                 reg660,
                 reg659,
                 reg658,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 reg651,
                 forvar650,
                 forvar649,
                 reg648,
                 reg647,
                 forvar644,
                 forvar642,
                 reg638,
                 reg637,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg640,
                 reg639,
                 forvar638,
                 forvar637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 forvar629,
                 forvar628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 forvar623,
                 forvar622,
                 reg621,
                 reg620,
                 reg619,
                 forvar618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg613,
                 reg612,
                 forvar611,
                 forvar610,
                 reg611,
                 forvar608,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 reg606,
                 wire605,
                 (1'h0)};
  assign wire605 = $signed($unsigned({((8'had) ^ wire604)}));
  always
    @(posedge clk) begin
      if ((8'hb0))
        begin
          if ({(~|((^~(8'ha9)) << (wire601 ? wire602 : wire602)))})
            begin
              if (wire605[(4'ha):(2'h2)])
                begin
                  if ((~^wire605[(4'hc):(2'h2)]))
                    begin
                      reg606 <= wire603[(3'h4):(2'h3)];
                      reg607 <= (wire602 + wire605[(3'h6):(3'h5)]);
                      reg608 <= $signed((reg607 ?
                          {wire603[(1'h0):(1'h0)]} : $unsigned(wire602[(4'he):(3'h4)])));
                      reg609 <= $signed(wire604);
                    end
                  else
                    begin
                      reg606 <= ((~^(wire603 ?
                              reg607[(1'h1):(1'h0)] : (^~(8'h9e)))) ?
                          (reg607 > (&$unsigned(wire604))) : ((^{reg606}) ?
                              wire605[(3'h7):(2'h2)] : $signed((|wire601))));
                    end
                  reg610 <= ((^{$signed(reg607)}) << $unsigned({wire601[(3'h7):(2'h2)]}));
                end
              else
                begin
                  if (reg607[(2'h2):(1'h1)])
                    begin
                      reg606 <= wire605;
                      reg607 <= (-reg606);
                    end
                  else
                    begin
                      reg606 <= reg606;
                      reg607 <= {wire603};
                    end
                  for (forvar608 = (1'h0); (forvar608 < (2'h3)); forvar608 = (forvar608 + (1'h1)))
                    begin
                      reg609 <= $signed(($signed($unsigned(wire603)) ?
                          $signed((reg606 <= wire605)) : $signed((reg609 ?
                              reg608 : wire605))));
                    end
                  reg610 <= $signed(($unsigned((!reg608)) ?
                      $unsigned($signed(reg608)) : $unsigned((reg609 ?
                          (8'hab) : reg608))));
                end
              reg611 <= $unsigned($unsigned(({reg609} * (reg608 ?
                  wire604 : reg609))));
            end
          else
            begin
              if ({$signed((^~wire604[(3'h6):(2'h2)]))})
                begin
                  reg606 <= reg606;
                  if ((((-(!wire604)) > $unsigned(reg610)) ?
                      $unsigned(((reg609 <<< wire603) ?
                          $signed(wire604) : (~|reg609))) : reg607[(3'h6):(3'h6)]))
                    begin
                      reg607 <= wire604;
                      reg608 <= reg610;
                      reg609 <= (~^(wire602 ?
                          ((^reg609) ?
                              reg607[(1'h1):(1'h0)] : (wire602 << reg607)) : $unsigned((forvar608 ?
                              reg606 : wire601))));
                    end
                  else
                    begin
                      reg607 <= reg610[(1'h0):(1'h0)];
                      reg608 <= (8'hae);
                      reg609 <= ($unsigned($signed((~reg608))) ^ $unsigned((((8'hb8) ?
                          wire605 : wire603) << (wire603 ?
                          (8'ha8) : wire605))));
                    end
                end
              else
                begin
                  if (wire604)
                    begin
                      reg606 <= $unsigned(((~|$signed(wire605)) ?
                          ($unsigned((8'h9d)) ?
                              reg607[(2'h2):(1'h1)] : $unsigned(reg608)) : reg606));
                      reg607 <= (!((&reg610) ?
                          $signed({wire603}) : {reg608[(2'h2):(1'h0)]}));
                    end
                  else
                    begin
                      reg606 <= ((8'h9e) && (($signed(forvar608) ?
                              reg606 : (reg609 >= reg607)) ?
                          (~|(wire601 ?
                              reg611 : wire601)) : $signed((~|(8'hae)))));
                      reg607 <= ({{(reg610 <<< reg611)}} * (wire603[(2'h3):(2'h3)] ?
                          reg610[(1'h1):(1'h1)] : $unsigned(reg606[(1'h0):(1'h0)])));
                      reg608 <= ((((reg610 ? wire603 : reg607) ?
                              $unsigned(reg606) : (forvar608 ?
                                  wire603 : wire605)) + ({(8'hb5)} ?
                              (wire601 ? wire602 : reg607) : {reg606})) ?
                          (!(|reg606)) : ((reg611[(1'h1):(1'h0)] ?
                              {(8'hb3)} : wire603[(2'h3):(2'h2)]) == (-(reg610 ?
                              reg606 : reg610))));
                      reg609 <= (~(+($signed(wire603) > (+wire603))));
                    end
                end
              for (forvar610 = (1'h0); (forvar610 < (1'h1)); forvar610 = (forvar610 + (1'h1)))
                begin
                  for (forvar611 = (1'h0); (forvar611 < (1'h0)); forvar611 = (forvar611 + (1'h1)))
                    begin
                      reg612 <= (~^$unsigned(($signed(wire602) ?
                          $unsigned(reg609) : $unsigned(reg610))));
                      reg613 <= wire603;
                      reg614 <= (((forvar608 ?
                                  (reg610 - forvar610) : $unsigned(forvar611)) ?
                              $signed((^reg611)) : wire601) ?
                          (8'h9d) : {$unsigned((reg613 >> reg606))});
                      reg615 <= (&(((reg611 == reg612) ?
                              $unsigned(forvar610) : $unsigned(reg611)) ?
                          reg613[(4'ha):(1'h1)] : reg608[(2'h2):(1'h0)]));
                    end
                  reg616 <= (wire602 < $unsigned($signed(reg612)));
                  reg617 <= (&wire605[(4'hf):(3'h5)]);
                  for (forvar618 = (1'h0); (forvar618 < (2'h2)); forvar618 = (forvar618 + (1'h1)))
                    begin
                      reg619 <= $signed((~^$signed((reg615 ?
                          reg615 : forvar608))));
                      reg620 <= reg612;
                      reg621 <= wire602[(4'h8):(2'h3)];
                    end
                end
            end
          for (forvar622 = (1'h0); (forvar622 < (1'h1)); forvar622 = (forvar622 + (1'h1)))
            begin
              if ($unsigned(((+forvar622) ? (^~(&(8'hac))) : (8'haf))))
                begin
                  for (forvar623 = (1'h0); (forvar623 < (2'h2)); forvar623 = (forvar623 + (1'h1)))
                    begin
                      reg624 <= $signed($unsigned($signed((reg617 >>> (8'ha6)))));
                      reg625 <= $signed(wire605);
                      reg626 <= $signed((+$unsigned(wire603[(3'h4):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar623 = (1'h0); (forvar623 < (1'h0)); forvar623 = (forvar623 + (1'h1)))
                    begin
                      reg624 <= wire602;
                    end
                  reg625 <= $unsigned((^~$unsigned(reg613)));
                  if ((+wire603[(2'h2):(2'h2)]))
                    begin
                      reg626 <= (({(reg610 ? forvar623 : reg624)} ?
                              reg609[(3'h5):(1'h0)] : forvar623[(1'h1):(1'h1)]) ?
                          (($signed(reg608) ?
                              (-forvar618) : (forvar608 ?
                                  reg621 : reg625)) & $signed(reg613)) : $unsigned(((^wire603) ~^ $unsigned(forvar618))));
                      reg627 <= $unsigned(reg624[(4'he):(4'h9)]);
                    end
                  else
                    begin
                      reg626 <= ((~^(~|(-reg606))) ?
                          ((!forvar611[(3'h5):(1'h0)]) * $unsigned((^reg613))) : $signed(((reg626 ?
                              wire603 : reg612) ^~ (reg610 >>> (8'hb9)))));
                      reg627 <= $signed($signed($unsigned($unsigned(reg617))));
                    end
                end
              for (forvar628 = (1'h0); (forvar628 < (1'h1)); forvar628 = (forvar628 + (1'h1)))
                begin
                  for (forvar629 = (1'h0); (forvar629 < (1'h0)); forvar629 = (forvar629 + (1'h1)))
                    begin
                      reg630 <= forvar611[(2'h2):(1'h1)];
                      reg631 <= reg624[(3'h6):(3'h4)];
                    end
                  reg632 <= (^($signed((reg627 && reg615)) ?
                      $unsigned($signed(reg615)) : ($unsigned((8'hb0)) >>> (reg611 ?
                          reg617 : (8'hb3)))));
                  reg633 <= (reg626 ?
                      ($signed(((8'haf) > wire604)) >> $signed(reg610[(1'h1):(1'h0)])) : $unsigned($unsigned((-reg631))));
                  if ((|(($signed(reg606) || reg621[(3'h5):(3'h5)]) || ((reg627 ?
                      reg624 : reg613) + ((8'ha0) ? (8'h9f) : forvar610)))))
                    begin
                      reg634 <= reg627[(2'h3):(2'h2)];
                      reg635 <= {$unsigned({$signed(forvar628)})};
                      reg636 <= ($unsigned($unsigned($unsigned(reg608))) >>> reg614[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg634 <= (^~reg610);
                      reg635 <= reg625[(4'h9):(3'h6)];
                      reg636 <= $unsigned(reg620);
                    end
                end
            end
          if ((($signed((forvar610 ~^ reg619)) < wire604) ?
              $unsigned($signed(forvar610[(1'h0):(1'h0)])) : (reg631[(1'h0):(1'h0)] ?
                  $unsigned($signed(forvar608)) : ($signed(reg619) << reg630))))
            begin
              for (forvar637 = (1'h0); (forvar637 < (1'h1)); forvar637 = (forvar637 + (1'h1)))
                begin
                  for (forvar638 = (1'h0); (forvar638 < (2'h2)); forvar638 = (forvar638 + (1'h1)))
                    begin
                      reg639 <= forvar611[(2'h2):(1'h0)];
                      reg640 <= (&($signed((!reg613)) | forvar628[(1'h0):(1'h0)]));
                      reg641 <= (~^reg624);
                    end
                  reg642 <= wire601;
                  reg643 <= {$signed($unsigned({(8'had)}))};
                  if ((|reg631[(3'h5):(2'h2)]))
                    begin
                      reg644 <= reg608;
                    end
                  else
                    begin
                      reg644 <= forvar622;
                      reg645 <= (reg643 ? forvar608[(1'h1):(1'h0)] : reg617);
                      reg646 <= (^$unsigned({forvar611[(1'h1):(1'h1)]}));
                    end
                end
            end
          else
            begin
              reg637 <= reg646;
              if ((^~((~$unsigned(reg619)) && $unsigned($signed((8'hae))))))
                begin
                  if (reg612)
                    begin
                      reg638 <= reg621;
                      reg639 <= $signed(reg636[(2'h3):(2'h2)]);
                      reg640 <= ((reg640[(4'h8):(3'h4)] <<< ((reg640 - reg627) ?
                              (forvar623 << forvar637) : (reg608 && reg625))) ?
                          (~(reg624[(4'h9):(1'h0)] ?
                              (forvar637 ?
                                  wire602 : reg645) : wire604[(4'h8):(3'h4)])) : ({$unsigned(reg613)} ?
                              (~&((8'hb4) <<< forvar610)) : reg615));
                      reg641 <= reg626[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg638 <= $unsigned($unsigned((reg608[(3'h5):(2'h2)] ?
                          (wire601 ? reg639 : reg621) : ((8'hb3) ?
                              forvar638 : forvar610))));
                      reg639 <= reg625[(4'h8):(1'h0)];
                      reg640 <= $signed((((reg638 ? reg639 : (8'hb8)) ?
                              (~forvar637) : (forvar611 | (8'ha0))) ?
                          reg630 : $unsigned($signed(forvar637))));
                    end
                  for (forvar642 = (1'h0); (forvar642 < (1'h1)); forvar642 = (forvar642 + (1'h1)))
                    begin
                      reg643 <= reg621[(3'h6):(3'h5)];
                    end
                  for (forvar644 = (1'h0); (forvar644 < (2'h2)); forvar644 = (forvar644 + (1'h1)))
                    begin
                      reg645 <= ($signed($unsigned(forvar628[(4'h8):(4'h8)])) ?
                          $signed((~|(reg627 ?
                              (8'hb2) : wire605))) : (-$unsigned((|wire602))));
                      reg646 <= $signed($signed(($unsigned(reg638) ?
                          (^reg609) : $unsigned(reg607))));
                      reg647 <= wire601[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  if ({wire603})
                    begin
                      reg638 <= {{$unsigned((reg612 * reg640))}};
                      reg639 <= ($signed(reg631) ^ (((~reg646) ?
                          $unsigned(forvar629) : (wire605 ?
                              reg641 : reg626)) << ((8'ha5) != $unsigned(reg635))));
                    end
                  else
                    begin
                      reg638 <= reg627;
                      reg639 <= (8'h9e);
                      reg640 <= ((($signed(reg636) ?
                              $signed(forvar642) : (forvar618 >> reg645)) >> ((~^forvar618) >> $unsigned(forvar629))) ?
                          ($unsigned((reg642 ? reg639 : reg612)) ?
                              $unsigned({(8'hb1)}) : reg635) : $unsigned((~|reg616)));
                      reg641 <= (!(~&$unsigned((-reg609))));
                    end
                  for (forvar642 = (1'h0); (forvar642 < (1'h0)); forvar642 = (forvar642 + (1'h1)))
                    begin
                      reg643 <= reg615;
                      reg644 <= $signed($unsigned((+reg621[(1'h1):(1'h0)])));
                    end
                  if (($signed(($signed(forvar623) ?
                      $signed((8'h9c)) : $signed(reg619))) >>> $unsigned({(reg644 ?
                          reg614 : reg630)})))
                    begin
                      reg645 <= reg625;
                    end
                  else
                    begin
                      reg645 <= reg642;
                    end
                  if ((($unsigned(reg631) ?
                      $unsigned((reg616 ?
                          (8'hb9) : reg613)) : $unsigned(forvar608)) - (|{$unsigned(reg635)})))
                    begin
                      reg646 <= $signed({(reg621 ?
                              ((8'hb4) ? reg624 : forvar644) : (forvar608 ?
                                  (8'hb4) : reg609))});
                    end
                  else
                    begin
                      reg646 <= reg606[(1'h0):(1'h0)];
                      reg647 <= {((reg624 ^~ $unsigned(forvar610)) ?
                              ((reg624 ? (8'hb0) : (8'haf)) ?
                                  (reg644 ? reg642 : reg620) : ((8'hb5) ?
                                      reg611 : reg617)) : $signed($unsigned(reg620)))};
                      reg648 <= $signed({(|{wire602})});
                    end
                end
              for (forvar649 = (1'h0); (forvar649 < (2'h3)); forvar649 = (forvar649 + (1'h1)))
                begin
                  for (forvar650 = (1'h0); (forvar650 < (2'h2)); forvar650 = (forvar650 + (1'h1)))
                    begin
                      reg651 <= (~forvar644);
                      reg652 <= forvar644;
                      reg653 <= reg647[(4'ha):(3'h6)];
                    end
                  if (forvar638)
                    begin
                      reg654 <= (+(~&forvar649));
                      reg655 <= reg608;
                      reg656 <= $unsigned(reg638[(4'ha):(3'h7)]);
                      reg657 <= ($unsigned((~^(reg641 == reg610))) ?
                          (~^(~&(reg625 ? reg654 : reg644))) : ((~(reg645 ?
                              reg619 : reg612)) || $unsigned(reg641)));
                    end
                  else
                    begin
                      reg654 <= (forvar650[(4'hb):(4'hb)] ?
                          (~|($unsigned((8'hb1)) ?
                              reg632[(2'h2):(1'h0)] : reg631[(1'h0):(1'h0)])) : (reg640[(1'h0):(1'h0)] ?
                              reg617 : $unsigned($unsigned(reg652))));
                      reg655 <= (reg640 < (reg608[(3'h6):(2'h2)] ?
                          $signed(reg632[(1'h0):(1'h0)]) : reg608[(1'h1):(1'h0)]));
                      reg656 <= (forvar611[(3'h4):(1'h1)] ?
                          (wire603[(2'h2):(1'h1)] ^~ {$unsigned(reg620)}) : forvar650);
                    end
                end
              if (reg633[(4'hc):(4'h8)])
                begin
                  if (($signed(reg645[(4'hf):(4'h8)]) ?
                      ($unsigned((^~reg654)) + $signed(reg647[(2'h2):(1'h1)])) : $signed($signed($signed(reg657)))))
                    begin
                      reg658 <= ((&$unsigned((reg627 == reg652))) ?
                          (reg644 ?
                              (+forvar650) : $unsigned((~|forvar611))) : {wire605});
                      reg659 <= reg616[(4'hb):(4'h8)];
                    end
                  else
                    begin
                      reg658 <= ((~(8'hb5)) >= {((~&reg625) == (forvar637 ?
                              wire604 : (8'had)))});
                    end
                end
              else
                begin
                  reg658 <= $unsigned($unsigned($signed((reg632 * forvar628))));
                end
            end
          if ($unsigned(reg659))
            begin
              reg660 <= ({(reg610 >> (~&wire605))} ?
                  $signed(reg657) : (|(~^$unsigned((8'ha0)))));
              for (forvar661 = (1'h0); (forvar661 < (1'h0)); forvar661 = (forvar661 + (1'h1)))
                begin
                  if ((~&forvar650))
                    begin
                      reg662 <= (8'ha3);
                      reg663 <= $unsigned((|((^reg642) ?
                          (reg643 || reg648) : $signed(reg621))));
                    end
                  else
                    begin
                      reg662 <= (^~(((~|reg636) ?
                          (8'ha7) : (~reg615)) ^~ {(reg657 >> reg655)}));
                      reg663 <= (($unsigned({(8'ha4)}) == reg611) - $unsigned(((~|reg660) ?
                          (reg657 ? reg654 : reg647) : (^reg646))));
                    end
                  for (forvar664 = (1'h0); (forvar664 < (1'h1)); forvar664 = (forvar664 + (1'h1)))
                    begin
                      reg665 <= (!reg625);
                    end
                end
              if ($unsigned(($signed((^forvar629)) <<< ($signed(forvar611) ?
                  reg619 : (forvar661 | reg655)))))
                begin
                  for (forvar666 = (1'h0); (forvar666 < (2'h2)); forvar666 = (forvar666 + (1'h1)))
                    begin
                      reg667 <= reg619[(3'h7):(3'h5)];
                      reg668 <= forvar642;
                      reg669 <= {reg615};
                      reg670 <= $signed({reg660});
                    end
                  reg671 <= reg660;
                  for (forvar672 = (1'h0); (forvar672 < (1'h0)); forvar672 = (forvar672 + (1'h1)))
                    begin
                      reg673 <= reg665[(4'h9):(3'h7)];
                      reg674 <= $signed($signed(wire603[(2'h3):(1'h0)]));
                      reg675 <= ((-(&(^(8'hb0)))) << $signed(reg658));
                    end
                end
              else
                begin
                  reg666 <= (reg670 ? forvar644[(1'h1):(1'h0)] : (~reg627));
                  if (($signed(({reg620} ?
                      $signed((8'ha5)) : ((8'haf) != forvar661))) || $unsigned((reg639[(2'h2):(1'h1)] ?
                      (reg670 ^~ reg611) : {reg624}))))
                    begin
                      reg667 <= reg653;
                    end
                  else
                    begin
                      reg667 <= $signed(reg632[(3'h4):(1'h0)]);
                      reg668 <= (8'ha3);
                      reg669 <= $unsigned({((reg639 ? forvar628 : reg648) ?
                              reg657[(1'h0):(1'h0)] : $signed(reg646))});
                      reg670 <= (({(forvar628 ?
                              reg633 : reg626)} <<< $unsigned((reg675 >>> forvar672))) <= (^($signed(reg671) ^~ reg674[(1'h0):(1'h0)])));
                    end
                  for (forvar671 = (1'h0); (forvar671 < (1'h0)); forvar671 = (forvar671 + (1'h1)))
                    begin
                      reg672 <= (-(~^$unsigned({forvar666})));
                      reg673 <= (~^(((&reg665) ?
                          $signed(reg631) : $unsigned(forvar628)) == forvar622));
                      reg674 <= ((8'hb5) >>> (&{(^reg646)}));
                      reg675 <= $unsigned((|(^~reg665[(4'ha):(3'h7)])));
                    end
                end
            end
          else
            begin
              for (forvar660 = (1'h0); (forvar660 < (1'h0)); forvar660 = (forvar660 + (1'h1)))
                begin
                  for (forvar661 = (1'h0); (forvar661 < (2'h2)); forvar661 = (forvar661 + (1'h1)))
                    begin
                      reg662 <= (!reg611[(2'h2):(2'h2)]);
                      reg663 <= (~^((8'hb5) & ((forvar650 < forvar623) ?
                          reg636 : {(8'h9f)})));
                      reg664 <= $signed(reg669);
                    end
                end
              for (forvar665 = (1'h0); (forvar665 < (2'h3)); forvar665 = (forvar665 + (1'h1)))
                begin
                  for (forvar666 = (1'h0); (forvar666 < (2'h2)); forvar666 = (forvar666 + (1'h1)))
                    begin
                      reg667 <= $unsigned((+(+$signed(reg636))));
                      reg668 <= {(!reg653[(3'h4):(1'h0)])};
                    end
                  for (forvar669 = (1'h0); (forvar669 < (1'h0)); forvar669 = (forvar669 + (1'h1)))
                    begin
                      reg670 <= ($signed(($signed((8'hba)) ?
                          (reg673 ?
                              reg624 : reg668) : (forvar629 ^~ (8'hb4)))) && reg638[(2'h2):(1'h1)]);
                      reg671 <= forvar664[(3'h4):(2'h3)];
                    end
                  reg672 <= {(reg666[(1'h0):(1'h0)] ?
                          $unsigned($unsigned(reg634)) : $unsigned(reg660[(3'h5):(1'h1)]))};
                  for (forvar673 = (1'h0); (forvar673 < (2'h3)); forvar673 = (forvar673 + (1'h1)))
                    begin
                      reg674 <= $unsigned({$signed((reg633 ^~ reg641))});
                    end
                end
            end
        end
      else
        begin
          for (forvar606 = (1'h0); (forvar606 < (2'h3)); forvar606 = (forvar606 + (1'h1)))
            begin
              if (($unsigned(reg656) >= {(reg655[(1'h1):(1'h0)] ?
                      (|reg675) : reg660[(3'h5):(3'h5)])}))
                begin
                  for (forvar607 = (1'h0); (forvar607 < (2'h3)); forvar607 = (forvar607 + (1'h1)))
                    begin
                      reg608 <= reg634;
                      reg609 <= $signed(wire604[(4'hf):(3'h7)]);
                    end
                  for (forvar610 = (1'h0); (forvar610 < (2'h2)); forvar610 = (forvar610 + (1'h1)))
                    begin
                      reg611 <= ($signed((reg668 << (forvar669 << (8'hac)))) && $unsigned($unsigned(reg647[(1'h1):(1'h0)])));
                    end
                  for (forvar612 = (1'h0); (forvar612 < (2'h3)); forvar612 = (forvar612 + (1'h1)))
                    begin
                      reg613 <= $signed((~($signed(reg615) >>> forvar606[(3'h5):(1'h1)])));
                      reg614 <= $unsigned((reg666 ?
                          reg675[(4'ha):(3'h4)] : ($signed(reg627) ?
                              (8'ha2) : (reg625 ? forvar650 : reg664))));
                    end
                  for (forvar615 = (1'h0); (forvar615 < (1'h0)); forvar615 = (forvar615 + (1'h1)))
                    begin
                      reg616 <= reg613[(3'h7):(3'h7)];
                      reg617 <= (($signed((reg608 ?
                              reg667 : forvar607)) < {(reg624 ?
                                  forvar644 : reg636)}) ?
                          ($signed(((8'ha0) << reg652)) && ((reg653 | wire604) ^ (forvar669 ?
                              reg610 : forvar666))) : $signed($unsigned({reg648})));
                      reg618 <= ($unsigned((-(forvar610 ~^ forvar615))) - (^~((-reg621) ?
                          $unsigned(reg663) : (reg635 + reg645))));
                      reg619 <= ((($unsigned((8'hac)) & $unsigned(reg672)) ^ $unsigned($unsigned(reg657))) >>> (reg670[(3'h7):(3'h5)] ?
                          (&$signed(reg610)) : ($signed(reg630) ?
                              (forvar611 == forvar644) : $unsigned((8'ha6)))));
                    end
                end
              else
                begin
                  if (((($signed(forvar623) >= $signed(reg618)) && reg609[(2'h3):(2'h3)]) > $unsigned($unsigned((&reg665)))))
                    begin
                      reg607 <= (reg665 ? reg658 : reg630);
                      reg608 <= (8'hb4);
                      reg609 <= reg666;
                      reg610 <= $signed({($signed(reg647) < forvar622)});
                    end
                  else
                    begin
                      reg607 <= {($unsigned($unsigned(forvar637)) <<< ($unsigned(reg616) ?
                              (reg640 ? reg619 : forvar638) : (forvar615 ?
                                  (8'hb1) : reg642)))};
                      reg608 <= (~$signed((8'hb7)));
                    end
                  if ($unsigned(reg636[(4'hc):(2'h3)]))
                    begin
                      reg611 <= (~$unsigned((^reg613[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg611 <= ((8'hb2) ? reg675 : wire601[(2'h2):(1'h0)]);
                      reg612 <= forvar661[(2'h3):(2'h3)];
                      reg613 <= forvar644[(3'h5):(3'h4)];
                    end
                  if (reg630[(1'h0):(1'h0)])
                    begin
                      reg614 <= ((forvar642[(4'hb):(3'h4)] ?
                              $unsigned((forvar607 ?
                                  (8'hab) : (8'h9f))) : (!forvar669[(1'h0):(1'h0)])) ?
                          $unsigned($unsigned((forvar660 == (8'had)))) : (|$unsigned($unsigned(reg656))));
                      reg615 <= ($unsigned((8'h9f)) != reg651[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg614 <= reg653[(2'h2):(1'h0)];
                      reg615 <= {(~|$unsigned((reg645 || reg657)))};
                      reg616 <= wire604;
                    end
                  for (forvar617 = (1'h0); (forvar617 < (1'h1)); forvar617 = (forvar617 + (1'h1)))
                    begin
                      reg618 <= $signed($unsigned($signed(reg657[(1'h0):(1'h0)])));
                      reg619 <= (~^$unsigned((forvar664 ?
                          $unsigned(forvar629) : (reg640 > (8'hb4)))));
                    end
                end
              for (forvar620 = (1'h0); (forvar620 < (1'h0)); forvar620 = (forvar620 + (1'h1)))
                begin
                  if ({((~&(+forvar617)) ?
                          {(8'hb8)} : ({wire601} - $unsigned(reg647)))})
                    begin
                      reg621 <= $unsigned(forvar617[(1'h0):(1'h0)]);
                      reg622 <= ((((~&reg631) && (reg613 < reg606)) != (reg613 == $signed(wire603))) ?
                          (!reg614[(4'hc):(4'ha)]) : $signed($signed(reg624)));
                      reg623 <= (forvar669[(3'h4):(3'h4)] ?
                          $unsigned((~&$unsigned(reg614))) : $signed(wire602[(4'hd):(3'h4)]));
                      reg624 <= ((|$signed($signed(reg654))) * reg635[(4'h9):(4'h8)]);
                    end
                  else
                    begin
                      reg621 <= reg615[(3'h4):(1'h0)];
                      reg622 <= forvar650[(2'h2):(1'h1)];
                      reg623 <= $unsigned(reg652);
                      reg624 <= {$unsigned((~|(forvar644 ?
                              forvar622 : forvar671)))};
                    end
                  if ($signed(reg658[(4'hb):(1'h1)]))
                    begin
                      reg625 <= reg643;
                    end
                  else
                    begin
                      reg625 <= reg674;
                      reg626 <= (~|{$signed($unsigned((8'hb1)))});
                    end
                end
              if (((&(+(|forvar615))) + {(reg663 ^ (+wire605))}))
                begin
                  for (forvar627 = (1'h0); (forvar627 < (2'h2)); forvar627 = (forvar627 + (1'h1)))
                    begin
                      reg628 <= $signed(($signed((forvar638 >= forvar617)) > $signed({reg608})));
                      reg629 <= {(|$signed($unsigned(reg616)))};
                      reg630 <= $signed(($signed((reg673 ? reg634 : (8'hb3))) ?
                          ({forvar627} ?
                              reg668[(2'h3):(2'h3)] : (reg632 >= forvar618)) : $unsigned($signed(forvar644))));
                      reg631 <= reg666;
                    end
                  if ({reg642})
                    begin
                      reg632 <= $unsigned($signed(forvar665));
                      reg633 <= reg624;
                      reg634 <= (8'hb8);
                    end
                  else
                    begin
                      reg632 <= wire602;
                      reg633 <= $signed(forvar642);
                      reg634 <= reg607[(4'ha):(1'h1)];
                      reg635 <= $signed((~&({reg641} ~^ (reg657 || reg673))));
                    end
                end
              else
                begin
                  for (forvar627 = (1'h0); (forvar627 < (2'h3)); forvar627 = (forvar627 + (1'h1)))
                    begin
                      reg628 <= {reg674[(2'h3):(2'h3)]};
                      reg629 <= reg675[(1'h1):(1'h1)];
                      reg630 <= $unsigned(forvar612[(3'h5):(3'h5)]);
                    end
                  for (forvar631 = (1'h0); (forvar631 < (2'h2)); forvar631 = (forvar631 + (1'h1)))
                    begin
                      reg632 <= reg660;
                      reg633 <= reg671;
                      reg634 <= reg611[(2'h2):(1'h0)];
                      reg635 <= $signed($unsigned(reg662[(2'h3):(1'h1)]));
                    end
                  if ((&{(~&forvar642[(3'h7):(3'h7)])}))
                    begin
                      reg636 <= reg638[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg636 <= ($signed((((8'haf) ?
                              forvar649 : reg631) - forvar672)) ?
                          reg625 : ($unsigned($signed(forvar649)) ?
                              forvar660 : forvar627));
                    end
                  if (forvar618[(5'h10):(2'h3)])
                    begin
                      reg637 <= ($unsigned(forvar660) ?
                          {((reg607 != reg629) ?
                                  $signed(reg675) : $unsigned(reg632))} : (forvar617[(1'h1):(1'h0)] > {$signed(forvar637)}));
                      reg638 <= $unsigned(($unsigned((+(8'hba))) ?
                          (~(reg638 ^~ (8'ha0))) : $signed((8'ha5))));
                    end
                  else
                    begin
                      reg637 <= ({reg665} >= (reg655[(2'h2):(1'h0)] ?
                          forvar664 : $unsigned($signed((8'h9d)))));
                    end
                end
              for (forvar639 = (1'h0); (forvar639 < (1'h0)); forvar639 = (forvar639 + (1'h1)))
                begin
                  reg640 <= $unsigned((($signed((8'h9d)) ?
                      reg606[(1'h0):(1'h0)] : $signed(forvar665)) >>> ((8'ha2) << reg622)));
                  for (forvar641 = (1'h0); (forvar641 < (2'h3)); forvar641 = (forvar641 + (1'h1)))
                    begin
                      reg642 <= ($unsigned(reg634) > $unsigned($unsigned($unsigned(wire605))));
                      reg643 <= reg612;
                      reg644 <= $unsigned((&(forvar612 > (^reg615))));
                    end
                end
            end
          if ($unsigned($signed($unsigned($unsigned((8'ha6))))))
            begin
              if (reg637)
                begin
                  if ((~^(|$unsigned((forvar664 >> forvar644)))))
                    begin
                      reg645 <= ({$unsigned($unsigned(forvar622))} & $unsigned(({reg662} - (8'hb6))));
                      reg646 <= (($unsigned($unsigned(reg655)) ?
                          {(~^forvar610)} : (8'ha3)) ~^ $signed((^$unsigned(forvar644))));
                      reg647 <= $unsigned((forvar639 ?
                          $signed(reg641[(2'h3):(2'h2)]) : reg642[(4'hf):(2'h2)]));
                    end
                  else
                    begin
                      reg645 <= (-forvar608);
                      reg646 <= ($unsigned(((reg641 ?
                          forvar622 : forvar606) == (~|forvar660))) || {(reg644 > forvar649)});
                    end
                  if ((+((|(forvar629 ~^ reg635)) || (~&(~^reg665)))))
                    begin
                      reg648 <= reg632;
                      reg649 <= $unsigned($unsigned($signed($unsigned(reg653))));
                      reg650 <= (8'hab);
                      reg651 <= (!reg667[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg648 <= wire602[(3'h7):(3'h6)];
                    end
                  for (forvar652 = (1'h0); (forvar652 < (2'h3)); forvar652 = (forvar652 + (1'h1)))
                    begin
                      reg653 <= reg617;
                    end
                  for (forvar654 = (1'h0); (forvar654 < (1'h1)); forvar654 = (forvar654 + (1'h1)))
                    begin
                      reg655 <= (^$unsigned(($signed((8'h9e)) != {reg652})));
                      reg656 <= ($unsigned(reg667[(4'hd):(4'h9)]) ^ (reg674 ^ $unsigned(reg620)));
                      reg657 <= (~reg621);
                    end
                end
              else
                begin
                  if (((((&forvar665) ?
                          ((8'haa) > wire605) : (~|reg636)) + (~^(reg618 ?
                          reg671 : (8'hb4)))) ?
                      {forvar673} : wire605[(3'h5):(2'h2)]))
                    begin
                      reg645 <= (~^(((reg607 ? reg652 : reg656) ?
                          reg672[(3'h4):(1'h1)] : (forvar628 ?
                              (8'ha3) : reg641)) == forvar623[(3'h7):(3'h5)]));
                      reg646 <= $unsigned($signed({(8'ha5)}));
                    end
                  else
                    begin
                      reg645 <= reg640;
                      reg646 <= reg612;
                      reg647 <= (~&(-((reg639 ~^ reg655) ? reg643 : {reg618})));
                    end
                  for (forvar648 = (1'h0); (forvar648 < (1'h0)); forvar648 = (forvar648 + (1'h1)))
                    begin
                      reg649 <= (~|(!forvar661));
                    end
                  for (forvar650 = (1'h0); (forvar650 < (1'h1)); forvar650 = (forvar650 + (1'h1)))
                    begin
                      reg651 <= (^$signed(reg627));
                      reg652 <= ($signed(wire603[(2'h3):(2'h2)]) ?
                          $unsigned(((reg614 ?
                              reg665 : (8'hba)) << reg631)) : forvar661[(1'h1):(1'h1)]);
                      reg653 <= {(reg657[(1'h1):(1'h0)] && $unsigned((reg610 ?
                              reg656 : (8'had))))};
                      reg654 <= $signed({((~reg664) ^ reg673[(3'h5):(1'h0)])});
                    end
                  reg655 <= $signed($signed(forvar610[(2'h3):(1'h1)]));
                end
              reg658 <= (~&(&{(-reg640)}));
            end
          else
            begin
              if ((reg632 ?
                  (+reg667[(4'hf):(4'hb)]) : $signed((forvar649[(2'h3):(1'h1)] == (reg615 - reg609)))))
                begin
                  for (forvar645 = (1'h0); (forvar645 < (2'h3)); forvar645 = (forvar645 + (1'h1)))
                    begin
                      reg646 <= forvar628[(3'h4):(3'h4)];
                      reg647 <= (~&reg624[(2'h2):(2'h2)]);
                      reg648 <= (forvar641 ? forvar631 : (~|reg606));
                      reg649 <= ((^~$signed(((8'haf) <= reg631))) | (forvar652[(3'h6):(3'h4)] + (~reg653[(1'h1):(1'h1)])));
                    end
                  if (reg628)
                    begin
                      reg650 <= $unsigned(forvar639[(1'h0):(1'h0)]);
                      reg651 <= ((((~&reg614) ?
                              $signed(reg611) : wire602[(4'ha):(3'h6)]) ?
                          $signed($unsigned((8'hb1))) : reg674) ~^ ((reg656[(3'h4):(2'h2)] == {reg651}) ?
                          $signed((-reg672)) : ($unsigned((8'ha4)) && $unsigned(forvar669))));
                      reg652 <= ($unsigned($unsigned((reg652 > reg641))) & $signed($unsigned($unsigned(reg623))));
                    end
                  else
                    begin
                      reg650 <= forvar669[(2'h3):(1'h1)];
                      reg651 <= (reg625[(3'h5):(3'h4)] ?
                          $signed(reg630) : {reg624[(1'h1):(1'h0)]});
                      reg652 <= $unsigned({{$unsigned(reg653)}});
                    end
                  for (forvar653 = (1'h0); (forvar653 < (1'h0)); forvar653 = (forvar653 + (1'h1)))
                    begin
                      reg654 <= (-$signed(((^~wire601) <= (forvar629 | reg666))));
                      reg655 <= reg608;
                    end
                end
              else
                begin
                  for (forvar645 = (1'h0); (forvar645 < (2'h3)); forvar645 = (forvar645 + (1'h1)))
                    begin
                      reg646 <= $unsigned($signed(reg656));
                      reg647 <= $unsigned((((&forvar606) ?
                              $signed(forvar666) : $signed(forvar649)) ?
                          (+$unsigned(forvar628)) : reg606[(1'h0):(1'h0)]));
                      reg648 <= $signed((((reg669 <<< (8'hb0)) >> (8'ha7)) ?
                          reg615 : $unsigned($signed(reg657))));
                      reg649 <= $signed((|($signed(forvar607) + reg628)));
                    end
                  for (forvar650 = (1'h0); (forvar650 < (2'h3)); forvar650 = (forvar650 + (1'h1)))
                    begin
                      reg651 <= (^reg611[(1'h0):(1'h0)]);
                    end
                end
            end
          for (forvar659 = (1'h0); (forvar659 < (1'h1)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 <= reg668;
              for (forvar661 = (1'h0); (forvar661 < (2'h2)); forvar661 = (forvar661 + (1'h1)))
                begin
                  if (((($unsigned(reg668) ?
                      $signed(reg618) : (reg617 ?
                          reg609 : reg658)) ~^ (((8'hb2) ?
                      reg628 : reg632) << {reg649})) ^ $signed($signed(reg633[(4'he):(1'h1)]))))
                    begin
                      reg662 <= (reg674[(1'h0):(1'h0)] > (((forvar653 ^ forvar615) ~^ (8'hb4)) ?
                          (((8'ha4) * reg666) > forvar644) : $signed((^~(8'ha3)))));
                      reg663 <= (({(forvar660 ?
                              (8'ha8) : reg626)} == reg664[(1'h0):(1'h0)]) << (!($signed(reg647) ?
                          reg654[(1'h0):(1'h0)] : reg627[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg662 <= forvar618;
                      reg663 <= {((~$unsigned(reg610)) > (forvar637 <<< (forvar659 == reg628)))};
                      reg664 <= reg650[(2'h3):(1'h1)];
                      reg665 <= $unsigned(forvar639[(3'h5):(2'h2)]);
                    end
                  if ((8'hb2))
                    begin
                      reg666 <= (reg655[(1'h0):(1'h0)] ?
                          $signed((wire605[(3'h4):(3'h4)] ^ {(8'haf)})) : reg646);
                      reg667 <= forvar622[(3'h4):(2'h2)];
                      reg668 <= $signed($signed(reg611[(1'h0):(1'h0)]));
                      reg669 <= $signed((^$signed((reg672 || reg631))));
                    end
                  else
                    begin
                      reg666 <= ($signed((+$unsigned((8'hb6)))) ?
                          (($signed(forvar671) ? forvar618 : {(8'hb9)}) ?
                              (^~$unsigned(reg621)) : $unsigned((!forvar611))) : (({reg659} - reg655) ?
                              (forvar631 ?
                                  $signed(reg651) : (reg619 ?
                                      reg645 : reg632)) : $unsigned({wire601})));
                      reg667 <= (^(8'hac));
                      reg668 <= (~{$signed($unsigned(reg629))});
                      reg669 <= (&$unsigned((~((8'hb6) == reg613))));
                    end
                  for (forvar670 = (1'h0); (forvar670 < (1'h0)); forvar670 = (forvar670 + (1'h1)))
                    begin
                      reg671 <= $unsigned((($unsigned(reg616) == $unsigned(reg675)) * forvar607));
                      reg672 <= ((reg631 ?
                              reg659[(3'h6):(2'h3)] : reg620[(3'h5):(2'h3)]) ?
                          (($signed(reg639) ?
                              reg629 : (8'hb1)) == {$signed(reg619)}) : $unsigned($signed(reg642[(2'h2):(1'h1)])));
                    end
                  if (forvar639)
                    begin
                      reg673 <= ((forvar666[(4'h8):(2'h3)] ?
                              {$signed(reg659)} : $signed($signed((8'hb4)))) ?
                          ((~wire604) >> (~&reg631)) : ($unsigned(reg671[(1'h0):(1'h0)]) ^ {((8'h9e) ?
                                  reg634 : forvar644)}));
                      reg674 <= {reg609[(3'h5):(2'h3)]};
                      reg675 <= $signed((~|$unsigned((reg639 & forvar659))));
                    end
                  else
                    begin
                      reg673 <= (!($signed(reg652) ?
                          $signed((^~forvar610)) : $signed((!reg664))));
                    end
                end
            end
          for (forvar676 = (1'h0); (forvar676 < (1'h0)); forvar676 = (forvar676 + (1'h1)))
            begin
              if ({($signed((!forvar672)) >>> $unsigned((&forvar649)))})
                begin
                  if ($unsigned(reg647))
                    begin
                      reg677 <= (reg654 ?
                          forvar659[(4'hb):(4'h9)] : {(^reg670)});
                      reg678 <= (reg672 ?
                          forvar638 : $signed(((~&forvar653) ^ (reg669 ?
                              reg630 : reg621))));
                      reg679 <= $signed(reg648[(3'h5):(1'h0)]);
                      reg680 <= reg678[(3'h6):(3'h6)];
                    end
                  else
                    begin
                      reg677 <= $unsigned(((!reg643) >> (reg619[(5'h10):(4'he)] >> ((8'hb0) ?
                          reg634 : wire601))));
                    end
                  for (forvar681 = (1'h0); (forvar681 < (2'h3)); forvar681 = (forvar681 + (1'h1)))
                    begin
                      reg682 <= (($unsigned(forvar644[(2'h3):(2'h3)]) >> (((8'ha8) + (8'ha6)) ?
                              {reg672} : (reg665 ^~ reg615))) ?
                          $unsigned({(~|forvar660)}) : $unsigned(forvar653[(3'h7):(3'h5)]));
                      reg683 <= $unsigned({(reg644[(2'h2):(1'h0)] ^~ reg655)});
                      reg684 <= (~|$unsigned($unsigned(((8'hac) ?
                          reg617 : (8'ha4)))));
                      reg685 <= ($unsigned(reg608[(4'ha):(3'h7)]) ?
                          $signed($signed((!reg653))) : forvar661);
                    end
                end
              else
                begin
                  reg677 <= ({$signed(forvar612)} & (8'ha8));
                  if ((((reg674 ?
                              ((8'hae) ?
                                  reg606 : (8'hba)) : $signed(forvar620)) ?
                          (|((8'hb7) < reg627)) : {$unsigned((8'ha0))}) ?
                      reg660 : {(reg606 ?
                              {forvar617} : (forvar638 ? reg608 : reg622))}))
                    begin
                      reg678 <= {(forvar676 >> (~&reg614))};
                      reg679 <= ($unsigned((reg622[(1'h0):(1'h0)] <= $signed(forvar628))) <= {((reg614 ?
                                  reg680 : reg654) ?
                              $unsigned(reg629) : reg638)});
                    end
                  else
                    begin
                      reg678 <= reg620;
                      reg679 <= reg626[(4'he):(4'he)];
                    end
                  reg680 <= (~((|forvar660) > $unsigned(((8'ha3) & reg642))));
                  if ((8'ha4))
                    begin
                      reg681 <= (~|($signed(reg669[(4'ha):(4'h8)]) ?
                          {(forvar620 ? forvar610 : reg606)} : {(~^reg683)}));
                      reg682 <= $unsigned(({$unsigned((8'ha4))} <<< reg658[(4'hf):(4'h9)]));
                    end
                  else
                    begin
                      reg681 <= $unsigned({$unsigned({forvar673})});
                      reg682 <= (-$unsigned(((~forvar666) ?
                          (forvar659 ?
                              forvar610 : reg615) : $signed((8'hb9)))));
                    end
                end
            end
        end
      for (forvar686 = (1'h0); (forvar686 < (2'h2)); forvar686 = (forvar686 + (1'h1)))
        begin
          for (forvar687 = (1'h0); (forvar687 < (1'h1)); forvar687 = (forvar687 + (1'h1)))
            begin
              if (forvar607)
                begin
                  if (((reg627[(3'h5):(3'h4)] <<< reg624) * reg672))
                    begin
                      reg688 <= (~&reg672);
                      reg689 <= reg611;
                    end
                  else
                    begin
                      reg688 <= $unsigned(($unsigned((|reg656)) << {forvar648}));
                      reg689 <= (reg619 >> forvar641[(1'h0):(1'h0)]);
                    end
                  for (forvar690 = (1'h0); (forvar690 < (1'h0)); forvar690 = (forvar690 + (1'h1)))
                    begin
                      reg691 <= reg617;
                      reg692 <= (wire605 ?
                          (-((forvar659 < (8'h9f)) ?
                              (^reg630) : $signed(forvar654))) : ({forvar664} ^~ ((reg643 > reg667) ?
                              (forvar607 ?
                                  reg644 : reg617) : reg610[(1'h1):(1'h0)])));
                      reg693 <= (forvar660 && (|{(reg634 ? wire603 : reg634)}));
                    end
                end
              else
                begin
                  reg688 <= ({$unsigned(reg630)} ?
                      reg632[(1'h1):(1'h1)] : {((forvar686 + forvar631) ?
                              ((8'ha8) >= reg656) : $unsigned(reg618))});
                  reg689 <= ($signed((~^(reg647 ? reg679 : forvar669))) ?
                      {(reg655[(2'h2):(2'h2)] ?
                              (~|forvar686) : {reg629})} : (($signed(reg666) ?
                              ((8'ha6) ? forvar648 : (8'hb3)) : (+reg640)) ?
                          {reg635[(4'hc):(2'h3)]} : reg610[(3'h5):(3'h4)]));
                end
            end
          for (forvar694 = (1'h0); (forvar694 < (1'h1)); forvar694 = (forvar694 + (1'h1)))
            begin
              for (forvar695 = (1'h0); (forvar695 < (1'h1)); forvar695 = (forvar695 + (1'h1)))
                begin
                  for (forvar696 = (1'h0); (forvar696 < (2'h2)); forvar696 = (forvar696 + (1'h1)))
                    begin
                      reg697 <= (8'hb5);
                      reg698 <= forvar627;
                    end
                end
            end
          for (forvar699 = (1'h0); (forvar699 < (1'h0)); forvar699 = (forvar699 + (1'h1)))
            begin
              if (forvar623)
                begin
                  if ((($signed((forvar699 ?
                          forvar673 : reg614)) <= reg650[(2'h3):(1'h0)]) ?
                      (~|{(forvar669 ? forvar670 : (8'hac))}) : reg692))
                    begin
                      reg700 <= ($unsigned($unsigned($unsigned((8'hab)))) ?
                          (((~^(8'h9d)) >= {reg691}) ?
                              ((^(8'ha0)) ?
                                  $unsigned((8'hb3)) : $unsigned(reg670)) : $signed((8'hb9))) : (+wire603[(1'h0):(1'h0)]));
                      reg701 <= ({reg659} ?
                          $unsigned(($unsigned(reg678) * ((8'h9e) ?
                              reg654 : reg632))) : forvar673);
                    end
                  else
                    begin
                      reg700 <= {($unsigned(reg684) ?
                              {{forvar690}} : reg678[(2'h2):(2'h2)])};
                      reg701 <= reg692[(4'hc):(3'h7)];
                      reg702 <= (reg682[(2'h2):(2'h2)] + (^reg614));
                      reg703 <= (((~|forvar665) ?
                              $unsigned((reg672 ? reg628 : reg642)) : reg641) ?
                          (&{((8'ha1) ?
                                  reg633 : forvar696)}) : ($unsigned(reg663) ?
                              reg647[(3'h5):(1'h0)] : (~reg685[(3'h4):(2'h2)])));
                    end
                  reg704 <= reg616[(4'he):(4'h8)];
                end
              else
                begin
                  if (wire603[(1'h1):(1'h0)])
                    begin
                      reg700 <= $unsigned((reg634[(2'h2):(2'h2)] == $unsigned((~^reg617))));
                    end
                  else
                    begin
                      reg700 <= $unsigned((~(~|(|(8'had)))));
                      reg701 <= {$signed($unsigned(forvar612[(3'h4):(1'h0)]))};
                      reg702 <= $signed(($unsigned((+reg659)) ?
                          ((&reg643) ?
                              $unsigned(reg634) : (forvar660 ?
                                  reg684 : forvar649)) : (^(~&forvar645))));
                    end
                  if (((!(~|reg632)) <= $unsigned($signed((forvar617 || forvar629)))))
                    begin
                      reg703 <= (~forvar676);
                      reg704 <= ((^$unsigned((reg644 ?
                          forvar617 : forvar608))) <<< {reg698[(4'hb):(3'h4)]});
                    end
                  else
                    begin
                      reg703 <= reg612;
                      reg704 <= ($signed($signed(forvar642[(3'h5):(2'h2)])) ?
                          (&(^reg689)) : reg682[(1'h1):(1'h1)]);
                    end
                  for (forvar705 = (1'h0); (forvar705 < (1'h0)); forvar705 = (forvar705 + (1'h1)))
                    begin
                      reg706 <= (reg652[(2'h2):(1'h0)] | reg637);
                    end
                  for (forvar707 = (1'h0); (forvar707 < (1'h1)); forvar707 = (forvar707 + (1'h1)))
                    begin
                      reg708 <= (reg644 ?
                          ($signed({forvar650}) ?
                              (&{forvar669}) : reg645) : reg631);
                      reg709 <= $unsigned((&forvar617));
                    end
                end
              if ({($unsigned((~&wire602)) ^ reg632)})
                begin
                  if ($signed(forvar652[(3'h5):(3'h5)]))
                    begin
                      reg710 <= ($signed((8'ha4)) >> ((!reg701) ?
                          forvar659 : reg653));
                      reg711 <= forvar654[(1'h1):(1'h1)];
                      reg712 <= $signed(forvar642[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg710 <= (^((+reg626[(2'h2):(2'h2)]) ?
                          {{forvar690}} : reg683));
                    end
                  for (forvar713 = (1'h0); (forvar713 < (1'h1)); forvar713 = (forvar713 + (1'h1)))
                    begin
                      reg714 <= forvar659;
                      reg715 <= ((reg703[(4'he):(3'h6)] ?
                          $signed(reg621[(3'h6):(2'h2)]) : (reg700 ^~ (^~reg655))) + (^~((&(8'ha0)) ?
                          (!forvar694) : forvar648[(2'h2):(1'h1)])));
                      reg716 <= (($signed($unsigned(forvar644)) ?
                              (+(reg640 ?
                                  forvar659 : forvar618)) : (((8'h9c) > forvar690) ?
                                  (reg644 ?
                                      reg691 : (8'ha1)) : $signed(reg706))) ?
                          forvar699[(2'h2):(1'h1)] : reg654[(3'h4):(1'h0)]);
                      reg717 <= $signed($unsigned((forvar645[(4'hb):(4'h9)] ?
                          (reg611 ? (8'h9c) : forvar650) : forvar707)));
                    end
                  if ($unsigned($unsigned($unsigned({(8'had)}))))
                    begin
                      reg718 <= $signed($signed($unsigned((reg610 > reg658))));
                    end
                  else
                    begin
                      reg718 <= (~^((!(reg692 ? reg666 : reg703)) ?
                          $signed((reg675 ~^ reg700)) : (reg652[(2'h2):(1'h0)] ?
                              $unsigned((8'hac)) : $signed(reg630))));
                      reg719 <= reg662[(3'h4):(1'h1)];
                      reg720 <= (((8'ha8) >= ({reg652} ?
                              $signed(reg649) : (~&reg683))) ?
                          $unsigned(forvar618) : (^~{reg665}));
                      reg721 <= $signed($unsigned(reg718[(2'h3):(2'h2)]));
                    end
                end
              else
                begin
                  reg710 <= $unsigned((|({reg704} ?
                      reg700 : (reg689 > reg701))));
                  reg711 <= reg613;
                end
            end
        end
      for (forvar722 = (1'h0); (forvar722 < (1'h1)); forvar722 = (forvar722 + (1'h1)))
        begin
          for (forvar723 = (1'h0); (forvar723 < (2'h3)); forvar723 = (forvar723 + (1'h1)))
            begin
              if ($signed((reg614 ? (^wire605) : (~^reg697[(5'h10):(5'h10)]))))
                begin
                  if ($unsigned(reg652[(1'h0):(1'h0)]))
                    begin
                      reg724 <= reg680;
                      reg725 <= $unsigned((^$signed(reg619)));
                    end
                  else
                    begin
                      reg724 <= $signed(({{forvar681}} ?
                          (~|(reg670 && forvar696)) : $unsigned($signed(reg619))));
                      reg725 <= (+$signed((reg671[(2'h2):(1'h0)] ?
                          (!wire603) : reg697[(2'h3):(1'h0)])));
                      reg726 <= $unsigned(reg701);
                    end
                end
              else
                begin
                  if (reg626[(4'hb):(4'hb)])
                    begin
                      reg724 <= forvar612[(3'h4):(2'h3)];
                      reg725 <= ($signed($unsigned(reg638[(4'hb):(1'h0)])) ?
                          $unsigned((+(reg716 ?
                              forvar620 : (8'h9c)))) : $signed($unsigned((~|reg658))));
                      reg726 <= reg623[(1'h1):(1'h1)];
                      reg727 <= ($unsigned((^(8'hac))) ?
                          ($signed($unsigned(forvar671)) > (|$unsigned(reg634))) : {(~&(|reg688))});
                    end
                  else
                    begin
                      reg724 <= $unsigned((~&(forvar627[(4'hd):(1'h0)] ?
                          $signed(reg606) : reg709)));
                      reg725 <= $signed(($signed(reg630) ?
                          ($signed(forvar665) ?
                              (reg668 ?
                                  (8'hb5) : reg656) : (8'hba)) : ($unsigned(reg664) >>> forvar699[(2'h3):(2'h3)])));
                      reg726 <= (+forvar705);
                    end
                  for (forvar728 = (1'h0); (forvar728 < (1'h0)); forvar728 = (forvar728 + (1'h1)))
                    begin
                      reg729 <= reg725;
                    end
                  reg730 <= $signed(forvar654[(5'h10):(2'h3)]);
                  if ($unsigned((+$unsigned(reg727))))
                    begin
                      reg731 <= (reg654 ?
                          reg645[(4'hd):(4'h8)] : $signed(forvar669[(1'h0):(1'h0)]));
                      reg732 <= (-($signed((~forvar607)) ?
                          (~reg641) : (8'ha6)));
                      reg733 <= ($signed($unsigned((^(8'ha8)))) ?
                          forvar681 : (+((forvar665 ? (8'ha0) : forvar694) ?
                              (reg637 ? reg611 : forvar686) : (~^reg708))));
                      reg734 <= forvar707[(4'hf):(4'h8)];
                    end
                  else
                    begin
                      reg731 <= (&$signed({(!reg703)}));
                      reg732 <= {(($signed(forvar649) ?
                                  $unsigned(reg649) : ((8'ha3) ~^ reg688)) ?
                              (forvar699 ?
                                  (forvar606 + reg709) : reg642) : reg673[(4'h9):(3'h4)])};
                      reg733 <= {(8'ha7)};
                    end
                end
              reg735 <= $signed(forvar615);
              if (forvar707)
                begin
                  if (((reg718 ?
                      ((reg684 ? forvar653 : reg620) * (reg709 ?
                          wire605 : reg633)) : (+(reg716 & reg629))) ^ (reg629[(4'hb):(2'h2)] > forvar722[(3'h7):(3'h5)])))
                    begin
                      reg736 <= reg667;
                      reg737 <= {(&((forvar649 ~^ forvar695) ?
                              $unsigned(forvar681) : forvar629))};
                    end
                  else
                    begin
                      reg736 <= (~&forvar618[(3'h4):(3'h4)]);
                      reg737 <= $signed($signed((~|$signed(forvar631))));
                    end
                  if (($unsigned({$unsigned(forvar671)}) - $unsigned(reg662)))
                    begin
                      reg738 <= $unsigned((^$unsigned(((8'hb3) >= forvar694))));
                      reg739 <= (reg727[(3'h6):(3'h6)] - reg637);
                      reg740 <= ((8'hab) ^~ $unsigned(($signed((8'ha9)) & $signed(reg674))));
                    end
                  else
                    begin
                      reg738 <= (reg625 ?
                          forvar652[(3'h4):(1'h0)] : $unsigned($signed((^~reg670))));
                      reg739 <= (({reg719[(3'h6):(1'h1)]} <= $signed($signed((8'hb6)))) ?
                          (((^reg685) * reg648[(1'h0):(1'h0)]) != (reg609 ?
                              (reg644 ?
                                  reg607 : (8'h9d)) : $signed(reg731))) : forvar650);
                      reg740 <= (~^$unsigned($unsigned((forvar645 == reg692))));
                    end
                  if ($signed($unsigned(forvar623)))
                    begin
                      reg741 <= wire602;
                      reg742 <= $signed(((forvar639[(3'h6):(3'h4)] ?
                              (reg663 >>> forvar661) : $unsigned(forvar612)) ?
                          {$unsigned(reg685)} : ($unsigned(forvar671) >> {reg706})));
                      reg743 <= (^($unsigned((forvar673 && forvar687)) ?
                          (((8'hb4) ~^ reg626) ?
                              $unsigned(forvar669) : (+forvar610)) : {(8'hb2)}));
                      reg744 <= (~&reg637[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg741 <= (8'ha3);
                      reg742 <= forvar690;
                    end
                end
              else
                begin
                  for (forvar736 = (1'h0); (forvar736 < (1'h1)); forvar736 = (forvar736 + (1'h1)))
                    begin
                      reg737 <= (($signed(((8'ha8) ? reg677 : forvar696)) ?
                              forvar713 : (reg709 ?
                                  (8'ha4) : (reg618 ? reg636 : reg688))) ?
                          reg608 : (8'haa));
                      reg738 <= reg679;
                      reg739 <= ($unsigned(reg610[(2'h3):(1'h0)]) == $signed($unsigned(forvar722[(4'hc):(4'hc)])));
                      reg740 <= (($unsigned(reg655[(1'h0):(1'h0)]) ?
                          $signed($signed((8'ha6))) : $signed(reg726[(2'h2):(1'h0)])) ^~ ($signed($unsigned(forvar664)) < forvar611));
                    end
                  for (forvar741 = (1'h0); (forvar741 < (2'h3)); forvar741 = (forvar741 + (1'h1)))
                    begin
                      reg742 <= $signed(((8'hb3) - ($unsigned((8'ha2)) ?
                          (forvar637 ^ wire603) : forvar649)));
                    end
                  if (((!{(forvar644 ? reg732 : (8'ha0))}) ?
                      (~$signed(forvar649)) : ((forvar612 ~^ forvar687[(3'h4):(2'h3)]) >>> reg621[(3'h6):(1'h1)])))
                    begin
                      reg743 <= $signed($unsigned(reg708));
                    end
                  else
                    begin
                      reg743 <= $signed(reg730[(2'h2):(2'h2)]);
                      reg744 <= $unsigned(($unsigned($signed(forvar671)) | ($unsigned(forvar653) & {forvar652})));
                      reg745 <= reg612;
                      reg746 <= reg649;
                    end
                  if (reg628)
                    begin
                      reg747 <= ((^~$signed((8'hae))) ?
                          forvar664[(2'h3):(1'h0)] : reg632[(2'h2):(1'h1)]);
                      reg748 <= $unsigned(($unsigned(reg679[(3'h4):(1'h0)]) ?
                          ({(8'hba)} ?
                              forvar615[(3'h7):(2'h2)] : (reg702 ?
                                  reg732 : reg621)) : forvar669));
                    end
                  else
                    begin
                      reg747 <= forvar741;
                      reg748 <= ($unsigned(reg607) >>> {((reg634 ?
                              forvar631 : forvar615) != $signed((8'ha0)))});
                    end
                end
              reg749 <= reg738[(3'h5):(2'h3)];
            end
          for (forvar750 = (1'h0); (forvar750 < (2'h3)); forvar750 = (forvar750 + (1'h1)))
            begin
              if ({$unsigned({reg727[(3'h7):(2'h2)]})})
                begin
                  reg751 <= $unsigned(reg691);
                  if ((~|(!(~|{forvar648}))))
                    begin
                      reg752 <= reg647[(4'hb):(3'h6)];
                      reg753 <= reg649;
                    end
                  else
                    begin
                      reg752 <= (^~(&((-reg643) ?
                          $unsigned(reg711) : $unsigned(reg674))));
                      reg753 <= $unsigned((reg715[(4'hb):(4'h9)] | $unsigned($signed(reg735))));
                      reg754 <= ($signed(forvar615[(3'h7):(3'h6)]) ?
                          forvar606 : {$signed($signed(reg631))});
                    end
                end
              else
                begin
                  if ($unsigned((-$unsigned((forvar660 ? reg651 : forvar728)))))
                    begin
                      reg751 <= reg660;
                    end
                  else
                    begin
                      reg751 <= {forvar707};
                      reg752 <= reg692;
                    end
                  if (((!$unsigned($unsigned((8'ha0)))) ?
                      (forvar653 ?
                          (&forvar606[(1'h0):(1'h0)]) : (reg674[(1'h1):(1'h1)] ?
                              forvar669 : (^reg675))) : $unsigned(($signed(reg631) >>> (~forvar648)))))
                    begin
                      reg753 <= reg669;
                      reg754 <= forvar637[(3'h5):(3'h4)];
                      reg755 <= forvar659;
                    end
                  else
                    begin
                      reg753 <= reg734[(3'h5):(3'h5)];
                      reg754 <= $signed(($signed((^(8'hb5))) ?
                          ((~^reg710) << forvar638[(3'h6):(1'h0)]) : ((forvar681 || reg652) ?
                              (8'ha3) : $unsigned(reg680))));
                      reg755 <= forvar722;
                      reg756 <= $signed(reg727);
                    end
                end
              for (forvar757 = (1'h0); (forvar757 < (1'h1)); forvar757 = (forvar757 + (1'h1)))
                begin
                  if ($unsigned((((^reg624) <= reg747) < reg737[(2'h3):(1'h1)])))
                    begin
                      reg758 <= reg714;
                      reg759 <= $signed($unsigned(($unsigned(reg617) ?
                          reg647 : (~reg620))));
                      reg760 <= forvar694;
                      reg761 <= ($signed((forvar661[(2'h2):(1'h0)] > (+reg734))) ?
                          forvar615[(1'h0):(1'h0)] : reg698[(4'h9):(3'h7)]);
                    end
                  else
                    begin
                      reg758 <= (reg609 <<< {{forvar736[(1'h0):(1'h0)]}});
                      reg759 <= (~$unsigned($unsigned((forvar654 ?
                          wire605 : reg613))));
                      reg760 <= forvar648[(2'h3):(2'h2)];
                    end
                  for (forvar762 = (1'h0); (forvar762 < (1'h1)); forvar762 = (forvar762 + (1'h1)))
                    begin
                      reg763 <= (8'hac);
                      reg764 <= (reg618 <<< (~$signed(reg693)));
                    end
                end
              if ((^~(reg731 ?
                  (^$unsigned(forvar631)) : reg657[(2'h2):(1'h1)])))
                begin
                  for (forvar765 = (1'h0); (forvar765 < (2'h2)); forvar765 = (forvar765 + (1'h1)))
                    begin
                      reg766 <= (^~(-$unsigned((forvar606 || reg756))));
                      reg767 <= $unsigned(((reg749[(1'h1):(1'h0)] != (~(8'h9d))) ?
                          (~|((8'ha9) & reg619)) : {forvar681[(3'h5):(3'h5)]}));
                      reg768 <= {(~^$signed((reg682 < forvar608)))};
                    end
                end
              else
                begin
                  reg765 <= (8'ha1);
                  if ($unsigned($unsigned((~^(~^forvar681)))))
                    begin
                      reg766 <= forvar653[(1'h0):(1'h0)];
                      reg767 <= (^~($unsigned($unsigned(forvar670)) ?
                          ((forvar622 ?
                              forvar722 : forvar762) == reg731[(1'h1):(1'h1)]) : (forvar631[(4'h9):(4'h9)] ?
                              reg611[(1'h1):(1'h1)] : $signed(reg719))));
                      reg768 <= ((!$unsigned((forvar705 ?
                          reg747 : (8'h9f)))) - reg746[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg766 <= wire603[(3'h4):(2'h3)];
                    end
                end
              if ((({reg683[(1'h1):(1'h1)]} ?
                  $signed($signed(reg745)) : forvar750[(4'h9):(3'h5)]) + ($signed((!reg646)) ?
                  (-$signed((8'had))) : ((~|reg645) ?
                      $unsigned(forvar707) : reg659[(3'h4):(1'h0)]))))
                begin
                  for (forvar769 = (1'h0); (forvar769 < (2'h2)); forvar769 = (forvar769 + (1'h1)))
                    begin
                      reg770 <= reg625[(1'h1):(1'h1)];
                      reg771 <= (|{((reg636 <= reg613) ?
                              $signed(reg615) : forvar615)});
                      reg772 <= ((!forvar695) ?
                          forvar673 : (^~$signed({forvar672})));
                    end
                  if (forvar627)
                    begin
                      reg773 <= (+($unsigned((~|forvar661)) && (wire605[(4'hb):(2'h2)] - ((8'ha4) ?
                          reg748 : reg724))));
                    end
                  else
                    begin
                      reg773 <= reg685;
                      reg774 <= (forvar620 ?
                          {forvar606[(2'h3):(1'h1)]} : reg680[(4'hb):(2'h3)]);
                      reg775 <= reg640;
                      reg776 <= (forvar617[(2'h3):(2'h3)] >= $signed($signed(((8'had) ?
                          reg681 : reg630))));
                    end
                  reg777 <= $unsigned((+reg741));
                end
              else
                begin
                  if ($signed($unsigned(((8'hb9) ?
                      reg751[(1'h0):(1'h0)] : {reg655}))))
                    begin
                      reg769 <= $unsigned((forvar671 ?
                          reg774[(2'h2):(1'h1)] : {(reg655 && (8'hb4))}));
                    end
                  else
                    begin
                      reg769 <= (^~forvar644);
                    end
                  for (forvar770 = (1'h0); (forvar770 < (2'h3)); forvar770 = (forvar770 + (1'h1)))
                    begin
                      reg771 <= reg727[(3'h5):(3'h4)];
                      reg772 <= (-$signed(($signed(forvar641) == forvar672)));
                      reg773 <= reg666[(1'h1):(1'h1)];
                    end
                end
            end
        end
      reg778 <= forvar650;
    end
  assign wire779 = (^~reg761[(2'h2):(1'h0)]);
  assign wire780 = (reg759 >>> forvar650);
  assign wire781 = {reg712};
  assign wire782 = ((forvar606[(1'h0):(1'h0)] != ({reg716} + reg708)) == (8'hb8));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1515
#( parameter param1646 = ((8'hb2) | (((8'ha5) < ((8'hb6) >= (8'hae))) ? (((8'ha5) >>> (8'hb9)) ? (8'h9d) : ((8'haf) ^~ (8'ha1))) : (((8'ha3) ? (8'ha1) : (8'ha8)) ? (^(8'h9d)) : {(8'h9c)}))) )
(y, clk, wire1520, wire1519, wire1518, wire1517, wire1516);
  output wire [(32'h4f5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'he):(1'h0)] wire1520;
  input wire signed [(2'h2):(1'h0)] wire1519;
  input wire [(3'h5):(1'h0)] wire1518;
  input wire signed [(5'h10):(1'h0)] wire1517;
  input wire signed [(4'hf):(1'h0)] wire1516;
  wire signed [(4'h9):(1'h0)] wire1645;
  wire signed [(4'hc):(1'h0)] wire1644;
  reg signed [(3'h4):(1'h0)] reg1643 = (1'h0);
  reg [(4'hd):(1'h0)] reg1544 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1541 = (1'h0);
  reg [(3'h6):(1'h0)] reg1539 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1536 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1535 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1528 = (1'h0);
  reg [(4'h8):(1'h0)] reg1530 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1642 = (1'h0);
  reg [(5'h10):(1'h0)] reg1641 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1640 = (1'h0);
  reg [(2'h2):(1'h0)] reg1639 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1638 = (1'h0);
  reg [(3'h5):(1'h0)] reg1636 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1635 = (1'h0);
  reg [(3'h4):(1'h0)] reg1637 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1636 = (1'h0);
  reg [(4'h8):(1'h0)] reg1635 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1632 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1631 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1629 = (1'h0);
  reg [(4'hd):(1'h0)] reg1634 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1633 = (1'h0);
  reg [(5'h10):(1'h0)] reg1632 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1631 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1630 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1629 = (1'h0);
  reg [(4'hc):(1'h0)] reg1628 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1627 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1621 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1619 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1627 = (1'h0);
  reg [(2'h2):(1'h0)] reg1626 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1625 = (1'h0);
  reg [(4'hb):(1'h0)] reg1624 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1623 = (1'h0);
  reg [(5'h10):(1'h0)] reg1622 = (1'h0);
  reg [(4'hb):(1'h0)] reg1621 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1620 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1619 = (1'h0);
  reg [(3'h7):(1'h0)] reg1618 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1617 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1616 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1615 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1614 = (1'h0);
  reg [(3'h4):(1'h0)] reg1613 = (1'h0);
  reg [(3'h7):(1'h0)] reg1612 = (1'h0);
  reg [(4'he):(1'h0)] forvar1611 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1610 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1609 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1608 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1607 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1606 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1605 = (1'h0);
  reg [(3'h7):(1'h0)] reg1604 = (1'h0);
  reg [(4'h8):(1'h0)] reg1603 = (1'h0);
  reg [(4'he):(1'h0)] forvar1602 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1601 = (1'h0);
  reg [(2'h3):(1'h0)] reg1600 = (1'h0);
  reg [(3'h6):(1'h0)] reg1599 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1598 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1597 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1596 = (1'h0);
  reg [(2'h3):(1'h0)] reg1595 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1594 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1593 = (1'h0);
  reg [(4'hf):(1'h0)] reg1592 = (1'h0);
  reg [(4'he):(1'h0)] forvar1591 = (1'h0);
  reg [(4'hf):(1'h0)] reg1591 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1590 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1589 = (1'h0);
  reg [(4'h9):(1'h0)] reg1588 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1587 = (1'h0);
  reg [(3'h7):(1'h0)] reg1586 = (1'h0);
  reg [(3'h4):(1'h0)] reg1585 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1584 = (1'h0);
  reg [(3'h5):(1'h0)] reg1583 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1582 = (1'h0);
  reg [(4'he):(1'h0)] reg1581 = (1'h0);
  reg [(4'hd):(1'h0)] reg1580 = (1'h0);
  reg [(4'hf):(1'h0)] reg1579 = (1'h0);
  reg [(4'h8):(1'h0)] reg1578 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1577 = (1'h0);
  reg [(4'ha):(1'h0)] reg1576 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1575 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1565 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1563 = (1'h0);
  reg [(4'hc):(1'h0)] reg1574 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1573 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1572 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1571 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1570 = (1'h0);
  reg [(4'h8):(1'h0)] reg1569 = (1'h0);
  reg [(4'h9):(1'h0)] reg1568 = (1'h0);
  reg [(3'h6):(1'h0)] reg1567 = (1'h0);
  reg [(4'h9):(1'h0)] reg1566 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1565 = (1'h0);
  reg [(3'h7):(1'h0)] reg1564 = (1'h0);
  reg [(4'h9):(1'h0)] reg1563 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1562 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1561 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1560 = (1'h0);
  reg [(4'h8):(1'h0)] reg1559 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1558 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1557 = (1'h0);
  reg [(4'h8):(1'h0)] reg1556 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1555 = (1'h0);
  reg [(2'h3):(1'h0)] reg1554 = (1'h0);
  reg [(5'h10):(1'h0)] reg1553 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1552 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1551 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1550 = (1'h0);
  reg [(3'h7):(1'h0)] reg1549 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1548 = (1'h0);
  reg [(4'hb):(1'h0)] reg1547 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1546 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1545 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1544 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1543 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1542 = (1'h0);
  reg [(4'ha):(1'h0)] reg1541 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1540 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1539 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1538 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1537 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1536 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1535 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1534 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1533 = (1'h0);
  reg [(3'h6):(1'h0)] reg1532 = (1'h0);
  reg [(3'h7):(1'h0)] reg1531 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1530 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1529 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1528 = (1'h0);
  wire [(3'h4):(1'h0)] wire1527;
  reg [(4'ha):(1'h0)] reg1526 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1525 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1524 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1523 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1522 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1521 = (1'h0);
  assign y = {wire1645,
                 wire1644,
                 reg1643,
                 reg1544,
                 forvar1541,
                 reg1539,
                 forvar1536,
                 forvar1535,
                 reg1528,
                 reg1530,
                 reg1642,
                 reg1641,
                 reg1640,
                 reg1639,
                 forvar1638,
                 reg1636,
                 forvar1635,
                 reg1637,
                 forvar1636,
                 reg1635,
                 forvar1632,
                 reg1631,
                 reg1629,
                 reg1634,
                 reg1633,
                 reg1632,
                 forvar1631,
                 reg1630,
                 forvar1629,
                 reg1628,
                 forvar1627,
                 forvar1621,
                 forvar1619,
                 reg1627,
                 reg1626,
                 reg1625,
                 reg1624,
                 forvar1623,
                 reg1622,
                 reg1621,
                 reg1620,
                 reg1619,
                 reg1618,
                 reg1617,
                 forvar1616,
                 reg1615,
                 forvar1614,
                 reg1613,
                 reg1612,
                 forvar1611,
                 reg1610,
                 forvar1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1603,
                 forvar1602,
                 forvar1601,
                 reg1600,
                 reg1599,
                 forvar1598,
                 reg1597,
                 reg1596,
                 reg1595,
                 reg1594,
                 reg1593,
                 reg1592,
                 forvar1591,
                 reg1591,
                 reg1590,
                 reg1589,
                 reg1588,
                 forvar1587,
                 reg1586,
                 reg1585,
                 reg1584,
                 reg1583,
                 forvar1582,
                 reg1581,
                 reg1580,
                 reg1579,
                 reg1578,
                 forvar1577,
                 reg1576,
                 forvar1575,
                 reg1565,
                 forvar1563,
                 reg1574,
                 reg1573,
                 reg1572,
                 reg1571,
                 forvar1570,
                 reg1569,
                 reg1568,
                 reg1567,
                 reg1566,
                 forvar1565,
                 reg1564,
                 reg1563,
                 forvar1562,
                 reg1561,
                 forvar1560,
                 reg1559,
                 forvar1558,
                 reg1557,
                 reg1556,
                 forvar1555,
                 reg1554,
                 reg1553,
                 reg1552,
                 reg1551,
                 forvar1550,
                 reg1549,
                 forvar1548,
                 reg1547,
                 reg1546,
                 reg1545,
                 forvar1544,
                 reg1543,
                 reg1542,
                 reg1541,
                 forvar1540,
                 forvar1539,
                 reg1538,
                 reg1537,
                 reg1536,
                 reg1535,
                 reg1534,
                 reg1533,
                 reg1532,
                 reg1531,
                 forvar1530,
                 forvar1529,
                 forvar1528,
                 wire1527,
                 reg1526,
                 reg1525,
                 reg1524,
                 forvar1523,
                 forvar1522,
                 forvar1521,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1521 = (1'h0); (forvar1521 < (2'h2)); forvar1521 = (forvar1521 + (1'h1)))
        begin
          for (forvar1522 = (1'h0); (forvar1522 < (2'h2)); forvar1522 = (forvar1522 + (1'h1)))
            begin
              for (forvar1523 = (1'h0); (forvar1523 < (1'h0)); forvar1523 = (forvar1523 + (1'h1)))
                begin
                  if ($unsigned(((wire1520 ?
                      wire1517 : (wire1517 & wire1519)) ^ ((forvar1523 + wire1517) >>> ((8'ha8) + (8'hab))))))
                    begin
                      reg1524 <= $unsigned((wire1519[(2'h2):(2'h2)] ?
                          $signed(wire1520[(4'hb):(3'h7)]) : $signed($unsigned(wire1520))));
                      reg1525 <= (~$unsigned(reg1524[(4'ha):(4'ha)]));
                    end
                  else
                    begin
                      reg1524 <= ((~&wire1520[(1'h1):(1'h1)]) ?
                          wire1517 : reg1525);
                      reg1525 <= (&forvar1521[(2'h2):(1'h1)]);
                      reg1526 <= forvar1522[(4'h9):(2'h2)];
                    end
                end
            end
        end
    end
  assign wire1527 = (^wire1518);
  always
    @(posedge clk) begin
      if ((~|($signed(reg1525[(1'h0):(1'h0)]) - $signed((~wire1518)))))
        begin
          for (forvar1528 = (1'h0); (forvar1528 < (2'h2)); forvar1528 = (forvar1528 + (1'h1)))
            begin
              for (forvar1529 = (1'h0); (forvar1529 < (1'h1)); forvar1529 = (forvar1529 + (1'h1)))
                begin
                  for (forvar1530 = (1'h0); (forvar1530 < (2'h2)); forvar1530 = (forvar1530 + (1'h1)))
                    begin
                      reg1531 <= (8'hae);
                      reg1532 <= wire1516[(4'hf):(1'h1)];
                      reg1533 <= (~(~reg1531[(2'h2):(1'h1)]));
                      reg1534 <= forvar1523;
                    end
                  if ($signed(reg1525[(4'hd):(4'hd)]))
                    begin
                      reg1535 <= (~&(($unsigned(reg1525) ?
                              (!reg1533) : reg1524) ?
                          ($unsigned((8'hb2)) >>> {reg1533}) : {$signed(reg1531)}));
                      reg1536 <= {$signed(((reg1534 - (8'hab)) ?
                              {reg1534} : reg1525[(4'h9):(4'h8)]))};
                      reg1537 <= (!$signed(((forvar1530 != forvar1529) ?
                          (reg1534 ? (8'ha0) : reg1535) : $signed(reg1531))));
                      reg1538 <= (~^(^~$signed(((8'hb1) ~^ forvar1522))));
                    end
                  else
                    begin
                      reg1535 <= (+$unsigned((~^(wire1516 ?
                          (8'ha9) : reg1525))));
                    end
                end
              for (forvar1539 = (1'h0); (forvar1539 < (2'h2)); forvar1539 = (forvar1539 + (1'h1)))
                begin
                  for (forvar1540 = (1'h0); (forvar1540 < (2'h2)); forvar1540 = (forvar1540 + (1'h1)))
                    begin
                      reg1541 <= ($unsigned((8'haf)) ?
                          (-({reg1538} ?
                              $unsigned(reg1531) : {wire1517})) : ((^{forvar1530}) + (^~{(8'h9c)})));
                      reg1542 <= $signed(reg1526[(1'h1):(1'h1)]);
                      reg1543 <= $signed(wire1518[(3'h4):(1'h1)]);
                    end
                  for (forvar1544 = (1'h0); (forvar1544 < (2'h3)); forvar1544 = (forvar1544 + (1'h1)))
                    begin
                      reg1545 <= ((~|($unsigned(wire1517) <<< (wire1517 ~^ reg1525))) && {((!wire1516) ~^ $unsigned(forvar1521))});
                      reg1546 <= ((-reg1538[(1'h0):(1'h0)]) ?
                          forvar1529 : ($signed($signed(forvar1529)) ?
                              $unsigned($signed(reg1526)) : wire1517));
                    end
                end
              if ((forvar1522[(4'h9):(1'h0)] ?
                  ((^forvar1540[(2'h3):(2'h2)]) && {{wire1519}}) : (reg1541[(2'h2):(1'h1)] ?
                      ((forvar1528 << (8'had)) << (!forvar1523)) : ((~&reg1532) ?
                          (8'ha0) : $unsigned(reg1546)))))
                begin
                  reg1547 <= $unsigned(((^$signed(reg1538)) ?
                      ($unsigned(reg1533) * $signed((8'ha3))) : ((reg1533 == reg1534) ?
                          $signed(wire1519) : {reg1524})));
                end
              else
                begin
                  reg1547 <= $signed($signed(($unsigned(reg1531) && $signed(reg1538))));
                  for (forvar1548 = (1'h0); (forvar1548 < (2'h3)); forvar1548 = (forvar1548 + (1'h1)))
                    begin
                      reg1549 <= $signed({reg1547});
                    end
                  for (forvar1550 = (1'h0); (forvar1550 < (1'h0)); forvar1550 = (forvar1550 + (1'h1)))
                    begin
                      reg1551 <= forvar1544[(3'h4):(2'h3)];
                      reg1552 <= forvar1530[(4'h8):(1'h0)];
                      reg1553 <= $signed($unsigned((reg1533 ?
                          reg1546[(2'h3):(1'h1)] : (forvar1530 >>> (8'hae)))));
                      reg1554 <= $signed(reg1552[(3'h4):(2'h3)]);
                    end
                  for (forvar1555 = (1'h0); (forvar1555 < (1'h1)); forvar1555 = (forvar1555 + (1'h1)))
                    begin
                      reg1556 <= $signed($signed(reg1526));
                      reg1557 <= (8'hb7);
                    end
                end
              for (forvar1558 = (1'h0); (forvar1558 < (1'h1)); forvar1558 = (forvar1558 + (1'h1)))
                begin
                  reg1559 <= ((+(~&$signed((8'hb4)))) - wire1519[(2'h2):(2'h2)]);
                  for (forvar1560 = (1'h0); (forvar1560 < (2'h3)); forvar1560 = (forvar1560 + (1'h1)))
                    begin
                      reg1561 <= {(^(reg1552[(3'h4):(3'h4)] ?
                              forvar1544[(4'ha):(4'h9)] : (reg1534 < (8'haf))))};
                    end
                end
            end
          for (forvar1562 = (1'h0); (forvar1562 < (2'h3)); forvar1562 = (forvar1562 + (1'h1)))
            begin
              if ((reg1536[(3'h6):(3'h6)] >= reg1538[(1'h0):(1'h0)]))
                begin
                  if ((reg1535 ?
                      $unsigned({(reg1526 == wire1517)}) : $unsigned(({reg1552} ?
                          reg1554 : (^reg1546)))))
                    begin
                      reg1563 <= $unsigned((~&reg1551));
                    end
                  else
                    begin
                      reg1563 <= forvar1562[(1'h1):(1'h0)];
                      reg1564 <= {$unsigned(({reg1552} ?
                              ((8'hb4) ?
                                  reg1534 : reg1556) : reg1543[(3'h4):(1'h0)]))};
                    end
                  for (forvar1565 = (1'h0); (forvar1565 < (1'h0)); forvar1565 = (forvar1565 + (1'h1)))
                    begin
                      reg1566 <= {{$unsigned(reg1557)}};
                      reg1567 <= reg1536;
                      reg1568 <= $unsigned((+(&reg1551)));
                      reg1569 <= ((reg1546[(1'h1):(1'h0)] ?
                              reg1537 : forvar1521) ?
                          (~(forvar1550 && reg1545)) : $unsigned({(8'ha1)}));
                    end
                  for (forvar1570 = (1'h0); (forvar1570 < (1'h0)); forvar1570 = (forvar1570 + (1'h1)))
                    begin
                      reg1571 <= $signed(reg1564[(3'h7):(2'h3)]);
                      reg1572 <= (~forvar1570[(4'h8):(4'h8)]);
                      reg1573 <= (~&($unsigned((forvar1562 ?
                          reg1561 : forvar1544)) + ((reg1551 ?
                          wire1519 : wire1517) - forvar1565)));
                      reg1574 <= reg1524;
                    end
                end
              else
                begin
                  for (forvar1563 = (1'h0); (forvar1563 < (2'h3)); forvar1563 = (forvar1563 + (1'h1)))
                    begin
                      reg1564 <= ($unsigned((+$unsigned(reg1559))) ?
                          reg1567[(3'h4):(3'h4)] : $unsigned($signed((forvar1539 ?
                              reg1525 : reg1572))));
                      reg1565 <= {(($unsigned((8'had)) <<< (reg1572 ?
                                  (8'hac) : forvar1523)) ?
                              reg1531 : wire1520)};
                      reg1566 <= ((forvar1528 < {{(8'h9e)}}) ?
                          (8'hb6) : reg1557[(1'h1):(1'h0)]);
                      reg1567 <= (+$signed(reg1553));
                    end
                end
              for (forvar1575 = (1'h0); (forvar1575 < (2'h3)); forvar1575 = (forvar1575 + (1'h1)))
                begin
                  reg1576 <= $signed($unsigned($signed((&(8'h9c)))));
                  for (forvar1577 = (1'h0); (forvar1577 < (2'h2)); forvar1577 = (forvar1577 + (1'h1)))
                    begin
                      reg1578 <= reg1552[(2'h2):(2'h2)];
                      reg1579 <= (({(forvar1558 ?
                                  reg1559 : (8'h9d))} * forvar1521) ?
                          reg1561 : $signed(($signed(forvar1570) ?
                              reg1559 : reg1526)));
                      reg1580 <= reg1578;
                      reg1581 <= (!$signed(reg1532[(2'h2):(1'h1)]));
                    end
                  for (forvar1582 = (1'h0); (forvar1582 < (2'h3)); forvar1582 = (forvar1582 + (1'h1)))
                    begin
                      reg1583 <= $unsigned({$unsigned($unsigned(reg1541))});
                      reg1584 <= $signed({($signed(wire1518) ?
                              (forvar1528 ?
                                  reg1564 : reg1573) : (reg1572 | forvar1563))});
                      reg1585 <= (~$unsigned($unsigned({forvar1522})));
                      reg1586 <= (&($unsigned((-forvar1582)) >= $unsigned((reg1573 ?
                          forvar1548 : forvar1570))));
                    end
                  for (forvar1587 = (1'h0); (forvar1587 < (1'h0)); forvar1587 = (forvar1587 + (1'h1)))
                    begin
                      reg1588 <= (&{(&$unsigned(reg1586))});
                      reg1589 <= (^~(~&((wire1516 == reg1542) ?
                          (reg1546 ^~ reg1564) : ((8'hb5) ?
                              forvar1530 : reg1574))));
                    end
                end
              reg1590 <= (^reg1578);
              if (reg1571)
                begin
                  reg1591 <= wire1519[(1'h0):(1'h0)];
                end
              else
                begin
                  for (forvar1591 = (1'h0); (forvar1591 < (2'h2)); forvar1591 = (forvar1591 + (1'h1)))
                    begin
                      reg1592 <= reg1533[(2'h3):(2'h3)];
                      reg1593 <= reg1579;
                      reg1594 <= $unsigned({($signed(forvar1544) != $unsigned(forvar1560))});
                    end
                  if ((reg1589[(3'h6):(2'h2)] + $signed((&{reg1532}))))
                    begin
                      reg1595 <= ((8'haf) ? {reg1553[(3'h4):(3'h4)]} : reg1567);
                      reg1596 <= (($signed($unsigned(wire1527)) ?
                          reg1567 : ((~^reg1572) <<< (reg1583 ?
                              forvar1560 : reg1557))) ^~ (^~$unsigned(forvar1539)));
                      reg1597 <= (((reg1576[(3'h4):(2'h2)] ?
                              ((8'haf) < wire1516) : $unsigned(forvar1544)) ?
                          ($unsigned(forvar1570) - ((8'h9d) >= (8'ha5))) : (~(reg1542 ?
                              reg1557 : reg1594))) || ((~|$signed((8'hb4))) ?
                          $unsigned($unsigned(reg1589)) : reg1537[(3'h7):(3'h5)]));
                    end
                  else
                    begin
                      reg1595 <= (((8'hb6) - (!(reg1541 ?
                          forvar1587 : (8'ha2)))) ^~ (8'ha0));
                    end
                  for (forvar1598 = (1'h0); (forvar1598 < (1'h1)); forvar1598 = (forvar1598 + (1'h1)))
                    begin
                      reg1599 <= ((reg1572 ?
                          $unsigned($unsigned(reg1541)) : $signed((8'haa))) != ((|$signed(reg1538)) ^~ $signed({reg1531})));
                      reg1600 <= reg1536;
                    end
                end
            end
          for (forvar1601 = (1'h0); (forvar1601 < (2'h2)); forvar1601 = (forvar1601 + (1'h1)))
            begin
              if (forvar1522[(3'h7):(3'h5)])
                begin
                  for (forvar1602 = (1'h0); (forvar1602 < (1'h0)); forvar1602 = (forvar1602 + (1'h1)))
                    begin
                      reg1603 <= ({({(8'ha7)} > (forvar1602 ~^ reg1535))} != $unsigned((forvar1539[(2'h2):(2'h2)] >= ((8'hb0) ?
                          reg1546 : wire1518))));
                      reg1604 <= (|reg1533);
                    end
                  reg1605 <= (~^(8'hb8));
                end
              else
                begin
                  for (forvar1602 = (1'h0); (forvar1602 < (1'h1)); forvar1602 = (forvar1602 + (1'h1)))
                    begin
                      reg1603 <= forvar1540;
                    end
                  if (forvar1523)
                    begin
                      reg1604 <= reg1590[(4'hb):(2'h2)];
                    end
                  else
                    begin
                      reg1604 <= (forvar1598[(4'h9):(2'h2)] ?
                          reg1605[(1'h0):(1'h0)] : reg1592[(4'hc):(4'h8)]);
                      reg1605 <= reg1573;
                      reg1606 <= $unsigned($signed((reg1597 ^~ reg1553)));
                    end
                  reg1607 <= (reg1545[(2'h2):(1'h0)] ?
                      (~reg1571[(4'hb):(3'h5)]) : $signed(reg1559[(3'h5):(2'h3)]));
                  reg1608 <= reg1545[(4'h8):(3'h7)];
                end
              for (forvar1609 = (1'h0); (forvar1609 < (2'h3)); forvar1609 = (forvar1609 + (1'h1)))
                begin
                  reg1610 <= ((~|{$signed(reg1531)}) ?
                      reg1561 : ((-reg1542) ?
                          $unsigned($unsigned(reg1604)) : ((reg1596 ?
                                  reg1574 : reg1534) ?
                              reg1525 : $unsigned((8'ha3)))));
                  for (forvar1611 = (1'h0); (forvar1611 < (2'h3)); forvar1611 = (forvar1611 + (1'h1)))
                    begin
                      reg1612 <= $unsigned(((8'hba) <<< $unsigned($signed(reg1572))));
                      reg1613 <= {(^~(8'hb5))};
                    end
                  for (forvar1614 = (1'h0); (forvar1614 < (2'h3)); forvar1614 = (forvar1614 + (1'h1)))
                    begin
                      reg1615 <= forvar1602[(2'h3):(1'h1)];
                    end
                  for (forvar1616 = (1'h0); (forvar1616 < (1'h1)); forvar1616 = (forvar1616 + (1'h1)))
                    begin
                      reg1617 <= {(-{forvar1540[(2'h2):(1'h1)]})};
                      reg1618 <= $unsigned((~&$unsigned((reg1566 ?
                          reg1547 : forvar1528))));
                    end
                end
            end
          if (reg1546[(2'h3):(2'h2)])
            begin
              if (reg1542[(1'h1):(1'h1)])
                begin
                  if (reg1594[(3'h4):(1'h0)])
                    begin
                      reg1619 <= $signed($signed({reg1591[(3'h7):(3'h4)]}));
                      reg1620 <= (~|($unsigned($unsigned((8'ha6))) ?
                          (~^reg1543[(2'h3):(1'h0)]) : forvar1550[(1'h1):(1'h1)]));
                      reg1621 <= {({(reg1584 ? reg1546 : reg1589)} ?
                              {((8'haf) >>> (8'hb8))} : forvar1544)};
                      reg1622 <= forvar1602;
                    end
                  else
                    begin
                      reg1619 <= reg1563;
                    end
                  for (forvar1623 = (1'h0); (forvar1623 < (1'h1)); forvar1623 = (forvar1623 + (1'h1)))
                    begin
                      reg1624 <= reg1551;
                      reg1625 <= $signed(forvar1562[(1'h1):(1'h0)]);
                      reg1626 <= (((&(8'hae)) ?
                          {(~&reg1556)} : ($signed(forvar1598) ?
                              reg1531 : (&reg1589))) ^ reg1535[(3'h6):(2'h2)]);
                    end
                  reg1627 <= reg1536;
                end
              else
                begin
                  for (forvar1619 = (1'h0); (forvar1619 < (2'h3)); forvar1619 = (forvar1619 + (1'h1)))
                    begin
                      reg1620 <= (8'h9e);
                      reg1621 <= (~|{reg1524});
                      reg1622 <= reg1556;
                    end
                end
            end
          else
            begin
              for (forvar1619 = (1'h0); (forvar1619 < (2'h2)); forvar1619 = (forvar1619 + (1'h1)))
                begin
                  reg1620 <= {(^~(-$signed(forvar1528)))};
                  for (forvar1621 = (1'h0); (forvar1621 < (1'h0)); forvar1621 = (forvar1621 + (1'h1)))
                    begin
                      reg1622 <= ($unsigned((!forvar1529[(2'h2):(1'h0)])) ?
                          reg1534 : $signed(reg1618[(1'h1):(1'h1)]));
                    end
                  for (forvar1623 = (1'h0); (forvar1623 < (2'h2)); forvar1623 = (forvar1623 + (1'h1)))
                    begin
                      reg1624 <= $unsigned(forvar1540);
                      reg1625 <= (8'had);
                      reg1626 <= ({forvar1587[(1'h1):(1'h1)]} - {((-forvar1591) ?
                              (~&reg1627) : (reg1590 ? (8'hb6) : reg1567))});
                    end
                end
              if (forvar1611)
                begin
                  for (forvar1627 = (1'h0); (forvar1627 < (1'h0)); forvar1627 = (forvar1627 + (1'h1)))
                    begin
                      reg1628 <= $signed((($signed(reg1556) ?
                          $signed(reg1556) : $unsigned((8'ha5))) != $unsigned($signed(reg1537))));
                    end
                  for (forvar1629 = (1'h0); (forvar1629 < (1'h0)); forvar1629 = (forvar1629 + (1'h1)))
                    begin
                      reg1630 <= (+forvar1616);
                    end
                  for (forvar1631 = (1'h0); (forvar1631 < (1'h0)); forvar1631 = (forvar1631 + (1'h1)))
                    begin
                      reg1632 <= reg1624;
                      reg1633 <= reg1551;
                      reg1634 <= (|(+reg1524));
                    end
                end
              else
                begin
                  for (forvar1627 = (1'h0); (forvar1627 < (2'h3)); forvar1627 = (forvar1627 + (1'h1)))
                    begin
                      reg1628 <= reg1524;
                      reg1629 <= (($unsigned(reg1574) ?
                          ((reg1605 ?
                              wire1516 : reg1585) <<< reg1576) : ($signed(reg1626) ?
                              reg1600 : $unsigned(reg1564))) ~^ $signed(reg1588));
                      reg1630 <= {{((reg1588 || reg1561) ?
                                  wire1527 : $unsigned((8'hac)))}};
                    end
                  if (reg1589)
                    begin
                      reg1631 <= (+{{reg1605}});
                    end
                  else
                    begin
                      reg1631 <= (~{reg1591});
                    end
                  for (forvar1632 = (1'h0); (forvar1632 < (2'h3)); forvar1632 = (forvar1632 + (1'h1)))
                    begin
                      reg1633 <= (8'ha5);
                    end
                end
              if ((^~((((8'hb8) ? reg1547 : (8'hb1)) ?
                      $signed((8'ha5)) : $signed(forvar1555)) ?
                  $signed($unsigned(reg1525)) : ((^reg1617) == (&reg1571)))))
                begin
                  reg1635 <= $signed(($signed((~&reg1621)) | (&reg1632[(3'h7):(2'h3)])));
                  for (forvar1636 = (1'h0); (forvar1636 < (1'h0)); forvar1636 = (forvar1636 + (1'h1)))
                    begin
                      reg1637 <= (~&(-$signed((reg1561 ? (8'ha8) : reg1531))));
                    end
                end
              else
                begin
                  for (forvar1635 = (1'h0); (forvar1635 < (1'h0)); forvar1635 = (forvar1635 + (1'h1)))
                    begin
                      reg1636 <= $unsigned({(~|forvar1636)});
                    end
                end
              for (forvar1638 = (1'h0); (forvar1638 < (1'h1)); forvar1638 = (forvar1638 + (1'h1)))
                begin
                  if ($signed(reg1536[(3'h5):(3'h4)]))
                    begin
                      reg1639 <= (^(!(forvar1587[(3'h4):(2'h2)] - ((8'hb9) + forvar1555))));
                      reg1640 <= $signed((|forvar1522[(3'h4):(1'h1)]));
                      reg1641 <= forvar1523[(4'h9):(2'h3)];
                      reg1642 <= (+reg1607);
                    end
                  else
                    begin
                      reg1639 <= (($unsigned({(8'ha3)}) && reg1585[(2'h2):(1'h1)]) ?
                          (reg1543 >= reg1563[(3'h5):(1'h0)]) : ($signed((reg1641 ^ forvar1627)) ?
                              reg1526[(4'h8):(1'h1)] : $signed(((8'ha5) ?
                                  reg1606 : reg1545))));
                      reg1640 <= (reg1536 <= {(^~reg1567[(3'h4):(2'h3)])});
                      reg1641 <= (8'hb9);
                    end
                end
            end
        end
      else
        begin
          if ({reg1592})
            begin
              for (forvar1528 = (1'h0); (forvar1528 < (1'h1)); forvar1528 = (forvar1528 + (1'h1)))
                begin
                  for (forvar1529 = (1'h0); (forvar1529 < (1'h0)); forvar1529 = (forvar1529 + (1'h1)))
                    begin
                      reg1530 <= $unsigned($signed((~|(reg1606 > (8'ha6)))));
                      reg1531 <= {reg1579[(4'hd):(1'h0)]};
                      reg1532 <= reg1564[(2'h3):(1'h0)];
                    end
                end
            end
          else
            begin
              reg1528 <= (!($signed((reg1612 ?
                  wire1516 : reg1627)) << (forvar1621[(3'h4):(3'h4)] ?
                  reg1642 : $unsigned(forvar1522))));
              for (forvar1529 = (1'h0); (forvar1529 < (1'h0)); forvar1529 = (forvar1529 + (1'h1)))
                begin
                  for (forvar1530 = (1'h0); (forvar1530 < (1'h0)); forvar1530 = (forvar1530 + (1'h1)))
                    begin
                      reg1531 <= $unsigned($signed(($unsigned(reg1552) <<< $unsigned(reg1603))));
                      reg1532 <= {((^(reg1543 ^ reg1573)) ?
                              (8'hab) : $signed($signed(reg1542)))};
                      reg1533 <= $unsigned((((&reg1605) ?
                          reg1573[(1'h0):(1'h0)] : reg1642[(2'h2):(1'h0)]) >> $signed(reg1633)));
                      reg1534 <= reg1603[(4'h8):(1'h1)];
                    end
                end
              for (forvar1535 = (1'h0); (forvar1535 < (1'h1)); forvar1535 = (forvar1535 + (1'h1)))
                begin
                  for (forvar1536 = (1'h0); (forvar1536 < (2'h2)); forvar1536 = (forvar1536 + (1'h1)))
                    begin
                      reg1537 <= (&reg1589);
                      reg1538 <= ((!((!reg1566) ? (8'ha9) : (+forvar1565))) ?
                          reg1568[(3'h7):(2'h3)] : $unsigned({(&reg1637)}));
                      reg1539 <= {($signed((^~reg1622)) ?
                              (forvar1627 < (reg1551 ~^ reg1557)) : $signed(((8'ha0) ?
                                  reg1596 : reg1552)))};
                    end
                end
              for (forvar1540 = (1'h0); (forvar1540 < (2'h2)); forvar1540 = (forvar1540 + (1'h1)))
                begin
                  for (forvar1541 = (1'h0); (forvar1541 < (1'h1)); forvar1541 = (forvar1541 + (1'h1)))
                    begin
                      reg1542 <= forvar1529;
                      reg1543 <= ({{(forvar1611 ? reg1547 : reg1607)}} ?
                          ($unsigned($unsigned(reg1634)) ?
                              reg1583 : $unsigned((reg1629 ?
                                  wire1518 : reg1590))) : $signed(((8'hb8) ?
                              reg1568 : (forvar1629 <<< forvar1611))));
                    end
                  if ((^~$signed($unsigned(reg1563))))
                    begin
                      reg1544 <= (~&forvar1548[(2'h3):(2'h3)]);
                      reg1545 <= $signed((8'hb2));
                      reg1546 <= (($unsigned((forvar1558 ?
                          reg1576 : forvar1563)) & {(reg1613 && reg1599)}) & (reg1627[(2'h3):(1'h1)] ?
                          $unsigned($unsigned(reg1636)) : $signed($signed(forvar1522))));
                      reg1547 <= reg1534[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1544 <= reg1554;
                      reg1545 <= reg1593;
                      reg1546 <= {$unsigned($signed((reg1595 || reg1566)))};
                    end
                end
            end
        end
      reg1643 <= $unsigned($unsigned($unsigned($unsigned(reg1531))));
    end
  assign wire1644 = ($signed(($unsigned((8'hac)) >>> (reg1630 ?
                        reg1542 : reg1626))) < (^~(wire1520 ?
                        ((8'hb2) != reg1639) : reg1573)));
  assign wire1645 = (~&reg1583);
endmodule
