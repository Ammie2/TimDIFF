module top
#( parameter param151 = (((((~&(8'hbc)) ? ((8'had) ? (8'ha4) : (7'h44)) : ((8'hb4) * (7'h41))) > (8'hb2)) ? {((|(8'hab)) && (-(7'h43)))} : ({((8'h9e) ^ (7'h43))} ? (((8'ha1) ? (8'ha1) : (8'hb5)) ? ((8'hb4) + (8'ha0)) : {(8'hb3)}) : {{(8'ha9)}, ((7'h40) ? (8'hb7) : (8'hb2))})) ? ((~((~&(7'h40)) ? ((8'hba) ? (8'ha6) : (8'h9c)) : (+(8'hb3)))) || (({(8'ha7)} >>> (~&(8'hae))) ? {((8'hb1) <<< (8'hb6)), ((8'hbd) ? (8'hbd) : (8'ha4))} : ((8'hb4) ? ((8'hb5) ^ (8'ha5)) : ((8'hb1) ? (8'hb6) : (8'hbc))))) : (&(((-(8'ha5)) ? (~|(8'hbf)) : {(8'ha5), (8'hb9)}) ~^ (((8'hba) ? (7'h40) : (7'h42)) < ((8'had) ~^ (8'h9c)))))) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h285):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire3;
  input wire [(5'h15):(1'h0)] wire2;
  input wire [(5'h13):(1'h0)] wire1;
  input wire [(5'h14):(1'h0)] wire0;
  wire [(5'h12):(1'h0)] wire150;
  wire signed [(4'hb):(1'h0)] wire149;
  wire [(5'h11):(1'h0)] wire148;
  wire signed [(3'h5):(1'h0)] wire146;
  wire signed [(2'h2):(1'h0)] wire145;
  wire signed [(5'h14):(1'h0)] wire144;
  wire signed [(4'ha):(1'h0)] wire77;
  wire [(5'h14):(1'h0)] wire6;
  wire signed [(5'h13):(1'h0)] wire5;
  wire signed [(5'h11):(1'h0)] wire4;
  wire [(5'h14):(1'h0)] wire79;
  reg signed [(4'h8):(1'h0)] reg80 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg81 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg82 = (1'h0);
  reg [(5'h13):(1'h0)] reg83 = (1'h0);
  reg [(5'h13):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg86 = (1'h0);
  reg [(4'hf):(1'h0)] reg87 = (1'h0);
  reg [(5'h10):(1'h0)] reg88 = (1'h0);
  reg signed [(4'he):(1'h0)] reg89 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg90 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg91 = (1'h0);
  reg [(5'h15):(1'h0)] reg92 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg93 = (1'h0);
  wire [(5'h14):(1'h0)] wire94;
  reg [(3'h7):(1'h0)] reg95 = (1'h0);
  reg [(4'h9):(1'h0)] reg96 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg97 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg98 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg100 = (1'h0);
  reg [(3'h4):(1'h0)] reg101 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg102 = (1'h0);
  reg [(4'ha):(1'h0)] reg103 = (1'h0);
  reg [(5'h10):(1'h0)] reg104 = (1'h0);
  reg [(5'h13):(1'h0)] reg105 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg106 = (1'h0);
  reg [(3'h4):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg108 = (1'h0);
  reg [(5'h12):(1'h0)] reg109 = (1'h0);
  reg [(5'h14):(1'h0)] reg110 = (1'h0);
  reg [(5'h15):(1'h0)] reg111 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg112 = (1'h0);
  reg [(5'h11):(1'h0)] reg113 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire139;
  wire signed [(4'hf):(1'h0)] wire141;
  wire [(4'hd):(1'h0)] wire142;
  assign y = {wire150,
                 wire149,
                 wire148,
                 wire146,
                 wire145,
                 wire144,
                 wire77,
                 wire6,
                 wire5,
                 wire4,
                 wire79,
                 reg80,
                 reg81,
                 reg82,
                 reg83,
                 reg84,
                 reg85,
                 reg86,
                 reg87,
                 reg88,
                 reg89,
                 reg90,
                 reg91,
                 reg92,
                 reg93,
                 wire94,
                 reg95,
                 reg96,
                 reg97,
                 reg98,
                 reg99,
                 reg100,
                 reg101,
                 reg102,
                 reg103,
                 reg104,
                 reg105,
                 reg106,
                 reg107,
                 reg108,
                 reg109,
                 reg110,
                 reg111,
                 reg112,
                 reg113,
                 wire139,
                 wire141,
                 wire142,
                 (1'h0)};
  assign wire4 = {wire2};
  assign wire5 = (wire4[(1'h0):(1'h0)] ? $signed(wire4) : wire3);
  assign wire6 = ((~(^(wire1 ? wire3[(4'ha):(1'h1)] : wire5))) ^~ (wire5 ?
                     {((wire1 ?
                             (8'ha7) : wire0) > $unsigned(wire3))} : ({$signed(wire1),
                             (wire3 == wire0)} ?
                         wire1 : (~^wire1))));
  module7 modinst78 (.wire12(wire0), .wire9(wire1), .y(wire77), .clk(clk), .wire11(wire6), .wire10(wire5), .wire8(wire4));
  assign wire79 = (~|wire6);
  always
    @(posedge clk) begin
      reg80 <= $signed((($signed(wire0[(5'h10):(3'h6)]) & (wire79 <= $signed(wire5))) ?
          {$signed((wire77 <= wire77)),
              $unsigned($signed(wire79))} : (((wire79 ^ wire5) ?
              wire6[(1'h1):(1'h0)] : ((8'hbd) ?
                  wire0 : wire5)) * $signed(((8'ha7) ? wire1 : wire6)))));
      reg81 <= (8'hb4);
      reg82 <= wire77[(4'h9):(3'h7)];
      if (wire5)
        begin
          reg83 <= ($signed(wire5) > ((8'hb3) ?
              wire2 : {((reg81 ~^ (8'ha6)) ?
                      reg80[(4'h8):(4'h8)] : (reg81 ? wire0 : wire3))}));
          reg84 <= reg81[(3'h4):(3'h4)];
          if ((-wire0))
            begin
              reg85 <= ((reg82 ?
                  $signed(($unsigned(wire4) ?
                      (~&wire79) : $unsigned(wire4))) : ($unsigned((+reg82)) ?
                      $unsigned(reg80[(3'h7):(3'h6)]) : $unsigned((^~wire3)))) >> $unsigned(reg84[(4'ha):(3'h6)]));
              reg86 <= ((reg80 <= (($signed(wire6) <<< (8'hae)) << $unsigned($signed(reg85)))) >= reg81[(4'hb):(1'h0)]);
              reg87 <= wire3;
              reg88 <= $signed(reg80);
            end
          else
            begin
              reg85 <= ($signed((wire1 > ((~^wire79) & ((8'ha2) ?
                      wire77 : (8'haa))))) ?
                  ({$signed((8'hb4))} >= $unsigned((8'h9d))) : (~$signed($signed($signed(reg80)))));
              reg86 <= wire77[(2'h2):(2'h2)];
            end
          if (reg80)
            begin
              reg89 <= reg82[(3'h7):(2'h2)];
              reg90 <= $unsigned({$unsigned($unsigned(reg88)), (~&wire77)});
              reg91 <= $signed((|$unsigned(wire4[(3'h5):(2'h3)])));
              reg92 <= $unsigned(({reg88[(4'h8):(3'h4)],
                  ($unsigned(wire4) ? (!wire6) : wire2)} || (reg84 ?
                  ((wire79 ?
                      reg91 : reg80) && $unsigned(reg84)) : (~|$signed((8'ha5))))));
            end
          else
            begin
              reg89 <= $signed($unsigned(reg83[(2'h3):(1'h0)]));
              reg90 <= $unsigned(wire6[(3'h5):(2'h3)]);
              reg91 <= $signed((((~^reg92) ?
                  reg89 : $unsigned($unsigned(wire1))) || $unsigned(reg84)));
              reg92 <= ((($signed({reg88}) ?
                          (|$signed(wire0)) : wire0[(5'h12):(1'h1)]) ?
                      {{(^reg81)}} : ($unsigned(reg88) ? reg82 : (~|reg81))) ?
                  reg91[(3'h5):(1'h1)] : ($unsigned({reg81, $signed(reg80)}) ?
                      reg86[(4'h9):(1'h0)] : $unsigned(($signed(reg84) ?
                          (reg82 || wire4) : {wire0, wire79}))));
            end
          reg93 <= (8'hb3);
        end
      else
        begin
          reg83 <= $unsigned((~|{wire6[(4'hc):(4'hc)], $unsigned(reg93)}));
          if ($unsigned(($unsigned((~$unsigned(wire1))) ?
              $unsigned(($signed(wire0) != (reg89 ?
                  reg81 : (8'hac)))) : (-wire4))))
            begin
              reg84 <= (+(((|wire79) ~^ {(reg87 ^ wire5),
                  {reg87}}) + $unsigned(wire6[(3'h4):(2'h2)])));
              reg85 <= reg90[(4'ha):(4'ha)];
              reg86 <= $signed($signed((~|$signed($unsigned(wire4)))));
            end
          else
            begin
              reg84 <= reg89;
              reg85 <= {(^~wire1[(4'hc):(4'hc)]),
                  (((reg91 != $signed(wire1)) << ((reg86 ? reg92 : reg91) ?
                      (reg86 ?
                          wire1 : reg86) : $signed(reg86))) + $unsigned((|reg80)))};
              reg86 <= (reg84 >>> reg91);
              reg87 <= (wire6[(4'hd):(3'h4)] ?
                  {reg88, $signed(reg86[(4'h9):(1'h0)])} : reg85);
            end
          reg88 <= (reg91 ? wire3[(4'h9):(3'h5)] : (|{reg86}));
          reg89 <= {wire5[(5'h12):(3'h7)],
              (wire1[(4'h8):(4'h8)] ?
                  (((8'h9d) ? $unsigned(reg80) : wire5) ?
                      $signed(((8'hb1) - (8'hb7))) : reg88[(3'h4):(2'h3)]) : ((wire79 ^ (reg90 ^~ (8'hbc))) + $signed(wire1[(1'h1):(1'h0)])))};
        end
    end
  assign wire94 = $signed($unsigned(($unsigned(reg92) | $signed(reg88[(1'h1):(1'h1)]))));
  always
    @(posedge clk) begin
      reg95 <= ((((8'ha6) ? wire0 : {(reg93 ? reg86 : reg83)}) - ((!(wire94 ?
                  reg88 : (8'ha5))) ?
              ($unsigned(reg87) ?
                  reg89[(4'h9):(3'h5)] : {(7'h44)}) : wire94[(4'hd):(3'h4)])) ?
          (-(reg81 ? wire0[(5'h13):(5'h10)] : reg81)) : $unsigned({(!((8'h9d) ?
                  reg86 : wire6))}));
      reg96 <= {$signed((wire77 ?
              $unsigned((reg87 != wire5)) : $signed((wire6 ?
                  (8'hbb) : reg86)))),
          reg80};
      if (reg93)
        begin
          reg97 <= (($signed(((wire3 <= reg82) ?
                  reg89 : $signed(wire79))) - reg87[(1'h0):(1'h0)]) ?
              ($signed(($signed(reg83) <= (reg87 ?
                  reg95 : reg82))) >= wire6) : (({(wire5 ?
                          wire94 : reg93)} <<< (|(reg93 ? (8'hac) : (8'hac)))) ?
                  {(~&(reg95 ? wire77 : reg96))} : (~&(~^{(8'hb1)}))));
          reg98 <= $unsigned((&{$signed($unsigned(wire0)),
              wire3[(4'hf):(4'he)]}));
        end
      else
        begin
          if ($signed({$signed(((wire3 <<< reg93) <= (reg98 ? reg93 : wire2))),
              (wire5[(3'h5):(2'h2)] ? {(8'ha1)} : $signed($signed(reg90)))}))
            begin
              reg97 <= (~|wire4);
              reg98 <= wire4[(3'h7):(3'h7)];
              reg99 <= {(reg93[(1'h1):(1'h0)] || reg95[(2'h2):(2'h2)])};
              reg100 <= $signed(reg90[(3'h6):(2'h2)]);
              reg101 <= $unsigned(({reg97, reg88} ?
                  $unsigned($unsigned((~|reg99))) : $unsigned((wire77[(1'h1):(1'h1)] ?
                      (^reg82) : wire1))));
            end
          else
            begin
              reg97 <= {({((-reg86) - (reg90 >> wire4)),
                      (reg86[(1'h0):(1'h0)] ^~ $signed(reg88))} * reg82),
                  (+($unsigned((-wire5)) ? {wire6, reg97} : (!(~wire5))))};
              reg98 <= ((-(+($signed(reg89) ~^ (wire79 && reg80)))) * (~^(8'hbf)));
              reg99 <= (+$signed(($signed(wire2) ?
                  (wire4 ?
                      {reg100,
                          reg100} : (wire6 || reg85)) : (reg82 && reg88))));
              reg100 <= $unsigned($signed(($unsigned($signed(wire1)) ?
                  (wire79[(2'h3):(2'h2)] + $signed(reg82)) : ($unsigned((8'ha0)) < (8'ha1)))));
              reg101 <= reg95[(1'h1):(1'h0)];
            end
          reg102 <= ((-{((~|reg81) ?
                      (reg91 ? (8'hb6) : wire6) : (~&(8'ha2)))}) ?
              ($signed((!reg96)) ?
                  $signed({$signed((8'hbb)),
                      (reg98 ? reg86 : wire2)}) : ($signed($signed((8'hae))) ?
                      $unsigned((~^reg101)) : $signed(reg89[(3'h5):(1'h0)]))) : (8'h9c));
          if (reg84)
            begin
              reg103 <= reg99;
            end
          else
            begin
              reg103 <= $unsigned((~^reg102[(1'h0):(1'h0)]));
              reg104 <= $signed({wire6[(5'h13):(5'h11)]});
              reg105 <= $unsigned((~|(^~reg103[(4'h9):(4'h8)])));
              reg106 <= reg98;
            end
          reg107 <= (~|(($unsigned($signed(reg104)) ?
              (~^(8'hac)) : reg104[(2'h3):(1'h1)]) ^~ $signed($signed(reg105[(4'ha):(3'h7)]))));
          reg108 <= (wire0[(5'h10):(3'h6)] - (((+reg91[(3'h7):(2'h3)]) > reg98[(3'h5):(3'h4)]) ?
              $unsigned($unsigned($unsigned(reg86))) : {$signed(wire5),
                  reg92}));
        end
      if (reg101)
        begin
          reg109 <= $signed((~|(-(+reg103[(4'h8):(1'h1)]))));
          reg110 <= $signed((~^(~&(+reg98[(4'hd):(4'h8)]))));
        end
      else
        begin
          if ((^~(~&$unsigned(($signed(reg104) >>> wire5)))))
            begin
              reg109 <= reg90[(3'h7):(2'h3)];
            end
          else
            begin
              reg109 <= (~((8'h9d) <= reg102));
              reg110 <= (-reg80[(4'h8):(2'h2)]);
            end
          reg111 <= ({$unsigned((wire77[(2'h2):(2'h2)] ^~ $unsigned(wire3))),
                  $unsigned((^reg91[(2'h3):(1'h0)]))} ?
              (reg83[(5'h10):(4'hb)] <= reg106) : reg104[(3'h6):(1'h0)]);
          reg112 <= (&(reg104 + (reg108[(4'he):(3'h7)] <= (reg105[(4'hb):(4'ha)] ?
              (reg93 ? reg96 : wire4) : (reg97 << reg80)))));
        end
      reg113 <= $signed(reg111);
    end
  module114 modinst140 (wire139, clk, reg89, reg111, reg88, wire2);
  assign wire141 = {((reg97 >= $signed($unsigned(reg100))) >> wire6[(1'h0):(1'h0)])};
  module19 modinst143 (.clk(clk), .wire24(wire4), .wire20(reg86), .wire21(reg110), .y(wire142), .wire22(reg113), .wire23(reg103));
  assign wire144 = reg81;
  assign wire145 = reg103;
  module114 modinst147 (.y(wire146), .wire115(reg92), .wire116(reg104), .wire117(reg109), .clk(clk), .wire118(reg110));
  assign wire148 = {(|reg80)};
  assign wire149 = (($signed($signed($signed(reg95))) << ((~$unsigned(reg99)) ?
                       (wire142[(3'h5):(2'h3)] >> reg83[(4'he):(3'h5)]) : reg112[(2'h2):(2'h2)])) | (reg113 >> $signed($unsigned(reg98[(4'hd):(2'h3)]))));
  assign wire150 = ($unsigned((wire148 < reg91)) ?
                       (|$unsigned($unsigned((|(8'hae))))) : wire94);
endmodule

module module114
#( parameter param138 = ({({{(8'haf), (8'hb6)}, ((8'hb5) ? (8'hbc) : (8'h9e))} ? (+(-(7'h42))) : {(~^(8'hbc)), {(8'hbc), (8'hb0)}}), ((~^(|(8'hbd))) && {{(8'h9e)}})} ^~ ((((~&(8'ha4)) * ((8'had) == (8'ha4))) ? ((8'ha3) ? {(8'ha3)} : {(8'ha6), (8'hb0)}) : (^~(~|(7'h41)))) << ((^~(^~(8'hb9))) ? {{(8'h9c), (8'ha6)}, ((7'h40) > (8'hb8))} : (((8'ha5) ? (8'hab) : (8'hb2)) & ((7'h43) ? (8'haa) : (8'hbd)))))) )
(y, clk, wire118, wire117, wire116, wire115);
  output wire [(32'h40):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire118;
  input wire signed [(5'h11):(1'h0)] wire117;
  input wire [(5'h10):(1'h0)] wire116;
  input wire signed [(5'h15):(1'h0)] wire115;
  wire [(4'hd):(1'h0)] wire137;
  wire signed [(4'hc):(1'h0)] wire136;
  wire [(5'h15):(1'h0)] wire135;
  wire signed [(5'h11):(1'h0)] wire133;
  assign y = {wire137, wire136, wire135, wire133, (1'h0)};
  module119 modinst134 (wire133, clk, wire115, wire116, wire117, wire118, (8'ha5));
  assign wire135 = (~(({(^wire133), (wire115 << wire116)} ?
                       (~&(wire115 ?
                           wire118 : wire115)) : $unsigned((wire115 ~^ wire118))) == (wire116 ?
                       $unsigned({wire118, wire116}) : wire118)));
  assign wire136 = $signed({wire117,
                       {wire116[(4'h9):(4'h8)], $unsigned(wire115)}});
  assign wire137 = $unsigned(wire135);
endmodule

module module7
#( parameter param76 = (((+(8'ha5)) ^~ {{((7'h43) ^~ (8'ha0)), (+(8'hb8))}, ((|(8'ha5)) ? ((8'hac) * (8'hbc)) : ((7'h40) ? (8'ha5) : (8'hbe)))}) ? (8'ha2) : (~{(~&((8'hb8) ? (8'had) : (8'ha2)))})) )
(y, clk, wire8, wire9, wire10, wire11, wire12);
  output wire [(32'h107):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire8;
  input wire signed [(4'h8):(1'h0)] wire9;
  input wire [(5'h13):(1'h0)] wire10;
  input wire [(5'h14):(1'h0)] wire11;
  input wire signed [(5'h14):(1'h0)] wire12;
  wire [(4'hc):(1'h0)] wire75;
  wire [(5'h10):(1'h0)] wire74;
  wire [(5'h14):(1'h0)] wire73;
  wire signed [(5'h11):(1'h0)] wire72;
  wire [(4'h8):(1'h0)] wire71;
  wire signed [(5'h13):(1'h0)] wire69;
  reg signed [(4'h8):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg54 = (1'h0);
  wire [(5'h15):(1'h0)] wire53;
  wire [(3'h7):(1'h0)] wire52;
  wire signed [(4'hd):(1'h0)] wire51;
  wire [(3'h5):(1'h0)] wire50;
  reg [(3'h4):(1'h0)] reg49 = (1'h0);
  wire [(4'hd):(1'h0)] wire13;
  wire [(2'h3):(1'h0)] wire14;
  wire signed [(5'h11):(1'h0)] wire15;
  wire [(5'h11):(1'h0)] wire16;
  wire [(5'h10):(1'h0)] wire17;
  wire [(5'h14):(1'h0)] wire18;
  wire signed [(5'h15):(1'h0)] wire47;
  assign y = {wire75,
                 wire74,
                 wire73,
                 wire72,
                 wire71,
                 wire69,
                 reg55,
                 reg54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 reg49,
                 wire13,
                 wire14,
                 wire15,
                 wire16,
                 wire17,
                 wire18,
                 wire47,
                 (1'h0)};
  assign wire13 = wire11[(1'h0):(1'h0)];
  assign wire14 = wire9[(2'h3):(1'h0)];
  assign wire15 = $signed(($unsigned((|(wire10 && wire8))) ?
                      wire9 : (^$signed({wire9, wire10}))));
  assign wire16 = (&$signed(wire9));
  assign wire17 = ($signed($unsigned($signed((+wire12)))) ^ wire15[(3'h5):(2'h3)]);
  assign wire18 = $signed((wire17 << (!((wire16 ? wire10 : wire16) ^~ (wire10 ?
                      wire14 : wire8)))));
  module19 modinst48 (wire47, clk, wire16, wire17, wire15, wire11, wire10);
  always
    @(posedge clk) begin
      reg49 <= $signed($signed(wire16[(3'h4):(2'h2)]));
    end
  assign wire50 = $unsigned($signed(($signed(wire12) ?
                      ((wire18 ? wire17 : wire10) ?
                          (~wire9) : wire8) : (~&(wire16 >>> wire18)))));
  assign wire51 = $unsigned(wire14[(2'h2):(1'h0)]);
  assign wire52 = $unsigned((~^wire9));
  assign wire53 = wire16;
  always
    @(posedge clk) begin
      reg54 <= $unsigned($unsigned(($signed((~^reg49)) + $signed($signed(wire15)))));
      reg55 <= {wire13,
          ($unsigned(wire17) ?
              (wire14 ^ (wire16 >>> (wire53 ?
                  wire13 : wire12))) : (&wire47[(4'h9):(3'h4)]))};
    end
  module56 modinst70 (wire69, clk, wire16, wire52, wire47, wire53);
  assign wire71 = reg54;
  assign wire72 = {$unsigned(($unsigned((~^wire10)) + wire15))};
  assign wire73 = (+(&((-(-wire51)) >> $signed($unsigned(wire8)))));
  assign wire74 = {wire16[(3'h4):(2'h2)], $unsigned(wire10)};
  assign wire75 = ((~^wire17) <<< (^$signed(wire69)));
endmodule

module module56
#( parameter param67 = ((((8'h9f) ? {((8'h9d) == (8'ha4)), ((8'hbc) >= (8'hbe))} : ({(7'h41)} >>> ((8'hbc) << (8'hbb)))) ^~ (&({(8'hbd)} ? (|(8'h9f)) : ((8'ha9) ? (8'hb9) : (8'hb6))))) ? (((!(8'hb0)) == {((8'hb1) ? (8'ha0) : (8'ha4)), (~&(8'ha5))}) ? (^~{((8'hbe) ? (8'h9c) : (8'hbd))}) : ((~&(^~(8'haf))) == ((&(8'hb8)) <= ((8'hb7) >> (8'hb9))))) : (!(8'ha8)))
, parameter param68 = ((((|(!param67)) ? (~&(!param67)) : ((param67 ? param67 : param67) ? param67 : (param67 ? param67 : param67))) == ({(param67 ? param67 : param67)} ? (param67 || ((8'h9d) <<< param67)) : ((param67 >> param67) >> param67))) + param67) )
(y, clk, wire60, wire59, wire58, wire57);
  output wire [(32'h4e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire60;
  input wire signed [(3'h7):(1'h0)] wire59;
  input wire signed [(5'h15):(1'h0)] wire58;
  input wire [(2'h2):(1'h0)] wire57;
  wire signed [(5'h12):(1'h0)] wire66;
  wire [(5'h10):(1'h0)] wire65;
  wire signed [(4'h9):(1'h0)] wire64;
  wire [(5'h11):(1'h0)] wire63;
  wire signed [(3'h5):(1'h0)] wire62;
  wire signed [(4'hc):(1'h0)] wire61;
  assign y = {wire66, wire65, wire64, wire63, wire62, wire61, (1'h0)};
  assign wire61 = ($signed($signed($unsigned((wire60 || wire58)))) ^~ $unsigned((~|(wire59 <= {wire59}))));
  assign wire62 = $unsigned($unsigned(wire60[(3'h4):(2'h3)]));
  assign wire63 = (wire58 || $signed($signed(((~wire57) != (~wire61)))));
  assign wire64 = (($unsigned(wire60) << $signed(((8'ha1) ?
                      (wire61 > wire58) : (-wire62)))) ^~ $signed((wire60 ?
                      ((~^wire60) <<< (^~(8'hb4))) : (8'hb2))));
  assign wire65 = $signed(wire57[(1'h0):(1'h0)]);
  assign wire66 = ({(^wire65[(3'h4):(1'h1)])} + wire62);
endmodule

module module19  (y, clk, wire24, wire23, wire22, wire21, wire20);
  output wire [(32'hf6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire24;
  input wire signed [(4'ha):(1'h0)] wire23;
  input wire signed [(5'h11):(1'h0)] wire22;
  input wire [(5'h14):(1'h0)] wire21;
  input wire signed [(5'h13):(1'h0)] wire20;
  reg [(4'h9):(1'h0)] reg46 = (1'h0);
  reg [(4'hb):(1'h0)] reg45 = (1'h0);
  reg [(3'h4):(1'h0)] reg44 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg43 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg42 = (1'h0);
  reg [(3'h7):(1'h0)] reg41 = (1'h0);
  reg [(3'h7):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg39 = (1'h0);
  reg [(5'h12):(1'h0)] reg38 = (1'h0);
  wire [(3'h4):(1'h0)] wire37;
  wire signed [(5'h10):(1'h0)] wire36;
  wire signed [(4'hf):(1'h0)] wire35;
  wire signed [(4'h8):(1'h0)] wire34;
  wire [(3'h7):(1'h0)] wire33;
  wire signed [(2'h2):(1'h0)] wire32;
  reg signed [(5'h15):(1'h0)] reg31 = (1'h0);
  reg [(4'ha):(1'h0)] reg30 = (1'h0);
  reg [(4'hc):(1'h0)] reg29 = (1'h0);
  reg [(3'h7):(1'h0)] reg28 = (1'h0);
  reg [(5'h10):(1'h0)] reg27 = (1'h0);
  reg [(5'h14):(1'h0)] reg26 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire25;
  assign y = {reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 wire37,
                 wire36,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 wire25,
                 (1'h0)};
  assign wire25 = $unsigned($signed(wire22[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      reg26 <= wire21;
      reg27 <= wire24;
      reg28 <= (^$unsigned((^~reg26)));
      reg29 <= $unsigned((&$signed(wire20[(3'h5):(2'h2)])));
    end
  always
    @(posedge clk) begin
      reg30 <= $unsigned((wire24[(2'h3):(2'h3)] ?
          (^(reg27[(4'hc):(3'h7)] <= (reg29 == wire23))) : $unsigned($signed($signed(wire23)))));
      reg31 <= ((wire23 ?
          reg26 : wire23[(3'h7):(1'h1)]) && $unsigned(wire21[(4'hf):(4'ha)]));
    end
  assign wire32 = wire25;
  assign wire33 = (^(reg30[(4'h9):(4'h9)] >> (8'hbb)));
  assign wire34 = reg27;
  assign wire35 = (+reg26[(3'h4):(3'h4)]);
  assign wire36 = (|wire21[(4'h8):(1'h1)]);
  assign wire37 = reg31;
  always
    @(posedge clk) begin
      reg38 <= {{wire33}};
      reg39 <= $signed({({wire22, {wire36}} ?
              (|wire33) : wire25[(1'h1):(1'h1)]),
          (^wire24[(4'he):(4'h9)])});
      if ($unsigned(wire36[(3'h5):(1'h0)]))
        begin
          if ((((wire21[(4'hd):(3'h4)] ?
                  ((reg28 < reg38) >> wire35[(3'h4):(1'h0)]) : $unsigned($unsigned(wire23))) & reg28) ?
              ((reg39[(4'hf):(4'hf)] ?
                      (|((8'ha7) ? wire20 : reg30)) : $unsigned((~|wire32))) ?
                  reg30 : $signed(((&reg29) ?
                      $signed((8'hb5)) : $signed((8'ha9))))) : (($unsigned(wire25) * reg38[(2'h2):(1'h1)]) - $unsigned((8'ha8)))))
            begin
              reg40 <= $signed($signed(wire23));
            end
          else
            begin
              reg40 <= (wire22[(1'h0):(1'h0)] ?
                  ($signed((-$unsigned(reg26))) + (~(reg27 ?
                      {(8'hba)} : wire21[(4'he):(4'hd)]))) : $unsigned(reg29[(2'h3):(1'h1)]));
              reg41 <= {(wire33 != {wire32[(1'h0):(1'h0)],
                      (reg39 > (reg29 && wire36))}),
                  {$signed(wire33),
                      $signed((wire35 ? (~&(8'hbe)) : ((8'hbe) * reg38)))}};
            end
        end
      else
        begin
          reg40 <= (wire32[(2'h2):(2'h2)] == $unsigned($signed((wire25[(2'h3):(1'h1)] ?
              (reg27 == wire25) : (wire37 ? reg29 : (8'hb9))))));
        end
      reg42 <= (((8'hbf) != (~&$unsigned(((8'ha8) ?
          reg39 : reg26)))) <= (~|{{reg29, (wire22 || wire23)}}));
      reg43 <= (reg39 != $signed((!($signed(reg42) <= $signed(reg31)))));
    end
  always
    @(posedge clk) begin
      reg44 <= (reg27 & $signed((reg26 ~^ {$signed(reg29), {wire36, reg27}})));
      reg45 <= wire23;
      reg46 <= (-(8'hb4));
    end
endmodule

module module119  (y, clk, wire124, wire123, wire122, wire121, wire120);
  output wire [(32'h59):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire124;
  input wire [(5'h10):(1'h0)] wire123;
  input wire signed [(5'h11):(1'h0)] wire122;
  input wire signed [(4'hd):(1'h0)] wire121;
  input wire [(5'h15):(1'h0)] wire120;
  wire signed [(2'h2):(1'h0)] wire132;
  wire signed [(4'he):(1'h0)] wire131;
  wire [(5'h10):(1'h0)] wire130;
  wire signed [(4'hf):(1'h0)] wire129;
  wire signed [(2'h3):(1'h0)] wire128;
  reg signed [(5'h15):(1'h0)] reg127 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg126 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire125;
  assign y = {wire132,
                 wire131,
                 wire130,
                 wire129,
                 wire128,
                 reg127,
                 reg126,
                 wire125,
                 (1'h0)};
  assign wire125 = (wire120 & ((($signed(wire124) >= (wire124 + wire120)) ?
                           ($signed(wire121) ?
                               wire121[(4'hb):(4'h8)] : $unsigned(wire124)) : $signed(wire121[(3'h4):(2'h3)])) ?
                       ($signed(wire122) + (8'hb1)) : {$signed((^wire121))}));
  always
    @(posedge clk) begin
      reg126 <= wire120;
      reg127 <= (($signed((wire123 && (~&wire121))) ?
          {{$signed((8'haa))},
              wire123} : (-((^reg126) & reg126[(2'h2):(1'h1)]))) && $signed(wire124));
    end
  assign wire128 = reg127[(2'h2):(1'h1)];
  assign wire129 = {reg127,
                       $unsigned((($unsigned(reg127) ?
                           (8'ha1) : (^~wire124)) ^~ wire122[(3'h4):(1'h1)]))};
  assign wire130 = $unsigned(wire120);
  assign wire131 = $signed((wire121 ?
                       wire123 : (^$unsigned($signed(wire121)))));
  assign wire132 = {(($signed(wire120) == (((8'hb0) <= wire131) >>> (wire121 ^ wire129))) <= (wire123 ?
                           $signed(wire125[(3'h6):(1'h1)]) : wire123))};
endmodule