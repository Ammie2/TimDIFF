(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param7783 = (^~(-(((8'hb9) & (8'ha9)) ? {(8'ha4)} : {(8'hb8)}))))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h6e6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire3;
  input wire signed [(4'h8):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire1;
  input wire [(5'h10):(1'h0)] wire0;
  wire signed [(3'h4):(1'h0)] wire7782;
  reg signed [(3'h4):(1'h0)] forvar7769 = (1'h0);
  reg [(4'ha):(1'h0)] reg7768 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7764 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7761 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7766 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7765 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7762 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7760 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7756 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7755 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7754 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar7749 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7746 = (1'h0);
  reg [(3'h7):(1'h0)] forvar7744 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7780 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7777 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7781 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7780 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7779 = (1'h0);
  reg [(5'h10):(1'h0)] reg7778 = (1'h0);
  reg [(5'h10):(1'h0)] reg7777 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7776 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7775 = (1'h0);
  reg [(4'h8):(1'h0)] reg7774 = (1'h0);
  reg [(2'h3):(1'h0)] reg7773 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7772 = (1'h0);
  reg [(3'h7):(1'h0)] reg7771 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7770 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7770 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7769 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7768 = (1'h0);
  reg [(4'ha):(1'h0)] reg7767 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7766 = (1'h0);
  reg [(4'he):(1'h0)] reg7765 = (1'h0);
  reg [(4'ha):(1'h0)] reg7764 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7763 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7762 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7761 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7760 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7759 = (1'h0);
  reg [(4'hf):(1'h0)] reg7758 = (1'h0);
  reg [(5'h10):(1'h0)] reg7757 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7756 = (1'h0);
  reg [(3'h6):(1'h0)] reg7755 = (1'h0);
  reg [(4'h9):(1'h0)] forvar7748 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7754 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7753 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7752 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7751 = (1'h0);
  reg [(3'h5):(1'h0)] reg7750 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7749 = (1'h0);
  reg [(3'h4):(1'h0)] reg7748 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7747 = (1'h0);
  reg [(3'h5):(1'h0)] forvar7746 = (1'h0);
  reg [(3'h5):(1'h0)] forvar7745 = (1'h0);
  reg [(2'h3):(1'h0)] reg7744 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7629 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7743 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7742 = (1'h0);
  reg [(4'hb):(1'h0)] reg7741 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7740 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7739 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7738 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7737 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7736 = (1'h0);
  reg [(3'h7):(1'h0)] reg7735 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar7734 = (1'h0);
  reg [(4'hb):(1'h0)] reg7733 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7732 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7731 = (1'h0);
  reg [(4'he):(1'h0)] reg7730 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7729 = (1'h0);
  reg [(4'hf):(1'h0)] reg7728 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7727 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7726 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7725 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7724 = (1'h0);
  reg [(4'he):(1'h0)] reg7723 = (1'h0);
  reg [(4'h8):(1'h0)] reg7722 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7721 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7720 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7719 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7718 = (1'h0);
  reg [(4'hc):(1'h0)] reg7717 = (1'h0);
  reg [(4'hc):(1'h0)] reg7716 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7715 = (1'h0);
  reg [(3'h7):(1'h0)] reg7714 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7713 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7712 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7711 = (1'h0);
  reg [(2'h2):(1'h0)] forvar7710 = (1'h0);
  reg [(2'h3):(1'h0)] reg7709 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7708 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7707 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7706 = (1'h0);
  reg [(2'h2):(1'h0)] reg7705 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7704 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7703 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7702 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7701 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7700 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7699 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7698 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7697 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7696 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7695 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7686 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7683 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7682 = (1'h0);
  reg [(4'hc):(1'h0)] reg7694 = (1'h0);
  reg [(4'hd):(1'h0)] reg7693 = (1'h0);
  reg [(3'h7):(1'h0)] reg7692 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7691 = (1'h0);
  reg [(3'h5):(1'h0)] reg7690 = (1'h0);
  reg [(4'hb):(1'h0)] reg7689 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7688 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7687 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar7686 = (1'h0);
  reg [(2'h3):(1'h0)] reg7685 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7684 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7683 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7682 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7681 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7680 = (1'h0);
  reg [(4'he):(1'h0)] reg7679 = (1'h0);
  reg [(3'h7):(1'h0)] reg7678 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7677 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7674 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7672 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7670 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7668 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7667 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7665 = (1'h0);
  reg [(5'h10):(1'h0)] reg7677 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7676 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7675 = (1'h0);
  reg [(5'h10):(1'h0)] reg7674 = (1'h0);
  reg [(4'h9):(1'h0)] reg7673 = (1'h0);
  reg [(3'h5):(1'h0)] forvar7672 = (1'h0);
  reg [(4'h8):(1'h0)] reg7671 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7670 = (1'h0);
  reg [(4'h9):(1'h0)] reg7669 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7668 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7667 = (1'h0);
  reg [(3'h7):(1'h0)] reg7666 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7665 = (1'h0);
  reg [(2'h2):(1'h0)] reg7664 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7663 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7662 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7661 = (1'h0);
  reg [(5'h10):(1'h0)] forvar7633 = (1'h0);
  reg [(4'hf):(1'h0)] reg7632 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7630 = (1'h0);
  reg [(5'h10):(1'h0)] reg7660 = (1'h0);
  reg [(4'ha):(1'h0)] reg7659 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7658 = (1'h0);
  reg [(2'h3):(1'h0)] reg7657 = (1'h0);
  reg [(4'hb):(1'h0)] reg7656 = (1'h0);
  reg [(4'hb):(1'h0)] reg7655 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7654 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar7653 = (1'h0);
  reg [(4'h8):(1'h0)] reg7652 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7651 = (1'h0);
  reg [(3'h6):(1'h0)] reg7650 = (1'h0);
  reg [(4'hd):(1'h0)] reg7649 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7648 = (1'h0);
  reg [(4'he):(1'h0)] reg7647 = (1'h0);
  reg [(5'h10):(1'h0)] reg7643 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7640 = (1'h0);
  reg [(4'ha):(1'h0)] reg7646 = (1'h0);
  reg [(4'hd):(1'h0)] reg7645 = (1'h0);
  reg [(2'h3):(1'h0)] reg7644 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7643 = (1'h0);
  reg [(4'hf):(1'h0)] reg7642 = (1'h0);
  reg [(3'h6):(1'h0)] reg7641 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7640 = (1'h0);
  reg [(3'h5):(1'h0)] reg7639 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7638 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7637 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7636 = (1'h0);
  reg [(5'h10):(1'h0)] reg7635 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7634 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7633 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7632 = (1'h0);
  reg [(4'hd):(1'h0)] reg7631 = (1'h0);
  reg [(3'h6):(1'h0)] reg7630 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7629 = (1'h0);
  wire [(2'h2):(1'h0)] wire7628;
  reg [(3'h4):(1'h0)] reg7627 = (1'h0);
  wire [(4'h8):(1'h0)] wire7625;
  wire signed [(3'h6):(1'h0)] wire618;
  wire [(4'ha):(1'h0)] wire5;
  wire [(5'h10):(1'h0)] wire4;
  assign y = {wire7782,
                 forvar7769,
                 reg7768,
                 forvar7764,
                 forvar7761,
                 reg7766,
                 forvar7765,
                 forvar7762,
                 reg7760,
                 reg7756,
                 forvar7755,
                 forvar7754,
                 forvar7749,
                 reg7746,
                 forvar7744,
                 reg7780,
                 forvar7777,
                 reg7781,
                 forvar7780,
                 reg7779,
                 reg7778,
                 reg7777,
                 reg7776,
                 reg7775,
                 reg7774,
                 reg7773,
                 forvar7772,
                 reg7771,
                 forvar7770,
                 reg7770,
                 reg7769,
                 forvar7768,
                 reg7767,
                 forvar7766,
                 reg7765,
                 reg7764,
                 reg7763,
                 reg7762,
                 reg7761,
                 forvar7760,
                 reg7759,
                 reg7758,
                 reg7757,
                 forvar7756,
                 reg7755,
                 forvar7748,
                 reg7754,
                 reg7753,
                 reg7752,
                 reg7751,
                 reg7750,
                 reg7749,
                 reg7748,
                 reg7747,
                 forvar7746,
                 forvar7745,
                 reg7744,
                 reg7629,
                 reg7743,
                 reg7742,
                 reg7741,
                 forvar7740,
                 reg7739,
                 reg7738,
                 reg7737,
                 forvar7736,
                 reg7735,
                 forvar7734,
                 reg7733,
                 reg7732,
                 reg7731,
                 reg7730,
                 forvar7729,
                 reg7728,
                 reg7727,
                 reg7726,
                 reg7725,
                 forvar7724,
                 reg7723,
                 reg7722,
                 reg7721,
                 reg7720,
                 reg7719,
                 reg7718,
                 reg7717,
                 reg7716,
                 reg7715,
                 reg7714,
                 forvar7713,
                 reg7712,
                 forvar7711,
                 forvar7710,
                 reg7709,
                 reg7708,
                 forvar7707,
                 reg7706,
                 reg7705,
                 forvar7704,
                 reg7703,
                 reg7702,
                 reg7701,
                 reg7700,
                 forvar7699,
                 forvar7698,
                 reg7697,
                 reg7696,
                 forvar7695,
                 reg7686,
                 forvar7683,
                 reg7682,
                 reg7694,
                 reg7693,
                 reg7692,
                 reg7691,
                 reg7690,
                 reg7689,
                 reg7688,
                 reg7687,
                 forvar7686,
                 reg7685,
                 reg7684,
                 reg7683,
                 forvar7682,
                 reg7681,
                 reg7680,
                 reg7679,
                 reg7678,
                 forvar7677,
                 forvar7674,
                 reg7672,
                 forvar7670,
                 reg7668,
                 reg7667,
                 forvar7665,
                 reg7677,
                 reg7676,
                 reg7675,
                 reg7674,
                 reg7673,
                 forvar7672,
                 reg7671,
                 reg7670,
                 reg7669,
                 forvar7668,
                 forvar7667,
                 reg7666,
                 reg7665,
                 reg7664,
                 reg7663,
                 reg7662,
                 forvar7661,
                 forvar7633,
                 reg7632,
                 forvar7630,
                 reg7660,
                 reg7659,
                 reg7658,
                 reg7657,
                 reg7656,
                 reg7655,
                 forvar7654,
                 forvar7653,
                 reg7652,
                 forvar7651,
                 reg7650,
                 reg7649,
                 reg7648,
                 reg7647,
                 reg7643,
                 forvar7640,
                 reg7646,
                 reg7645,
                 reg7644,
                 forvar7643,
                 reg7642,
                 reg7641,
                 reg7640,
                 reg7639,
                 reg7638,
                 reg7637,
                 reg7636,
                 reg7635,
                 reg7634,
                 reg7633,
                 forvar7632,
                 reg7631,
                 reg7630,
                 forvar7629,
                 wire7628,
                 reg7627,
                 wire7625,
                 wire618,
                 wire5,
                 wire4,
                 (1'h0)};
  assign wire4 = (-$signed((!((8'hb9) ? wire1 : wire3))));
  assign wire5 = wire1[(1'h1):(1'h1)];
  module6 modinst619 (wire618, clk, wire4, wire3, wire1, wire5);
  module620 modinst7626 (wire7625, clk, wire4, wire0, wire3, wire1);
  always
    @(posedge clk) begin
      reg7627 <= (~(~$unsigned((^~wire618))));
    end
  assign wire7628 = wire2[(3'h4):(2'h2)];
  always
    @(posedge clk) begin
      if (($signed(($unsigned(wire618) == wire618[(1'h1):(1'h0)])) * wire7625))
        begin
          if ((^~$unsigned($signed((wire0 ? wire0 : wire0)))))
            begin
              for (forvar7629 = (1'h0); (forvar7629 < (2'h3)); forvar7629 = (forvar7629 + (1'h1)))
                begin
                  if ($unsigned(forvar7629))
                    begin
                      reg7630 <= ((!(~|wire2[(4'h8):(3'h4)])) <= {(reg7627[(2'h3):(2'h3)] || $signed(wire2))});
                      reg7631 <= (wire7625[(3'h5):(1'h0)] ?
                          $signed($unsigned({(8'h9f)})) : (~^((reg7630 ?
                              wire2 : wire0) > wire1)));
                    end
                  else
                    begin
                      reg7630 <= $unsigned((($signed((8'hab)) ~^ (reg7631 >>> forvar7629)) | wire618[(1'h0):(1'h0)]));
                      reg7631 <= ((|wire4) ?
                          ((~^wire4[(4'hf):(3'h5)]) ?
                              (~&$unsigned(reg7630)) : $signed(wire7625[(1'h0):(1'h0)])) : {wire4});
                    end
                  for (forvar7632 = (1'h0); (forvar7632 < (1'h0)); forvar7632 = (forvar7632 + (1'h1)))
                    begin
                      reg7633 <= forvar7632;
                      reg7634 <= $unsigned((~^((wire4 * wire618) >>> (~|reg7627))));
                    end
                  reg7635 <= $unsigned($unsigned((^(+reg7627))));
                  if (wire2)
                    begin
                      reg7636 <= (reg7635[(4'h9):(4'h9)] ?
                          (!(8'hb0)) : reg7631[(2'h2):(1'h0)]);
                      reg7637 <= {((|(reg7634 ?
                              (8'hae) : reg7636)) > wire5[(3'h7):(3'h4)])};
                    end
                  else
                    begin
                      reg7636 <= {((8'hb8) - $unsigned(reg7637[(1'h1):(1'h1)]))};
                      reg7637 <= wire5;
                      reg7638 <= (-$unsigned({{reg7633}}));
                      reg7639 <= $signed((((|forvar7629) >= (wire618 && (8'hb0))) ?
                          forvar7632[(1'h1):(1'h0)] : ((reg7633 >> reg7637) <= wire7628[(1'h1):(1'h0)])));
                    end
                end
              if ((^~$signed($signed({forvar7629}))))
                begin
                  if (reg7631[(3'h4):(1'h1)])
                    begin
                      reg7640 <= (&($signed((&reg7635)) <= $signed({wire5})));
                      reg7641 <= $unsigned((~(-forvar7632)));
                      reg7642 <= $unsigned((wire7625 || reg7627[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg7640 <= {reg7641};
                      reg7641 <= ($signed((+$signed((8'hb5)))) <= wire0);
                    end
                  for (forvar7643 = (1'h0); (forvar7643 < (2'h3)); forvar7643 = (forvar7643 + (1'h1)))
                    begin
                      reg7644 <= ($signed((reg7635 ?
                          {wire2} : wire2[(2'h3):(2'h3)])) ^ (-$unsigned(reg7634[(2'h2):(2'h2)])));
                      reg7645 <= $unsigned({(~|(~^wire7625))});
                      reg7646 <= forvar7643[(3'h6):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar7640 = (1'h0); (forvar7640 < (1'h1)); forvar7640 = (forvar7640 + (1'h1)))
                    begin
                      reg7641 <= $signed(forvar7643);
                    end
                  if ($unsigned((|($unsigned(wire1) - ((8'hb0) + wire7628)))))
                    begin
                      reg7642 <= ((({wire3} != (wire1 ?
                          reg7639 : reg7637)) ^ wire4[(2'h2):(1'h1)]) * ($signed(reg7646[(2'h2):(2'h2)]) * forvar7632[(2'h2):(2'h2)]));
                      reg7643 <= forvar7632[(1'h1):(1'h0)];
                      reg7644 <= {$unsigned(wire7625)};
                      reg7645 <= $signed($unsigned($signed(reg7630)));
                    end
                  else
                    begin
                      reg7642 <= {$signed(reg7644[(1'h1):(1'h0)])};
                      reg7643 <= wire618;
                      reg7644 <= reg7646[(4'ha):(1'h0)];
                    end
                  reg7646 <= (((8'hb0) ? reg7630[(3'h5):(2'h3)] : wire7628) ?
                      wire3 : $signed(((+wire0) ?
                          $unsigned((8'hb7)) : {(8'h9d)})));
                  if ((+reg7641[(1'h1):(1'h1)]))
                    begin
                      reg7647 <= ({$unsigned(reg7643[(1'h1):(1'h1)])} > $signed(((reg7634 ?
                              wire2 : wire618) ?
                          $signed((8'haa)) : reg7644)));
                      reg7648 <= ({reg7642[(1'h0):(1'h0)]} > reg7646);
                      reg7649 <= (^reg7646);
                      reg7650 <= (~^$unsigned(((reg7636 ?
                          reg7627 : reg7638) ~^ (reg7647 && (8'hab)))));
                    end
                  else
                    begin
                      reg7647 <= (+$signed($signed($signed(wire4))));
                      reg7648 <= $unsigned($unsigned(wire7625[(3'h7):(2'h3)]));
                      reg7649 <= $unsigned(wire5);
                    end
                end
              for (forvar7651 = (1'h0); (forvar7651 < (2'h2)); forvar7651 = (forvar7651 + (1'h1)))
                begin
                  if ($unsigned($signed($unsigned($signed((8'had))))))
                    begin
                      reg7652 <= (~$signed($unsigned((&reg7633))));
                    end
                  else
                    begin
                      reg7652 <= reg7649[(3'h7):(3'h5)];
                    end
                end
              for (forvar7653 = (1'h0); (forvar7653 < (2'h3)); forvar7653 = (forvar7653 + (1'h1)))
                begin
                  for (forvar7654 = (1'h0); (forvar7654 < (1'h0)); forvar7654 = (forvar7654 + (1'h1)))
                    begin
                      reg7655 <= forvar7654;
                      reg7656 <= reg7630;
                    end
                  if ($unsigned((~(|((8'h9c) ? reg7646 : forvar7632)))))
                    begin
                      reg7657 <= $signed(reg7635);
                      reg7658 <= (8'hb0);
                    end
                  else
                    begin
                      reg7657 <= (forvar7632 | (reg7631 || wire0[(3'h7):(2'h3)]));
                      reg7658 <= $signed((reg7658 + $unsigned(forvar7654[(3'h7):(1'h0)])));
                      reg7659 <= $unsigned($signed(wire618));
                      reg7660 <= (!$signed(((wire3 ^~ wire0) ?
                          $signed(reg7656) : (wire7625 | (8'had)))));
                    end
                end
            end
          else
            begin
              for (forvar7629 = (1'h0); (forvar7629 < (1'h1)); forvar7629 = (forvar7629 + (1'h1)))
                begin
                  for (forvar7630 = (1'h0); (forvar7630 < (1'h0)); forvar7630 = (forvar7630 + (1'h1)))
                    begin
                      reg7631 <= $unsigned((^(~(~|wire7625))));
                    end
                  reg7632 <= (^~forvar7653[(4'ha):(1'h1)]);
                  for (forvar7633 = (1'h0); (forvar7633 < (2'h2)); forvar7633 = (forvar7633 + (1'h1)))
                    begin
                      reg7634 <= reg7645[(3'h4):(1'h1)];
                      reg7635 <= ((-reg7659) ?
                          reg7639 : (($unsigned(reg7660) ?
                              (reg7637 ? forvar7633 : forvar7654) : (reg7659 ?
                                  reg7627 : (8'hac))) * reg7656[(3'h4):(2'h2)]));
                      reg7636 <= wire618[(1'h0):(1'h0)];
                    end
                  if (($unsigned(wire618) + $unsigned($signed(forvar7654[(3'h5):(3'h4)]))))
                    begin
                      reg7637 <= (((reg7638 ?
                              $unsigned(forvar7629) : (forvar7632 ?
                                  reg7638 : wire4)) ?
                          {forvar7654[(3'h5):(3'h5)]} : ((reg7642 + (8'ha4)) | $unsigned(reg7641))) <<< (({forvar7653} ?
                          reg7657[(2'h3):(1'h0)] : reg7656[(3'h6):(3'h4)]) - (reg7632[(4'hc):(4'ha)] >= (^~wire0))));
                      reg7638 <= $signed((-((reg7648 ? reg7660 : forvar7651) ?
                          (&(8'h9c)) : (wire2 < forvar7653))));
                      reg7639 <= forvar7640[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg7637 <= {{(&$unsigned(wire4))}};
                      reg7638 <= $signed((((reg7655 ?
                          reg7645 : reg7656) || (8'hac)) ^~ $unsigned(reg7647[(3'h5):(1'h1)])));
                    end
                end
              for (forvar7640 = (1'h0); (forvar7640 < (1'h0)); forvar7640 = (forvar7640 + (1'h1)))
                begin
                  reg7641 <= ($signed((reg7638[(1'h0):(1'h0)] ?
                      reg7639 : {reg7643})) >>> ({((8'hab) ? reg7644 : wire0)} ?
                      reg7649 : $signed($unsigned(reg7642))));
                end
            end
          if (({$signed((reg7646 ?
                  reg7641 : forvar7633))} < $signed($unsigned(reg7642[(4'ha):(2'h2)]))))
            begin
              for (forvar7661 = (1'h0); (forvar7661 < (1'h0)); forvar7661 = (forvar7661 + (1'h1)))
                begin
                  reg7662 <= ((8'hba) == reg7644);
                  if (({wire3[(4'hb):(3'h4)]} - reg7655[(4'hb):(3'h4)]))
                    begin
                      reg7663 <= $signed({$signed($signed(wire4))});
                    end
                  else
                    begin
                      reg7663 <= forvar7629;
                      reg7664 <= (8'ha8);
                      reg7665 <= {$signed(reg7641[(1'h1):(1'h0)])};
                    end
                  reg7666 <= forvar7630;
                end
              for (forvar7667 = (1'h0); (forvar7667 < (2'h2)); forvar7667 = (forvar7667 + (1'h1)))
                begin
                  for (forvar7668 = (1'h0); (forvar7668 < (2'h2)); forvar7668 = (forvar7668 + (1'h1)))
                    begin
                      reg7669 <= (-reg7652);
                      reg7670 <= forvar7667;
                      reg7671 <= reg7670[(2'h2):(2'h2)];
                    end
                  for (forvar7672 = (1'h0); (forvar7672 < (1'h1)); forvar7672 = (forvar7672 + (1'h1)))
                    begin
                      reg7673 <= $signed(({$unsigned(reg7634)} ?
                          reg7657[(2'h2):(1'h1)] : (reg7630 ?
                              $signed(reg7660) : $signed(wire5))));
                      reg7674 <= {(~^reg7647)};
                    end
                  if ((($signed((^~reg7630)) <<< (^{reg7655})) != reg7658[(1'h0):(1'h0)]))
                    begin
                      reg7675 <= {$signed($signed((forvar7668 ?
                              reg7635 : reg7650)))};
                    end
                  else
                    begin
                      reg7675 <= (-$signed(forvar7632[(2'h2):(1'h0)]));
                      reg7676 <= {((~^reg7673) ?
                              $signed(((8'ha5) ?
                                  (8'h9c) : wire1)) : ($signed(reg7647) ?
                                  (~|forvar7661) : $unsigned(reg7640)))};
                    end
                end
              reg7677 <= ($unsigned(reg7674) ~^ (~reg7632[(4'hf):(1'h0)]));
            end
          else
            begin
              if ({($unsigned($unsigned(reg7665)) ^ (reg7647 && ((8'hba) >>> reg7656)))})
                begin
                  for (forvar7661 = (1'h0); (forvar7661 < (1'h1)); forvar7661 = (forvar7661 + (1'h1)))
                    begin
                      reg7662 <= reg7643;
                      reg7663 <= ((+((forvar7667 ? reg7675 : wire5) ?
                          reg7670 : reg7666[(1'h1):(1'h0)])) ^ reg7655[(3'h5):(2'h2)]);
                      reg7664 <= (wire7628 ?
                          (~^forvar7654) : (+($unsigned(wire1) ?
                              $unsigned(wire4) : (8'haf))));
                    end
                  for (forvar7665 = (1'h0); (forvar7665 < (1'h0)); forvar7665 = (forvar7665 + (1'h1)))
                    begin
                      reg7666 <= reg7648[(4'hd):(4'hb)];
                      reg7667 <= $unsigned(forvar7651);
                      reg7668 <= (^~{$signed(forvar7668)});
                      reg7669 <= forvar7672[(2'h2):(2'h2)];
                    end
                  for (forvar7670 = (1'h0); (forvar7670 < (1'h0)); forvar7670 = (forvar7670 + (1'h1)))
                    begin
                      reg7671 <= $unsigned({($unsigned(reg7673) << (8'ha9))});
                      reg7672 <= $unsigned(forvar7653);
                      reg7673 <= ($signed(((reg7676 ? forvar7672 : reg7677) ?
                          (reg7656 << reg7663) : forvar7670[(1'h1):(1'h0)])) != $signed((~^(~^forvar7640))));
                    end
                end
              else
                begin
                  for (forvar7661 = (1'h0); (forvar7661 < (2'h2)); forvar7661 = (forvar7661 + (1'h1)))
                    begin
                      reg7662 <= ({(reg7670[(1'h1):(1'h1)] & reg7655[(3'h6):(2'h3)])} ?
                          $unsigned($unsigned($unsigned((8'hb3)))) : {({forvar7665} ?
                                  wire7625[(2'h3):(2'h2)] : (forvar7643 - reg7656))});
                    end
                end
              for (forvar7674 = (1'h0); (forvar7674 < (1'h0)); forvar7674 = (forvar7674 + (1'h1)))
                begin
                  if ($unsigned((({reg7658} ?
                      (reg7666 ? (8'ha9) : wire5) : (reg7636 ?
                          reg7666 : reg7630)) <= $signed({reg7647}))))
                    begin
                      reg7675 <= forvar7632[(1'h0):(1'h0)];
                      reg7676 <= $signed(reg7650[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg7675 <= reg7667;
                      reg7676 <= forvar7640;
                    end
                end
              if (reg7662)
                begin
                  for (forvar7677 = (1'h0); (forvar7677 < (1'h0)); forvar7677 = (forvar7677 + (1'h1)))
                    begin
                      reg7678 <= $signed(reg7631);
                      reg7679 <= ($signed(((+reg7669) ?
                              (8'hac) : forvar7668[(3'h7):(3'h6)])) ?
                          ((+forvar7667[(4'h9):(1'h0)]) != (-reg7633)) : forvar7630[(1'h0):(1'h0)]);
                      reg7680 <= ((forvar7674[(2'h3):(1'h0)] || reg7643) || $unsigned((reg7669 >>> (reg7668 * reg7633))));
                      reg7681 <= (-$unsigned({(reg7639 ^ reg7678)}));
                    end
                  for (forvar7682 = (1'h0); (forvar7682 < (2'h3)); forvar7682 = (forvar7682 + (1'h1)))
                    begin
                      reg7683 <= (~|{reg7662});
                      reg7684 <= $unsigned($signed(reg7663));
                      reg7685 <= reg7667[(1'h0):(1'h0)];
                    end
                  for (forvar7686 = (1'h0); (forvar7686 < (2'h3)); forvar7686 = (forvar7686 + (1'h1)))
                    begin
                      reg7687 <= (reg7671 * (($signed(reg7655) | $unsigned(reg7643)) ~^ reg7666[(1'h1):(1'h1)]));
                      reg7688 <= (forvar7643 ?
                          (-((reg7646 <= reg7680) * (wire5 ?
                              reg7641 : reg7652))) : reg7638[(3'h6):(2'h2)]);
                      reg7689 <= (8'ha0);
                      reg7690 <= (wire4 ? (~reg7649) : {$unsigned(forvar7654)});
                    end
                  if ($unsigned(({(-forvar7651)} >> {(|reg7645)})))
                    begin
                      reg7691 <= reg7673;
                      reg7692 <= forvar7670[(1'h1):(1'h1)];
                      reg7693 <= forvar7653[(4'hc):(2'h3)];
                      reg7694 <= {$unsigned(({(8'hb7)} ?
                              (!forvar7670) : $signed(reg7688)))};
                    end
                  else
                    begin
                      reg7691 <= (({$unsigned(reg7627)} ~^ $unsigned($unsigned(wire7628))) >>> (8'haa));
                      reg7692 <= $signed(reg7655[(1'h1):(1'h1)]);
                      reg7693 <= ((~^reg7663) ?
                          (8'h9c) : ((~$signed(wire618)) ?
                              reg7681[(3'h7):(1'h0)] : {reg7684[(3'h5):(2'h3)]}));
                      reg7694 <= (8'ha7);
                    end
                end
              else
                begin
                  for (forvar7677 = (1'h0); (forvar7677 < (1'h1)); forvar7677 = (forvar7677 + (1'h1)))
                    begin
                      reg7678 <= $unsigned(($signed($signed(reg7672)) ?
                          (8'hb4) : ((reg7639 ? reg7670 : forvar7643) ?
                              $signed(wire1) : $unsigned(reg7671))));
                      reg7679 <= reg7648;
                      reg7680 <= reg7633;
                    end
                  if ($unsigned($signed($unsigned($unsigned(reg7694)))))
                    begin
                      reg7681 <= $unsigned(forvar7661);
                      reg7682 <= (8'hb8);
                    end
                  else
                    begin
                      reg7681 <= forvar7667;
                      reg7682 <= (($unsigned(reg7669[(3'h4):(3'h4)]) ?
                          $signed($signed(forvar7670)) : (reg7630[(1'h0):(1'h0)] || $unsigned(reg7687))) != (reg7633 < reg7656[(3'h4):(1'h1)]));
                    end
                  for (forvar7683 = (1'h0); (forvar7683 < (1'h1)); forvar7683 = (forvar7683 + (1'h1)))
                    begin
                      reg7684 <= $signed((^({reg7656} | (wire4 ?
                          reg7647 : reg7638))));
                    end
                  if ($unsigned((reg7650[(3'h4):(2'h3)] >= $signed((~|reg7637)))))
                    begin
                      reg7685 <= (~|{$signed((reg7690 * reg7631))});
                      reg7686 <= (8'hb2);
                      reg7687 <= reg7638;
                    end
                  else
                    begin
                      reg7685 <= (reg7650[(3'h6):(2'h3)] ?
                          $signed($unsigned((8'ha3))) : ((~&$signed(forvar7670)) ?
                              {(8'hb0)} : $unsigned((reg7641 ?
                                  reg7677 : reg7676))));
                      reg7686 <= reg7637;
                      reg7687 <= reg7633;
                      reg7688 <= $signed($unsigned(reg7669[(4'h8):(3'h7)]));
                    end
                end
              for (forvar7695 = (1'h0); (forvar7695 < (1'h1)); forvar7695 = (forvar7695 + (1'h1)))
                begin
                  reg7696 <= $unsigned(reg7694);
                  reg7697 <= $unsigned($signed((!(reg7687 ?
                      reg7676 : (8'hab)))));
                end
            end
          for (forvar7698 = (1'h0); (forvar7698 < (2'h2)); forvar7698 = (forvar7698 + (1'h1)))
            begin
              for (forvar7699 = (1'h0); (forvar7699 < (1'h1)); forvar7699 = (forvar7699 + (1'h1)))
                begin
                  if ($signed(($unsigned((~^wire4)) ?
                      (~^(~forvar7683)) : ($signed(forvar7667) * $unsigned(reg7631)))))
                    begin
                      reg7700 <= $unsigned(wire5);
                      reg7701 <= ($signed(reg7650) < reg7667[(4'hf):(4'hb)]);
                      reg7702 <= (((-(forvar7629 ?
                              reg7671 : wire618)) ^ forvar7661[(1'h0):(1'h0)]) ?
                          ((wire618[(1'h0):(1'h0)] << $unsigned(reg7669)) ?
                              $signed((~&forvar7677)) : ((reg7674 + wire7625) >> {reg7627})) : (~&({reg7660} < (-forvar7686))));
                      reg7703 <= ($unsigned(($signed(reg7631) ?
                              (|reg7679) : reg7632)) ?
                          $unsigned(((8'hb2) ?
                              (8'ha6) : forvar7683)) : forvar7640[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg7700 <= (8'ha0);
                      reg7701 <= {(($unsigned(reg7679) ?
                              (-(8'h9f)) : (reg7702 ?
                                  reg7648 : wire3)) || ((^~reg7700) ?
                              (forvar7677 ?
                                  (8'had) : forvar7672) : (reg7678 > reg7645)))};
                    end
                  for (forvar7704 = (1'h0); (forvar7704 < (2'h3)); forvar7704 = (forvar7704 + (1'h1)))
                    begin
                      reg7705 <= (~(reg7650 & ($signed(reg7637) >= ((8'hb6) ?
                          reg7650 : forvar7653))));
                      reg7706 <= ($unsigned($signed(((8'hb2) || forvar7632))) | ((reg7664 ?
                              reg7627 : reg7646[(1'h1):(1'h1)]) ?
                          (~|$signed((8'hb7))) : {$signed(reg7627)}));
                    end
                  for (forvar7707 = (1'h0); (forvar7707 < (1'h0)); forvar7707 = (forvar7707 + (1'h1)))
                    begin
                      reg7708 <= (forvar7704 - forvar7683);
                      reg7709 <= reg7676;
                    end
                end
              for (forvar7710 = (1'h0); (forvar7710 < (1'h0)); forvar7710 = (forvar7710 + (1'h1)))
                begin
                  for (forvar7711 = (1'h0); (forvar7711 < (2'h3)); forvar7711 = (forvar7711 + (1'h1)))
                    begin
                      reg7712 <= $unsigned((forvar7710[(2'h2):(1'h0)] ?
                          $unsigned(reg7659) : ((-forvar7695) & (reg7667 == reg7632))));
                    end
                  for (forvar7713 = (1'h0); (forvar7713 < (1'h0)); forvar7713 = (forvar7713 + (1'h1)))
                    begin
                      reg7714 <= $unsigned(((~(reg7657 ?
                          forvar7668 : reg7636)) * forvar7632));
                      reg7715 <= (8'haa);
                      reg7716 <= wire2;
                    end
                  if (((^~((forvar7668 ?
                          forvar7704 : reg7697) - $unsigned(wire7628))) ?
                      forvar7672 : wire2[(1'h0):(1'h0)]))
                    begin
                      reg7717 <= $signed(reg7639[(3'h5):(2'h3)]);
                      reg7718 <= ($signed((-$signed(reg7659))) & reg7641);
                    end
                  else
                    begin
                      reg7717 <= (8'ha4);
                      reg7718 <= forvar7713;
                      reg7719 <= {{(forvar7661 ?
                                  forvar7668[(3'h6):(3'h5)] : ((8'hac) ?
                                      reg7639 : reg7635))}};
                      reg7720 <= (^(reg7655 & $signed((reg7712 != reg7627))));
                    end
                  if (($unsigned(reg7691) >>> reg7678))
                    begin
                      reg7721 <= reg7666;
                    end
                  else
                    begin
                      reg7721 <= ($signed(reg7697) <<< ($signed({reg7676}) >= $unsigned($unsigned((8'haa)))));
                      reg7722 <= $signed({$unsigned({reg7685})});
                    end
                end
              reg7723 <= reg7670;
              for (forvar7724 = (1'h0); (forvar7724 < (1'h1)); forvar7724 = (forvar7724 + (1'h1)))
                begin
                  if (reg7632)
                    begin
                      reg7725 <= {($unsigned($unsigned(reg7657)) ?
                              $signed((~^forvar7699)) : $unsigned($unsigned(reg7630)))};
                      reg7726 <= (reg7702[(4'hb):(1'h1)] >= ($unsigned((-reg7714)) == reg7646[(2'h2):(1'h1)]));
                      reg7727 <= $unsigned(((~&reg7701[(3'h6):(1'h1)]) ?
                          (reg7687[(2'h2):(2'h2)] | wire1[(4'hc):(4'ha)]) : ((|reg7663) ?
                              $unsigned((8'ha4)) : (forvar7686 ?
                                  (8'hb6) : reg7673))));
                    end
                  else
                    begin
                      reg7725 <= (~forvar7698);
                      reg7726 <= reg7664[(1'h0):(1'h0)];
                    end
                end
            end
          if (forvar7710)
            begin
              reg7728 <= $unsigned($unsigned(($unsigned(reg7656) ?
                  (reg7668 <<< reg7647) : ((8'h9d) + reg7655))));
              for (forvar7729 = (1'h0); (forvar7729 < (1'h1)); forvar7729 = (forvar7729 + (1'h1)))
                begin
                  reg7730 <= {{(8'hba)}};
                  if ((+{forvar7677[(4'hc):(3'h5)]}))
                    begin
                      reg7731 <= (reg7680[(3'h6):(2'h2)] ?
                          (!(&(!reg7697))) : (8'hae));
                      reg7732 <= ($unsigned(forvar7668[(3'h4):(2'h3)]) ~^ wire7625);
                      reg7733 <= reg7716;
                    end
                  else
                    begin
                      reg7731 <= {(forvar7640 ?
                              $signed($signed(forvar7665)) : reg7703)};
                      reg7732 <= ($unsigned({reg7720}) ^ $unsigned({(forvar7711 >= reg7725)}));
                      reg7733 <= reg7637[(1'h1):(1'h0)];
                    end
                  for (forvar7734 = (1'h0); (forvar7734 < (2'h3)); forvar7734 = (forvar7734 + (1'h1)))
                    begin
                      reg7735 <= (+(reg7722[(3'h5):(3'h5)] ?
                          reg7631 : reg7730[(3'h4):(3'h4)]));
                    end
                end
              for (forvar7736 = (1'h0); (forvar7736 < (1'h1)); forvar7736 = (forvar7736 + (1'h1)))
                begin
                  if (reg7643)
                    begin
                      reg7737 <= ($unsigned($unsigned($signed(reg7672))) ?
                          ($signed((|reg7674)) ?
                              (forvar7654[(4'h8):(2'h3)] >> $unsigned(forvar7668)) : (reg7689[(3'h4):(1'h0)] ?
                                  forvar7698[(1'h0):(1'h0)] : reg7683[(1'h0):(1'h0)])) : $unsigned((~(&forvar7670))));
                    end
                  else
                    begin
                      reg7737 <= reg7648;
                      reg7738 <= $signed((&$unsigned(((8'hb2) | reg7687))));
                      reg7739 <= $signed((~|$signed($unsigned(reg7722))));
                    end
                  for (forvar7740 = (1'h0); (forvar7740 < (2'h3)); forvar7740 = (forvar7740 + (1'h1)))
                    begin
                      reg7741 <= {$signed(reg7730[(1'h0):(1'h0)])};
                      reg7742 <= {forvar7661};
                      reg7743 <= (wire0[(4'hb):(4'h8)] ?
                          (8'hb6) : reg7650[(2'h2):(1'h0)]);
                    end
                end
            end
          else
            begin
              reg7728 <= ((~^$unsigned($signed(reg7668))) ?
                  $unsigned((!(~|(8'hba)))) : $unsigned((^~(+(8'hba)))));
            end
        end
      else
        begin
          reg7629 <= reg7718[(3'h4):(3'h4)];
          for (forvar7630 = (1'h0); (forvar7630 < (1'h0)); forvar7630 = (forvar7630 + (1'h1)))
            begin
              reg7631 <= reg7685[(2'h2):(1'h0)];
            end
        end
      if (reg7677)
        begin
          reg7744 <= forvar7710[(2'h2):(1'h1)];
          for (forvar7745 = (1'h0); (forvar7745 < (2'h2)); forvar7745 = (forvar7745 + (1'h1)))
            begin
              if ((forvar7740 ? reg7721 : {$unsigned((^~wire0))}))
                begin
                  for (forvar7746 = (1'h0); (forvar7746 < (1'h0)); forvar7746 = (forvar7746 + (1'h1)))
                    begin
                      reg7747 <= $unsigned({forvar7632});
                      reg7748 <= (reg7685 <= reg7637[(2'h3):(1'h1)]);
                      reg7749 <= $signed(($signed(reg7723[(3'h5):(1'h1)]) * reg7679));
                      reg7750 <= (wire0[(4'h8):(1'h0)] >= $unsigned({((8'hab) <<< reg7714)}));
                    end
                  if ($unsigned($signed(((forvar7632 ?
                      (8'haf) : reg7658) ^ forvar7710))))
                    begin
                      reg7751 <= $signed((($unsigned((8'h9d)) >> reg7659[(4'h9):(3'h4)]) && {{forvar7670}}));
                      reg7752 <= forvar7667;
                    end
                  else
                    begin
                      reg7751 <= reg7693;
                      reg7752 <= $signed(reg7725);
                      reg7753 <= $signed($unsigned($unsigned((reg7631 ?
                          reg7639 : (8'hb3)))));
                    end
                  reg7754 <= {reg7633[(2'h3):(1'h0)]};
                end
              else
                begin
                  for (forvar7746 = (1'h0); (forvar7746 < (2'h3)); forvar7746 = (forvar7746 + (1'h1)))
                    begin
                      reg7747 <= $signed($signed(forvar7736[(4'h9):(3'h6)]));
                    end
                  for (forvar7748 = (1'h0); (forvar7748 < (1'h1)); forvar7748 = (forvar7748 + (1'h1)))
                    begin
                      reg7749 <= ($signed((-wire4[(2'h3):(1'h0)])) + $unsigned(($signed(reg7662) ?
                          $unsigned(reg7672) : reg7662[(2'h3):(2'h2)])));
                      reg7750 <= $signed(((^~reg7658) ?
                          $unsigned(forvar7653) : ($unsigned(forvar7686) - reg7679)));
                    end
                end
              reg7755 <= (forvar7674 < $signed(({forvar7713} ^~ reg7728[(3'h4):(2'h2)])));
              if ($unsigned($unsigned((|((8'ha2) == forvar7740)))))
                begin
                  for (forvar7756 = (1'h0); (forvar7756 < (1'h0)); forvar7756 = (forvar7756 + (1'h1)))
                    begin
                      reg7757 <= ((((reg7689 ? reg7631 : reg7631) ?
                              {reg7749} : (reg7700 <<< reg7655)) >>> $signed(reg7676[(2'h2):(2'h2)])) ?
                          (&$signed((~|forvar7668))) : reg7744[(2'h2):(2'h2)]);
                      reg7758 <= $unsigned(($unsigned((&reg7693)) ?
                          $unsigned($unsigned(reg7675)) : $signed(reg7712)));
                      reg7759 <= (({(reg7739 ?
                                  reg7681 : reg7749)} > $unsigned(reg7674)) ?
                          ((+forvar7698) & (reg7682[(3'h7):(2'h3)] >= wire2[(3'h4):(3'h4)])) : reg7633);
                    end
                  for (forvar7760 = (1'h0); (forvar7760 < (2'h3)); forvar7760 = (forvar7760 + (1'h1)))
                    begin
                      reg7761 <= $unsigned((!{forvar7643}));
                      reg7762 <= $unsigned(reg7723);
                    end
                end
              else
                begin
                  for (forvar7756 = (1'h0); (forvar7756 < (1'h1)); forvar7756 = (forvar7756 + (1'h1)))
                    begin
                      reg7757 <= {reg7685[(2'h3):(1'h0)]};
                      reg7758 <= ((forvar7734 < (&(~^reg7663))) ?
                          reg7739[(4'hb):(2'h2)] : $unsigned($signed((reg7741 | forvar7629))));
                    end
                  reg7759 <= (^~$unsigned((forvar7710[(1'h0):(1'h0)] ?
                      $signed(forvar7748) : {reg7754})));
                  for (forvar7760 = (1'h0); (forvar7760 < (2'h2)); forvar7760 = (forvar7760 + (1'h1)))
                    begin
                      reg7761 <= ($signed(((reg7725 > forvar7677) != (~&(8'hb5)))) >>> reg7751);
                      reg7762 <= forvar7724;
                      reg7763 <= {{{(reg7757 ? forvar7630 : reg7741)}}};
                      reg7764 <= $signed($signed((^(reg7709 ?
                          reg7640 : forvar7686))));
                    end
                end
              reg7765 <= ($signed((~|(~|reg7735))) ~^ reg7712);
            end
          for (forvar7766 = (1'h0); (forvar7766 < (1'h1)); forvar7766 = (forvar7766 + (1'h1)))
            begin
              if (reg7758[(1'h0):(1'h0)])
                begin
                  if ($signed((8'hb0)))
                    begin
                      reg7767 <= (reg7634[(2'h3):(1'h0)] ?
                          ((~&(8'hb7)) ?
                              wire0 : reg7754[(4'h9):(3'h6)]) : ($signed((-reg7670)) >>> $unsigned($signed(reg7721))));
                    end
                  else
                    begin
                      reg7767 <= $signed(({$unsigned(reg7644)} ?
                          ((reg7678 != reg7705) == forvar7711) : (+(reg7742 ?
                              wire3 : forvar7674))));
                    end
                  for (forvar7768 = (1'h0); (forvar7768 < (1'h0)); forvar7768 = (forvar7768 + (1'h1)))
                    begin
                      reg7769 <= (^~reg7636);
                      reg7770 <= (!$unsigned({{(8'hb6)}}));
                    end
                end
              else
                begin
                  reg7767 <= ((reg7694 ? reg7639 : (!$unsigned(forvar7653))) ?
                      reg7753[(2'h2):(1'h1)] : ($unsigned((forvar7683 >= reg7681)) ?
                          {(reg7770 >> forvar7668)} : reg7685[(1'h0):(1'h0)]));
                  for (forvar7768 = (1'h0); (forvar7768 < (2'h3)); forvar7768 = (forvar7768 + (1'h1)))
                    begin
                      reg7769 <= (+$unsigned(reg7757[(1'h1):(1'h0)]));
                    end
                  for (forvar7770 = (1'h0); (forvar7770 < (2'h2)); forvar7770 = (forvar7770 + (1'h1)))
                    begin
                      reg7771 <= $unsigned((reg7665 ?
                          wire3[(3'h7):(3'h7)] : $signed($unsigned((8'hb8)))));
                    end
                  for (forvar7772 = (1'h0); (forvar7772 < (2'h3)); forvar7772 = (forvar7772 + (1'h1)))
                    begin
                      reg7773 <= wire0;
                    end
                end
              if (reg7685[(1'h0):(1'h0)])
                begin
                  reg7774 <= $signed(reg7656);
                  if (reg7774[(2'h2):(2'h2)])
                    begin
                      reg7775 <= $signed((^~{$signed(reg7627)}));
                      reg7776 <= $signed((~|(-$unsigned(wire3))));
                      reg7777 <= (forvar7748[(3'h4):(1'h1)] ?
                          (8'ha7) : $signed(reg7750[(2'h3):(2'h2)]));
                      reg7778 <= ((~|reg7663) ?
                          forvar7695 : (reg7657 & ((|reg7753) - $signed(forvar7640))));
                    end
                  else
                    begin
                      reg7775 <= (({$signed(reg7747)} ?
                          $unsigned($unsigned(reg7752)) : $unsigned((reg7652 ?
                              reg7721 : reg7751))) * (^~(^~(^~reg7731))));
                      reg7776 <= ($signed($signed($unsigned(reg7662))) ?
                          (~(forvar7729 ? {reg7679} : reg7677)) : ((!(reg7700 ?
                              reg7749 : reg7763)) + reg7733));
                      reg7777 <= ($unsigned(forvar7686[(4'hc):(2'h3)]) ?
                          $signed((!(&reg7749))) : reg7726[(4'h8):(1'h0)]);
                      reg7778 <= reg7761;
                    end
                  reg7779 <= $unsigned(forvar7677);
                  for (forvar7780 = (1'h0); (forvar7780 < (2'h2)); forvar7780 = (forvar7780 + (1'h1)))
                    begin
                      reg7781 <= ((reg7655[(1'h0):(1'h0)] ?
                          (8'haf) : reg7629) + {{$unsigned(reg7648)}});
                    end
                end
              else
                begin
                  if (forvar7713)
                    begin
                      reg7774 <= $signed($signed(reg7667[(4'ha):(1'h0)]));
                      reg7775 <= forvar7710;
                      reg7776 <= (^(($unsigned(forvar7729) ?
                          $signed(reg7720) : (wire4 ?
                              reg7715 : forvar7661)) | $signed((8'haf))));
                    end
                  else
                    begin
                      reg7774 <= (8'h9c);
                      reg7775 <= reg7721[(4'h8):(4'h8)];
                    end
                  for (forvar7777 = (1'h0); (forvar7777 < (1'h1)); forvar7777 = (forvar7777 + (1'h1)))
                    begin
                      reg7778 <= (reg7774 ?
                          reg7672[(4'h9):(1'h0)] : $unsigned($signed((~(8'ha9)))));
                      reg7779 <= forvar7683[(3'h7):(3'h5)];
                      reg7780 <= (|(reg7678[(3'h7):(3'h7)] ?
                          $unsigned((reg7748 || reg7764)) : $signed(reg7776)));
                      reg7781 <= $unsigned((($unsigned((8'ha0)) ?
                          $signed(reg7735) : $signed(forvar7746)) <= (&(reg7672 ?
                          forvar7667 : reg7679))));
                    end
                end
            end
        end
      else
        begin
          for (forvar7744 = (1'h0); (forvar7744 < (1'h1)); forvar7744 = (forvar7744 + (1'h1)))
            begin
              for (forvar7745 = (1'h0); (forvar7745 < (2'h3)); forvar7745 = (forvar7745 + (1'h1)))
                begin
                  if (reg7629[(1'h0):(1'h0)])
                    begin
                      reg7746 <= reg7776[(2'h2):(2'h2)];
                      reg7747 <= ($signed($signed($signed(wire7628))) ?
                          $unsigned((8'haf)) : $signed(forvar7632[(1'h0):(1'h0)]));
                      reg7748 <= (~|(reg7688[(2'h2):(1'h1)] ?
                          $signed({forvar7768}) : ({reg7658} ?
                              (forvar7713 * reg7780) : reg7683)));
                    end
                  else
                    begin
                      reg7746 <= $unsigned(forvar7744[(1'h0):(1'h0)]);
                      reg7747 <= $signed(($unsigned(reg7769) ?
                          {(~|forvar7629)} : ($signed(reg7639) + (8'ha2))));
                      reg7748 <= (-(($signed(reg7644) ?
                              $signed(reg7631) : (~|reg7738)) ?
                          ((^~reg7629) ?
                              (reg7753 | wire618) : $signed(reg7683)) : $signed((|forvar7695))));
                    end
                  for (forvar7749 = (1'h0); (forvar7749 < (1'h1)); forvar7749 = (forvar7749 + (1'h1)))
                    begin
                      reg7750 <= $signed((forvar7654 >> $unsigned({forvar7770})));
                    end
                  if (reg7690[(2'h2):(2'h2)])
                    begin
                      reg7751 <= (((reg7721 - (8'hb8)) + (!(reg7731 ?
                              reg7680 : (8'h9f)))) ?
                          reg7754 : $unsigned($signed(((8'hac) << wire5))));
                      reg7752 <= forvar7736;
                      reg7753 <= (&$unsigned(($signed((8'h9f)) >= forvar7734)));
                    end
                  else
                    begin
                      reg7751 <= reg7636[(2'h2):(2'h2)];
                    end
                end
            end
          for (forvar7754 = (1'h0); (forvar7754 < (2'h2)); forvar7754 = (forvar7754 + (1'h1)))
            begin
              for (forvar7755 = (1'h0); (forvar7755 < (2'h3)); forvar7755 = (forvar7755 + (1'h1)))
                begin
                  if ($signed((((~&reg7629) ?
                          (reg7686 ?
                              (8'ha8) : forvar7746) : reg7649[(4'h9):(3'h6)]) ?
                      reg7696[(1'h1):(1'h1)] : $unsigned($signed(reg7738)))))
                    begin
                      reg7756 <= $unsigned((($signed((8'hb7)) ?
                              $signed((8'ha4)) : (forvar7748 ~^ (8'had))) ?
                          ({reg7776} ?
                              (reg7680 > reg7753) : $unsigned((8'hab))) : $unsigned((reg7763 != (8'hb0)))));
                    end
                  else
                    begin
                      reg7756 <= (&$unsigned($unsigned((8'h9f))));
                      reg7757 <= (~({reg7747} ?
                          forvar7686 : (~|((8'h9f) ? forvar7665 : reg7738))));
                    end
                  reg7758 <= (($signed(reg7657) ?
                          {reg7638[(1'h1):(1'h1)]} : $unsigned($unsigned(reg7756))) ?
                      ($signed((&forvar7749)) <<< reg7678) : {$signed($signed(reg7677))});
                  if ($signed({reg7780[(2'h2):(2'h2)]}))
                    begin
                      reg7759 <= (reg7687 ?
                          $signed({$signed(reg7716)}) : $unsigned({(|(8'ha7))}));
                    end
                  else
                    begin
                      reg7759 <= reg7731;
                      reg7760 <= reg7636;
                    end
                end
              if ((({$unsigned((8'hb3))} | reg7696[(2'h2):(1'h1)]) ?
                  (^($signed(reg7663) * $signed(forvar7754))) : forvar7756))
                begin
                  reg7761 <= wire3[(3'h4):(2'h3)];
                  for (forvar7762 = (1'h0); (forvar7762 < (2'h2)); forvar7762 = (forvar7762 + (1'h1)))
                    begin
                      reg7763 <= $signed({((-reg7683) ?
                              forvar7661[(1'h1):(1'h1)] : $signed(reg7777))});
                      reg7764 <= (((forvar7632[(1'h1):(1'h1)] ?
                              forvar7736 : $signed((8'h9c))) || $signed(forvar7643)) ?
                          ((reg7759 ?
                              {reg7627} : reg7781[(1'h0):(1'h0)]) <= reg7686) : $signed($unsigned((reg7744 - reg7662))));
                    end
                  for (forvar7765 = (1'h0); (forvar7765 < (1'h0)); forvar7765 = (forvar7765 + (1'h1)))
                    begin
                      reg7766 <= $signed($signed($unsigned((8'hb7))));
                    end
                  reg7767 <= reg7747;
                end
              else
                begin
                  for (forvar7761 = (1'h0); (forvar7761 < (2'h3)); forvar7761 = (forvar7761 + (1'h1)))
                    begin
                      reg7762 <= reg7779[(2'h3):(2'h2)];
                      reg7763 <= $unsigned(($unsigned($unsigned(reg7737)) + $unsigned(reg7752)));
                    end
                  for (forvar7764 = (1'h0); (forvar7764 < (2'h2)); forvar7764 = (forvar7764 + (1'h1)))
                    begin
                      reg7765 <= reg7780[(1'h0):(1'h0)];
                      reg7766 <= reg7669[(3'h7):(1'h0)];
                      reg7767 <= (8'hb9);
                      reg7768 <= reg7722[(3'h6):(3'h6)];
                    end
                end
              for (forvar7769 = (1'h0); (forvar7769 < (1'h1)); forvar7769 = (forvar7769 + (1'h1)))
                begin
                  for (forvar7770 = (1'h0); (forvar7770 < (2'h3)); forvar7770 = (forvar7770 + (1'h1)))
                    begin
                      reg7771 <= reg7731;
                    end
                  for (forvar7772 = (1'h0); (forvar7772 < (2'h2)); forvar7772 = (forvar7772 + (1'h1)))
                    begin
                      reg7773 <= $signed((reg7684[(3'h5):(3'h5)] * ($unsigned(forvar7670) >= $unsigned(reg7635))));
                      reg7774 <= forvar7654[(2'h2):(2'h2)];
                      reg7775 <= reg7667;
                    end
                end
            end
        end
    end
  assign wire7782 = (forvar7672 || $signed((^~(reg7647 ? reg7759 : (8'ha3)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module620  (y, clk, wire624, wire623, wire622, wire621);
  output wire [(32'ha47):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire624;
  input wire [(4'hc):(1'h0)] wire623;
  input wire signed [(2'h3):(1'h0)] wire622;
  input wire [(3'h5):(1'h0)] wire621;
  wire [(4'h8):(1'h0)] wire7624;
  reg signed [(3'h6):(1'h0)] reg7623 = (1'h0);
  reg [(3'h7):(1'h0)] reg7619 = (1'h0);
  reg [(2'h3):(1'h0)] reg7622 = (1'h0);
  reg [(4'h8):(1'h0)] reg7621 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7620 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar7619 = (1'h0);
  reg [(5'h10):(1'h0)] reg7618 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7617 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7616 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7615 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7614 = (1'h0);
  reg [(3'h4):(1'h0)] reg7613 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7612 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7611 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7610 = (1'h0);
  reg [(3'h6):(1'h0)] forvar7609 = (1'h0);
  reg [(3'h4):(1'h0)] reg7608 = (1'h0);
  reg [(4'hd):(1'h0)] reg7607 = (1'h0);
  reg [(2'h2):(1'h0)] reg7606 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7605 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7604 = (1'h0);
  reg [(2'h3):(1'h0)] reg7603 = (1'h0);
  reg [(4'h9):(1'h0)] reg7602 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar7601 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7600 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7599 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7598 = (1'h0);
  reg [(4'ha):(1'h0)] reg7597 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7596 = (1'h0);
  reg [(4'hd):(1'h0)] reg7595 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7594 = (1'h0);
  reg [(5'h10):(1'h0)] reg7593 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7592 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7591 = (1'h0);
  reg [(3'h6):(1'h0)] reg7590 = (1'h0);
  reg [(4'ha):(1'h0)] reg7589 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7587 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7582 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7577 = (1'h0);
  reg [(3'h5):(1'h0)] reg7576 = (1'h0);
  reg [(3'h6):(1'h0)] reg7585 = (1'h0);
  reg [(4'hd):(1'h0)] reg7588 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7587 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7586 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7585 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7584 = (1'h0);
  reg [(4'hd):(1'h0)] reg7583 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7582 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7581 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7580 = (1'h0);
  reg [(4'hb):(1'h0)] reg7579 = (1'h0);
  reg [(4'h8):(1'h0)] reg7578 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7577 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar7576 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7575 = (1'h0);
  reg [(5'h10):(1'h0)] forvar7574 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7573 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7572 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7571 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar7570 = (1'h0);
  reg [(4'hd):(1'h0)] reg7569 = (1'h0);
  reg [(5'h10):(1'h0)] reg7568 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7567 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7566 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7565 = (1'h0);
  reg [(4'hf):(1'h0)] reg7564 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7563 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7562 = (1'h0);
  reg [(3'h4):(1'h0)] reg7561 = (1'h0);
  reg [(3'h7):(1'h0)] reg7560 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7559 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7558 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7557 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7556 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7555 = (1'h0);
  reg [(4'hb):(1'h0)] reg7554 = (1'h0);
  reg [(2'h3):(1'h0)] reg7553 = (1'h0);
  reg [(3'h4):(1'h0)] reg7552 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7551 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7550 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7549 = (1'h0);
  reg [(4'hc):(1'h0)] reg7548 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7547 = (1'h0);
  reg [(3'h5):(1'h0)] forvar7546 = (1'h0);
  reg [(2'h2):(1'h0)] reg7546 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7545 = (1'h0);
  reg [(4'ha):(1'h0)] forvar7543 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7539 = (1'h0);
  reg [(3'h5):(1'h0)] reg7544 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7543 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7542 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7541 = (1'h0);
  reg [(4'h9):(1'h0)] reg7540 = (1'h0);
  reg [(3'h6):(1'h0)] reg7539 = (1'h0);
  reg [(4'hd):(1'h0)] reg7538 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7537 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7536 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7531 = (1'h0);
  reg [(3'h5):(1'h0)] reg7535 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7534 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7533 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7532 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7531 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7530 = (1'h0);
  reg [(4'hd):(1'h0)] reg7529 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7528 = (1'h0);
  reg [(4'ha):(1'h0)] reg7527 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7526 = (1'h0);
  reg [(4'hf):(1'h0)] reg7525 = (1'h0);
  reg [(4'ha):(1'h0)] reg7524 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7523 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7522 = (1'h0);
  reg [(4'hb):(1'h0)] reg7521 = (1'h0);
  reg [(4'hc):(1'h0)] reg7520 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7519 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7518 = (1'h0);
  reg [(4'h9):(1'h0)] reg7517 = (1'h0);
  reg [(4'ha):(1'h0)] reg7516 = (1'h0);
  reg [(4'hc):(1'h0)] reg7515 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7514 = (1'h0);
  reg [(4'he):(1'h0)] reg7513 = (1'h0);
  reg [(3'h5):(1'h0)] reg7512 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7511 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7510 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7509 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7508 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7507 = (1'h0);
  reg [(4'ha):(1'h0)] reg7506 = (1'h0);
  reg [(5'h10):(1'h0)] reg7505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7504 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7503 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7502 = (1'h0);
  reg [(4'h9):(1'h0)] reg7501 = (1'h0);
  reg [(3'h7):(1'h0)] reg7500 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7493 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7499 = (1'h0);
  reg [(4'hc):(1'h0)] reg7498 = (1'h0);
  reg [(4'hd):(1'h0)] reg7497 = (1'h0);
  reg [(4'hc):(1'h0)] reg7496 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7495 = (1'h0);
  reg [(4'he):(1'h0)] reg7494 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7493 = (1'h0);
  reg [(4'hb):(1'h0)] reg7492 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7491 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7490 = (1'h0);
  reg [(3'h5):(1'h0)] reg7489 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7488 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7487 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7486 = (1'h0);
  reg [(4'ha):(1'h0)] reg7485 = (1'h0);
  reg [(4'he):(1'h0)] reg7484 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7483 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7482 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7481 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7480 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar7479 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7478 = (1'h0);
  reg [(3'h5):(1'h0)] forvar7477 = (1'h0);
  reg [(4'he):(1'h0)] forvar7454 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7449 = (1'h0);
  reg [(3'h6):(1'h0)] forvar7446 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7443 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7442 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7440 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7441 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7438 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7437 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7436 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7476 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar7475 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7474 = (1'h0);
  reg [(5'h10):(1'h0)] reg7466 = (1'h0);
  reg [(4'hf):(1'h0)] reg7473 = (1'h0);
  reg [(4'hb):(1'h0)] reg7472 = (1'h0);
  reg [(3'h6):(1'h0)] reg7471 = (1'h0);
  reg [(5'h10):(1'h0)] forvar7470 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7469 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7468 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7467 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7466 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7465 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7464 = (1'h0);
  reg [(4'h9):(1'h0)] reg7462 = (1'h0);
  reg [(3'h4):(1'h0)] reg7461 = (1'h0);
  reg [(3'h6):(1'h0)] reg7456 = (1'h0);
  reg [(4'he):(1'h0)] reg7457 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7450 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7448 = (1'h0);
  reg [(3'h4):(1'h0)] reg7445 = (1'h0);
  reg [(3'h4):(1'h0)] reg7463 = (1'h0);
  reg [(4'ha):(1'h0)] forvar7462 = (1'h0);
  reg [(3'h7):(1'h0)] forvar7461 = (1'h0);
  reg [(4'hb):(1'h0)] reg7460 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7459 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7458 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar7457 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7456 = (1'h0);
  reg [(3'h7):(1'h0)] reg7455 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7454 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7453 = (1'h0);
  reg [(4'he):(1'h0)] reg7452 = (1'h0);
  reg [(4'ha):(1'h0)] reg7451 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7450 = (1'h0);
  reg [(4'hd):(1'h0)] reg7449 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7448 = (1'h0);
  reg [(3'h7):(1'h0)] reg7447 = (1'h0);
  reg [(5'h10):(1'h0)] reg7446 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7445 = (1'h0);
  reg [(2'h3):(1'h0)] reg7444 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7443 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7442 = (1'h0);
  reg [(4'hb):(1'h0)] reg7441 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7440 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7439 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7438 = (1'h0);
  reg [(3'h7):(1'h0)] forvar7437 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7436 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire7435;
  wire signed [(4'hf):(1'h0)] wire7433;
  wire signed [(4'he):(1'h0)] wire7432;
  wire signed [(3'h5):(1'h0)] wire7431;
  wire [(2'h2):(1'h0)] wire7430;
  wire signed [(4'hf):(1'h0)] wire7429;
  wire [(4'hb):(1'h0)] wire7427;
  reg signed [(4'h8):(1'h0)] forvar643 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg642 = (1'h0);
  reg [(3'h5):(1'h0)] forvar639 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg638 = (1'h0);
  reg [(4'he):(1'h0)] reg637 = (1'h0);
  reg [(4'he):(1'h0)] forvar636 = (1'h0);
  reg [(3'h5):(1'h0)] reg672 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar671 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg667 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg674 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg673 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar672 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg671 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg670 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg669 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg668 = (1'h0);
  reg [(4'hc):(1'h0)] forvar667 = (1'h0);
  reg [(3'h7):(1'h0)] reg666 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg665 = (1'h0);
  reg [(3'h4):(1'h0)] reg664 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg663 = (1'h0);
  reg [(4'hf):(1'h0)] forvar662 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg661 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg660 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar659 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg658 = (1'h0);
  reg [(3'h7):(1'h0)] reg651 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar648 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar644 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg657 = (1'h0);
  reg [(4'he):(1'h0)] reg656 = (1'h0);
  reg [(5'h10):(1'h0)] reg655 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar654 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg653 = (1'h0);
  reg signed [(4'he):(1'h0)] reg652 = (1'h0);
  reg [(4'h8):(1'h0)] forvar651 = (1'h0);
  reg [(4'hf):(1'h0)] reg650 = (1'h0);
  reg [(2'h2):(1'h0)] reg649 = (1'h0);
  reg [(5'h10):(1'h0)] reg648 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg647 = (1'h0);
  reg [(3'h7):(1'h0)] reg646 = (1'h0);
  reg [(3'h4):(1'h0)] reg645 = (1'h0);
  reg [(4'h9):(1'h0)] reg644 = (1'h0);
  reg [(4'hd):(1'h0)] reg643 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar642 = (1'h0);
  reg [(3'h4):(1'h0)] reg641 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg640 = (1'h0);
  reg [(4'hd):(1'h0)] reg639 = (1'h0);
  reg [(4'ha):(1'h0)] forvar638 = (1'h0);
  reg [(3'h6):(1'h0)] forvar637 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg635 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar632 = (1'h0);
  reg [(4'hd):(1'h0)] reg636 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar635 = (1'h0);
  reg [(4'hb):(1'h0)] reg634 = (1'h0);
  reg [(2'h3):(1'h0)] reg633 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg632 = (1'h0);
  reg [(3'h6):(1'h0)] forvar631 = (1'h0);
  wire [(4'hc):(1'h0)] wire630;
  wire [(3'h6):(1'h0)] wire629;
  wire signed [(3'h4):(1'h0)] wire628;
  wire signed [(4'ha):(1'h0)] wire627;
  wire [(4'ha):(1'h0)] wire626;
  wire [(4'hb):(1'h0)] wire625;
  assign y = {wire7624,
                 reg7623,
                 reg7619,
                 reg7622,
                 reg7621,
                 reg7620,
                 forvar7619,
                 reg7618,
                 forvar7617,
                 reg7616,
                 reg7615,
                 reg7614,
                 reg7613,
                 reg7612,
                 reg7611,
                 reg7610,
                 forvar7609,
                 reg7608,
                 reg7607,
                 reg7606,
                 forvar7605,
                 reg7604,
                 reg7603,
                 reg7602,
                 forvar7601,
                 forvar7600,
                 forvar7599,
                 forvar7598,
                 reg7597,
                 forvar7596,
                 reg7595,
                 reg7594,
                 reg7593,
                 reg7592,
                 reg7591,
                 reg7590,
                 reg7589,
                 forvar7587,
                 forvar7582,
                 reg7577,
                 reg7576,
                 reg7585,
                 reg7588,
                 reg7587,
                 reg7586,
                 forvar7585,
                 reg7584,
                 reg7583,
                 reg7582,
                 reg7581,
                 reg7580,
                 reg7579,
                 reg7578,
                 forvar7577,
                 forvar7576,
                 reg7575,
                 forvar7574,
                 reg7573,
                 reg7572,
                 reg7571,
                 forvar7570,
                 reg7569,
                 reg7568,
                 reg7567,
                 reg7566,
                 forvar7565,
                 reg7564,
                 reg7563,
                 reg7562,
                 reg7561,
                 reg7560,
                 reg7559,
                 forvar7558,
                 forvar7557,
                 reg7556,
                 forvar7555,
                 reg7554,
                 reg7553,
                 reg7552,
                 forvar7551,
                 reg7550,
                 reg7549,
                 reg7548,
                 reg7547,
                 forvar7546,
                 reg7546,
                 reg7545,
                 forvar7543,
                 forvar7539,
                 reg7544,
                 reg7543,
                 reg7542,
                 reg7541,
                 reg7540,
                 reg7539,
                 reg7538,
                 reg7537,
                 reg7536,
                 reg7531,
                 reg7535,
                 reg7534,
                 reg7533,
                 reg7532,
                 forvar7531,
                 forvar7530,
                 reg7529,
                 forvar7528,
                 reg7527,
                 reg7526,
                 reg7525,
                 reg7524,
                 forvar7523,
                 forvar7522,
                 reg7521,
                 reg7520,
                 forvar7519,
                 reg7518,
                 reg7517,
                 reg7516,
                 reg7515,
                 forvar7514,
                 reg7513,
                 reg7512,
                 reg7511,
                 reg7510,
                 reg7509,
                 forvar7508,
                 forvar7507,
                 reg7506,
                 reg7505,
                 reg7504,
                 reg7503,
                 reg7502,
                 reg7501,
                 reg7500,
                 reg7493,
                 reg7499,
                 reg7498,
                 reg7497,
                 reg7496,
                 reg7495,
                 reg7494,
                 forvar7493,
                 reg7492,
                 reg7491,
                 forvar7490,
                 reg7489,
                 forvar7488,
                 forvar7487,
                 reg7486,
                 reg7485,
                 reg7484,
                 reg7483,
                 forvar7482,
                 reg7481,
                 reg7480,
                 forvar7479,
                 forvar7478,
                 forvar7477,
                 forvar7454,
                 forvar7449,
                 forvar7446,
                 reg7443,
                 forvar7442,
                 forvar7440,
                 forvar7441,
                 forvar7438,
                 reg7437,
                 reg7436,
                 reg7476,
                 forvar7475,
                 reg7474,
                 reg7466,
                 reg7473,
                 reg7472,
                 reg7471,
                 forvar7470,
                 reg7469,
                 reg7468,
                 reg7467,
                 forvar7466,
                 reg7465,
                 reg7464,
                 reg7462,
                 reg7461,
                 reg7456,
                 reg7457,
                 reg7450,
                 forvar7448,
                 reg7445,
                 reg7463,
                 forvar7462,
                 forvar7461,
                 reg7460,
                 reg7459,
                 reg7458,
                 forvar7457,
                 forvar7456,
                 reg7455,
                 reg7454,
                 reg7453,
                 reg7452,
                 reg7451,
                 forvar7450,
                 reg7449,
                 reg7448,
                 reg7447,
                 reg7446,
                 forvar7445,
                 reg7444,
                 forvar7443,
                 reg7442,
                 reg7441,
                 reg7440,
                 reg7439,
                 reg7438,
                 forvar7437,
                 forvar7436,
                 wire7435,
                 wire7433,
                 wire7432,
                 wire7431,
                 wire7430,
                 wire7429,
                 wire7427,
                 forvar643,
                 reg642,
                 forvar639,
                 reg638,
                 reg637,
                 forvar636,
                 reg672,
                 forvar671,
                 reg667,
                 reg674,
                 reg673,
                 forvar672,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 forvar667,
                 reg666,
                 reg665,
                 reg664,
                 reg663,
                 forvar662,
                 reg661,
                 reg660,
                 forvar659,
                 reg658,
                 reg651,
                 forvar648,
                 forvar644,
                 reg657,
                 reg656,
                 reg655,
                 forvar654,
                 reg653,
                 reg652,
                 forvar651,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 forvar642,
                 reg641,
                 reg640,
                 reg639,
                 forvar638,
                 forvar637,
                 reg635,
                 forvar632,
                 reg636,
                 forvar635,
                 reg634,
                 reg633,
                 reg632,
                 forvar631,
                 wire630,
                 wire629,
                 wire628,
                 wire627,
                 wire626,
                 wire625,
                 (1'h0)};
  assign wire625 = {wire622};
  assign wire626 = (^~wire625);
  assign wire627 = wire622;
  assign wire628 = ({wire625[(4'hb):(1'h1)]} ?
                       (($signed(wire625) ? (|wire627) : wire623) ?
                           $unsigned(wire622[(1'h0):(1'h0)]) : (wire626 ?
                               $signed(wire622) : (^wire625))) : wire624[(1'h0):(1'h0)]);
  assign wire629 = $signed(($signed($unsigned(wire621)) ?
                       (wire623[(3'h7):(3'h6)] ?
                           {wire626} : wire622) : (&((8'hb2) ?
                           wire625 : wire621))));
  assign wire630 = wire621;
  always
    @(posedge clk) begin
      if ($signed(wire623[(4'hb):(2'h3)]))
        begin
          for (forvar631 = (1'h0); (forvar631 < (2'h3)); forvar631 = (forvar631 + (1'h1)))
            begin
              if ((|{$signed((wire629 ? wire622 : wire623))}))
                begin
                  if ((+((wire621[(1'h0):(1'h0)] ?
                      wire625 : wire623[(4'h9):(4'h8)]) ^ (((8'hb8) + wire629) ?
                      ((8'haa) > forvar631) : forvar631[(2'h3):(1'h0)]))))
                    begin
                      reg632 <= $signed($signed($signed(wire629)));
                      reg633 <= (8'ha6);
                    end
                  else
                    begin
                      reg632 <= (!$signed((!$signed(wire621))));
                      reg633 <= $signed(wire627[(4'h8):(3'h6)]);
                      reg634 <= $signed((+wire626));
                    end
                  for (forvar635 = (1'h0); (forvar635 < (1'h0)); forvar635 = (forvar635 + (1'h1)))
                    begin
                      reg636 <= ({$unsigned($signed(wire629))} | $unsigned($signed((wire623 ?
                          wire626 : wire629))));
                    end
                end
              else
                begin
                  for (forvar632 = (1'h0); (forvar632 < (1'h1)); forvar632 = (forvar632 + (1'h1)))
                    begin
                      reg633 <= $signed($unsigned($unsigned(wire623)));
                      reg634 <= forvar632[(2'h3):(2'h2)];
                      reg635 <= $unsigned(forvar635);
                    end
                end
              for (forvar637 = (1'h0); (forvar637 < (1'h1)); forvar637 = (forvar637 + (1'h1)))
                begin
                  for (forvar638 = (1'h0); (forvar638 < (1'h1)); forvar638 = (forvar638 + (1'h1)))
                    begin
                      reg639 <= (!$signed($unsigned(((8'ha5) ^~ reg634))));
                      reg640 <= (wire622[(1'h1):(1'h1)] ? wire624 : wire622);
                      reg641 <= reg639;
                    end
                  for (forvar642 = (1'h0); (forvar642 < (2'h3)); forvar642 = (forvar642 + (1'h1)))
                    begin
                      reg643 <= reg634[(3'h7):(1'h1)];
                    end
                end
              if ($unsigned($unsigned(wire621[(1'h1):(1'h1)])))
                begin
                  if ($signed(wire625[(3'h7):(2'h3)]))
                    begin
                      reg644 <= $signed($signed($signed(((8'ha8) & forvar638))));
                      reg645 <= (8'hb8);
                    end
                  else
                    begin
                      reg644 <= ($unsigned((|(reg632 ? reg633 : wire623))) ?
                          reg634[(1'h1):(1'h1)] : {(^$unsigned(forvar635))});
                      reg645 <= forvar637;
                      reg646 <= ($unsigned(forvar631) >= reg645);
                      reg647 <= $unsigned(reg635[(2'h2):(1'h1)]);
                    end
                  if ({forvar638[(4'h9):(2'h2)]})
                    begin
                      reg648 <= (~&wire627[(3'h5):(2'h3)]);
                      reg649 <= wire625;
                      reg650 <= $unsigned(((wire628[(1'h1):(1'h1)] <= $unsigned(reg639)) ?
                          $signed($signed(forvar642)) : forvar637[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg648 <= reg639[(3'h7):(3'h5)];
                    end
                  for (forvar651 = (1'h0); (forvar651 < (1'h0)); forvar651 = (forvar651 + (1'h1)))
                    begin
                      reg652 <= reg643;
                      reg653 <= $signed(reg641);
                    end
                  for (forvar654 = (1'h0); (forvar654 < (2'h2)); forvar654 = (forvar654 + (1'h1)))
                    begin
                      reg655 <= forvar635[(3'h6):(1'h0)];
                      reg656 <= (~|reg640[(3'h4):(1'h0)]);
                      reg657 <= reg633[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar644 = (1'h0); (forvar644 < (2'h3)); forvar644 = (forvar644 + (1'h1)))
                    begin
                      reg645 <= reg657[(3'h6):(3'h4)];
                      reg646 <= wire626;
                      reg647 <= reg646[(2'h3):(1'h1)];
                    end
                  for (forvar648 = (1'h0); (forvar648 < (2'h3)); forvar648 = (forvar648 + (1'h1)))
                    begin
                      reg649 <= $signed(forvar651);
                      reg650 <= (|(+reg635[(1'h1):(1'h1)]));
                    end
                  reg651 <= reg655[(4'h8):(1'h1)];
                end
              reg658 <= reg634;
            end
          for (forvar659 = (1'h0); (forvar659 < (2'h3)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 <= forvar637;
              reg661 <= (-$unsigned(($unsigned(forvar642) != wire630[(4'hb):(4'ha)])));
              if ($signed((^wire629)))
                begin
                  for (forvar662 = (1'h0); (forvar662 < (1'h0)); forvar662 = (forvar662 + (1'h1)))
                    begin
                      reg663 <= $signed(reg639[(3'h6):(2'h3)]);
                      reg664 <= $signed($unsigned((forvar659[(3'h6):(2'h3)] ?
                          reg653[(2'h3):(1'h1)] : (wire623 ?
                              reg646 : (8'ha6)))));
                      reg665 <= ($unsigned({(^forvar659)}) ?
                          $signed(((^(8'had)) ?
                              $unsigned(wire627) : ((8'hab) ?
                                  (8'hb9) : forvar642))) : reg633[(2'h3):(2'h2)]);
                      reg666 <= reg634;
                    end
                  for (forvar667 = (1'h0); (forvar667 < (1'h0)); forvar667 = (forvar667 + (1'h1)))
                    begin
                      reg668 <= $signed({$unsigned($signed(forvar638))});
                      reg669 <= $signed($unsigned((~&{wire626})));
                    end
                  if (reg658[(4'ha):(4'ha)])
                    begin
                      reg670 <= $unsigned((~^{(+forvar662)}));
                      reg671 <= (!($signed(reg664[(1'h1):(1'h0)]) >>> reg635[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg670 <= $unsigned(reg668);
                    end
                  for (forvar672 = (1'h0); (forvar672 < (1'h1)); forvar672 = (forvar672 + (1'h1)))
                    begin
                      reg673 <= ($unsigned(reg643) ?
                          reg643[(4'hd):(3'h7)] : $unsigned((reg660 ?
                              reg641 : (reg636 << (8'hba)))));
                      reg674 <= (+$signed(reg640[(2'h2):(1'h1)]));
                    end
                end
              else
                begin
                  for (forvar662 = (1'h0); (forvar662 < (2'h3)); forvar662 = (forvar662 + (1'h1)))
                    begin
                      reg663 <= ((8'ha4) ~^ ($signed((reg634 && reg635)) | reg652[(4'h8):(3'h7)]));
                      reg664 <= (($signed(reg644[(3'h4):(3'h4)]) ?
                              ((|forvar631) == reg646) : reg632[(1'h1):(1'h1)]) ?
                          wire627[(4'ha):(3'h6)] : {reg641[(3'h4):(2'h2)]});
                      reg665 <= ((|$signed((&forvar662))) || $unsigned((reg656[(1'h0):(1'h0)] ?
                          (+reg640) : $signed(forvar638))));
                    end
                  if ($signed((~&$unsigned($unsigned(reg660)))))
                    begin
                      reg666 <= forvar642;
                    end
                  else
                    begin
                      reg666 <= ($signed(forvar631) * {{$unsigned(wire626)}});
                      reg667 <= (reg651[(1'h1):(1'h0)] ?
                          (+(^~(reg632 ?
                              reg669 : reg673))) : $unsigned(reg669[(2'h3):(2'h2)]));
                      reg668 <= ((!(~&$unsigned(reg645))) ^~ (forvar659 || $unsigned((reg668 <<< (8'ha6)))));
                      reg669 <= (8'ha7);
                    end
                  reg670 <= (~(&reg671[(4'hb):(4'h9)]));
                  for (forvar671 = (1'h0); (forvar671 < (1'h1)); forvar671 = (forvar671 + (1'h1)))
                    begin
                      reg672 <= $signed(reg673[(1'h0):(1'h0)]);
                      reg673 <= {wire623};
                      reg674 <= ((wire625 ~^ reg634[(1'h0):(1'h0)]) ?
                          ($signed((reg672 >> (8'hb3))) - wire623) : reg667[(2'h2):(2'h2)]);
                    end
                end
            end
        end
      else
        begin
          for (forvar631 = (1'h0); (forvar631 < (1'h0)); forvar631 = (forvar631 + (1'h1)))
            begin
              if (($unsigned({(^forvar651)}) ?
                  forvar672[(3'h4):(1'h0)] : reg663))
                begin
                  if ((({(reg666 + (8'ha2))} ?
                      {(reg673 & wire625)} : {(forvar651 ?
                              reg668 : reg673)}) && reg669))
                    begin
                      reg632 <= reg667[(2'h2):(2'h2)];
                      reg633 <= wire626[(4'h8):(1'h0)];
                      reg634 <= ($signed(reg636) << forvar638[(3'h5):(3'h5)]);
                      reg635 <= $unsigned($signed(reg661[(3'h7):(1'h1)]));
                    end
                  else
                    begin
                      reg632 <= {($signed($unsigned(reg634)) <= ((forvar651 | forvar635) || (~|(8'ha5))))};
                      reg633 <= (8'ha3);
                      reg634 <= wire623[(3'h6):(1'h0)];
                    end
                  for (forvar636 = (1'h0); (forvar636 < (2'h3)); forvar636 = (forvar636 + (1'h1)))
                    begin
                      reg637 <= (reg672 >> (reg632 ?
                          $unsigned((+reg653)) : reg653));
                      reg638 <= $signed(reg650);
                    end
                  for (forvar639 = (1'h0); (forvar639 < (2'h3)); forvar639 = (forvar639 + (1'h1)))
                    begin
                      reg640 <= $signed(($unsigned(reg661[(4'ha):(2'h2)]) | {$signed(forvar671)}));
                      reg641 <= reg671;
                      reg642 <= forvar632[(3'h6):(2'h3)];
                    end
                  for (forvar643 = (1'h0); (forvar643 < (2'h2)); forvar643 = (forvar643 + (1'h1)))
                    begin
                      reg644 <= wire623;
                      reg645 <= reg643[(4'hc):(1'h0)];
                      reg646 <= $signed(($signed((!reg674)) >>> ($unsigned(wire625) ?
                          {reg660} : (wire623 ? forvar637 : reg655))));
                      reg647 <= forvar644[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  if ($unsigned((forvar671[(1'h1):(1'h0)] != (8'ha7))))
                    begin
                      reg632 <= reg647;
                    end
                  else
                    begin
                      reg632 <= reg645[(2'h3):(1'h1)];
                    end
                end
              reg648 <= $unsigned((~^wire626[(3'h5):(2'h2)]));
            end
        end
    end
  module675 modinst7428 (wire7427, clk, forvar635, forvar659, forvar662, reg637);
  assign wire7429 = ((&forvar671[(3'h5):(3'h4)]) << ((8'h9c) ?
                        ((reg637 ? reg632 : reg656) ?
                            forvar638 : $unsigned((8'ha2))) : (~&(wire624 ^ reg663))));
  assign wire7430 = {$signed($signed((reg636 ? reg644 : (8'ha4))))};
  assign wire7431 = (^(((forvar632 & forvar635) ?
                            reg652[(4'h9):(3'h7)] : forvar639) ?
                        ((|reg636) ?
                            forvar631[(3'h4):(2'h2)] : {wire629}) : $signed($signed((8'ha2)))));
  assign wire7432 = {{$signed((wire630 >> forvar648))}};
  module4572 modinst7434 (.wire4574(reg656), .y(wire7433), .clk(clk), .wire4575(reg641), .wire4573(forvar635), .wire4576(reg651));
  assign wire7435 = $signed((($signed(forvar662) ?
                            $signed(reg661) : $signed(reg663)) ?
                        ($unsigned(reg668) >= (~|reg660)) : $unsigned({wire7429})));
  always
    @(posedge clk) begin
      if ($signed($unsigned(reg638[(3'h6):(3'h4)])))
        begin
          for (forvar7436 = (1'h0); (forvar7436 < (2'h2)); forvar7436 = (forvar7436 + (1'h1)))
            begin
              for (forvar7437 = (1'h0); (forvar7437 < (1'h0)); forvar7437 = (forvar7437 + (1'h1)))
                begin
                  if (reg672)
                    begin
                      reg7438 <= forvar635[(3'h4):(3'h4)];
                      reg7439 <= (&({forvar637} ?
                          $signed((forvar644 ?
                              reg636 : (8'hb3))) : (|$signed(reg664))));
                      reg7440 <= reg657[(4'h9):(4'h8)];
                      reg7441 <= (^(reg646[(1'h1):(1'h0)] ?
                          reg637[(4'h9):(1'h1)] : $unsigned((reg647 ?
                              forvar671 : reg637))));
                    end
                  else
                    begin
                      reg7438 <= (-(reg7440[(4'h9):(1'h0)] && (reg656 >= {reg663})));
                      reg7439 <= (reg655[(3'h6):(3'h6)] ?
                          (!(reg671[(3'h5):(2'h2)] > (reg649 ?
                              forvar662 : (8'hb6)))) : (~&(+(forvar636 >>> wire7430))));
                    end
                end
              reg7442 <= $unsigned(wire624);
              for (forvar7443 = (1'h0); (forvar7443 < (2'h3)); forvar7443 = (forvar7443 + (1'h1)))
                begin
                  reg7444 <= (8'h9e);
                end
            end
          if ((8'hb1))
            begin
              for (forvar7445 = (1'h0); (forvar7445 < (1'h1)); forvar7445 = (forvar7445 + (1'h1)))
                begin
                  if (reg632)
                    begin
                      reg7446 <= ((^{$unsigned(wire7431)}) == forvar672[(4'hc):(2'h2)]);
                      reg7447 <= ((reg667 != (((8'hb8) <<< forvar667) - (forvar637 ~^ wire7427))) * $unsigned((~|(8'ha8))));
                      reg7448 <= $unsigned(($signed($signed(forvar659)) >>> (8'haf)));
                      reg7449 <= ($unsigned(((reg646 ?
                              wire7427 : (8'hb6)) >> (reg668 ?
                              wire7433 : reg7446))) ?
                          reg7438 : (reg669[(1'h1):(1'h0)] ?
                              (reg661 <= (-(8'hb5))) : $signed((wire7429 | reg640))));
                    end
                  else
                    begin
                      reg7446 <= reg658[(4'ha):(4'ha)];
                      reg7447 <= {{(~|$unsigned(reg672))}};
                      reg7448 <= {$unsigned((^(reg632 ? (8'hb3) : forvar672)))};
                    end
                  for (forvar7450 = (1'h0); (forvar7450 < (1'h1)); forvar7450 = (forvar7450 + (1'h1)))
                    begin
                      reg7451 <= reg632;
                    end
                  if (($signed($unsigned(reg634[(3'h7):(2'h2)])) ?
                      ($unsigned($signed(reg7441)) * $signed((reg667 ?
                          forvar639 : reg7444))) : {reg664}))
                    begin
                      reg7452 <= (reg666[(3'h4):(1'h1)] || $signed($signed($unsigned((8'ha7)))));
                      reg7453 <= reg673[(1'h0):(1'h0)];
                      reg7454 <= $signed((~&($unsigned(forvar7443) ^ (^(8'ha1)))));
                      reg7455 <= reg7440;
                    end
                  else
                    begin
                      reg7452 <= reg668[(3'h6):(3'h5)];
                      reg7453 <= ((|(~|(^reg663))) ?
                          (reg663[(1'h0):(1'h0)] ?
                              ((reg639 ? forvar7445 : reg646) ?
                                  {forvar632} : reg657[(4'h9):(1'h0)]) : reg661[(4'ha):(2'h3)]) : $signed(((~&forvar7443) ?
                              {forvar7443} : reg657)));
                    end
                end
              for (forvar7456 = (1'h0); (forvar7456 < (1'h1)); forvar7456 = (forvar7456 + (1'h1)))
                begin
                  for (forvar7457 = (1'h0); (forvar7457 < (1'h0)); forvar7457 = (forvar7457 + (1'h1)))
                    begin
                      reg7458 <= ((((forvar642 >> wire622) ?
                          (reg7452 && (8'hb1)) : $unsigned(reg7440)) ^ (|(reg649 > reg652))) + reg658[(3'h7):(1'h1)]);
                      reg7459 <= $unsigned((!forvar631[(1'h0):(1'h0)]));
                      reg7460 <= ((($unsigned(wire630) - $signed(reg7442)) & reg664[(1'h1):(1'h1)]) ?
                          ($signed(wire621[(1'h1):(1'h0)]) ?
                              ($signed((8'ha8)) ?
                                  $unsigned(reg643) : forvar7456[(3'h4):(2'h2)]) : (((8'hab) ?
                                      reg635 : reg645) ?
                                  reg7446 : reg660)) : ($signed((reg664 ?
                                  forvar639 : (8'had))) ?
                              (!(^forvar662)) : ((reg633 ?
                                  reg633 : reg646) > forvar672[(3'h7):(2'h3)])));
                    end
                end
              for (forvar7461 = (1'h0); (forvar7461 < (2'h2)); forvar7461 = (forvar7461 + (1'h1)))
                begin
                  for (forvar7462 = (1'h0); (forvar7462 < (1'h1)); forvar7462 = (forvar7462 + (1'h1)))
                    begin
                      reg7463 <= forvar7437;
                    end
                end
            end
          else
            begin
              if ($signed(((&(reg666 ^ (8'ha7))) ?
                  $unsigned($signed(wire630)) : (^~(forvar7436 != reg642)))))
                begin
                  if (((({(8'h9d)} && $signed((8'hb5))) ?
                      $unsigned($unsigned(wire625)) : $unsigned((forvar637 ?
                          forvar643 : forvar648))) & {$signed((&forvar648))}))
                    begin
                      reg7445 <= (reg633 ?
                          $unsigned(((~&wire7435) <= (-reg658))) : (&reg7440));
                      reg7446 <= reg7451[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg7445 <= ($signed(reg7452) ~^ (8'ha0));
                      reg7446 <= $signed($unsigned(((reg656 * reg655) + (reg7458 * reg660))));
                      reg7447 <= ($signed(reg7438[(4'h9):(4'h8)]) == $signed(reg7463));
                    end
                  for (forvar7448 = (1'h0); (forvar7448 < (1'h0)); forvar7448 = (forvar7448 + (1'h1)))
                    begin
                      reg7449 <= (($unsigned((-forvar7448)) ?
                              ((reg7455 | wire623) ^ (wire628 ?
                                  wire7430 : forvar7457)) : (reg7441[(2'h3):(2'h3)] ?
                                  (~reg649) : (reg668 == (8'ha4)))) ?
                          {(^$signed(reg656))} : reg7451[(3'h5):(3'h4)]);
                    end
                end
              else
                begin
                  for (forvar7445 = (1'h0); (forvar7445 < (1'h0)); forvar7445 = (forvar7445 + (1'h1)))
                    begin
                      reg7446 <= (~reg650);
                      reg7447 <= $unsigned(forvar643[(4'h8):(3'h5)]);
                      reg7448 <= $signed($unsigned($unsigned($unsigned(reg7441))));
                      reg7449 <= (forvar651[(1'h1):(1'h1)] ?
                          $signed($unsigned(forvar632)) : $signed(reg656[(3'h5):(3'h5)]));
                    end
                  if ($signed(((~|((8'h9d) ? reg668 : wire7429)) ?
                      $unsigned(reg7445) : (-$unsigned(forvar7436)))))
                    begin
                      reg7450 <= (!forvar654[(3'h5):(2'h2)]);
                      reg7451 <= (~(!$signed(wire621[(2'h3):(1'h0)])));
                    end
                  else
                    begin
                      reg7450 <= {wire7432};
                      reg7451 <= (($signed({reg7463}) == reg673[(2'h3):(1'h0)]) ?
                          reg652[(4'he):(4'ha)] : $signed($signed(forvar636[(3'h4):(1'h1)])));
                    end
                  if ($unsigned($signed({{(8'hae)}})))
                    begin
                      reg7452 <= ((^~(~^wire624[(3'h7):(3'h5)])) ?
                          (!(~^{reg646})) : $signed($unsigned(wire625[(4'h9):(3'h5)])));
                      reg7453 <= {reg666[(1'h1):(1'h0)]};
                      reg7454 <= forvar7450[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg7452 <= (($unsigned(reg672) ?
                          $signed((|reg7459)) : $unsigned($unsigned(reg656))) > $unsigned((wire629 ?
                          (reg7447 ~^ reg661) : {(8'ha7)})));
                      reg7453 <= ({$unsigned(forvar639)} ?
                          ((~^$signed((8'hb9))) ?
                              $unsigned(reg7438[(4'ha):(3'h6)]) : ((forvar635 < reg7450) ^~ $unsigned(wire7435))) : $signed($signed((8'haf))));
                      reg7454 <= forvar644[(1'h0):(1'h0)];
                    end
                end
              reg7455 <= ($unsigned({reg647[(3'h7):(3'h4)]}) ?
                  reg7446 : $signed(((8'ha6) <<< (~|reg7454))));
              if ((&($unsigned((+reg7460)) ?
                  reg636[(3'h4):(2'h2)] : $unsigned($unsigned((8'hb1))))))
                begin
                  for (forvar7456 = (1'h0); (forvar7456 < (1'h1)); forvar7456 = (forvar7456 + (1'h1)))
                    begin
                      reg7457 <= wire630;
                      reg7458 <= ((+(!(!reg7450))) >> $unsigned(($signed(forvar639) ?
                          {reg641} : (reg637 && forvar667))));
                    end
                end
              else
                begin
                  reg7456 <= $signed((8'haf));
                  reg7457 <= (~|reg633[(1'h1):(1'h1)]);
                  if ($unsigned(reg7454))
                    begin
                      reg7458 <= (!(~^(reg7457[(3'h5):(3'h5)] ?
                          $unsigned(forvar7437) : wire629[(3'h6):(3'h4)])));
                      reg7459 <= {((&reg7448[(1'h1):(1'h0)]) && $unsigned((reg647 && reg7451)))};
                      reg7460 <= reg673[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg7458 <= $signed(({{(8'ha6)}} ?
                          $unsigned({reg7457}) : $unsigned(wire629)));
                      reg7459 <= (reg664 == (8'ha0));
                    end
                  if ($signed(((~^(^(8'hb5))) >= (reg660[(3'h5):(3'h5)] ?
                      $signed(forvar7448) : ((8'hab) ? reg639 : reg635)))))
                    begin
                      reg7461 <= reg649;
                    end
                  else
                    begin
                      reg7461 <= reg7444;
                    end
                end
              if ((forvar671[(1'h1):(1'h0)] ^ {(reg7439[(2'h2):(2'h2)] >= reg644[(1'h0):(1'h0)])}))
                begin
                  if (((8'hb9) < $signed($signed((wire622 ?
                      reg7438 : reg7452)))))
                    begin
                      reg7462 <= reg663;
                      reg7463 <= (~(~(|forvar632[(3'h4):(3'h4)])));
                      reg7464 <= ($signed(forvar7461[(3'h5):(2'h2)]) || ({forvar7461} ?
                          $signed((wire7429 < forvar671)) : reg660[(1'h0):(1'h0)]));
                      reg7465 <= {((reg7446[(3'h7):(1'h0)] ?
                                  $signed(forvar672) : forvar667[(3'h5):(1'h0)]) ?
                              reg7458[(2'h2):(2'h2)] : $unsigned(reg7459[(2'h3):(2'h3)]))};
                    end
                  else
                    begin
                      reg7462 <= $unsigned(($unsigned((forvar7436 < reg7455)) == $signed(reg660[(3'h4):(2'h3)])));
                    end
                  for (forvar7466 = (1'h0); (forvar7466 < (2'h2)); forvar7466 = (forvar7466 + (1'h1)))
                    begin
                      reg7467 <= (forvar638 ?
                          ($signed(reg7457) - ((reg634 ?
                              reg7465 : forvar642) != (reg634 != wire623))) : forvar651[(1'h0):(1'h0)]);
                      reg7468 <= (forvar7466 || ((reg7460 > (reg7440 >> forvar662)) ?
                          (~$unsigned(forvar637)) : forvar7448[(2'h2):(1'h0)]));
                    end
                  reg7469 <= (~|$unsigned({(8'ha3)}));
                  for (forvar7470 = (1'h0); (forvar7470 < (1'h0)); forvar7470 = (forvar7470 + (1'h1)))
                    begin
                      reg7471 <= (forvar7450 ?
                          $unsigned($unsigned((8'ha3))) : (((forvar7462 & reg636) ?
                              (^~reg668) : (~&wire7433)) <<< (|reg651)));
                      reg7472 <= $signed(($signed(((8'hb5) | reg637)) >> ((8'ha9) ?
                          $signed(reg673) : (reg670 ? wire7429 : wire7433))));
                      reg7473 <= (|(((reg652 ?
                              reg7444 : forvar7457) >> (reg656 ?
                              reg7447 : reg641)) ?
                          $unsigned(forvar7443[(4'hd):(3'h7)]) : (reg7444 <= $unsigned(reg672))));
                    end
                end
              else
                begin
                  for (forvar7462 = (1'h0); (forvar7462 < (2'h2)); forvar7462 = (forvar7462 + (1'h1)))
                    begin
                      reg7463 <= ($unsigned({$signed(forvar7443)}) ?
                          reg7461[(2'h2):(2'h2)] : $unsigned({$unsigned(reg633)}));
                      reg7464 <= (forvar7456 ?
                          (|{(forvar667 ^ reg656)}) : (((reg7473 ?
                                  reg7450 : reg7458) + (reg7438 > reg670)) ?
                              $signed($unsigned((8'hab))) : reg658));
                      reg7465 <= (+$signed({{reg7446}}));
                    end
                  if ((($signed((&forvar672)) == (&(reg650 | (8'hb1)))) ?
                      reg650[(3'h6):(1'h1)] : (({forvar643} | {forvar672}) >> (&(8'hb4)))))
                    begin
                      reg7466 <= (~&(^~($signed(reg642) ?
                          $unsigned(reg643) : reg652)));
                      reg7467 <= $signed({($signed(wire626) + (reg643 <<< reg7458))});
                      reg7468 <= {(^~{$unsigned(reg647)})};
                      reg7469 <= {$signed(((+reg7447) ?
                              $signed(reg661) : forvar639[(3'h4):(1'h1)]))};
                    end
                  else
                    begin
                      reg7466 <= ($signed((8'hb5)) ?
                          ({$unsigned(forvar7462)} >= reg657) : reg653);
                      reg7467 <= (wire7433 ^ $signed((8'haf)));
                      reg7468 <= (~&$unsigned(((reg644 || reg7463) << reg7466)));
                      reg7469 <= $unsigned($signed(reg656[(4'ha):(4'h9)]));
                    end
                  for (forvar7470 = (1'h0); (forvar7470 < (1'h0)); forvar7470 = (forvar7470 + (1'h1)))
                    begin
                      reg7471 <= (8'hb7);
                      reg7472 <= reg7469;
                      reg7473 <= $unsigned($signed($unsigned(reg672)));
                      reg7474 <= (8'had);
                    end
                  for (forvar7475 = (1'h0); (forvar7475 < (2'h3)); forvar7475 = (forvar7475 + (1'h1)))
                    begin
                      reg7476 <= reg635;
                    end
                end
            end
        end
      else
        begin
          if ($signed({$unsigned(((8'hb0) ? forvar7436 : (8'h9c)))}))
            begin
              if (reg636[(4'h9):(2'h2)])
                begin
                  if (reg656)
                    begin
                      reg7436 <= (^~wire7435);
                      reg7437 <= (8'ha7);
                    end
                  else
                    begin
                      reg7436 <= $signed(reg666);
                      reg7437 <= reg637;
                    end
                end
              else
                begin
                  if (forvar637[(1'h1):(1'h0)])
                    begin
                      reg7436 <= (-$signed($signed((reg634 ?
                          reg666 : reg647))));
                      reg7437 <= (($unsigned($unsigned(reg7466)) ?
                              (|{reg7456}) : (+(forvar671 + forvar7462))) ?
                          (~^((reg7452 ?
                              reg7454 : reg644) ~^ reg632[(3'h4):(2'h2)])) : (~^forvar7462));
                    end
                  else
                    begin
                      reg7436 <= {(~^reg7461)};
                    end
                  for (forvar7438 = (1'h0); (forvar7438 < (1'h0)); forvar7438 = (forvar7438 + (1'h1)))
                    begin
                      reg7439 <= forvar651[(2'h2):(1'h1)];
                      reg7440 <= reg638;
                    end
                end
              for (forvar7441 = (1'h0); (forvar7441 < (1'h1)); forvar7441 = (forvar7441 + (1'h1)))
                begin
                  reg7442 <= forvar7445;
                end
              for (forvar7443 = (1'h0); (forvar7443 < (1'h0)); forvar7443 = (forvar7443 + (1'h1)))
                begin
                  reg7444 <= ((+$signed($signed(reg7440))) ~^ ($unsigned(forvar7462) && {(^reg645)}));
                  if ((((((8'hb1) ? reg7460 : wire627) ^ (~^(8'hb1))) ?
                      $signed(reg674[(2'h2):(1'h0)]) : ($unsigned(wire7431) && ((8'hb1) ^~ (8'hb0)))) != (reg7451[(1'h0):(1'h0)] ?
                      (reg7437 > (reg7469 >>> reg674)) : $unsigned({(8'hb7)}))))
                    begin
                      reg7445 <= $signed((8'hb1));
                      reg7446 <= forvar671;
                    end
                  else
                    begin
                      reg7445 <= reg632[(3'h5):(2'h3)];
                      reg7446 <= reg7448[(4'hb):(4'hb)];
                      reg7447 <= {$unsigned($unsigned((|(8'ha3))))};
                    end
                  for (forvar7448 = (1'h0); (forvar7448 < (1'h1)); forvar7448 = (forvar7448 + (1'h1)))
                    begin
                      reg7449 <= wire629[(1'h0):(1'h0)];
                      reg7450 <= ($unsigned(reg666) > $signed($signed(wire7432[(4'ha):(2'h2)])));
                      reg7451 <= (~|((reg7453[(3'h7):(2'h2)] ?
                          $unsigned(forvar639) : forvar635[(3'h6):(1'h0)]) >= reg656[(2'h3):(2'h3)]));
                    end
                  reg7452 <= wire7429[(4'hf):(4'he)];
                end
            end
          else
            begin
              if ($signed(reg7439[(1'h0):(1'h0)]))
                begin
                  if ((($unsigned($signed(reg7449)) >>> {(reg7457 ?
                          reg641 : forvar643)}) ~^ $unsigned((!reg7449))))
                    begin
                      reg7436 <= $unsigned($signed(reg7442[(2'h3):(2'h3)]));
                      reg7437 <= $unsigned($unsigned((~|reg652[(3'h6):(3'h4)])));
                      reg7438 <= forvar7443[(4'h9):(1'h1)];
                      reg7439 <= reg634;
                    end
                  else
                    begin
                      reg7436 <= (reg643[(1'h1):(1'h0)] ?
                          (-(~^{reg7442})) : (((reg637 || reg650) <= reg7451[(1'h0):(1'h0)]) * wire7433));
                      reg7437 <= $unsigned($signed($signed($unsigned(reg7437))));
                      reg7438 <= reg7476[(4'h8):(3'h4)];
                      reg7439 <= ((&($signed(reg632) >>> $unsigned(forvar638))) ?
                          $signed((-(^~forvar7457))) : forvar662[(4'hd):(1'h1)]);
                    end
                  for (forvar7440 = (1'h0); (forvar7440 < (2'h2)); forvar7440 = (forvar7440 + (1'h1)))
                    begin
                      reg7441 <= ((~^(^$signed(reg640))) * reg665);
                    end
                  for (forvar7442 = (1'h0); (forvar7442 < (2'h3)); forvar7442 = (forvar7442 + (1'h1)))
                    begin
                      reg7443 <= (reg669 ?
                          $signed(($signed(forvar7450) * (forvar671 ?
                              reg638 : forvar639))) : {(((8'ha5) ~^ reg7436) ?
                                  (forvar7442 + reg7450) : (reg7455 ?
                                      (8'ha4) : (8'hac)))});
                      reg7444 <= $unsigned($unsigned(((forvar7448 >>> reg7476) == $unsigned(reg7439))));
                      reg7445 <= $unsigned($signed($signed(reg7476[(2'h3):(2'h3)])));
                    end
                end
              else
                begin
                  for (forvar7436 = (1'h0); (forvar7436 < (2'h2)); forvar7436 = (forvar7436 + (1'h1)))
                    begin
                      reg7437 <= $unsigned({$unsigned(reg7456)});
                      reg7438 <= reg656;
                      reg7439 <= {{$signed({(8'hb3)})}};
                      reg7440 <= ($unsigned(reg668[(2'h3):(1'h1)]) | (^~{(-reg657)}));
                    end
                end
              for (forvar7446 = (1'h0); (forvar7446 < (1'h1)); forvar7446 = (forvar7446 + (1'h1)))
                begin
                  reg7447 <= (((&$signed(reg650)) > {$unsigned(forvar648)}) == ((~&$signed(reg7467)) > reg7441));
                end
              reg7448 <= {(($unsigned(reg653) ?
                          $unsigned(reg639) : (forvar7436 >> reg7464)) ?
                      $unsigned($unsigned(forvar7446)) : {forvar7448[(2'h3):(1'h1)]})};
              for (forvar7449 = (1'h0); (forvar7449 < (2'h2)); forvar7449 = (forvar7449 + (1'h1)))
                begin
                  if ({((8'hb1) ?
                          $unsigned((|(8'ha4))) : (!$unsigned((8'hb8))))})
                    begin
                      reg7450 <= ({reg7437} ?
                          (forvar7436[(2'h3):(1'h0)] ?
                              (&(~|forvar654)) : $signed((wire7427 ~^ forvar7437))) : $unsigned($signed(reg7466[(4'he):(1'h1)])));
                    end
                  else
                    begin
                      reg7450 <= ($signed(forvar635) && ($signed(reg638) ?
                          (^~$signed(wire627)) : reg669));
                      reg7451 <= reg637;
                      reg7452 <= ({({forvar635} ?
                              forvar648 : (reg661 ^~ forvar651))} + (8'had));
                      reg7453 <= reg7457[(4'hb):(4'h8)];
                    end
                  for (forvar7454 = (1'h0); (forvar7454 < (1'h0)); forvar7454 = (forvar7454 + (1'h1)))
                    begin
                      reg7455 <= reg650[(4'hf):(3'h7)];
                      reg7456 <= (+reg635);
                      reg7457 <= (~^reg638[(1'h0):(1'h0)]);
                    end
                end
            end
        end
      for (forvar7477 = (1'h0); (forvar7477 < (2'h2)); forvar7477 = (forvar7477 + (1'h1)))
        begin
          for (forvar7478 = (1'h0); (forvar7478 < (2'h2)); forvar7478 = (forvar7478 + (1'h1)))
            begin
              for (forvar7479 = (1'h0); (forvar7479 < (1'h1)); forvar7479 = (forvar7479 + (1'h1)))
                begin
                  if (reg7445)
                    begin
                      reg7480 <= $signed({$signed((reg644 ?
                              (8'ha0) : reg7465))});
                      reg7481 <= ((~&$signed((reg7474 ?
                          (8'ha9) : reg645))) <<< $signed(((~reg660) < (reg7476 ?
                          reg651 : wire621))));
                    end
                  else
                    begin
                      reg7480 <= (forvar7461 ?
                          ((~|(^reg661)) ?
                              (~reg671) : reg634[(3'h5):(2'h2)]) : reg7453);
                    end
                  for (forvar7482 = (1'h0); (forvar7482 < (1'h0)); forvar7482 = (forvar7482 + (1'h1)))
                    begin
                      reg7483 <= {({forvar7448[(2'h3):(2'h3)]} <= $unsigned($unsigned(forvar636)))};
                      reg7484 <= reg7436;
                      reg7485 <= ($unsigned($unsigned(reg7441[(4'hb):(4'h8)])) ^ reg7438[(1'h1):(1'h1)]);
                    end
                  reg7486 <= ((^((&forvar7446) == (reg7464 < forvar671))) ?
                      $unsigned($unsigned((~^reg7469))) : $signed((reg7461[(1'h0):(1'h0)] ?
                          $unsigned((8'hb5)) : (&forvar7441))));
                end
            end
        end
      for (forvar7487 = (1'h0); (forvar7487 < (2'h3)); forvar7487 = (forvar7487 + (1'h1)))
        begin
          for (forvar7488 = (1'h0); (forvar7488 < (1'h1)); forvar7488 = (forvar7488 + (1'h1)))
            begin
              reg7489 <= ($signed(reg7485[(3'h4):(2'h2)]) ?
                  (reg7446[(4'h8):(3'h5)] ?
                      reg7440[(4'hc):(4'h8)] : $unsigned((forvar7449 <= wire7431))) : {$unsigned(((8'ha4) ?
                          (8'hb1) : reg635))});
              if ((wire621[(2'h3):(2'h2)] ?
                  (^~reg640) : (~|{(reg7446 ? (8'hb6) : forvar7475)})))
                begin
                  for (forvar7490 = (1'h0); (forvar7490 < (2'h2)); forvar7490 = (forvar7490 + (1'h1)))
                    begin
                      reg7491 <= reg635[(3'h6):(1'h1)];
                      reg7492 <= $signed({forvar671[(1'h1):(1'h1)]});
                    end
                  for (forvar7493 = (1'h0); (forvar7493 < (1'h0)); forvar7493 = (forvar7493 + (1'h1)))
                    begin
                      reg7494 <= ((^~(forvar7446[(1'h1):(1'h0)] == (reg633 ?
                              forvar7493 : forvar7461))) ?
                          ({$signed(reg639)} ?
                              ($unsigned((8'ha7)) ?
                                  forvar7437 : $signed((8'ha0))) : $signed(((8'had) ?
                                  reg7486 : wire629))) : (reg635[(3'h4):(2'h2)] ?
                              $unsigned($unsigned(reg7468)) : ((~(8'ha3)) & forvar635[(4'hb):(3'h6)])));
                      reg7495 <= $signed(((8'hb6) > ((reg645 < reg7476) ?
                          (forvar7466 != wire624) : $signed(reg7469))));
                      reg7496 <= $unsigned((+(~{reg7447})));
                      reg7497 <= reg650;
                    end
                  if (reg7486)
                    begin
                      reg7498 <= forvar667[(4'h8):(1'h0)];
                      reg7499 <= $signed(($signed($unsigned((8'hb8))) ?
                          reg7472[(3'h7):(3'h5)] : reg7467));
                    end
                  else
                    begin
                      reg7498 <= reg7489;
                      reg7499 <= forvar644;
                    end
                end
              else
                begin
                  for (forvar7490 = (1'h0); (forvar7490 < (1'h1)); forvar7490 = (forvar7490 + (1'h1)))
                    begin
                      reg7491 <= ({($signed(reg641) ?
                                  $unsigned((8'ha1)) : reg7469[(2'h2):(1'h0)])} ?
                          ((-reg667[(1'h0):(1'h0)]) ?
                              (~&(forvar638 << (8'ha2))) : $signed((+(8'ha7)))) : reg7451);
                      reg7492 <= ({($unsigned(reg7483) != (-reg7461))} >>> $unsigned($signed(((8'ha4) >> wire7432))));
                      reg7493 <= reg7458[(4'h8):(3'h4)];
                      reg7494 <= reg7481[(4'he):(4'hc)];
                    end
                end
              if ({forvar7437[(3'h4):(3'h4)]})
                begin
                  reg7500 <= ($unsigned(((^~reg666) >= reg650[(3'h4):(2'h2)])) ~^ $unsigned((!$unsigned(forvar671))));
                  reg7501 <= reg643;
                  if ({wire7432})
                    begin
                      reg7502 <= reg7436;
                      reg7503 <= (^~$signed(reg7494));
                    end
                  else
                    begin
                      reg7502 <= reg640[(3'h7):(1'h0)];
                      reg7503 <= (&reg7484[(4'hc):(1'h1)]);
                      reg7504 <= reg669;
                      reg7505 <= $unsigned(reg7474[(4'ha):(4'h8)]);
                    end
                  reg7506 <= {$signed((reg7504[(4'h9):(1'h1)] ?
                          $signed(reg7505) : $unsigned((8'hb3))))};
                end
              else
                begin
                  if ((~^reg7461[(1'h1):(1'h0)]))
                    begin
                      reg7500 <= {((-{forvar642}) || reg672[(1'h1):(1'h0)])};
                    end
                  else
                    begin
                      reg7500 <= (($signed((^~forvar648)) - {$unsigned(reg645)}) == (reg7438[(4'h9):(1'h1)] ?
                          ((reg650 ?
                              reg7463 : (8'hb7)) == {forvar662}) : reg632[(3'h6):(2'h2)]));
                      reg7501 <= (~$unsigned($unsigned((forvar7438 ?
                          wire7431 : wire7429))));
                      reg7502 <= ((^~reg7497[(2'h2):(1'h0)]) ?
                          forvar637 : (forvar636 ?
                              forvar7438 : (+$unsigned(forvar672))));
                    end
                end
              for (forvar7507 = (1'h0); (forvar7507 < (1'h1)); forvar7507 = (forvar7507 + (1'h1)))
                begin
                  for (forvar7508 = (1'h0); (forvar7508 < (2'h2)); forvar7508 = (forvar7508 + (1'h1)))
                    begin
                      reg7509 <= {(!$unsigned((&reg7463)))};
                      reg7510 <= $unsigned(reg7501[(2'h3):(2'h2)]);
                      reg7511 <= $unsigned(reg7439);
                      reg7512 <= (8'h9d);
                    end
                  if (reg647)
                    begin
                      reg7513 <= {((forvar7441[(2'h3):(2'h2)] ?
                                  (forvar7436 | forvar638) : $signed(reg7459)) ?
                              ($unsigned((8'hb5)) ?
                                  reg7480[(3'h5):(2'h2)] : (forvar7477 ?
                                      reg7510 : reg648)) : ((forvar7438 ?
                                  reg7501 : reg7499) > reg7501[(3'h5):(3'h5)]))};
                    end
                  else
                    begin
                      reg7513 <= wire623;
                    end
                  for (forvar7514 = (1'h0); (forvar7514 < (2'h2)); forvar7514 = (forvar7514 + (1'h1)))
                    begin
                      reg7515 <= ((!$unsigned((+reg7460))) || $unsigned(({forvar7462} >> $signed(forvar662))));
                      reg7516 <= $unsigned(reg7510);
                      reg7517 <= reg7449;
                      reg7518 <= reg646[(2'h3):(1'h0)];
                    end
                end
            end
          for (forvar7519 = (1'h0); (forvar7519 < (2'h2)); forvar7519 = (forvar7519 + (1'h1)))
            begin
              reg7520 <= reg7438[(3'h4):(1'h1)];
              reg7521 <= (-(|$unsigned((-(8'haf)))));
              for (forvar7522 = (1'h0); (forvar7522 < (2'h3)); forvar7522 = (forvar7522 + (1'h1)))
                begin
                  for (forvar7523 = (1'h0); (forvar7523 < (1'h0)); forvar7523 = (forvar7523 + (1'h1)))
                    begin
                      reg7524 <= {{($unsigned(reg7484) ?
                                  forvar648[(1'h0):(1'h0)] : (reg7474 ?
                                      forvar7514 : wire626))}};
                      reg7525 <= (+((^forvar7437) ?
                          (~&reg7501[(1'h0):(1'h0)]) : wire7435[(1'h1):(1'h1)]));
                      reg7526 <= $signed($unsigned(reg7489));
                    end
                end
              reg7527 <= $unsigned(((~|$unsigned((8'hb2))) ?
                  ($signed(reg7451) ? reg646 : (~|forvar7475)) : (forvar636 ?
                      {forvar7445} : reg7509)));
            end
        end
      for (forvar7528 = (1'h0); (forvar7528 < (1'h0)); forvar7528 = (forvar7528 + (1'h1)))
        begin
          reg7529 <= (8'hb7);
          if (forvar7462[(2'h3):(2'h2)])
            begin
              for (forvar7530 = (1'h0); (forvar7530 < (2'h2)); forvar7530 = (forvar7530 + (1'h1)))
                begin
                  for (forvar7531 = (1'h0); (forvar7531 < (1'h0)); forvar7531 = (forvar7531 + (1'h1)))
                    begin
                      reg7532 <= (wire621 ?
                          reg651 : $signed(reg642[(1'h0):(1'h0)]));
                      reg7533 <= (~(reg637 || $unsigned((reg7483 ~^ reg667))));
                      reg7534 <= (reg7526 ?
                          ($unsigned($unsigned((8'ha6))) && {(forvar7456 <= reg633)}) : wire629[(3'h5):(2'h3)]);
                      reg7535 <= (~reg646);
                    end
                end
            end
          else
            begin
              for (forvar7530 = (1'h0); (forvar7530 < (1'h0)); forvar7530 = (forvar7530 + (1'h1)))
                begin
                  if ($signed($unsigned({((8'ha4) ? forvar7477 : (8'hb6))})))
                    begin
                      reg7531 <= ((forvar7479 <<< $unsigned((8'hba))) ?
                          reg7473 : ($unsigned($unsigned((8'ha6))) > $unsigned(forvar7479)));
                    end
                  else
                    begin
                      reg7531 <= (~|(8'h9e));
                      reg7532 <= forvar7482[(3'h6):(3'h6)];
                      reg7533 <= $unsigned({reg656});
                      reg7534 <= (+{(forvar636 <<< $signed(reg7436))});
                    end
                  if ((({(+forvar7522)} ?
                      forvar7522[(3'h5):(1'h1)] : forvar7479) != $signed((&$signed(reg638)))))
                    begin
                      reg7535 <= ($signed(((reg672 >> forvar7531) ^~ (wire7429 | reg7502))) - ({$unsigned(forvar7487)} ?
                          {$signed(reg639)} : forvar672));
                      reg7536 <= $signed(reg673);
                      reg7537 <= reg7480;
                      reg7538 <= (((reg635[(2'h3):(1'h0)] << $unsigned(reg7466)) + $signed(((8'hb2) > wire629))) == forvar7437[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg7535 <= $unsigned((reg7483[(2'h2):(2'h2)] ?
                          (^{reg7538}) : {reg643}));
                      reg7536 <= $signed($signed({wire624}));
                    end
                end
              if (reg7463)
                begin
                  reg7539 <= (-$unsigned((^(reg7468 > reg653))));
                  if (((&$signed((~|wire7430))) || $signed({(+reg651)})))
                    begin
                      reg7540 <= reg7489;
                      reg7541 <= ({$signed((reg7457 ? reg7459 : forvar7482))} ?
                          (forvar7454 != $unsigned((^forvar642))) : (($signed(reg651) >= $unsigned((8'h9d))) ?
                              reg7486 : ({reg7511} < reg7484[(4'hc):(3'h5)])));
                    end
                  else
                    begin
                      reg7540 <= reg7456;
                      reg7541 <= ($unsigned($unsigned((reg7455 * forvar7531))) ?
                          (reg7534[(2'h3):(2'h2)] ?
                              reg660[(3'h4):(3'h4)] : (~|(reg7453 ?
                                  wire625 : (8'hb9)))) : $unsigned($signed(reg7448)));
                      reg7542 <= $unsigned({((reg7500 ?
                              forvar648 : (8'ha5)) * ((8'hb0) && wire624))});
                    end
                  if (($signed({(&(8'ha3))}) ?
                      (forvar7438 * {(reg7446 ~^ forvar7531)}) : $unsigned((^reg635[(1'h1):(1'h0)]))))
                    begin
                      reg7543 <= $signed(wire7435[(2'h2):(2'h2)]);
                      reg7544 <= reg650;
                    end
                  else
                    begin
                      reg7543 <= forvar7531[(4'h8):(3'h7)];
                      reg7544 <= reg665[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar7539 = (1'h0); (forvar7539 < (2'h3)); forvar7539 = (forvar7539 + (1'h1)))
                    begin
                      reg7540 <= $unsigned(($signed($unsigned((8'h9e))) + (~&(8'hb1))));
                      reg7541 <= $signed($unsigned((&(forvar7450 < reg7543))));
                      reg7542 <= $unsigned($signed(forvar639[(2'h3):(2'h3)]));
                    end
                  for (forvar7543 = (1'h0); (forvar7543 < (1'h0)); forvar7543 = (forvar7543 + (1'h1)))
                    begin
                      reg7544 <= $signed((((reg7521 < wire624) + (^~reg7491)) + ((^reg634) << (8'haa))));
                      reg7545 <= (forvar7477 >= $unsigned(((^reg638) ^~ $unsigned(reg671))));
                    end
                end
            end
          if (($unsigned($signed($unsigned(reg671))) > ({{(8'ha6)}} || $unsigned((~|(8'h9e))))))
            begin
              reg7546 <= ({($signed(wire627) ?
                      forvar7448 : forvar7443[(4'hc):(2'h2)])} || ({$unsigned(reg7450)} ?
                  $signed(reg656) : (~(&forvar7530))));
            end
          else
            begin
              for (forvar7546 = (1'h0); (forvar7546 < (1'h0)); forvar7546 = (forvar7546 + (1'h1)))
                begin
                  if ((-reg7440[(1'h1):(1'h0)]))
                    begin
                      reg7547 <= $unsigned($unsigned($signed({(8'h9d)})));
                      reg7548 <= (($unsigned($signed(forvar7523)) ?
                              reg655[(3'h7):(2'h3)] : forvar7482) ?
                          {{reg651[(3'h7):(3'h7)]}} : ($unsigned($unsigned(reg7464)) <<< $signed($signed(reg7444))));
                      reg7549 <= reg7526;
                      reg7550 <= (reg7529[(1'h1):(1'h1)] >> (~|{reg7464[(3'h6):(1'h0)]}));
                    end
                  else
                    begin
                      reg7547 <= reg7544;
                      reg7548 <= (($signed($unsigned(reg7529)) ?
                          $unsigned((reg7529 > reg7512)) : reg7454) == (reg7509 ?
                          ((8'h9f) <<< ((8'h9f) >= reg7516)) : (~(^~reg7466))));
                      reg7549 <= (8'h9e);
                    end
                  for (forvar7551 = (1'h0); (forvar7551 < (1'h0)); forvar7551 = (forvar7551 + (1'h1)))
                    begin
                      reg7552 <= $unsigned(forvar7450[(2'h3):(2'h2)]);
                      reg7553 <= (((~&(!reg7513)) ?
                          forvar7446 : ($unsigned(reg644) ?
                              (reg7436 ?
                                  reg7459 : (8'hab)) : $signed(forvar671))) * reg645[(3'h4):(1'h1)]);
                    end
                  reg7554 <= $unsigned($signed($signed(reg7449[(2'h3):(1'h0)])));
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar7555 = (1'h0); (forvar7555 < (2'h2)); forvar7555 = (forvar7555 + (1'h1)))
        begin
          reg7556 <= $signed((|{forvar7523}));
          for (forvar7557 = (1'h0); (forvar7557 < (1'h1)); forvar7557 = (forvar7557 + (1'h1)))
            begin
              for (forvar7558 = (1'h0); (forvar7558 < (1'h0)); forvar7558 = (forvar7558 + (1'h1)))
                begin
                  reg7559 <= ($unsigned($unsigned(reg7442[(1'h0):(1'h0)])) | reg7496);
                  if (reg7467)
                    begin
                      reg7560 <= $signed((~forvar7482[(3'h4):(3'h4)]));
                    end
                  else
                    begin
                      reg7560 <= forvar7456;
                      reg7561 <= forvar642;
                      reg7562 <= forvar7557[(4'hc):(4'h8)];
                      reg7563 <= $signed($signed((forvar7443[(2'h2):(2'h2)] ?
                          (forvar7555 ? reg647 : reg7436) : $signed(reg635))));
                    end
                  reg7564 <= $signed((wire628[(2'h3):(1'h1)] < reg7546[(1'h0):(1'h0)]));
                end
              for (forvar7565 = (1'h0); (forvar7565 < (2'h2)); forvar7565 = (forvar7565 + (1'h1)))
                begin
                  if (({forvar7546[(1'h0):(1'h0)]} ?
                      reg7469[(1'h1):(1'h1)] : $unsigned((reg7513[(4'hb):(2'h3)] ?
                          (reg7447 ^ forvar7446) : reg7502[(2'h2):(2'h2)]))))
                    begin
                      reg7566 <= (~|reg670[(3'h4):(3'h4)]);
                      reg7567 <= (-$signed(((&(8'hb8)) << $signed(reg643))));
                      reg7568 <= forvar7528;
                      reg7569 <= (8'hb2);
                    end
                  else
                    begin
                      reg7566 <= $unsigned({$signed((8'haa))});
                      reg7567 <= (reg7568 ?
                          (~{(reg7510 || reg7493)}) : reg7484[(4'hb):(4'ha)]);
                    end
                  for (forvar7570 = (1'h0); (forvar7570 < (1'h0)); forvar7570 = (forvar7570 + (1'h1)))
                    begin
                      reg7571 <= wire629;
                      reg7572 <= $unsigned($unsigned((forvar7470 && (forvar7490 ?
                          forvar7470 : (8'hac)))));
                      reg7573 <= (|forvar648[(1'h0):(1'h0)]);
                    end
                end
            end
          if ((-wire626))
            begin
              for (forvar7574 = (1'h0); (forvar7574 < (1'h1)); forvar7574 = (forvar7574 + (1'h1)))
                begin
                  if ({forvar632[(2'h3):(2'h3)]})
                    begin
                      reg7575 <= (~&(&(^$signed(reg7560))));
                    end
                  else
                    begin
                      reg7575 <= reg7471[(1'h0):(1'h0)];
                    end
                end
              for (forvar7576 = (1'h0); (forvar7576 < (2'h2)); forvar7576 = (forvar7576 + (1'h1)))
                begin
                  for (forvar7577 = (1'h0); (forvar7577 < (1'h1)); forvar7577 = (forvar7577 + (1'h1)))
                    begin
                      reg7578 <= $signed($unsigned($signed($unsigned(forvar7457))));
                      reg7579 <= {((+$signed(reg7505)) - ((reg7527 ?
                              reg7493 : reg7575) == $signed(reg7521)))};
                      reg7580 <= (&($unsigned($signed(forvar7523)) || forvar7530));
                    end
                  if ((((8'ha4) ?
                      $unsigned(reg7543[(2'h3):(2'h3)]) : (reg7453[(3'h4):(2'h3)] || (~&reg643))) ~^ $signed((forvar7523 ?
                      $unsigned(reg671) : forvar7475[(3'h5):(2'h3)]))))
                    begin
                      reg7581 <= (reg7454[(1'h1):(1'h1)] && ($unsigned($unsigned(forvar7507)) * (reg7550 << (^reg7532))));
                    end
                  else
                    begin
                      reg7581 <= reg7469;
                      reg7582 <= (($unsigned({reg7498}) ?
                              ((|reg7567) ^~ forvar7479[(4'hc):(3'h5)]) : {{forvar7462}}) ?
                          (8'h9c) : $unsigned(reg7520));
                      reg7583 <= forvar7442;
                    end
                end
              reg7584 <= reg7506[(1'h0):(1'h0)];
              if ((+forvar7457[(3'h4):(2'h3)]))
                begin
                  for (forvar7585 = (1'h0); (forvar7585 < (2'h3)); forvar7585 = (forvar7585 + (1'h1)))
                    begin
                      reg7586 <= reg7543;
                    end
                  if (forvar672)
                    begin
                      reg7587 <= $signed((!(reg7439[(4'h9):(2'h2)] >= reg7552[(2'h3):(1'h0)])));
                      reg7588 <= ((-({reg7474} && $unsigned(reg7498))) != $unsigned({(8'hb8)}));
                    end
                  else
                    begin
                      reg7587 <= reg632;
                    end
                end
              else
                begin
                  if (($signed(forvar644) > (reg7436[(2'h2):(1'h1)] ?
                      forvar7437[(3'h4):(2'h2)] : $signed((forvar637 + reg7581)))))
                    begin
                      reg7585 <= forvar7456[(1'h0):(1'h0)];
                      reg7586 <= $signed(((+$signed(forvar7440)) ^ $signed({reg664})));
                      reg7587 <= (forvar7445[(1'h1):(1'h1)] | {((~^reg7493) ?
                              $unsigned(reg657) : wire7432[(4'he):(3'h7)])});
                      reg7588 <= ((!$unsigned(reg7554[(4'h8):(2'h3)])) - $signed(({forvar7457} * wire624[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg7585 <= (reg7493[(2'h2):(1'h1)] >> (wire7433[(1'h0):(1'h0)] * reg632[(3'h5):(3'h4)]));
                    end
                end
            end
          else
            begin
              for (forvar7574 = (1'h0); (forvar7574 < (2'h2)); forvar7574 = (forvar7574 + (1'h1)))
                begin
                  if ($unsigned((reg7459 ?
                      ((reg7492 + (8'h9d)) ?
                          reg667[(2'h3):(1'h0)] : $unsigned(reg7521)) : $signed((reg664 * reg7537)))))
                    begin
                      reg7575 <= $signed(($signed((-reg7449)) ^ {reg7562[(3'h6):(3'h5)]}));
                      reg7576 <= ((^~$unsigned((forvar7574 - (8'hb0)))) ?
                          reg640 : ((~^(!reg674)) ?
                              forvar671 : ((~&(8'ha2)) ?
                                  (+reg660) : $signed(forvar632))));
                      reg7577 <= ((((reg668 == reg632) > reg644[(4'h8):(3'h6)]) >>> $unsigned((+forvar7488))) ?
                          ({reg7496} ?
                              $unsigned((|(8'hac))) : (((8'had) * forvar7508) ?
                                  $unsigned(reg635) : (reg637 > forvar7441))) : ($unsigned((~^reg7498)) ?
                              $unsigned({reg7474}) : ($signed(reg7526) ?
                                  $signed((8'hb7)) : $unsigned(reg670))));
                    end
                  else
                    begin
                      reg7575 <= (((forvar7478 ?
                                  {reg7575} : forvar7488[(4'h9):(2'h3)]) ?
                              {((8'haa) > reg7545)} : forvar7475[(4'hb):(4'h8)]) ?
                          ($signed((reg7564 ? reg7440 : reg674)) ?
                              reg7587 : $signed((reg7529 ?
                                  forvar7531 : (8'h9c)))) : ((~^reg7568[(2'h3):(2'h3)]) < (reg7517 ?
                              {forvar7488} : $signed(forvar7477))));
                      reg7576 <= {(^~$signed($unsigned(reg7496)))};
                      reg7577 <= $unsigned((8'haa));
                      reg7578 <= wire628[(1'h1):(1'h0)];
                    end
                  if (($unsigned($unsigned({reg7540})) ~^ $signed(($unsigned(reg7527) != $unsigned(reg634)))))
                    begin
                      reg7579 <= reg657[(2'h3):(1'h1)];
                      reg7580 <= ((^~((~^reg7566) ?
                              forvar639[(2'h2):(1'h0)] : reg7461[(1'h0):(1'h0)])) ?
                          reg7575[(1'h1):(1'h0)] : reg649[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg7579 <= (reg7499 ?
                          reg7560 : forvar7470[(3'h4):(2'h3)]);
                      reg7580 <= forvar7576[(3'h5):(2'h2)];
                      reg7581 <= $signed($signed(($signed(wire628) ?
                          (reg7498 ? reg7460 : reg7499) : $unsigned(reg7464))));
                    end
                end
              for (forvar7582 = (1'h0); (forvar7582 < (2'h2)); forvar7582 = (forvar7582 + (1'h1)))
                begin
                  if ($unsigned($signed((~(8'hae)))))
                    begin
                      reg7583 <= reg7587;
                      reg7584 <= ((|$signed($signed(reg7545))) >> reg7550);
                      reg7585 <= reg668[(3'h4):(3'h4)];
                      reg7586 <= $signed($unsigned((reg652 < reg7450)));
                    end
                  else
                    begin
                      reg7583 <= reg7444;
                      reg7584 <= (~&({$signed((8'hb6))} <<< reg7584[(3'h6):(3'h5)]));
                      reg7585 <= {$signed(wire628[(1'h0):(1'h0)])};
                    end
                  for (forvar7587 = (1'h0); (forvar7587 < (1'h1)); forvar7587 = (forvar7587 + (1'h1)))
                    begin
                      reg7588 <= (8'h9c);
                      reg7589 <= $unsigned($signed($signed({forvar7438})));
                      reg7590 <= (&forvar7576);
                      reg7591 <= $signed({(((8'hab) ?
                              forvar7543 : reg7571) ^~ (forvar659 ?
                              forvar7440 : wire7430))});
                    end
                  reg7592 <= forvar7587;
                  if ($signed($unsigned(($unsigned(reg7548) ?
                      reg7547[(4'ha):(1'h0)] : (^reg7471)))))
                    begin
                      reg7593 <= $signed(reg7525);
                      reg7594 <= $unsigned($signed((-forvar7440)));
                      reg7595 <= $unsigned($unsigned((8'hac)));
                    end
                  else
                    begin
                      reg7593 <= $unsigned(reg7578);
                    end
                end
            end
          for (forvar7596 = (1'h0); (forvar7596 < (1'h0)); forvar7596 = (forvar7596 + (1'h1)))
            begin
              reg7597 <= $unsigned(((reg7455[(2'h2):(1'h0)] ~^ wire624) & $signed((+forvar7557))));
            end
        end
      for (forvar7598 = (1'h0); (forvar7598 < (2'h2)); forvar7598 = (forvar7598 + (1'h1)))
        begin
          for (forvar7599 = (1'h0); (forvar7599 < (2'h3)); forvar7599 = (forvar7599 + (1'h1)))
            begin
              for (forvar7600 = (1'h0); (forvar7600 < (1'h0)); forvar7600 = (forvar7600 + (1'h1)))
                begin
                  for (forvar7601 = (1'h0); (forvar7601 < (1'h0)); forvar7601 = (forvar7601 + (1'h1)))
                    begin
                      reg7602 <= forvar7599[(4'ha):(2'h2)];
                      reg7603 <= ($unsigned(reg632[(3'h4):(3'h4)]) + (($signed(reg7572) ?
                              (reg7540 ?
                                  reg7525 : reg7494) : $signed(wire622)) ?
                          reg7480 : ((+wire7429) ?
                              reg647 : (reg7554 || reg656))));
                      reg7604 <= (~&({(-forvar7546)} != ((^~(8'ha6)) ^~ (reg7456 + forvar7577))));
                    end
                  for (forvar7605 = (1'h0); (forvar7605 < (2'h3)); forvar7605 = (forvar7605 + (1'h1)))
                    begin
                      reg7606 <= ((wire624[(3'h6):(2'h3)] > (+reg7524[(3'h6):(2'h2)])) ?
                          $unsigned($unsigned($unsigned(reg653))) : (8'hb8));
                      reg7607 <= (^$signed(forvar635));
                      reg7608 <= ((($signed((8'hb4)) * forvar654) * $unsigned((forvar7438 > (8'ha9)))) ?
                          ($signed(reg7515[(3'h6):(2'h2)]) != $signed($signed((8'hac)))) : (reg7544[(3'h4):(2'h2)] + ((reg7512 ?
                                  forvar7546 : reg7448) ?
                              forvar7461[(3'h7):(2'h2)] : $signed(reg642))));
                    end
                  for (forvar7609 = (1'h0); (forvar7609 < (1'h0)); forvar7609 = (forvar7609 + (1'h1)))
                    begin
                      reg7610 <= $unsigned((-$unsigned(((8'ha3) ?
                          forvar7543 : (8'ha2)))));
                      reg7611 <= $signed((!(8'ha0)));
                      reg7612 <= reg7472[(3'h5):(1'h0)];
                    end
                  if ((reg7509[(2'h3):(1'h0)] ?
                      $unsigned((reg7503[(2'h2):(2'h2)] ?
                          (~^forvar7488) : (&reg7608))) : ($unsigned((forvar7479 > wire625)) < (8'hb5))))
                    begin
                      reg7613 <= reg7505[(3'h5):(3'h5)];
                      reg7614 <= (~forvar7576);
                      reg7615 <= (-(~&{$signed((8'h9e))}));
                    end
                  else
                    begin
                      reg7613 <= (reg7445 | ($signed(((8'ha1) ?
                          reg7503 : forvar7600)) <= $signed(forvar659)));
                      reg7614 <= (^forvar7600[(2'h3):(1'h1)]);
                      reg7615 <= reg7590[(2'h3):(2'h2)];
                      reg7616 <= (+(-($signed(forvar636) || $signed(reg7584))));
                    end
                end
              if ((^reg648))
                begin
                  for (forvar7617 = (1'h0); (forvar7617 < (2'h3)); forvar7617 = (forvar7617 + (1'h1)))
                    begin
                      reg7618 <= (&(((~|reg7584) ?
                          (^reg7444) : {reg673}) + $signed($unsigned(reg7503))));
                    end
                  for (forvar7619 = (1'h0); (forvar7619 < (1'h0)); forvar7619 = (forvar7619 + (1'h1)))
                    begin
                      reg7620 <= (reg7581[(2'h3):(2'h3)] ?
                          ((reg636[(4'hd):(3'h5)] == reg7580) ?
                              (|(~(8'ha7))) : reg7483[(1'h0):(1'h0)]) : wire629[(3'h4):(2'h2)]);
                      reg7621 <= forvar7466;
                      reg7622 <= reg7456[(3'h6):(3'h4)];
                    end
                end
              else
                begin
                  for (forvar7617 = (1'h0); (forvar7617 < (1'h0)); forvar7617 = (forvar7617 + (1'h1)))
                    begin
                      reg7618 <= reg7610[(1'h1):(1'h0)];
                      reg7619 <= reg7602;
                      reg7620 <= {reg7529[(4'h8):(4'h8)]};
                    end
                end
            end
          reg7623 <= $unsigned({reg7616[(4'ha):(3'h6)]});
        end
    end
  assign wire7624 = ($unsigned(reg7481[(3'h5):(2'h3)]) ?
                        $signed($signed(((8'ha9) || reg7542))) : reg7500);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module6
#( parameter param617 = ({(((8'hb4) ? (8'h9d) : (8'haf)) ? (!(8'ha5)) : ((8'hb2) > (8'hb6)))} & {(((8'ha9) >>> (8'ha9)) == (~(8'hb9)))}) )
(y, clk, wire7, wire8, wire9, wire10);
  output wire [(32'haa1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire7;
  input wire [(4'ha):(1'h0)] wire8;
  input wire [(4'hd):(1'h0)] wire9;
  input wire [(4'ha):(1'h0)] wire10;
  wire signed [(2'h2):(1'h0)] wire616;
  reg signed [(3'h6):(1'h0)] reg615 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg614 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg613 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar612 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg611 = (1'h0);
  reg [(3'h4):(1'h0)] reg610 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar609 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar608 = (1'h0);
  reg [(2'h2):(1'h0)] forvar607 = (1'h0);
  reg [(4'h9):(1'h0)] forvar606 = (1'h0);
  reg [(2'h2):(1'h0)] reg605 = (1'h0);
  reg signed [(4'he):(1'h0)] reg604 = (1'h0);
  reg [(4'h8):(1'h0)] reg603 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg602 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg601 = (1'h0);
  reg [(2'h3):(1'h0)] reg600 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar599 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg598 = (1'h0);
  reg [(2'h2):(1'h0)] reg597 = (1'h0);
  reg [(3'h4):(1'h0)] forvar596 = (1'h0);
  reg [(5'h10):(1'h0)] reg595 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg594 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg593 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg592 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar591 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar590 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar589 = (1'h0);
  reg [(2'h3):(1'h0)] reg588 = (1'h0);
  reg [(3'h5):(1'h0)] forvar587 = (1'h0);
  reg [(4'hc):(1'h0)] reg586 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg585 = (1'h0);
  reg [(4'hd):(1'h0)] reg584 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar583 = (1'h0);
  reg [(4'hf):(1'h0)] forvar582 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg581 = (1'h0);
  reg [(4'ha):(1'h0)] reg580 = (1'h0);
  reg [(3'h7):(1'h0)] reg579 = (1'h0);
  reg [(4'h9):(1'h0)] reg578 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar576 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg577 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg576 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg575 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar574 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg571 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg573 = (1'h0);
  reg [(3'h5):(1'h0)] reg572 = (1'h0);
  reg [(3'h7):(1'h0)] forvar571 = (1'h0);
  reg [(3'h7):(1'h0)] reg570 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg569 = (1'h0);
  reg [(4'hb):(1'h0)] reg568 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg567 = (1'h0);
  reg [(3'h7):(1'h0)] reg566 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg565 = (1'h0);
  reg [(4'hf):(1'h0)] forvar564 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar563 = (1'h0);
  reg [(5'h10):(1'h0)] reg560 = (1'h0);
  reg [(3'h5):(1'h0)] forvar557 = (1'h0);
  reg [(4'hc):(1'h0)] reg555 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg562 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg561 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar560 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg559 = (1'h0);
  reg [(4'hb):(1'h0)] reg558 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg557 = (1'h0);
  reg [(4'h9):(1'h0)] reg556 = (1'h0);
  reg [(3'h6):(1'h0)] forvar555 = (1'h0);
  reg signed [(4'he):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg553 = (1'h0);
  reg [(3'h7):(1'h0)] reg552 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg551 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar550 = (1'h0);
  reg [(4'ha):(1'h0)] reg549 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg548 = (1'h0);
  reg [(4'hb):(1'h0)] reg547 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar545 = (1'h0);
  reg [(4'hd):(1'h0)] forvar543 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg541 = (1'h0);
  reg [(4'hf):(1'h0)] forvar540 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg546 = (1'h0);
  reg [(3'h7):(1'h0)] reg545 = (1'h0);
  reg [(4'hd):(1'h0)] reg544 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg543 = (1'h0);
  reg [(4'ha):(1'h0)] reg542 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar541 = (1'h0);
  reg [(2'h2):(1'h0)] reg540 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg539 = (1'h0);
  reg [(3'h5):(1'h0)] reg538 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg537 = (1'h0);
  reg [(4'ha):(1'h0)] forvar536 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg535 = (1'h0);
  reg [(4'hd):(1'h0)] reg534 = (1'h0);
  reg [(3'h7):(1'h0)] reg533 = (1'h0);
  reg [(4'hf):(1'h0)] reg532 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar531 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar526 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg524 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar521 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg531 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg529 = (1'h0);
  reg [(4'hc):(1'h0)] reg528 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg527 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg526 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg525 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar524 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg523 = (1'h0);
  reg [(2'h3):(1'h0)] reg522 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg521 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg520 = (1'h0);
  reg [(3'h7):(1'h0)] reg519 = (1'h0);
  reg [(4'hb):(1'h0)] forvar516 = (1'h0);
  reg [(4'hc):(1'h0)] forvar510 = (1'h0);
  reg signed [(4'he):(1'h0)] reg518 = (1'h0);
  reg [(4'he):(1'h0)] reg517 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg516 = (1'h0);
  reg [(2'h2):(1'h0)] reg515 = (1'h0);
  reg [(4'hd):(1'h0)] reg514 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg513 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg511 = (1'h0);
  reg [(4'hc):(1'h0)] reg510 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar509 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar508 = (1'h0);
  wire [(3'h4):(1'h0)] wire506;
  wire [(4'hb):(1'h0)] wire337;
  reg [(4'hf):(1'h0)] reg336 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg335 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg334 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar333 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg332 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg331 = (1'h0);
  reg [(4'he):(1'h0)] reg330 = (1'h0);
  reg signed [(4'he):(1'h0)] reg329 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg328 = (1'h0);
  reg [(3'h4):(1'h0)] reg327 = (1'h0);
  reg [(4'h9):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg325 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar323 = (1'h0);
  reg [(4'hd):(1'h0)] forvar322 = (1'h0);
  reg [(3'h6):(1'h0)] reg321 = (1'h0);
  reg [(4'hc):(1'h0)] reg320 = (1'h0);
  reg [(4'ha):(1'h0)] reg319 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar318 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar317 = (1'h0);
  reg [(2'h3):(1'h0)] forvar316 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar311 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg310 = (1'h0);
  reg [(4'hd):(1'h0)] reg308 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar306 = (1'h0);
  reg [(4'he):(1'h0)] forvar304 = (1'h0);
  reg [(4'h9):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg315 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg314 = (1'h0);
  reg [(4'hb):(1'h0)] reg313 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar310 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg309 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar308 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar307 = (1'h0);
  reg [(3'h7):(1'h0)] reg302 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar299 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg297 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg306 = (1'h0);
  reg [(4'hb):(1'h0)] reg305 = (1'h0);
  reg [(2'h2):(1'h0)] reg304 = (1'h0);
  reg signed [(4'he):(1'h0)] reg303 = (1'h0);
  reg [(2'h2):(1'h0)] forvar302 = (1'h0);
  reg [(3'h7):(1'h0)] reg301 = (1'h0);
  reg signed [(4'he):(1'h0)] reg300 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg299 = (1'h0);
  reg [(2'h2):(1'h0)] reg298 = (1'h0);
  reg [(4'hd):(1'h0)] forvar297 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg296 = (1'h0);
  reg [(3'h5):(1'h0)] reg295 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar293 = (1'h0);
  reg [(3'h7):(1'h0)] forvar292 = (1'h0);
  reg [(4'ha):(1'h0)] reg291 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire290;
  reg signed [(4'he):(1'h0)] reg289 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar287 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg284 = (1'h0);
  reg [(3'h5):(1'h0)] reg288 = (1'h0);
  reg [(4'hd):(1'h0)] reg287 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg286 = (1'h0);
  reg [(4'hd):(1'h0)] reg285 = (1'h0);
  reg [(2'h2):(1'h0)] forvar284 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg283 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg281 = (1'h0);
  reg [(4'hd):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar279 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg277 = (1'h0);
  reg signed [(4'he):(1'h0)] reg276 = (1'h0);
  reg [(4'hd):(1'h0)] reg275 = (1'h0);
  reg [(3'h6):(1'h0)] reg274 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg273 = (1'h0);
  reg [(3'h4):(1'h0)] reg272 = (1'h0);
  reg [(5'h10):(1'h0)] reg271 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar270 = (1'h0);
  reg [(4'ha):(1'h0)] reg269 = (1'h0);
  reg [(4'hd):(1'h0)] forvar268 = (1'h0);
  reg [(5'h10):(1'h0)] forvar267 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg264 = (1'h0);
  reg [(4'h8):(1'h0)] forvar263 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar259 = (1'h0);
  reg [(2'h2):(1'h0)] reg258 = (1'h0);
  reg [(2'h3):(1'h0)] forvar254 = (1'h0);
  reg [(4'hf):(1'h0)] reg263 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg262 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar261 = (1'h0);
  reg [(4'h9):(1'h0)] reg260 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg259 = (1'h0);
  reg [(5'h10):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg257 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg256 = (1'h0);
  reg signed [(4'he):(1'h0)] reg255 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg254 = (1'h0);
  reg [(4'he):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar252 = (1'h0);
  reg [(4'h9):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg249 = (1'h0);
  reg [(4'he):(1'h0)] reg248 = (1'h0);
  reg [(4'ha):(1'h0)] forvar247 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar246 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar245 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar239 = (1'h0);
  reg [(4'hd):(1'h0)] forvar232 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar234 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg233 = (1'h0);
  reg [(4'he):(1'h0)] reg244 = (1'h0);
  reg [(3'h7):(1'h0)] reg243 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg241 = (1'h0);
  reg [(3'h7):(1'h0)] reg240 = (1'h0);
  reg [(4'h8):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg238 = (1'h0);
  reg [(2'h2):(1'h0)] reg237 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg236 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg234 = (1'h0);
  reg [(4'hb):(1'h0)] forvar233 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg232 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg210 = (1'h0);
  reg [(3'h4):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg230 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar229 = (1'h0);
  reg [(4'ha):(1'h0)] reg228 = (1'h0);
  reg [(4'hc):(1'h0)] reg227 = (1'h0);
  reg [(4'hc):(1'h0)] reg226 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg225 = (1'h0);
  reg [(4'hd):(1'h0)] forvar224 = (1'h0);
  reg [(3'h5):(1'h0)] forvar223 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg221 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg220 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg219 = (1'h0);
  reg [(4'h9):(1'h0)] forvar218 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg217 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar216 = (1'h0);
  reg [(5'h10):(1'h0)] reg215 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg214 = (1'h0);
  reg [(5'h10):(1'h0)] forvar213 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg212 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar211 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar210 = (1'h0);
  reg [(5'h10):(1'h0)] forvar209 = (1'h0);
  reg [(4'hd):(1'h0)] reg208 = (1'h0);
  wire [(3'h4):(1'h0)] wire11;
  wire signed [(4'hd):(1'h0)] wire12;
  wire signed [(4'he):(1'h0)] wire13;
  wire signed [(4'hc):(1'h0)] wire14;
  wire signed [(5'h10):(1'h0)] wire15;
  wire [(4'ha):(1'h0)] wire16;
  wire signed [(4'hc):(1'h0)] wire17;
  wire signed [(4'ha):(1'h0)] wire18;
  wire [(3'h5):(1'h0)] wire206;
  assign y = {wire616,
                 reg615,
                 reg614,
                 reg613,
                 forvar612,
                 reg611,
                 reg610,
                 forvar609,
                 forvar608,
                 forvar607,
                 forvar606,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 forvar599,
                 reg598,
                 reg597,
                 forvar596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 forvar591,
                 forvar590,
                 forvar589,
                 reg588,
                 forvar587,
                 reg586,
                 reg585,
                 reg584,
                 forvar583,
                 forvar582,
                 reg581,
                 reg580,
                 reg579,
                 reg578,
                 forvar576,
                 reg577,
                 reg576,
                 reg575,
                 forvar574,
                 reg571,
                 reg573,
                 reg572,
                 forvar571,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 forvar564,
                 forvar563,
                 reg560,
                 forvar557,
                 reg555,
                 reg562,
                 reg561,
                 forvar560,
                 reg559,
                 reg558,
                 reg557,
                 reg556,
                 forvar555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 forvar550,
                 reg549,
                 reg548,
                 reg547,
                 forvar545,
                 forvar543,
                 reg541,
                 forvar540,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 forvar541,
                 reg540,
                 reg539,
                 reg538,
                 reg537,
                 forvar536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 forvar531,
                 forvar526,
                 reg524,
                 forvar521,
                 reg531,
                 reg530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 forvar524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 forvar516,
                 forvar510,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 forvar509,
                 forvar508,
                 wire506,
                 wire337,
                 reg336,
                 reg335,
                 reg334,
                 forvar333,
                 reg332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 forvar323,
                 forvar322,
                 reg321,
                 reg320,
                 reg319,
                 forvar318,
                 forvar317,
                 forvar316,
                 forvar311,
                 reg310,
                 reg308,
                 reg307,
                 forvar306,
                 forvar304,
                 reg293,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 reg309,
                 forvar308,
                 forvar307,
                 reg302,
                 forvar299,
                 reg297,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 forvar302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 forvar297,
                 reg296,
                 reg295,
                 reg294,
                 forvar293,
                 forvar292,
                 reg291,
                 wire290,
                 reg289,
                 forvar287,
                 reg284,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 forvar284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 forvar279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 forvar270,
                 reg269,
                 forvar268,
                 forvar267,
                 reg266,
                 reg265,
                 reg264,
                 forvar263,
                 reg261,
                 forvar259,
                 reg258,
                 forvar254,
                 reg263,
                 reg262,
                 forvar261,
                 reg260,
                 reg259,
                 forvar258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 forvar252,
                 reg251,
                 reg250,
                 reg249,
                 reg248,
                 forvar247,
                 forvar246,
                 forvar245,
                 forvar239,
                 forvar232,
                 forvar234,
                 reg233,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 forvar233,
                 reg232,
                 reg210,
                 reg231,
                 reg230,
                 forvar229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 forvar224,
                 forvar223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 forvar218,
                 reg217,
                 forvar216,
                 reg215,
                 reg214,
                 forvar213,
                 reg212,
                 forvar211,
                 forvar210,
                 forvar209,
                 reg208,
                 wire11,
                 wire12,
                 wire13,
                 wire14,
                 wire15,
                 wire16,
                 wire17,
                 wire18,
                 wire206,
                 (1'h0)};
  assign wire11 = (~&$unsigned((((8'ha6) ? wire7 : (8'hb6)) ?
                      $signed(wire10) : (wire7 <<< (8'h9e)))));
  assign wire12 = (+$unsigned(wire10[(3'h6):(3'h5)]));
  assign wire13 = $unsigned($signed(((wire10 <= wire11) != (wire9 ~^ wire12))));
  assign wire14 = (~|$unsigned($signed({wire9})));
  assign wire15 = (+{(wire11 && (wire9 ? wire11 : (8'hb7)))});
  assign wire16 = ($signed((^$signed(wire11))) ?
                      wire13[(3'h4):(2'h3)] : (+{(wire10 ? (8'hb5) : wire9)}));
  assign wire17 = (~|wire8);
  assign wire18 = $signed(wire8[(4'ha):(3'h7)]);
  module19 modinst207 (wire206, clk, wire17, wire16, wire9, wire14, wire15);
  always
    @(posedge clk) begin
      reg208 <= wire17[(2'h3):(1'h0)];
      for (forvar209 = (1'h0); (forvar209 < (2'h2)); forvar209 = (forvar209 + (1'h1)))
        begin
          if (wire18[(1'h1):(1'h0)])
            begin
              for (forvar210 = (1'h0); (forvar210 < (2'h2)); forvar210 = (forvar210 + (1'h1)))
                begin
                  for (forvar211 = (1'h0); (forvar211 < (2'h3)); forvar211 = (forvar211 + (1'h1)))
                    begin
                      reg212 <= {wire11};
                    end
                  for (forvar213 = (1'h0); (forvar213 < (2'h3)); forvar213 = (forvar213 + (1'h1)))
                    begin
                      reg214 <= (~^(((wire18 ? wire12 : wire10) == wire15) ?
                          $unsigned((forvar211 && wire12)) : wire17[(4'h9):(4'h9)]));
                      reg215 <= ($unsigned(wire206[(1'h1):(1'h1)]) ?
                          wire17 : wire8);
                    end
                  for (forvar216 = (1'h0); (forvar216 < (1'h1)); forvar216 = (forvar216 + (1'h1)))
                    begin
                      reg217 <= (((|((8'haf) ?
                              wire12 : forvar210)) < (~&$unsigned(wire13))) ?
                          ((8'hb3) & (8'hb4)) : $signed(($signed((8'ha3)) == (8'ha0))));
                    end
                  for (forvar218 = (1'h0); (forvar218 < (2'h3)); forvar218 = (forvar218 + (1'h1)))
                    begin
                      reg219 <= ((&($unsigned(wire15) ?
                              ((8'hb3) ?
                                  forvar209 : wire9) : $signed(wire11))) ?
                          (~&(~|$unsigned((8'hb5)))) : (+(forvar211 ?
                              forvar218[(3'h4):(2'h2)] : wire12)));
                      reg220 <= $signed(wire9[(1'h1):(1'h1)]);
                      reg221 <= {$unsigned(forvar218)};
                    end
                end
              reg222 <= {wire17};
              for (forvar223 = (1'h0); (forvar223 < (2'h3)); forvar223 = (forvar223 + (1'h1)))
                begin
                  for (forvar224 = (1'h0); (forvar224 < (1'h1)); forvar224 = (forvar224 + (1'h1)))
                    begin
                      reg225 <= wire10;
                      reg226 <= $unsigned((wire14 ?
                          $signed(reg220[(2'h3):(1'h0)]) : forvar209[(4'hf):(3'h7)]));
                      reg227 <= $signed(reg215);
                      reg228 <= ({$unsigned($unsigned(wire9))} ?
                          $signed(((forvar223 && forvar211) || (!wire17))) : (+$unsigned($unsigned(forvar216))));
                    end
                end
              for (forvar229 = (1'h0); (forvar229 < (1'h0)); forvar229 = (forvar229 + (1'h1)))
                begin
                  reg230 <= (8'hb8);
                  reg231 <= $unsigned((forvar211 < $unsigned($signed(reg208))));
                end
            end
          else
            begin
              reg210 <= ($unsigned(($signed((8'h9c)) ?
                  {(8'hb9)} : forvar213)) | (((wire14 ? forvar229 : (8'ha5)) ?
                      (reg225 & reg215) : (reg221 ? wire7 : (8'ha7))) ?
                  wire9[(2'h3):(1'h0)] : $signed(wire13[(1'h1):(1'h0)])));
            end
          if ({(^reg208)})
            begin
              reg232 <= wire18[(1'h1):(1'h1)];
              if ($unsigned(forvar213))
                begin
                  for (forvar233 = (1'h0); (forvar233 < (2'h3)); forvar233 = (forvar233 + (1'h1)))
                    begin
                      reg234 <= {(wire17[(1'h0):(1'h0)] ?
                              $unsigned(reg231) : wire17)};
                      reg235 <= forvar229;
                      reg236 <= ($signed((|wire9)) | ($signed((8'hb1)) ?
                          $unsigned(wire206) : (wire18 != $signed(forvar229))));
                    end
                  if ((&($unsigned(reg222[(1'h0):(1'h0)]) ?
                      reg221 : (^(reg226 ? reg231 : forvar223)))))
                    begin
                      reg237 <= {reg226};
                    end
                  else
                    begin
                      reg237 <= $unsigned(((^reg219[(2'h2):(1'h1)]) ?
                          (((8'hba) ? wire17 : forvar218) ?
                              {forvar229} : (8'ha1)) : $unsigned({reg226})));
                      reg238 <= forvar210;
                      reg239 <= ($signed(((reg219 ?
                          wire11 : reg219) == (8'h9c))) && $signed(($unsigned(reg234) >= (^~reg235))));
                      reg240 <= reg208;
                    end
                  if ($signed(((!{(8'hab)}) ?
                      $signed($signed(reg217)) : $unsigned((reg234 | reg221)))))
                    begin
                      reg241 <= forvar213[(4'h8):(2'h2)];
                    end
                  else
                    begin
                      reg241 <= ($signed(wire15) ? wire18 : (8'ha0));
                      reg242 <= reg241;
                      reg243 <= ({wire8} >>> {$signed($unsigned((8'hb6)))});
                      reg244 <= (reg220 <= $signed(reg230));
                    end
                end
              else
                begin
                  reg233 <= ($unsigned((&$unsigned(reg228))) ?
                      forvar224[(2'h2):(1'h0)] : $signed((~^$unsigned(reg243))));
                  for (forvar234 = (1'h0); (forvar234 < (2'h2)); forvar234 = (forvar234 + (1'h1)))
                    begin
                      reg235 <= $unsigned((+((wire8 << reg212) ?
                          $unsigned(wire7) : (8'haf))));
                      reg236 <= wire15;
                      reg237 <= ($unsigned($signed($signed(wire18))) > $signed(((+(8'h9f)) ?
                          $signed(reg220) : reg233[(4'hc):(2'h3)])));
                    end
                end
            end
          else
            begin
              for (forvar232 = (1'h0); (forvar232 < (1'h0)); forvar232 = (forvar232 + (1'h1)))
                begin
                  if ((forvar223[(3'h5):(2'h3)] ?
                      forvar213[(1'h1):(1'h0)] : forvar224))
                    begin
                      reg233 <= reg210[(3'h4):(3'h4)];
                      reg234 <= (((8'h9c) ?
                          reg238[(2'h3):(1'h1)] : $unsigned((^wire14))) * {((forvar234 != forvar209) ?
                              (8'hb3) : reg239)});
                    end
                  else
                    begin
                      reg233 <= ($unsigned(reg234[(2'h3):(2'h2)]) ?
                          (+$unsigned((wire206 ?
                              reg244 : reg243))) : reg226[(4'hc):(3'h6)]);
                      reg234 <= (^$unsigned(({wire9} ?
                          $unsigned(reg244) : (reg234 ? reg232 : reg214))));
                      reg235 <= $signed({(reg214[(3'h6):(3'h5)] ?
                              (reg232 ?
                                  wire17 : reg228) : (wire15 != wire17))});
                    end
                  if ($signed($unsigned(((reg217 * forvar229) ?
                      (^reg243) : $unsigned((8'ha1))))))
                    begin
                      reg236 <= $unsigned((|(&((8'ha7) ? wire15 : (8'ha4)))));
                      reg237 <= (^$signed($signed((^reg221))));
                      reg238 <= $signed($signed(forvar211[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg236 <= $unsigned((~|((reg242 ?
                          reg238 : forvar213) && (wire17 ? reg212 : wire12))));
                      reg237 <= $unsigned($signed($signed($unsigned(forvar209))));
                      reg238 <= {$unsigned(wire10[(2'h3):(2'h2)])};
                    end
                  for (forvar239 = (1'h0); (forvar239 < (2'h2)); forvar239 = (forvar239 + (1'h1)))
                    begin
                      reg240 <= forvar233;
                      reg241 <= ((forvar229 ?
                          (wire11[(3'h4):(1'h1)] <<< (-wire18)) : ($signed((8'h9d)) > reg230)) & ($signed(forvar223) == (8'hb9)));
                      reg242 <= (reg225 ?
                          $unsigned((|((8'h9d) <<< reg233))) : ($unsigned(forvar229) ?
                              (~^{wire18}) : wire206));
                    end
                end
            end
          for (forvar245 = (1'h0); (forvar245 < (2'h2)); forvar245 = (forvar245 + (1'h1)))
            begin
              for (forvar246 = (1'h0); (forvar246 < (2'h3)); forvar246 = (forvar246 + (1'h1)))
                begin
                  for (forvar247 = (1'h0); (forvar247 < (2'h3)); forvar247 = (forvar247 + (1'h1)))
                    begin
                      reg248 <= (+$unsigned(forvar210));
                      reg249 <= {((~^(8'ha4)) == (~&(reg214 > (8'hba))))};
                      reg250 <= $unsigned(($signed($signed(reg215)) ~^ {$signed(reg243)}));
                      reg251 <= $signed(({(+(8'hb6))} ?
                          (~&reg228[(1'h1):(1'h1)]) : wire10[(3'h7):(3'h5)]));
                    end
                  for (forvar252 = (1'h0); (forvar252 < (2'h3)); forvar252 = (forvar252 + (1'h1)))
                    begin
                      reg253 <= forvar229[(3'h5):(1'h1)];
                    end
                end
              if ((~forvar247))
                begin
                  if (reg240[(2'h3):(1'h0)])
                    begin
                      reg254 <= reg212;
                      reg255 <= (reg249[(2'h3):(1'h0)] ?
                          wire16[(1'h0):(1'h0)] : (wire17[(4'ha):(4'h9)] ?
                              ({(8'hb8)} ?
                                  {reg240} : $signed(forvar218)) : {$unsigned(reg231)}));
                    end
                  else
                    begin
                      reg254 <= $signed($unsigned({$unsigned(wire9)}));
                      reg255 <= ({{{(8'ha6)}}} & forvar223[(2'h3):(1'h0)]);
                      reg256 <= ((reg254[(3'h6):(3'h5)] ~^ ((+reg214) ?
                              (8'hb3) : reg238[(3'h5):(1'h1)])) ?
                          (&$unsigned(forvar233[(4'h8):(1'h1)])) : forvar232);
                    end
                  reg257 <= {$unsigned(reg233)};
                  for (forvar258 = (1'h0); (forvar258 < (2'h3)); forvar258 = (forvar258 + (1'h1)))
                    begin
                      reg259 <= (+(((~^forvar232) >> reg241[(3'h4):(1'h1)]) >= (&reg228[(3'h6):(2'h2)])));
                      reg260 <= (!(reg232[(3'h6):(3'h4)] << ($signed(reg238) ?
                          ((8'h9e) ~^ (8'ha1)) : (|reg221))));
                    end
                  for (forvar261 = (1'h0); (forvar261 < (2'h3)); forvar261 = (forvar261 + (1'h1)))
                    begin
                      reg262 <= (8'ha0);
                      reg263 <= (!(-((reg242 ?
                          forvar223 : (8'hb6)) != $unsigned(forvar258))));
                    end
                end
              else
                begin
                  for (forvar254 = (1'h0); (forvar254 < (2'h2)); forvar254 = (forvar254 + (1'h1)))
                    begin
                      reg255 <= wire8;
                      reg256 <= $signed((reg260[(2'h3):(1'h0)] ?
                          ((reg237 + wire8) ?
                              (wire11 ?
                                  reg256 : reg262) : $signed(forvar246)) : (8'ha6)));
                      reg257 <= reg251[(1'h0):(1'h0)];
                    end
                  reg258 <= ((wire16 + $unsigned({reg220})) >= $signed($signed((~^wire206))));
                  for (forvar259 = (1'h0); (forvar259 < (1'h0)); forvar259 = (forvar259 + (1'h1)))
                    begin
                      reg260 <= (&forvar239[(1'h1):(1'h1)]);
                      reg261 <= $signed($unsigned($signed(((8'hb5) >>> reg256))));
                      reg262 <= (~&$unsigned($signed((reg258 ?
                          forvar252 : wire206))));
                    end
                  for (forvar263 = (1'h0); (forvar263 < (2'h2)); forvar263 = (forvar263 + (1'h1)))
                    begin
                      reg264 <= ((~&{reg227[(3'h4):(2'h3)]}) ^ $signed((|$unsigned(reg233))));
                      reg265 <= ((({forvar216} * (wire9 != reg258)) ^~ $unsigned($unsigned(reg254))) ?
                          reg226[(4'ha):(4'ha)] : (|$unsigned((~^reg214))));
                      reg266 <= $unsigned((&((-(8'h9d)) & $signed(wire206))));
                    end
                end
              for (forvar267 = (1'h0); (forvar267 < (2'h3)); forvar267 = (forvar267 + (1'h1)))
                begin
                  for (forvar268 = (1'h0); (forvar268 < (1'h0)); forvar268 = (forvar268 + (1'h1)))
                    begin
                      reg269 <= reg251[(3'h7):(3'h4)];
                    end
                  for (forvar270 = (1'h0); (forvar270 < (1'h0)); forvar270 = (forvar270 + (1'h1)))
                    begin
                      reg271 <= $unsigned(reg219);
                      reg272 <= wire8[(3'h7):(3'h4)];
                      reg273 <= reg265[(3'h4):(2'h2)];
                      reg274 <= wire8;
                    end
                  if ((($signed(forvar259[(5'h10):(4'h8)]) && (+reg264)) <<< reg254[(3'h4):(3'h4)]))
                    begin
                      reg275 <= $signed($unsigned(reg250[(4'hc):(3'h4)]));
                    end
                  else
                    begin
                      reg275 <= $unsigned(((((8'ha2) ? reg242 : reg222) ?
                          (forvar254 ?
                              reg248 : (8'ha6)) : $unsigned(forvar218)) - ((-reg249) | (^reg222))));
                      reg276 <= $signed($unsigned(($unsigned((8'ha6)) ?
                          $unsigned(reg208) : reg272)));
                    end
                  if (reg256)
                    begin
                      reg277 <= $signed(((reg215[(3'h4):(2'h2)] >>> {reg273}) ?
                          $unsigned($unsigned(forvar233)) : $signed(reg255[(4'hd):(4'hc)])));
                      reg278 <= (+wire7);
                    end
                  else
                    begin
                      reg277 <= forvar216[(3'h6):(1'h0)];
                    end
                end
            end
          for (forvar279 = (1'h0); (forvar279 < (1'h1)); forvar279 = (forvar279 + (1'h1)))
            begin
              if ({(reg232[(2'h3):(1'h0)] ?
                      (~|(reg249 >= (8'hab))) : $unsigned((forvar239 ?
                          forvar259 : forvar210)))})
                begin
                  if (forvar213)
                    begin
                      reg280 <= $signed((^~reg210));
                      reg281 <= ($signed(reg249[(2'h2):(1'h1)]) || reg278);
                      reg282 <= (!reg244[(4'hb):(3'h5)]);
                      reg283 <= ($signed(reg273) != (&(&$unsigned(reg273))));
                    end
                  else
                    begin
                      reg280 <= $signed(reg210[(1'h0):(1'h0)]);
                      reg281 <= forvar232;
                      reg282 <= ({$signed((wire16 ^~ (8'ha1)))} >>> reg259[(2'h2):(1'h1)]);
                      reg283 <= (wire9[(4'ha):(2'h3)] ? forvar229 : forvar261);
                    end
                  for (forvar284 = (1'h0); (forvar284 < (1'h0)); forvar284 = (forvar284 + (1'h1)))
                    begin
                      reg285 <= (^{reg258[(2'h2):(1'h1)]});
                      reg286 <= ($signed(($unsigned(reg248) >>> (forvar211 ?
                              wire12 : (8'ha9)))) ?
                          (!$signed((reg275 ?
                              reg237 : forvar224))) : (|wire8[(3'h6):(3'h5)]));
                      reg287 <= $signed($signed(reg253[(1'h1):(1'h1)]));
                      reg288 <= forvar213;
                    end
                end
              else
                begin
                  if ($signed(forvar259[(3'h4):(3'h4)]))
                    begin
                      reg280 <= reg210;
                      reg281 <= $unsigned($signed(reg272[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg280 <= {$unsigned((|(forvar268 ^ (8'ha1))))};
                    end
                  if ($signed($unsigned(((reg260 == (8'ha5)) ?
                      forvar211 : (forvar270 ? (8'ha4) : (8'hb1))))))
                    begin
                      reg282 <= forvar224[(3'h7):(3'h6)];
                      reg283 <= {forvar239};
                      reg284 <= reg251;
                    end
                  else
                    begin
                      reg282 <= ({$unsigned(((8'had) ? (8'hb6) : (8'h9d)))} ?
                          forvar263 : $unsigned($signed((~(8'h9c)))));
                    end
                  if ($unsigned(forvar213[(4'h9):(4'h9)]))
                    begin
                      reg285 <= $unsigned($signed({{(8'hac)}}));
                      reg286 <= (reg225 >= $signed(forvar229));
                    end
                  else
                    begin
                      reg285 <= (8'hb6);
                    end
                  for (forvar287 = (1'h0); (forvar287 < (1'h0)); forvar287 = (forvar287 + (1'h1)))
                    begin
                      reg288 <= $unsigned({$unsigned(((8'ha1) ?
                              (8'had) : forvar224))});
                    end
                end
              reg289 <= reg264[(2'h3):(1'h1)];
            end
        end
    end
  assign wire290 = wire14[(4'hc):(3'h4)];
  always
    @(posedge clk) begin
      reg291 <= (~&(($signed(forvar268) | (&wire16)) + {(8'had)}));
      if (($unsigned(reg232[(4'hb):(3'h4)]) + ($unsigned((reg265 ?
              wire9 : reg263)) ?
          forvar218[(4'h9):(3'h4)] : $unsigned($unsigned((8'hb4))))))
        begin
          for (forvar292 = (1'h0); (forvar292 < (1'h1)); forvar292 = (forvar292 + (1'h1)))
            begin
              if (reg239[(2'h2):(2'h2)])
                begin
                  for (forvar293 = (1'h0); (forvar293 < (1'h0)); forvar293 = (forvar293 + (1'h1)))
                    begin
                      reg294 <= forvar218[(3'h7):(3'h7)];
                      reg295 <= ({$unsigned(reg289[(1'h1):(1'h1)])} + (~|(&forvar252[(4'hf):(4'hc)])));
                      reg296 <= reg226[(2'h3):(2'h2)];
                    end
                  for (forvar297 = (1'h0); (forvar297 < (2'h3)); forvar297 = (forvar297 + (1'h1)))
                    begin
                      reg298 <= $unsigned($signed(({(8'hb5)} ?
                          (~|(8'h9c)) : (!forvar216))));
                      reg299 <= forvar216;
                      reg300 <= $unsigned((~&(8'hb1)));
                      reg301 <= (reg248 >>> forvar239[(3'h7):(3'h7)]);
                    end
                  for (forvar302 = (1'h0); (forvar302 < (1'h0)); forvar302 = (forvar302 + (1'h1)))
                    begin
                      reg303 <= ((((reg242 ?
                          reg227 : reg254) ^~ {reg212}) < $signed($signed(reg291))) || (forvar224[(3'h7):(1'h0)] << $signed(reg237[(1'h1):(1'h1)])));
                      reg304 <= reg227;
                      reg305 <= (-(reg261[(3'h6):(1'h1)] - $signed($signed(forvar224))));
                    end
                  reg306 <= reg277;
                end
              else
                begin
                  for (forvar293 = (1'h0); (forvar293 < (2'h2)); forvar293 = (forvar293 + (1'h1)))
                    begin
                      reg294 <= reg269[(4'h8):(2'h2)];
                      reg295 <= (({reg263[(4'h9):(1'h1)]} << ((forvar268 ?
                              reg232 : forvar287) ?
                          $unsigned(reg259) : forvar247[(2'h2):(2'h2)])) | ($unsigned(reg275[(3'h5):(3'h5)]) ?
                          forvar224[(4'hc):(2'h3)] : (+$signed(wire206))));
                    end
                  if ($signed($signed($signed(forvar246))))
                    begin
                      reg296 <= reg299;
                    end
                  else
                    begin
                      reg296 <= (-({$signed(forvar302)} ?
                          reg289 : ((^~forvar268) > {reg253})));
                      reg297 <= $signed((^~forvar267[(4'hb):(3'h6)]));
                      reg298 <= (({(8'ha9)} <= (8'hb4)) || $unsigned($signed(reg278[(3'h4):(1'h1)])));
                    end
                  for (forvar299 = (1'h0); (forvar299 < (1'h1)); forvar299 = (forvar299 + (1'h1)))
                    begin
                      reg300 <= ($unsigned(((&reg281) ?
                              $signed(reg212) : (!reg299))) ?
                          $signed(reg257[(4'ha):(2'h2)]) : forvar299[(3'h6):(2'h2)]);
                      reg301 <= forvar302[(1'h1):(1'h0)];
                    end
                  reg302 <= reg242;
                end
            end
          for (forvar307 = (1'h0); (forvar307 < (1'h1)); forvar307 = (forvar307 + (1'h1)))
            begin
              for (forvar308 = (1'h0); (forvar308 < (1'h1)); forvar308 = (forvar308 + (1'h1)))
                begin
                  reg309 <= reg251[(3'h7):(3'h6)];
                  for (forvar310 = (1'h0); (forvar310 < (1'h0)); forvar310 = (forvar310 + (1'h1)))
                    begin
                      reg311 <= ($unsigned((~(-reg255))) ?
                          (~(wire14 ?
                              (reg262 ~^ reg281) : ((8'ha6) ?
                                  reg239 : forvar263))) : reg297[(3'h4):(1'h0)]);
                      reg312 <= reg220;
                      reg313 <= ((^(+$signed(forvar234))) ?
                          (8'hb9) : (((8'hab) > (~reg242)) ?
                              reg269 : reg299[(1'h1):(1'h1)]));
                    end
                end
              reg314 <= reg236;
            end
          reg315 <= $unsigned((!((forvar299 == reg226) >= (~^reg222))));
        end
      else
        begin
          for (forvar292 = (1'h0); (forvar292 < (2'h3)); forvar292 = (forvar292 + (1'h1)))
            begin
              if ((($signed($unsigned((8'ha8))) ?
                      {forvar279} : ((^~reg305) ~^ ((8'hb1) != forvar252))) ?
                  $unsigned($signed($signed((8'hae)))) : $signed(reg288)))
                begin
                  if ($signed((~reg257[(3'h6):(3'h4)])))
                    begin
                      reg293 <= {forvar268};
                      reg294 <= $unsigned(($signed(reg299) ?
                          ((reg254 ? (8'h9e) : reg303) ?
                              $unsigned(reg227) : $unsigned(wire10)) : $signed((^~forvar223))));
                    end
                  else
                    begin
                      reg293 <= ((~|$unsigned({forvar211})) * $signed(((~reg222) ?
                          (8'ha9) : $unsigned(wire12))));
                      reg294 <= forvar234;
                      reg295 <= $unsigned(({(|reg231)} + ({reg271} != reg256[(1'h0):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar293 = (1'h0); (forvar293 < (1'h1)); forvar293 = (forvar293 + (1'h1)))
                    begin
                      reg294 <= forvar293;
                    end
                  reg295 <= ((+(((8'h9d) * reg239) ?
                      (~(8'hb2)) : reg285[(4'h8):(3'h7)])) | reg272[(1'h1):(1'h1)]);
                end
              reg296 <= $signed($unsigned(($unsigned(reg275) > forvar302[(1'h1):(1'h0)])));
            end
          if ((~^((+$unsigned(wire206)) + forvar258[(1'h0):(1'h0)])))
            begin
              for (forvar297 = (1'h0); (forvar297 < (2'h2)); forvar297 = (forvar297 + (1'h1)))
                begin
                  if ($signed((((|reg238) ?
                      (-(8'ha5)) : (~reg273)) >>> ((reg249 == reg255) ?
                      $unsigned(forvar308) : {(8'ha6)}))))
                    begin
                      reg298 <= forvar218;
                    end
                  else
                    begin
                      reg298 <= (((forvar245[(1'h0):(1'h0)] >>> reg251) <= $signed({reg289})) ^~ {forvar247});
                    end
                  if ({$unsigned({reg214[(3'h4):(1'h0)]})})
                    begin
                      reg299 <= {$signed((^reg249[(3'h4):(2'h2)]))};
                      reg300 <= $signed(reg234[(3'h6):(1'h0)]);
                      reg301 <= $unsigned($signed({(reg214 | (8'ha4))}));
                    end
                  else
                    begin
                      reg299 <= (forvar218 ^~ (&$unsigned({reg237})));
                      reg300 <= reg266[(1'h0):(1'h0)];
                    end
                end
              reg302 <= $unsigned((+(forvar302[(2'h2):(1'h1)] ?
                  reg250[(4'he):(3'h7)] : {reg305})));
            end
          else
            begin
              if ((reg315[(4'ha):(1'h0)] ? (|(8'hac)) : wire10))
                begin
                  for (forvar297 = (1'h0); (forvar297 < (2'h2)); forvar297 = (forvar297 + (1'h1)))
                    begin
                      reg298 <= ((((wire290 ? reg214 : forvar292) ?
                              (reg225 & forvar209) : ((8'hb9) ?
                                  forvar216 : reg303)) || $signed({reg231})) ?
                          wire16 : (reg278 ?
                              ($unsigned(reg254) ?
                                  reg291[(2'h2):(2'h2)] : $signed(reg263)) : forvar210));
                    end
                  if (reg215[(3'h6):(2'h2)])
                    begin
                      reg299 <= (|$signed($unsigned((wire15 >>> reg262))));
                      reg300 <= ($unsigned(forvar308[(1'h1):(1'h1)]) ?
                          $unsigned(reg284[(4'hd):(4'h9)]) : reg210);
                    end
                  else
                    begin
                      reg299 <= ({(~^(~&reg263))} ?
                          reg300[(4'hc):(2'h2)] : ({(~^forvar232)} ?
                              reg313 : forvar261));
                      reg300 <= ((8'h9d) + ((((8'hb4) ?
                          forvar232 : reg291) == $unsigned(reg273)) >= $unsigned($signed((8'hac)))));
                    end
                  if (reg249[(1'h0):(1'h0)])
                    begin
                      reg301 <= (&$signed((~((8'ha1) >> reg244))));
                      reg302 <= (reg243[(3'h7):(1'h0)] * forvar258);
                    end
                  else
                    begin
                      reg301 <= $signed(reg255);
                      reg302 <= $signed((~reg313[(1'h0):(1'h0)]));
                      reg303 <= (reg227[(3'h6):(2'h2)] ?
                          wire7[(3'h6):(2'h3)] : $unsigned((&$signed(forvar268))));
                    end
                end
              else
                begin
                  for (forvar297 = (1'h0); (forvar297 < (1'h0)); forvar297 = (forvar297 + (1'h1)))
                    begin
                      reg298 <= (8'hb2);
                      reg299 <= forvar293;
                      reg300 <= (^~$unsigned((~|{(8'hb9)})));
                      reg301 <= $unsigned(reg248);
                    end
                end
              for (forvar304 = (1'h0); (forvar304 < (1'h1)); forvar304 = (forvar304 + (1'h1)))
                begin
                  reg305 <= $unsigned($signed((wire12 | (reg215 ?
                      reg215 : forvar239))));
                  for (forvar306 = (1'h0); (forvar306 < (1'h0)); forvar306 = (forvar306 + (1'h1)))
                    begin
                      reg307 <= {(~&(|(reg314 ? reg217 : reg208)))};
                      reg308 <= (^$unsigned({$unsigned(reg241)}));
                      reg309 <= (&(|$signed((forvar284 | reg250))));
                      reg310 <= (forvar299 > $unsigned(((forvar232 ^~ forvar211) << (reg307 ?
                          forvar254 : reg215))));
                    end
                end
              if ((&$unsigned($signed(((8'ha2) & (8'h9d))))))
                begin
                  if ((wire12[(3'h4):(1'h1)] & $signed($signed(reg286[(3'h4):(1'h0)]))))
                    begin
                      reg311 <= (wire18[(3'h4):(1'h0)] ?
                          $signed($signed($signed(reg308))) : ($unsigned(reg309) < (|(forvar297 ?
                              reg274 : reg297))));
                      reg312 <= reg249[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg311 <= ((^~forvar268) | $signed(($signed(wire14) ~^ wire18)));
                      reg312 <= {($unsigned(reg275[(2'h3):(2'h2)]) != ((|reg275) ?
                              reg241 : reg311))};
                    end
                end
              else
                begin
                  for (forvar311 = (1'h0); (forvar311 < (1'h1)); forvar311 = (forvar311 + (1'h1)))
                    begin
                      reg312 <= $signed(forvar254);
                      reg313 <= $signed(reg301[(1'h1):(1'h0)]);
                      reg314 <= (reg295 ?
                          ($unsigned({(8'ha0)}) ?
                              reg275 : $signed((wire17 != (8'hba)))) : (~($signed(reg289) >> (forvar297 ~^ reg307))));
                      reg315 <= {(~&$unsigned($signed(forvar259)))};
                    end
                end
            end
          for (forvar316 = (1'h0); (forvar316 < (1'h1)); forvar316 = (forvar316 + (1'h1)))
            begin
              for (forvar317 = (1'h0); (forvar317 < (2'h2)); forvar317 = (forvar317 + (1'h1)))
                begin
                  for (forvar318 = (1'h0); (forvar318 < (1'h0)); forvar318 = (forvar318 + (1'h1)))
                    begin
                      reg319 <= (forvar229[(3'h5):(3'h4)] ?
                          forvar254[(1'h0):(1'h0)] : (8'hb5));
                      reg320 <= (((!reg232) && (-$unsigned(reg273))) ?
                          forvar223 : (!(-((8'hb1) ^ wire15))));
                      reg321 <= $signed(forvar267);
                    end
                end
              for (forvar322 = (1'h0); (forvar322 < (2'h2)); forvar322 = (forvar322 + (1'h1)))
                begin
                  for (forvar323 = (1'h0); (forvar323 < (1'h1)); forvar323 = (forvar323 + (1'h1)))
                    begin
                      reg324 <= $signed(($signed((reg293 ?
                          (8'ha5) : reg305)) <<< (|(|wire11))));
                      reg325 <= reg288[(2'h2):(1'h0)];
                    end
                  if (((({(8'ha7)} == (+(8'ha1))) ?
                      $signed($signed(reg269)) : {$unsigned(reg312)}) ^ ($signed((reg303 ?
                      (8'ha6) : reg315)) <<< $signed($unsigned(forvar210)))))
                    begin
                      reg326 <= $unsigned(reg238);
                      reg327 <= $unsigned((8'ha7));
                      reg328 <= $unsigned(reg308[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg326 <= reg277[(2'h2):(2'h2)];
                      reg327 <= (reg293[(3'h6):(3'h4)] - $unsigned($unsigned($unsigned(forvar259))));
                    end
                  if (((reg293 ?
                          $unsigned((|forvar304)) : reg215[(4'h8):(1'h0)]) ?
                      reg291 : forvar268))
                    begin
                      reg329 <= reg284;
                      reg330 <= reg222;
                      reg331 <= (~^$signed(reg260[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg329 <= (((^~(wire15 - reg264)) ^ $unsigned((wire290 ?
                              (8'ha3) : (8'h9d)))) ?
                          reg303[(4'h9):(3'h7)] : $signed(((reg278 >= forvar223) | reg264)));
                      reg330 <= $signed((reg248 ?
                          $unsigned((forvar316 - reg309)) : (~|(forvar317 >> forvar261))));
                    end
                end
              reg332 <= reg277;
              for (forvar333 = (1'h0); (forvar333 < (1'h1)); forvar333 = (forvar333 + (1'h1)))
                begin
                  if ({reg250})
                    begin
                      reg334 <= reg274;
                      reg335 <= (forvar223[(2'h3):(2'h3)] ?
                          ((forvar306[(2'h2):(1'h0)] ~^ (wire290 * forvar218)) > reg272) : {(~&reg324[(4'ha):(3'h5)])});
                      reg336 <= $unsigned($signed((8'h9f)));
                    end
                  else
                    begin
                      reg334 <= (~(|($unsigned((8'hb8)) ?
                          reg328 : reg298[(2'h2):(2'h2)])));
                      reg335 <= (forvar268[(2'h2):(2'h2)] ?
                          wire13[(4'h8):(2'h2)] : reg291);
                    end
                end
            end
        end
    end
  assign wire337 = $unsigned({$signed($unsigned((8'ha8)))});
  module338 modinst507 (wire506, clk, reg291, reg276, reg299, forvar258);
  always
    @(posedge clk) begin
      for (forvar508 = (1'h0); (forvar508 < (1'h0)); forvar508 = (forvar508 + (1'h1)))
        begin
          if ({$unsigned($signed((reg262 ? forvar247 : reg212)))})
            begin
              for (forvar509 = (1'h0); (forvar509 < (1'h1)); forvar509 = (forvar509 + (1'h1)))
                begin
                  if ((8'ha9))
                    begin
                      reg510 <= {({$signed((8'hb8))} >= (8'ha4))};
                      reg511 <= ((wire7 > reg334) && ($unsigned(reg325[(3'h7):(2'h2)]) ?
                          ((wire10 >> forvar229) || (forvar316 ?
                              reg243 : forvar318)) : $signed($unsigned(reg271))));
                      reg512 <= $signed(reg215);
                    end
                  else
                    begin
                      reg510 <= (!forvar299[(3'h4):(1'h0)]);
                      reg511 <= (^$unsigned(reg221[(1'h0):(1'h0)]));
                      reg512 <= forvar252;
                    end
                  reg513 <= reg238;
                  reg514 <= ((reg276 ?
                      (forvar258[(5'h10):(4'hd)] ?
                          (reg325 * reg295) : (~(8'hb4))) : reg256) == $signed($unsigned((forvar210 | reg230))));
                  if (reg335[(3'h5):(1'h1)])
                    begin
                      reg515 <= reg324[(3'h4):(2'h2)];
                      reg516 <= (((~^forvar293) || forvar254) ?
                          (&($unsigned((8'hb2)) ?
                              reg285[(4'ha):(4'h8)] : $signed(reg225))) : ($signed(wire11[(1'h0):(1'h0)]) && {$signed(reg286)}));
                      reg517 <= (wire506[(1'h0):(1'h0)] + (forvar229[(2'h3):(1'h0)] - ((reg312 ?
                              forvar293 : wire8) ?
                          (reg330 ?
                              forvar318 : reg514) : ((8'ha4) <= reg217))));
                      reg518 <= ($unsigned($signed((reg264 ^ reg308))) & ((((8'hb4) && reg230) ?
                              (reg264 ?
                                  forvar323 : (8'hac)) : (reg309 >= reg210)) ?
                          $signed((reg220 > (8'ha9))) : (~|(~^reg331))));
                    end
                  else
                    begin
                      reg515 <= $signed((^~(~|forvar245[(1'h0):(1'h0)])));
                      reg516 <= (wire506[(1'h1):(1'h1)] + $signed($unsigned($signed(reg242))));
                      reg517 <= forvar308;
                    end
                end
            end
          else
            begin
              for (forvar509 = (1'h0); (forvar509 < (1'h0)); forvar509 = (forvar509 + (1'h1)))
                begin
                  for (forvar510 = (1'h0); (forvar510 < (2'h3)); forvar510 = (forvar510 + (1'h1)))
                    begin
                      reg511 <= (~^reg300[(2'h2):(1'h1)]);
                      reg512 <= reg315;
                      reg513 <= ((wire17[(4'hc):(1'h1)] < (reg239 ?
                          $unsigned((8'hb1)) : $signed(reg236))) > {({(8'ha6)} ?
                              (forvar209 ^~ reg225) : (reg263 ~^ reg266))});
                      reg514 <= $unsigned((!reg321[(1'h1):(1'h1)]));
                    end
                  reg515 <= ($unsigned((8'ha9)) ?
                      wire9 : ($signed({forvar218}) ? reg321 : reg212));
                  for (forvar516 = (1'h0); (forvar516 < (1'h0)); forvar516 = (forvar516 + (1'h1)))
                    begin
                      reg517 <= $signed(((forvar304 ?
                          reg319[(2'h2):(1'h0)] : reg210[(2'h3):(2'h2)]) << reg233));
                      reg518 <= $signed($signed(((reg275 - reg259) ?
                          (forvar333 ?
                              reg298 : (8'h9f)) : $signed(forvar318))));
                      reg519 <= {{$unsigned(reg514[(1'h1):(1'h1)])}};
                      reg520 <= $unsigned($unsigned(reg214[(1'h0):(1'h0)]));
                    end
                end
              if ({$unsigned(((forvar210 ^~ (8'ha4)) - (forvar310 == reg282)))})
                begin
                  if ($signed($signed($signed(reg275))))
                    begin
                      reg521 <= (wire7[(3'h7):(3'h5)] ?
                          ($unsigned($unsigned(reg327)) ^ (^~reg329[(3'h6):(2'h2)])) : ((^(|forvar287)) & reg265[(1'h1):(1'h1)]));
                      reg522 <= $unsigned((|(~|(~&reg225))));
                      reg523 <= (forvar259[(1'h0):(1'h0)] ?
                          (8'hb1) : ((8'hb7) <<< (((8'ha2) < reg313) <<< (~^reg214))));
                    end
                  else
                    begin
                      reg521 <= {$unsigned(((8'hba) ?
                              (forvar299 ? reg263 : forvar232) : wire9))};
                      reg522 <= reg233[(4'hd):(4'hd)];
                    end
                  for (forvar524 = (1'h0); (forvar524 < (2'h2)); forvar524 = (forvar524 + (1'h1)))
                    begin
                      reg525 <= $signed(reg303);
                      reg526 <= reg320;
                      reg527 <= forvar213;
                    end
                  if (((-(^~{(8'hb7)})) ? reg313 : $signed((+$signed(reg255)))))
                    begin
                      reg528 <= $unsigned((+$signed(((8'hb7) - reg517))));
                    end
                  else
                    begin
                      reg528 <= ($unsigned(reg263) == wire11);
                      reg529 <= forvar239[(2'h3):(1'h1)];
                      reg530 <= wire15[(3'h6):(1'h0)];
                      reg531 <= $signed($signed((!$unsigned(reg320))));
                    end
                end
              else
                begin
                  for (forvar521 = (1'h0); (forvar521 < (2'h3)); forvar521 = (forvar521 + (1'h1)))
                    begin
                      reg522 <= (!reg283[(1'h1):(1'h1)]);
                      reg523 <= {forvar524};
                      reg524 <= ($unsigned(forvar297) ~^ reg215);
                      reg525 <= (~&reg222[(1'h0):(1'h0)]);
                    end
                  for (forvar526 = (1'h0); (forvar526 < (1'h0)); forvar526 = (forvar526 + (1'h1)))
                    begin
                      reg527 <= reg269;
                      reg528 <= ($unsigned($signed(reg294)) <<< ($unsigned((~&reg208)) ?
                          (~^$signed(forvar317)) : $unsigned(reg262[(1'h1):(1'h0)])));
                      reg529 <= (~&(($unsigned(reg249) ~^ $signed(reg293)) & {reg259}));
                      reg530 <= $signed(reg306[(2'h2):(2'h2)]);
                    end
                  for (forvar531 = (1'h0); (forvar531 < (2'h2)); forvar531 = (forvar531 + (1'h1)))
                    begin
                      reg532 <= (forvar316[(2'h3):(1'h1)] && (^forvar509));
                      reg533 <= (($unsigned(reg272[(2'h3):(2'h3)]) != (&reg217[(4'hb):(3'h5)])) ?
                          reg532[(4'hc):(3'h6)] : (8'h9e));
                      reg534 <= (($unsigned(reg529) ?
                              $signed(reg233) : ($unsigned(reg282) <<< reg286[(2'h2):(1'h0)])) ?
                          ((~&$unsigned(forvar323)) ?
                              forvar233 : (^$signed(reg516))) : reg300[(1'h0):(1'h0)]);
                      reg535 <= reg298;
                    end
                  for (forvar536 = (1'h0); (forvar536 < (2'h2)); forvar536 = (forvar536 + (1'h1)))
                    begin
                      reg537 <= $unsigned((-(((8'ha1) ?
                          reg255 : forvar224) ~^ (reg301 | forvar210))));
                      reg538 <= $unsigned({($signed(reg286) && {reg282})});
                      reg539 <= $unsigned($unsigned(((reg288 ?
                          wire17 : reg526) ^ $unsigned(reg520))));
                    end
                end
              if (reg259[(2'h3):(2'h3)])
                begin
                  reg540 <= (|reg276[(4'ha):(1'h1)]);
                  for (forvar541 = (1'h0); (forvar541 < (1'h0)); forvar541 = (forvar541 + (1'h1)))
                    begin
                      reg542 <= ((reg210 <<< $signed({forvar323})) >>> $unsigned(($signed(reg257) > reg513)));
                      reg543 <= reg542[(1'h1):(1'h0)];
                    end
                  if (reg532[(4'h9):(3'h5)])
                    begin
                      reg544 <= (forvar270 ?
                          $signed((+forvar239)) : $unsigned(reg215[(4'hb):(4'h8)]));
                      reg545 <= (forvar259[(3'h6):(3'h6)] ?
                          $signed($signed({reg263})) : (($unsigned(reg265) - (reg304 ^ reg313)) && {((8'h9e) >>> reg257)}));
                      reg546 <= (~$signed($signed($unsigned(reg253))));
                    end
                  else
                    begin
                      reg544 <= reg250;
                      reg545 <= ($unsigned((forvar254[(2'h2):(1'h1)] < {reg293})) >= ((reg517[(4'ha):(3'h4)] || $unsigned((8'h9e))) ^~ {wire337[(1'h1):(1'h0)]}));
                    end
                end
              else
                begin
                  for (forvar540 = (1'h0); (forvar540 < (2'h2)); forvar540 = (forvar540 + (1'h1)))
                    begin
                      reg541 <= ((~((8'hb1) ?
                          {reg296} : $unsigned(reg230))) - reg238);
                      reg542 <= reg324;
                    end
                  for (forvar543 = (1'h0); (forvar543 < (2'h2)); forvar543 = (forvar543 + (1'h1)))
                    begin
                      reg544 <= $signed({(~|$signed(reg276))});
                    end
                  for (forvar545 = (1'h0); (forvar545 < (2'h3)); forvar545 = (forvar545 + (1'h1)))
                    begin
                      reg546 <= reg244;
                      reg547 <= (forvar516 ?
                          (&reg271[(3'h4):(3'h4)]) : (8'h9e));
                      reg548 <= $signed((^~($signed(reg310) ?
                          $signed(wire18) : (forvar545 >> forvar211))));
                      reg549 <= (~^$signed((|(&reg319))));
                    end
                  for (forvar550 = (1'h0); (forvar550 < (2'h3)); forvar550 = (forvar550 + (1'h1)))
                    begin
                      reg551 <= reg547;
                      reg552 <= {reg255};
                      reg553 <= {$signed($unsigned({(8'ha1)}))};
                    end
                end
              reg554 <= {(({(8'hb1)} ? reg311 : $signed(reg312)) >= reg258)};
            end
          if ({reg238[(3'h5):(3'h5)]})
            begin
              for (forvar555 = (1'h0); (forvar555 < (1'h1)); forvar555 = (forvar555 + (1'h1)))
                begin
                  if ($signed($signed(forvar306[(3'h5):(3'h5)])))
                    begin
                      reg556 <= (({$unsigned(reg237)} ?
                          $unsigned(wire16) : $unsigned((~&(8'ha1)))) & $unsigned((8'h9d)));
                      reg557 <= (({(~|reg208)} ?
                              $unsigned(reg208) : ($signed(forvar254) ?
                                  $unsigned(reg301) : (forvar279 || reg551))) ?
                          (({reg324} ? $unsigned(reg214) : forvar317) ?
                              (wire15[(5'h10):(4'hf)] >= (reg524 - wire206)) : {(reg297 | reg237)}) : wire12);
                      reg558 <= {$unsigned({(reg280 ? reg303 : reg530)})};
                    end
                  else
                    begin
                      reg556 <= (($signed((-reg253)) ?
                          (^~reg543) : wire206[(1'h1):(1'h0)]) == reg336[(1'h1):(1'h0)]);
                      reg557 <= reg231[(3'h4):(2'h3)];
                      reg558 <= (8'hb7);
                      reg559 <= wire17[(3'h7):(2'h2)];
                    end
                  for (forvar560 = (1'h0); (forvar560 < (1'h1)); forvar560 = (forvar560 + (1'h1)))
                    begin
                      reg561 <= wire18[(1'h0):(1'h0)];
                      reg562 <= (-wire15);
                    end
                end
            end
          else
            begin
              if (forvar508[(4'he):(3'h6)])
                begin
                  if ((^reg243[(3'h7):(3'h7)]))
                    begin
                      reg555 <= $signed($signed(forvar311[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg555 <= $unsigned({(reg335 ?
                              (reg210 ~^ (8'hae)) : {forvar316})});
                      reg556 <= (~(8'haa));
                    end
                  for (forvar557 = (1'h0); (forvar557 < (1'h0)); forvar557 = (forvar557 + (1'h1)))
                    begin
                      reg558 <= (reg325 ?
                          ($signed((forvar247 ?
                              reg516 : forvar263)) + $signed({(8'ha1)})) : (($signed((8'haf)) >> $signed(reg271)) ?
                              (~|forvar279) : $unsigned((!reg528))));
                    end
                  if ($signed((~&$signed(((8'hb4) <<< wire17)))))
                    begin
                      reg559 <= ((8'ha4) ?
                          forvar252[(4'hc):(3'h5)] : $unsigned($signed($signed(forvar223))));
                      reg560 <= reg255[(3'h7):(1'h0)];
                      reg561 <= $unsigned(reg236[(3'h6):(3'h6)]);
                      reg562 <= forvar302;
                    end
                  else
                    begin
                      reg559 <= forvar279;
                      reg560 <= $unsigned((|(forvar555[(3'h4):(2'h3)] != (reg300 >> reg511))));
                      reg561 <= ($signed({(reg242 ?
                              reg250 : reg327)}) & $unsigned(((reg562 >>> reg557) ?
                          $unsigned((8'hb3)) : {reg302})));
                    end
                end
              else
                begin
                  for (forvar555 = (1'h0); (forvar555 < (2'h2)); forvar555 = (forvar555 + (1'h1)))
                    begin
                      reg556 <= {reg227};
                      reg557 <= $unsigned(reg519[(1'h0):(1'h0)]);
                      reg558 <= (!forvar218[(1'h1):(1'h0)]);
                    end
                  reg559 <= reg518[(1'h0):(1'h0)];
                end
            end
          for (forvar563 = (1'h0); (forvar563 < (1'h1)); forvar563 = (forvar563 + (1'h1)))
            begin
              if ($unsigned(reg230))
                begin
                  for (forvar564 = (1'h0); (forvar564 < (2'h2)); forvar564 = (forvar564 + (1'h1)))
                    begin
                      reg565 <= reg562;
                    end
                  reg566 <= (8'hb4);
                  if (forvar318[(1'h0):(1'h0)])
                    begin
                      reg567 <= {(~$signed((~^reg263)))};
                    end
                  else
                    begin
                      reg567 <= reg225;
                      reg568 <= {{(reg566 ~^ (forvar246 ?
                                  reg308 : forvar292))}};
                      reg569 <= (&(-($signed(forvar210) & (reg568 ?
                          reg250 : forvar310))));
                      reg570 <= ((({reg549} ?
                              forvar213[(4'h9):(3'h4)] : (~|reg568)) ?
                          (reg533[(3'h6):(2'h2)] ?
                              {reg528} : $unsigned((8'ha5))) : $unsigned(wire10[(1'h1):(1'h0)])) == reg248[(1'h0):(1'h0)]);
                    end
                  for (forvar571 = (1'h0); (forvar571 < (1'h1)); forvar571 = (forvar571 + (1'h1)))
                    begin
                      reg572 <= $unsigned((forvar246 & reg282[(3'h4):(2'h3)]));
                      reg573 <= (wire7 ?
                          reg219 : ($unsigned((|reg512)) >>> reg302));
                    end
                end
              else
                begin
                  for (forvar564 = (1'h0); (forvar564 < (1'h1)); forvar564 = (forvar564 + (1'h1)))
                    begin
                      reg565 <= $signed((^~(+$unsigned((8'h9e)))));
                      reg566 <= (forvar543 <= ((8'haf) + reg512));
                      reg567 <= (~^reg300);
                      reg568 <= ($signed(reg529) < ((~&$signed(reg520)) >> ((8'h9d) & $unsigned(reg234))));
                    end
                  reg569 <= reg235;
                  reg570 <= $signed((($signed(reg565) ?
                          $unsigned(reg332) : reg275[(2'h3):(2'h2)]) ?
                      $signed((~&wire13)) : ((reg541 ?
                          (8'hae) : reg313) >= $unsigned(reg525))));
                  if (reg559[(4'hf):(3'h4)])
                    begin
                      reg571 <= forvar247[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg571 <= (($unsigned((wire7 ? reg537 : forvar304)) ?
                              (~^$unsigned((8'hb6))) : (8'hac)) ?
                          forvar333[(4'ha):(3'h5)] : (-(reg526[(2'h3):(1'h0)] ?
                              $unsigned(forvar543) : (!forvar299))));
                      reg572 <= (reg297 <<< (((^~forvar232) ?
                              (reg324 ? (8'ha0) : reg569) : $unsigned(reg331)) ?
                          (^~(reg558 != reg266)) : (forvar536[(3'h4):(1'h1)] ?
                              $signed(forvar571) : reg548)));
                    end
                end
              if ({($unsigned((reg273 ? reg548 : reg565)) ?
                      (~&(~reg305)) : {reg537[(4'h8):(2'h3)]})})
                begin
                  for (forvar574 = (1'h0); (forvar574 < (1'h0)); forvar574 = (forvar574 + (1'h1)))
                    begin
                      reg575 <= $unsigned(reg291[(4'h9):(3'h6)]);
                      reg576 <= (^~($signed(reg299[(1'h0):(1'h0)]) ^~ ((~|reg568) + reg558[(4'h8):(2'h2)])));
                      reg577 <= ($unsigned(($signed(reg514) ?
                              (reg242 ?
                                  reg283 : forvar510) : $signed(reg554))) ?
                          $unsigned(((~reg327) ?
                              reg529[(4'h9):(3'h4)] : {reg327})) : (8'hb5));
                    end
                end
              else
                begin
                  for (forvar574 = (1'h0); (forvar574 < (2'h3)); forvar574 = (forvar574 + (1'h1)))
                    begin
                      reg575 <= (8'ha6);
                    end
                  for (forvar576 = (1'h0); (forvar576 < (2'h3)); forvar576 = (forvar576 + (1'h1)))
                    begin
                      reg577 <= ((forvar540 ?
                              forvar526 : forvar550[(3'h6):(3'h6)]) ?
                          {(8'hb0)} : $signed((reg253 ?
                              $unsigned(reg297) : ((8'hac) >= reg532))));
                      reg578 <= reg547[(3'h4):(3'h4)];
                      reg579 <= (forvar297[(4'hb):(1'h1)] || reg516);
                      reg580 <= $unsigned(forvar545);
                    end
                  reg581 <= {(8'hb5)};
                end
              for (forvar582 = (1'h0); (forvar582 < (2'h2)); forvar582 = (forvar582 + (1'h1)))
                begin
                  for (forvar583 = (1'h0); (forvar583 < (2'h3)); forvar583 = (forvar583 + (1'h1)))
                    begin
                      reg584 <= {(reg291 && $signed((forvar224 ?
                              reg236 : reg301)))};
                    end
                  reg585 <= ($signed((forvar287[(1'h0):(1'h0)] ?
                      reg549[(4'ha):(2'h3)] : (reg263 ?
                          wire10 : reg235))) > $signed(((reg560 * (8'h9f)) ?
                      reg561 : (reg559 ? reg523 : reg542))));
                end
            end
          reg586 <= reg511[(3'h4):(1'h0)];
        end
      for (forvar587 = (1'h0); (forvar587 < (1'h0)); forvar587 = (forvar587 + (1'h1)))
        begin
          reg588 <= (^(reg539[(2'h2):(1'h1)] & $unsigned($unsigned(forvar297))));
          for (forvar589 = (1'h0); (forvar589 < (1'h1)); forvar589 = (forvar589 + (1'h1)))
            begin
              for (forvar590 = (1'h0); (forvar590 < (2'h3)); forvar590 = (forvar590 + (1'h1)))
                begin
                  for (forvar591 = (1'h0); (forvar591 < (1'h0)); forvar591 = (forvar591 + (1'h1)))
                    begin
                      reg592 <= (reg303 > reg243);
                      reg593 <= forvar245;
                      reg594 <= reg217[(3'h5):(1'h1)];
                      reg595 <= (($unsigned((reg230 ? forvar297 : reg562)) ?
                              reg527[(4'h8):(3'h7)] : forvar224) ?
                          reg286 : {forvar587});
                    end
                  for (forvar596 = (1'h0); (forvar596 < (2'h3)); forvar596 = (forvar596 + (1'h1)))
                    begin
                      reg597 <= $unsigned(reg537);
                      reg598 <= (reg555 ?
                          (reg573[(4'hd):(3'h6)] <<< (&(^~reg283))) : ((reg265 ?
                                  (forvar509 * reg227) : reg299[(3'h6):(1'h0)]) ?
                              (((8'h9c) + reg315) > (reg576 | (8'hb7))) : $signed({forvar583})));
                    end
                  for (forvar599 = (1'h0); (forvar599 < (2'h3)); forvar599 = (forvar599 + (1'h1)))
                    begin
                      reg600 <= reg526;
                      reg601 <= $signed((((forvar245 ?
                              reg274 : reg332) + (~&reg237)) ?
                          forvar258 : ((forvar574 << forvar210) ?
                              (reg210 ? (8'ha4) : reg571) : (forvar599 ?
                                  reg528 : (8'ha3)))));
                      reg602 <= {$signed((~&reg579))};
                    end
                  if ((8'hb8))
                    begin
                      reg603 <= {forvar318[(1'h1):(1'h0)]};
                      reg604 <= forvar531;
                      reg605 <= ($unsigned(((reg521 ? (8'hb1) : reg249) ?
                              reg283[(3'h6):(3'h4)] : (^~reg308))) ?
                          (&(|(reg301 ?
                              reg553 : reg310))) : {$signed(reg282[(4'hb):(4'hb)])});
                    end
                  else
                    begin
                      reg603 <= reg580;
                      reg604 <= (~&((reg282 ?
                          $unsigned(reg567) : (~wire7)) >= ($signed(forvar267) ^~ $signed((8'hac)))));
                    end
                end
            end
        end
      for (forvar606 = (1'h0); (forvar606 < (1'h1)); forvar606 = (forvar606 + (1'h1)))
        begin
          for (forvar607 = (1'h0); (forvar607 < (2'h3)); forvar607 = (forvar607 + (1'h1)))
            begin
              for (forvar608 = (1'h0); (forvar608 < (1'h0)); forvar608 = (forvar608 + (1'h1)))
                begin
                  for (forvar609 = (1'h0); (forvar609 < (2'h3)); forvar609 = (forvar609 + (1'h1)))
                    begin
                      reg610 <= {{((reg261 ? reg533 : (8'hac)) ?
                                  $signed(reg539) : {reg518})}};
                      reg611 <= (reg573 ?
                          reg559[(4'h9):(3'h5)] : (reg274 ?
                              $signed((reg534 ?
                                  (8'ha7) : reg313)) : {{reg578}}));
                    end
                end
              for (forvar612 = (1'h0); (forvar612 < (1'h1)); forvar612 = (forvar612 + (1'h1)))
                begin
                  if (reg240)
                    begin
                      reg613 <= {($signed((|reg535)) <<< $unsigned({reg276}))};
                    end
                  else
                    begin
                      reg613 <= reg208;
                      reg614 <= {($signed((|(8'hb5))) ?
                              forvar574 : $unsigned(reg249))};
                      reg615 <= reg261[(2'h2):(2'h2)];
                    end
                end
            end
        end
    end
  assign wire616 = forvar311;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module338
#( parameter param505 = {((((8'hb5) ? (8'haa) : (8'hb2)) ? (~^(8'hb5)) : ((8'ha0) ? (8'ha1) : (8'hb4))) ? (8'hb7) : {(~(8'hb8))})} )
(y, clk, wire342, wire341, wire340, wire339);
  output wire [(32'h632):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire342;
  input wire [(4'he):(1'h0)] wire341;
  input wire [(2'h3):(1'h0)] wire340;
  input wire [(5'h10):(1'h0)] wire339;
  wire [(4'h8):(1'h0)] wire504;
  reg [(4'hb):(1'h0)] reg503 = (1'h0);
  reg [(4'h8):(1'h0)] reg502 = (1'h0);
  reg [(3'h6):(1'h0)] reg501 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar500 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg499 = (1'h0);
  reg [(3'h7):(1'h0)] reg498 = (1'h0);
  reg [(4'hb):(1'h0)] forvar497 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar496 = (1'h0);
  reg [(2'h2):(1'h0)] reg495 = (1'h0);
  reg [(5'h10):(1'h0)] reg494 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg493 = (1'h0);
  reg [(4'ha):(1'h0)] reg492 = (1'h0);
  reg [(4'he):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg490 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg489 = (1'h0);
  reg [(4'h9):(1'h0)] forvar487 = (1'h0);
  reg [(5'h10):(1'h0)] forvar485 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg488 = (1'h0);
  reg [(4'ha):(1'h0)] reg487 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg486 = (1'h0);
  reg [(4'ha):(1'h0)] reg485 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg484 = (1'h0);
  reg [(3'h4):(1'h0)] reg483 = (1'h0);
  reg [(3'h6):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg481 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar480 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar479 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg478 = (1'h0);
  reg [(4'he):(1'h0)] reg477 = (1'h0);
  reg [(4'h9):(1'h0)] reg476 = (1'h0);
  reg [(2'h3):(1'h0)] reg475 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar474 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg473 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar472 = (1'h0);
  reg [(3'h5):(1'h0)] reg471 = (1'h0);
  reg [(4'h8):(1'h0)] forvar470 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar469 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire468;
  wire signed [(2'h3):(1'h0)] wire467;
  reg signed [(2'h3):(1'h0)] reg466 = (1'h0);
  reg [(4'hc):(1'h0)] reg465 = (1'h0);
  reg [(4'he):(1'h0)] reg464 = (1'h0);
  reg [(4'ha):(1'h0)] forvar463 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg462 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg461 = (1'h0);
  reg [(4'hf):(1'h0)] reg460 = (1'h0);
  reg [(4'hb):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg458 = (1'h0);
  reg [(2'h3):(1'h0)] forvar457 = (1'h0);
  reg [(5'h10):(1'h0)] reg456 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg455 = (1'h0);
  reg [(4'h8):(1'h0)] reg454 = (1'h0);
  reg [(4'h9):(1'h0)] forvar453 = (1'h0);
  reg [(4'ha):(1'h0)] reg452 = (1'h0);
  reg [(4'hd):(1'h0)] reg451 = (1'h0);
  reg [(4'hc):(1'h0)] forvar450 = (1'h0);
  reg [(3'h7):(1'h0)] reg449 = (1'h0);
  reg [(4'he):(1'h0)] reg448 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg447 = (1'h0);
  reg [(3'h6):(1'h0)] reg446 = (1'h0);
  reg [(2'h2):(1'h0)] forvar445 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg444 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg443 = (1'h0);
  reg [(3'h7):(1'h0)] reg442 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg441 = (1'h0);
  reg [(4'hd):(1'h0)] forvar440 = (1'h0);
  reg [(2'h3):(1'h0)] forvar439 = (1'h0);
  reg [(4'he):(1'h0)] reg432 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar431 = (1'h0);
  reg [(4'hd):(1'h0)] reg427 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg438 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg436 = (1'h0);
  reg [(4'h9):(1'h0)] reg435 = (1'h0);
  reg [(4'hc):(1'h0)] reg434 = (1'h0);
  reg [(4'hb):(1'h0)] reg433 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar432 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg431 = (1'h0);
  reg [(2'h2):(1'h0)] reg430 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg429 = (1'h0);
  reg [(4'he):(1'h0)] reg428 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar427 = (1'h0);
  reg [(4'h9):(1'h0)] forvar426 = (1'h0);
  reg [(4'h9):(1'h0)] reg425 = (1'h0);
  reg [(3'h7):(1'h0)] reg424 = (1'h0);
  reg [(2'h2):(1'h0)] reg423 = (1'h0);
  reg [(4'ha):(1'h0)] reg422 = (1'h0);
  reg [(4'hc):(1'h0)] forvar421 = (1'h0);
  reg [(4'he):(1'h0)] reg420 = (1'h0);
  reg [(2'h2):(1'h0)] reg419 = (1'h0);
  reg [(4'he):(1'h0)] reg418 = (1'h0);
  reg [(4'h8):(1'h0)] reg417 = (1'h0);
  reg [(3'h4):(1'h0)] reg416 = (1'h0);
  reg [(3'h7):(1'h0)] forvar415 = (1'h0);
  reg [(4'h9):(1'h0)] reg414 = (1'h0);
  reg [(3'h7):(1'h0)] forvar413 = (1'h0);
  reg [(3'h7):(1'h0)] forvar405 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar402 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg407 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar404 = (1'h0);
  reg [(4'hc):(1'h0)] reg412 = (1'h0);
  reg [(4'ha):(1'h0)] reg411 = (1'h0);
  reg [(4'h8):(1'h0)] reg410 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg409 = (1'h0);
  reg [(4'ha):(1'h0)] reg408 = (1'h0);
  reg [(3'h6):(1'h0)] forvar407 = (1'h0);
  reg [(2'h2):(1'h0)] reg406 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg405 = (1'h0);
  reg [(4'h8):(1'h0)] reg404 = (1'h0);
  reg [(4'hd):(1'h0)] reg403 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg402 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar401 = (1'h0);
  reg [(3'h7):(1'h0)] forvar400 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar385 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar386 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg382 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar381 = (1'h0);
  reg [(3'h6):(1'h0)] forvar380 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg401 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg396 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar395 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar393 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg390 = (1'h0);
  reg [(2'h3):(1'h0)] forvar389 = (1'h0);
  reg [(3'h5):(1'h0)] forvar388 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg400 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg399 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg398 = (1'h0);
  reg [(4'ha):(1'h0)] reg397 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar396 = (1'h0);
  reg [(2'h2):(1'h0)] reg395 = (1'h0);
  reg [(4'hc):(1'h0)] reg394 = (1'h0);
  reg [(4'hd):(1'h0)] reg393 = (1'h0);
  reg [(4'hf):(1'h0)] reg392 = (1'h0);
  reg [(2'h3):(1'h0)] forvar391 = (1'h0);
  reg [(3'h4):(1'h0)] forvar390 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg389 = (1'h0);
  reg [(4'h9):(1'h0)] reg388 = (1'h0);
  reg [(5'h10):(1'h0)] reg387 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg386 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg385 = (1'h0);
  reg [(3'h6):(1'h0)] reg384 = (1'h0);
  reg [(2'h3):(1'h0)] reg383 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar382 = (1'h0);
  reg [(3'h5):(1'h0)] reg381 = (1'h0);
  reg [(4'h9):(1'h0)] reg380 = (1'h0);
  reg [(4'ha):(1'h0)] reg379 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar378 = (1'h0);
  reg [(3'h4):(1'h0)] forvar377 = (1'h0);
  reg [(4'hf):(1'h0)] reg376 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg375 = (1'h0);
  reg signed [(4'he):(1'h0)] reg374 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg373 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg372 = (1'h0);
  reg [(4'hc):(1'h0)] forvar371 = (1'h0);
  reg [(3'h5):(1'h0)] reg370 = (1'h0);
  reg [(2'h2):(1'h0)] reg369 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar368 = (1'h0);
  reg signed [(4'he):(1'h0)] reg367 = (1'h0);
  reg [(3'h7):(1'h0)] reg366 = (1'h0);
  reg [(4'ha):(1'h0)] reg365 = (1'h0);
  reg [(3'h7):(1'h0)] reg364 = (1'h0);
  reg [(2'h2):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar362 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar361 = (1'h0);
  reg [(3'h7):(1'h0)] reg360 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg359 = (1'h0);
  reg [(2'h2):(1'h0)] reg358 = (1'h0);
  reg [(4'he):(1'h0)] reg357 = (1'h0);
  reg [(4'he):(1'h0)] forvar356 = (1'h0);
  reg [(3'h4):(1'h0)] forvar355 = (1'h0);
  reg [(3'h4):(1'h0)] reg354 = (1'h0);
  reg [(4'he):(1'h0)] forvar353 = (1'h0);
  reg [(4'hb):(1'h0)] reg352 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg350 = (1'h0);
  reg [(3'h6):(1'h0)] reg349 = (1'h0);
  reg [(4'ha):(1'h0)] forvar348 = (1'h0);
  reg [(4'h9):(1'h0)] reg347 = (1'h0);
  reg [(2'h3):(1'h0)] forvar346 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar345 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar344 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar343 = (1'h0);
  assign y = {wire504,
                 reg503,
                 reg502,
                 reg501,
                 forvar500,
                 reg499,
                 reg498,
                 forvar497,
                 forvar496,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg490,
                 reg489,
                 forvar487,
                 forvar485,
                 reg488,
                 reg487,
                 reg486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 forvar480,
                 forvar479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 forvar474,
                 reg473,
                 forvar472,
                 reg471,
                 forvar470,
                 forvar469,
                 wire468,
                 wire467,
                 reg466,
                 reg465,
                 reg464,
                 forvar463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg458,
                 forvar457,
                 reg456,
                 reg455,
                 reg454,
                 forvar453,
                 reg452,
                 reg451,
                 forvar450,
                 reg449,
                 reg448,
                 reg447,
                 reg446,
                 forvar445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 forvar440,
                 forvar439,
                 reg432,
                 forvar431,
                 reg427,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 forvar432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 forvar427,
                 forvar426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 forvar421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 forvar415,
                 reg414,
                 forvar413,
                 forvar405,
                 forvar402,
                 reg407,
                 forvar404,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 forvar407,
                 reg406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 forvar401,
                 forvar400,
                 forvar385,
                 forvar386,
                 reg382,
                 forvar381,
                 forvar380,
                 reg401,
                 reg396,
                 forvar395,
                 forvar393,
                 reg391,
                 reg390,
                 forvar389,
                 forvar388,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 forvar396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 forvar391,
                 forvar390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 reg383,
                 forvar382,
                 reg381,
                 reg380,
                 reg379,
                 forvar378,
                 forvar377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 forvar371,
                 reg370,
                 reg369,
                 forvar368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 forvar362,
                 forvar361,
                 reg360,
                 reg359,
                 reg358,
                 reg357,
                 forvar356,
                 forvar355,
                 reg354,
                 forvar353,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 forvar348,
                 reg347,
                 forvar346,
                 forvar345,
                 forvar344,
                 forvar343,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar343 = (1'h0); (forvar343 < (1'h1)); forvar343 = (forvar343 + (1'h1)))
        begin
          for (forvar344 = (1'h0); (forvar344 < (2'h2)); forvar344 = (forvar344 + (1'h1)))
            begin
              for (forvar345 = (1'h0); (forvar345 < (2'h2)); forvar345 = (forvar345 + (1'h1)))
                begin
                  for (forvar346 = (1'h0); (forvar346 < (2'h2)); forvar346 = (forvar346 + (1'h1)))
                    begin
                      reg347 <= $unsigned({forvar345});
                    end
                end
              if ((+(reg347 ? $signed(reg347[(2'h3):(1'h1)]) : forvar343)))
                begin
                  for (forvar348 = (1'h0); (forvar348 < (1'h1)); forvar348 = (forvar348 + (1'h1)))
                    begin
                      reg349 <= $unsigned($signed($unsigned($unsigned((8'ha0)))));
                      reg350 <= $signed(wire339[(4'h9):(1'h1)]);
                      reg351 <= reg350[(2'h2):(2'h2)];
                      reg352 <= $signed((|forvar346[(2'h2):(2'h2)]));
                    end
                  for (forvar353 = (1'h0); (forvar353 < (1'h1)); forvar353 = (forvar353 + (1'h1)))
                    begin
                      reg354 <= reg349[(3'h5):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar348 = (1'h0); (forvar348 < (2'h3)); forvar348 = (forvar348 + (1'h1)))
                    begin
                      reg349 <= ($unsigned(reg347[(2'h3):(1'h0)]) - ($signed(wire342) ?
                          wire342 : $unsigned((forvar343 && forvar344))));
                      reg350 <= reg350[(4'h8):(1'h0)];
                    end
                end
              for (forvar355 = (1'h0); (forvar355 < (2'h2)); forvar355 = (forvar355 + (1'h1)))
                begin
                  for (forvar356 = (1'h0); (forvar356 < (1'h0)); forvar356 = (forvar356 + (1'h1)))
                    begin
                      reg357 <= {$unsigned($signed((!forvar355)))};
                      reg358 <= (($signed(forvar345[(3'h5):(2'h2)]) ?
                          reg347[(3'h5):(2'h3)] : (8'hb7)) ~^ ((~&(!(8'hb1))) ^ {reg357[(3'h4):(2'h2)]}));
                      reg359 <= reg352;
                    end
                end
            end
          reg360 <= forvar343[(2'h2):(1'h1)];
          for (forvar361 = (1'h0); (forvar361 < (1'h1)); forvar361 = (forvar361 + (1'h1)))
            begin
              if (forvar344[(2'h3):(2'h2)])
                begin
                  for (forvar362 = (1'h0); (forvar362 < (2'h2)); forvar362 = (forvar362 + (1'h1)))
                    begin
                      reg363 <= {(~|($unsigned(wire339) ?
                              $signed(forvar361) : {(8'haa)}))};
                    end
                end
              else
                begin
                  for (forvar362 = (1'h0); (forvar362 < (2'h3)); forvar362 = (forvar362 + (1'h1)))
                    begin
                      reg363 <= ($unsigned(($unsigned(reg351) ?
                          (~&forvar348) : $unsigned(reg359))) < reg347[(2'h2):(1'h1)]);
                      reg364 <= reg347[(4'h8):(3'h4)];
                      reg365 <= (reg354[(3'h4):(2'h3)] ?
                          (wire339[(2'h2):(1'h0)] == $unsigned(forvar355[(2'h3):(1'h0)])) : forvar345);
                      reg366 <= (~|{$signed((~|forvar362))});
                    end
                  reg367 <= (+(reg351[(1'h0):(1'h0)] ?
                      (forvar343 ?
                          (!reg360) : (8'hab)) : ($unsigned(reg366) || forvar348[(4'h9):(2'h2)])));
                  for (forvar368 = (1'h0); (forvar368 < (1'h0)); forvar368 = (forvar368 + (1'h1)))
                    begin
                      reg369 <= reg350;
                      reg370 <= ($signed(forvar361[(2'h2):(1'h1)]) ?
                          forvar346[(1'h1):(1'h0)] : (~|reg352));
                    end
                end
              for (forvar371 = (1'h0); (forvar371 < (1'h1)); forvar371 = (forvar371 + (1'h1)))
                begin
                  reg372 <= $signed(reg359[(3'h6):(3'h6)]);
                  if (forvar371)
                    begin
                      reg373 <= (reg350 ?
                          {(reg370[(2'h2):(1'h1)] ?
                                  (reg350 << reg357) : (wire342 ~^ forvar368))} : (!(((8'hb2) ?
                                  wire342 : (8'hae)) ?
                              (wire340 ?
                                  reg347 : wire341) : $signed(forvar353))));
                    end
                  else
                    begin
                      reg373 <= reg369[(1'h1):(1'h1)];
                      reg374 <= $unsigned(reg369[(1'h0):(1'h0)]);
                      reg375 <= $signed(reg374[(3'h4):(1'h1)]);
                    end
                  reg376 <= ($signed({(reg372 ? reg347 : wire339)}) ?
                      (-($signed(reg374) <<< reg375[(1'h0):(1'h0)])) : $signed((+$signed(reg365))));
                end
            end
        end
      if ((wire341 >= forvar343))
        begin
          for (forvar377 = (1'h0); (forvar377 < (1'h1)); forvar377 = (forvar377 + (1'h1)))
            begin
              for (forvar378 = (1'h0); (forvar378 < (1'h0)); forvar378 = (forvar378 + (1'h1)))
                begin
                  if (($signed((reg370[(1'h0):(1'h0)] >= (reg375 > (8'hac)))) ^~ ({reg347[(4'h8):(4'h8)]} ?
                      (~((8'hb1) >= reg376)) : $unsigned(reg347[(4'h8):(3'h7)]))))
                    begin
                      reg379 <= (8'ha3);
                      reg380 <= (($signed($signed(forvar355)) ?
                          ((reg354 ? reg367 : forvar348) ~^ (forvar344 ?
                              reg359 : (8'h9c))) : forvar371[(4'h8):(4'h8)]) <= (&((forvar353 * reg365) + $unsigned(reg358))));
                      reg381 <= reg380[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg379 <= {(^~({(8'hb9)} << wire340))};
                      reg380 <= (~|(!((reg354 ? reg358 : forvar344) ?
                          forvar353 : $signed((8'ha4)))));
                      reg381 <= (|(-(forvar343[(3'h6):(1'h1)] ?
                          $signed(wire342) : ((8'ha6) ?
                              forvar377 : forvar353))));
                    end
                  for (forvar382 = (1'h0); (forvar382 < (1'h1)); forvar382 = (forvar382 + (1'h1)))
                    begin
                      reg383 <= {({$signed(reg375)} ?
                              forvar356[(3'h5):(2'h2)] : ($unsigned(reg350) <= (reg347 ?
                                  reg352 : forvar355)))};
                      reg384 <= $unsigned($signed(((reg357 ?
                              reg376 : forvar371) ?
                          (~reg372) : (~&reg360))));
                    end
                  if (forvar348[(4'ha):(3'h5)])
                    begin
                      reg385 <= ({(~|(reg350 < reg347))} >>> (((~forvar353) ?
                              {reg351} : (reg367 ? wire341 : reg364)) ?
                          $signed(forvar382) : $unsigned($unsigned(forvar355))));
                      reg386 <= (~forvar361[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg385 <= ((~(~|(forvar382 ? reg385 : forvar368))) ?
                          $unsigned((~^$unsigned(forvar362))) : $unsigned($unsigned($signed(reg354))));
                    end
                  reg387 <= reg376[(3'h5):(3'h4)];
                end
            end
          if (reg349)
            begin
              reg388 <= $signed((forvar368 && $signed((!(8'h9c)))));
              reg389 <= ((~$unsigned(((8'hab) < reg350))) - {$unsigned(reg354[(1'h1):(1'h1)])});
              for (forvar390 = (1'h0); (forvar390 < (1'h1)); forvar390 = (forvar390 + (1'h1)))
                begin
                  for (forvar391 = (1'h0); (forvar391 < (1'h0)); forvar391 = (forvar391 + (1'h1)))
                    begin
                      reg392 <= (($unsigned({forvar344}) ^ ({forvar348} ?
                          (&reg367) : (forvar348 ?
                              reg384 : forvar378))) >= {reg373[(1'h0):(1'h0)]});
                      reg393 <= reg392;
                      reg394 <= (~$signed($unsigned((8'haa))));
                      reg395 <= (8'ha0);
                    end
                  for (forvar396 = (1'h0); (forvar396 < (1'h1)); forvar396 = (forvar396 + (1'h1)))
                    begin
                      reg397 <= $signed((reg393[(1'h0):(1'h0)] >> $signed(forvar390[(3'h4):(3'h4)])));
                      reg398 <= ((+reg357[(4'ha):(3'h6)]) ?
                          $signed(reg376[(2'h2):(1'h0)]) : forvar353[(1'h1):(1'h1)]);
                      reg399 <= reg350;
                    end
                  reg400 <= (($unsigned($signed(forvar362)) >>> (reg381 ?
                          (forvar353 ? reg394 : reg367) : forvar371)) ?
                      forvar396[(3'h6):(2'h3)] : $signed($unsigned($signed(reg373))));
                end
            end
          else
            begin
              for (forvar388 = (1'h0); (forvar388 < (1'h1)); forvar388 = (forvar388 + (1'h1)))
                begin
                  for (forvar389 = (1'h0); (forvar389 < (1'h1)); forvar389 = (forvar389 + (1'h1)))
                    begin
                      reg390 <= $signed((((forvar388 ? reg385 : forvar391) ?
                              (reg372 ?
                                  reg384 : wire342) : reg369[(1'h1):(1'h1)]) ?
                          wire341[(4'h8):(2'h3)] : $unsigned($unsigned(forvar355))));
                      reg391 <= {$signed((+{(8'hb1)}))};
                      reg392 <= $signed((^~((+forvar362) ?
                          $signed(forvar391) : {reg375})));
                    end
                  for (forvar393 = (1'h0); (forvar393 < (1'h1)); forvar393 = (forvar393 + (1'h1)))
                    begin
                      reg394 <= (+(&reg388[(2'h3):(2'h2)]));
                    end
                  for (forvar395 = (1'h0); (forvar395 < (2'h2)); forvar395 = (forvar395 + (1'h1)))
                    begin
                      reg396 <= (~^$signed(reg349[(3'h5):(1'h1)]));
                      reg397 <= (~&$unsigned($signed({reg373})));
                      reg398 <= ((($signed(forvar348) ?
                                  reg354[(2'h3):(1'h0)] : reg395) ?
                              ((8'hac) ? (8'ha4) : $signed(reg359)) : (8'ha4)) ?
                          ($unsigned((~^forvar393)) ?
                              ((!reg367) >= reg360[(2'h2):(1'h0)]) : (|(forvar393 * forvar396))) : reg392[(4'ha):(1'h0)]);
                      reg399 <= $signed(reg396);
                    end
                  if (reg380[(4'h8):(2'h2)])
                    begin
                      reg400 <= $unsigned((~&$unsigned((|reg376))));
                      reg401 <= $unsigned((^~wire341));
                    end
                  else
                    begin
                      reg400 <= $unsigned(((reg397[(4'h9):(3'h7)] ?
                          (forvar382 <<< forvar344) : $signed(forvar371)) && ($unsigned((8'ha7)) || forvar393)));
                      reg401 <= ({(8'hba)} & forvar390[(3'h4):(1'h1)]);
                    end
                end
            end
        end
      else
        begin
          if ($unsigned(forvar378))
            begin
              for (forvar377 = (1'h0); (forvar377 < (2'h3)); forvar377 = (forvar377 + (1'h1)))
                begin
                  for (forvar378 = (1'h0); (forvar378 < (1'h0)); forvar378 = (forvar378 + (1'h1)))
                    begin
                      reg379 <= $signed($unsigned(($signed(reg365) < $signed(reg360))));
                    end
                end
              for (forvar380 = (1'h0); (forvar380 < (2'h2)); forvar380 = (forvar380 + (1'h1)))
                begin
                  for (forvar381 = (1'h0); (forvar381 < (1'h1)); forvar381 = (forvar381 + (1'h1)))
                    begin
                      reg382 <= $unsigned($unsigned($unsigned({reg360})));
                      reg383 <= $signed(reg396[(2'h2):(2'h2)]);
                      reg384 <= reg360[(2'h2):(2'h2)];
                      reg385 <= (reg352 | $unsigned(({reg363} + $signed(forvar371))));
                    end
                  for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
                    begin
                      reg387 <= $unsigned(($unsigned($signed(forvar381)) + ((reg357 >> reg351) ?
                          (~|reg396) : $signed(forvar355))));
                    end
                end
              for (forvar388 = (1'h0); (forvar388 < (1'h1)); forvar388 = (forvar388 + (1'h1)))
                begin
                  for (forvar389 = (1'h0); (forvar389 < (1'h1)); forvar389 = (forvar389 + (1'h1)))
                    begin
                      reg390 <= forvar368[(1'h0):(1'h0)];
                      reg391 <= (((^$unsigned(reg358)) <= reg390) + reg392);
                    end
                end
              reg392 <= forvar391;
            end
          else
            begin
              for (forvar377 = (1'h0); (forvar377 < (2'h3)); forvar377 = (forvar377 + (1'h1)))
                begin
                  for (forvar378 = (1'h0); (forvar378 < (1'h0)); forvar378 = (forvar378 + (1'h1)))
                    begin
                      reg379 <= ((((reg388 && forvar391) != $unsigned(reg366)) ~^ (forvar371[(4'hb):(1'h0)] ?
                          (forvar393 ? reg383 : (8'hba)) : (reg390 ?
                              forvar343 : reg370))) >> reg381[(1'h0):(1'h0)]);
                      reg380 <= wire339;
                    end
                  if ((-(8'ha0)))
                    begin
                      reg381 <= reg396;
                      reg382 <= (^reg399[(1'h0):(1'h0)]);
                      reg383 <= (reg370 + (forvar386[(1'h0):(1'h0)] << ((forvar380 ?
                              reg389 : wire342) ?
                          (forvar389 - reg384) : $unsigned((8'hb0)))));
                      reg384 <= {(~(^$signed(reg381)))};
                    end
                  else
                    begin
                      reg381 <= reg385[(1'h1):(1'h0)];
                      reg382 <= {({(forvar381 == reg396)} == ($unsigned(reg366) <= (forvar396 ?
                              reg397 : wire340)))};
                    end
                  for (forvar385 = (1'h0); (forvar385 < (1'h0)); forvar385 = (forvar385 + (1'h1)))
                    begin
                      reg386 <= reg400[(1'h0):(1'h0)];
                      reg387 <= $signed(forvar382);
                    end
                end
              if (reg396)
                begin
                  for (forvar388 = (1'h0); (forvar388 < (2'h2)); forvar388 = (forvar388 + (1'h1)))
                    begin
                      reg389 <= $signed((reg359[(3'h6):(3'h6)] * $unsigned(reg383)));
                      reg390 <= forvar371[(4'ha):(3'h4)];
                    end
                  for (forvar391 = (1'h0); (forvar391 < (2'h3)); forvar391 = (forvar391 + (1'h1)))
                    begin
                      reg392 <= $unsigned($unsigned({(reg374 ?
                              (8'hb8) : (8'haf))}));
                      reg393 <= {forvar368[(1'h0):(1'h0)]};
                      reg394 <= (8'ha0);
                      reg395 <= $unsigned(reg363);
                    end
                  if ((wire342 ?
                      (reg365 >> (-(~|forvar382))) : $unsigned(forvar356[(4'he):(3'h5)])))
                    begin
                      reg396 <= (^$unsigned(($unsigned(forvar348) | (reg400 & reg401))));
                      reg397 <= (forvar378[(2'h3):(2'h3)] ?
                          (8'haa) : (forvar391[(1'h0):(1'h0)] != reg397[(4'h9):(3'h4)]));
                      reg398 <= ((+$signed(reg387[(4'he):(4'h9)])) <<< $unsigned($unsigned($unsigned(forvar391))));
                      reg399 <= $signed(($unsigned((wire341 ~^ (8'hb5))) && $unsigned(forvar362)));
                    end
                  else
                    begin
                      reg396 <= (-reg359);
                      reg397 <= ({{(~wire342)}} ?
                          (~^$unsigned(((8'haf) ?
                              reg349 : reg392))) : (reg394[(1'h0):(1'h0)] <= (8'ha0)));
                    end
                end
              else
                begin
                  if ((8'hb9))
                    begin
                      reg388 <= {reg383};
                      reg389 <= ($signed(reg354) || (reg365 ?
                          reg374 : $unsigned((reg365 ^~ reg385))));
                      reg390 <= (forvar388 << reg347);
                      reg391 <= (forvar344 ?
                          ((reg397 != (^~forvar344)) ?
                              ((reg347 ? reg379 : reg385) ?
                                  forvar353 : reg386) : $unsigned(reg369)) : (((8'ha1) ?
                              (reg375 ? reg397 : wire341) : (forvar353 ?
                                  wire340 : reg388)) || (8'ha9)));
                    end
                  else
                    begin
                      reg388 <= $unsigned(({$signed(reg354)} >>> ((~reg400) != reg363[(1'h1):(1'h0)])));
                      reg389 <= $unsigned($unsigned(((8'h9c) ^~ (reg390 ?
                          reg389 : wire340))));
                    end
                  if ($signed($signed($signed(((8'ha6) ? (8'ha0) : reg390)))))
                    begin
                      reg392 <= ($signed(reg358[(1'h1):(1'h1)]) ?
                          $signed((forvar361[(1'h0):(1'h0)] >> (reg394 ^ (8'hb2)))) : {$unsigned((|forvar389))});
                      reg393 <= (($signed((reg373 >= forvar381)) ?
                          $signed((reg391 >> (8'h9c))) : $signed(((8'haf) & (8'hba)))) >>> forvar353[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg392 <= (reg350 ?
                          (~|(~^(reg389 | forvar356))) : (reg369[(1'h1):(1'h0)] ?
                              ($signed(reg389) ?
                                  (8'hb1) : $signed(forvar386)) : {(reg376 | forvar346)}));
                      reg393 <= forvar368;
                      reg394 <= (($unsigned((forvar382 ? forvar395 : reg382)) ?
                          reg389[(2'h3):(2'h3)] : ({reg375} == reg352[(3'h6):(2'h3)])) << $signed($signed($signed(reg376))));
                    end
                  if (reg380)
                    begin
                      reg395 <= {{($signed(forvar356) >> $unsigned(forvar396))}};
                      reg396 <= (((8'hac) < $unsigned(reg381[(1'h1):(1'h1)])) ?
                          reg387[(1'h1):(1'h1)] : (forvar395 ?
                              $signed(forvar396) : (reg360 | $signed(reg367))));
                    end
                  else
                    begin
                      reg395 <= ($signed(reg350[(4'h9):(3'h7)]) >>> ($unsigned({(8'haf)}) > (reg395 ?
                          reg369[(1'h0):(1'h0)] : (forvar389 ?
                              reg390 : (8'haa)))));
                      reg396 <= $unsigned(((reg381[(3'h5):(3'h5)] ?
                              (forvar385 >= reg398) : $signed(reg393)) ?
                          $signed($unsigned(forvar353)) : ($unsigned(reg349) ?
                              reg388[(2'h3):(1'h0)] : $signed((8'hb9)))));
                      reg397 <= {forvar378};
                    end
                end
            end
          if ((((forvar348 ?
              {reg379} : wire339[(3'h7):(2'h3)]) <= {(~|reg385)}) > (reg351 ^ $unsigned((8'hb3)))))
            begin
              for (forvar400 = (1'h0); (forvar400 < (1'h1)); forvar400 = (forvar400 + (1'h1)))
                begin
                  for (forvar401 = (1'h0); (forvar401 < (2'h3)); forvar401 = (forvar401 + (1'h1)))
                    begin
                      reg402 <= (wire341[(4'hd):(2'h3)] ?
                          ((&(~^forvar380)) ?
                              $unsigned((forvar348 ^ forvar356)) : $unsigned(reg352)) : (reg350[(3'h4):(2'h2)] ?
                              $unsigned({reg385}) : (~(reg398 * reg384))));
                    end
                  if (forvar353[(2'h2):(1'h1)])
                    begin
                      reg403 <= $signed(reg384[(1'h0):(1'h0)]);
                      reg404 <= $signed(reg382);
                      reg405 <= $unsigned(((forvar346[(1'h1):(1'h1)] ?
                              (forvar361 ? (8'haa) : wire342) : (-reg350)) ?
                          ($unsigned(forvar385) ?
                              (forvar353 ?
                                  reg367 : reg404) : (reg347 ~^ forvar395)) : reg372[(3'h4):(1'h1)]));
                    end
                  else
                    begin
                      reg403 <= (&forvar356[(4'hd):(4'h9)]);
                      reg404 <= reg382[(1'h1):(1'h0)];
                    end
                  reg406 <= $signed($unsigned(forvar401));
                end
              for (forvar407 = (1'h0); (forvar407 < (1'h0)); forvar407 = (forvar407 + (1'h1)))
                begin
                  if (((+((!reg369) ?
                      {reg372} : forvar391[(1'h0):(1'h0)])) < reg372[(2'h3):(2'h2)]))
                    begin
                      reg408 <= {((~$signed((8'hab))) ?
                              $signed((forvar385 >> (8'hae))) : $signed(reg347))};
                      reg409 <= ($signed($unsigned((&forvar391))) ?
                          $signed($unsigned($signed(reg392))) : $signed(reg392));
                      reg410 <= ($signed($unsigned((reg370 >>> reg379))) >> (~reg376));
                      reg411 <= {$signed(($unsigned(reg385) ?
                              $signed(forvar348) : $unsigned(reg408)))};
                    end
                  else
                    begin
                      reg408 <= reg382;
                    end
                  reg412 <= $signed(reg389[(3'h4):(1'h0)]);
                end
            end
          else
            begin
              if ({$signed({(forvar371 || reg404)})})
                begin
                  for (forvar400 = (1'h0); (forvar400 < (1'h0)); forvar400 = (forvar400 + (1'h1)))
                    begin
                      reg401 <= (((+((8'h9e) * forvar368)) < $unsigned(reg383)) ^~ {forvar390});
                      reg402 <= forvar378;
                      reg403 <= (forvar385 & (((reg373 * reg357) ?
                          (forvar386 ?
                              reg365 : (8'haa)) : (~&reg412)) >= $unsigned((!reg370))));
                    end
                  for (forvar404 = (1'h0); (forvar404 < (1'h1)); forvar404 = (forvar404 + (1'h1)))
                    begin
                      reg405 <= (~(((forvar353 ?
                          reg354 : reg373) ~^ $signed(forvar388)) || ((+(8'hb6)) ^ $unsigned(reg347))));
                      reg406 <= reg388[(2'h3):(2'h3)];
                      reg407 <= (+(forvar356[(3'h5):(1'h1)] > ($unsigned(reg389) ?
                          $unsigned(forvar346) : reg370[(3'h5):(2'h3)])));
                      reg408 <= (~|reg411);
                    end
                end
              else
                begin
                  for (forvar400 = (1'h0); (forvar400 < (1'h1)); forvar400 = (forvar400 + (1'h1)))
                    begin
                      reg401 <= (reg352 ?
                          $unsigned(forvar389[(2'h2):(1'h0)]) : $signed(reg359[(3'h5):(3'h5)]));
                    end
                  for (forvar402 = (1'h0); (forvar402 < (2'h3)); forvar402 = (forvar402 + (1'h1)))
                    begin
                      reg403 <= (~|(reg379[(2'h3):(1'h1)] != reg354));
                      reg404 <= (+($unsigned((forvar385 ?
                          forvar395 : reg380)) != $signed(forvar401)));
                    end
                  for (forvar405 = (1'h0); (forvar405 < (2'h2)); forvar405 = (forvar405 + (1'h1)))
                    begin
                      reg406 <= $signed((^~(!$signed(forvar405))));
                      reg407 <= $signed($signed(((8'h9d) >> reg380[(4'h8):(3'h5)])));
                    end
                  reg408 <= (8'hb1);
                end
            end
          for (forvar413 = (1'h0); (forvar413 < (1'h1)); forvar413 = (forvar413 + (1'h1)))
            begin
              reg414 <= {({forvar345} - {(^wire339)})};
              for (forvar415 = (1'h0); (forvar415 < (2'h2)); forvar415 = (forvar415 + (1'h1)))
                begin
                  if (forvar404[(4'hb):(1'h1)])
                    begin
                      reg416 <= (~(reg390[(1'h1):(1'h0)] << reg408[(3'h5):(1'h1)]));
                      reg417 <= forvar388[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg416 <= $unsigned(reg395);
                    end
                  if ((forvar377 ?
                      (reg381 ?
                          reg360[(3'h6):(1'h0)] : $signed(forvar402)) : (-((-forvar396) ?
                          $signed(forvar345) : $signed(reg379)))))
                    begin
                      reg418 <= $signed($signed($signed($unsigned(reg367))));
                    end
                  else
                    begin
                      reg418 <= (reg407[(2'h2):(1'h0)] ?
                          forvar415[(2'h3):(1'h0)] : $unsigned(forvar402[(2'h3):(2'h2)]));
                      reg419 <= (~|((forvar371 < reg358[(2'h2):(1'h1)]) ?
                          forvar345[(4'h8):(1'h1)] : reg406[(1'h1):(1'h0)]));
                      reg420 <= reg350[(5'h10):(4'hf)];
                    end
                  for (forvar421 = (1'h0); (forvar421 < (2'h2)); forvar421 = (forvar421 + (1'h1)))
                    begin
                      reg422 <= $signed({$unsigned(reg372)});
                    end
                  if (($signed(($signed(forvar402) ^ $signed(reg375))) ?
                      $unsigned($signed((forvar390 ?
                          (8'hb0) : reg366))) : $unsigned(((wire341 != forvar393) - (reg350 ?
                          reg350 : reg404)))))
                    begin
                      reg423 <= $unsigned((((reg386 ~^ reg409) <<< reg351) ^~ $signed($signed(reg387))));
                      reg424 <= forvar401;
                      reg425 <= reg395[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg423 <= forvar348;
                    end
                end
            end
          for (forvar426 = (1'h0); (forvar426 < (2'h3)); forvar426 = (forvar426 + (1'h1)))
            begin
              if (forvar388[(3'h4):(3'h4)])
                begin
                  for (forvar427 = (1'h0); (forvar427 < (1'h0)); forvar427 = (forvar427 + (1'h1)))
                    begin
                      reg428 <= (~&(((reg393 ?
                          reg376 : forvar407) == $unsigned((8'ha0))) < $unsigned({reg365})));
                      reg429 <= $signed(reg358);
                      reg430 <= (~^reg410[(1'h1):(1'h0)]);
                      reg431 <= $signed((reg373[(3'h4):(2'h3)] + ({reg385} ?
                          $signed(forvar407) : $unsigned(reg392))));
                    end
                  for (forvar432 = (1'h0); (forvar432 < (2'h2)); forvar432 = (forvar432 + (1'h1)))
                    begin
                      reg433 <= (({(reg409 ? reg414 : (8'hba))} ?
                              ((reg385 ?
                                  wire340 : reg416) >>> $signed(reg367)) : $unsigned((reg393 ?
                                  reg384 : (8'ha9)))) ?
                          reg352 : (~^reg347[(4'h8):(3'h4)]));
                    end
                  if ({(reg414[(4'h8):(3'h5)] ?
                          ((forvar390 ?
                              reg373 : reg405) + reg360) : $signed((forvar381 ^~ forvar356)))})
                    begin
                      reg434 <= ((^~reg385[(3'h4):(1'h0)]) - (-reg405));
                    end
                  else
                    begin
                      reg434 <= ({((wire342 ~^ reg372) - reg388[(3'h7):(3'h7)])} ?
                          {($signed(reg397) || reg414)} : reg384[(1'h0):(1'h0)]);
                      reg435 <= ($signed(reg387) - (^~$unsigned((-wire339))));
                      reg436 <= reg384;
                    end
                  if ($unsigned($signed(({reg417} ?
                      $unsigned(reg395) : (!(8'haa))))))
                    begin
                      reg437 <= {reg382[(1'h0):(1'h0)]};
                    end
                  else
                    begin
                      reg437 <= reg383;
                      reg438 <= (($signed(reg405) ?
                              $signed(((8'haa) ?
                                  (8'haf) : (8'h9e))) : (-(forvar382 ?
                                  reg366 : (8'hac)))) ?
                          reg405 : forvar368);
                    end
                end
              else
                begin
                  if ((8'ha9))
                    begin
                      reg427 <= $signed($signed($signed(reg347[(1'h1):(1'h0)])));
                      reg428 <= {(^((forvar421 ^~ (8'hb2)) ?
                              $signed(forvar402) : reg390[(1'h1):(1'h1)]))};
                      reg429 <= $signed(forvar378[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg427 <= (reg417[(3'h7):(3'h4)] & $unsigned(forvar368));
                      reg428 <= $unsigned(((~|$signed(forvar386)) != (-reg352)));
                      reg429 <= (reg437 ?
                          $unsigned($unsigned(forvar388)) : {($signed((8'h9e)) ?
                                  reg363[(2'h2):(1'h0)] : $signed(reg412))});
                      reg430 <= ({$unsigned(reg360)} * {reg429});
                    end
                  for (forvar431 = (1'h0); (forvar431 < (1'h1)); forvar431 = (forvar431 + (1'h1)))
                    begin
                      reg432 <= forvar343;
                      reg433 <= (~^forvar388[(3'h5):(1'h0)]);
                    end
                end
              for (forvar439 = (1'h0); (forvar439 < (1'h0)); forvar439 = (forvar439 + (1'h1)))
                begin
                  for (forvar440 = (1'h0); (forvar440 < (2'h3)); forvar440 = (forvar440 + (1'h1)))
                    begin
                      reg441 <= reg405;
                      reg442 <= forvar396;
                      reg443 <= (reg437[(3'h5):(2'h2)] ?
                          $unsigned($signed(reg402)) : {$unsigned($signed(forvar431))});
                      reg444 <= forvar413[(2'h3):(1'h0)];
                    end
                  for (forvar445 = (1'h0); (forvar445 < (1'h0)); forvar445 = (forvar445 + (1'h1)))
                    begin
                      reg446 <= reg354[(1'h1):(1'h0)];
                      reg447 <= $unsigned(($unsigned($unsigned(reg408)) ~^ ((reg397 ~^ reg391) ^ {forvar388})));
                      reg448 <= (8'ha5);
                      reg449 <= $unsigned((-((|wire340) ?
                          reg447[(2'h3):(2'h3)] : (reg406 ? reg360 : reg409))));
                    end
                  for (forvar450 = (1'h0); (forvar450 < (2'h3)); forvar450 = (forvar450 + (1'h1)))
                    begin
                      reg451 <= (~^$unsigned($unsigned(reg357)));
                      reg452 <= ($signed(((forvar388 && reg357) <= reg406[(1'h1):(1'h1)])) ?
                          $signed(forvar445) : {{reg382[(2'h3):(1'h1)]}});
                    end
                end
              for (forvar453 = (1'h0); (forvar453 < (2'h2)); forvar453 = (forvar453 + (1'h1)))
                begin
                  if ({(&{(forvar382 ? forvar362 : forvar361)})})
                    begin
                      reg454 <= reg411[(1'h1):(1'h1)];
                      reg455 <= reg429;
                      reg456 <= ((~forvar377[(1'h0):(1'h0)]) < $signed($unsigned(reg425)));
                    end
                  else
                    begin
                      reg454 <= (~^reg423[(1'h0):(1'h0)]);
                    end
                  for (forvar457 = (1'h0); (forvar457 < (1'h1)); forvar457 = (forvar457 + (1'h1)))
                    begin
                      reg458 <= $signed({reg456[(4'hb):(2'h3)]});
                      reg459 <= reg388;
                      reg460 <= ((&(^~(reg432 | reg397))) ?
                          reg410 : (~reg418[(4'he):(3'h7)]));
                      reg461 <= $unsigned($unsigned(({reg364} ?
                          (!reg347) : (forvar457 ? forvar355 : reg458))));
                    end
                  reg462 <= reg460[(2'h3):(1'h1)];
                  for (forvar463 = (1'h0); (forvar463 < (1'h1)); forvar463 = (forvar463 + (1'h1)))
                    begin
                      reg464 <= forvar463;
                      reg465 <= reg458[(3'h4):(1'h0)];
                      reg466 <= $unsigned((($unsigned((8'ha9)) < reg411) ?
                          {{reg350}} : ($signed(reg412) ^~ $signed((8'had)))));
                    end
                end
            end
        end
    end
  assign wire467 = $unsigned(reg444);
  assign wire468 = (~|$unsigned(reg454));
  always
    @(posedge clk) begin
      for (forvar469 = (1'h0); (forvar469 < (2'h3)); forvar469 = (forvar469 + (1'h1)))
        begin
          for (forvar470 = (1'h0); (forvar470 < (1'h0)); forvar470 = (forvar470 + (1'h1)))
            begin
              if ((8'haa))
                begin
                  reg471 <= $unsigned(wire468);
                end
              else
                begin
                  if ($unsigned(forvar381[(1'h0):(1'h0)]))
                    begin
                      reg471 <= $unsigned((reg444 - (~&(&reg349))));
                    end
                  else
                    begin
                      reg471 <= ($signed(forvar415[(2'h2):(2'h2)]) ?
                          forvar344 : $signed((^{reg409})));
                    end
                end
            end
          for (forvar472 = (1'h0); (forvar472 < (2'h3)); forvar472 = (forvar472 + (1'h1)))
            begin
              reg473 <= reg358;
              for (forvar474 = (1'h0); (forvar474 < (2'h2)); forvar474 = (forvar474 + (1'h1)))
                begin
                  if (({($unsigned((8'ha8)) ?
                          (forvar421 || reg399) : (reg434 ^~ forvar407))} ^~ (^$signed(wire339[(3'h6):(1'h1)]))))
                    begin
                      reg475 <= ((reg458 >= $unsigned((-forvar426))) << {reg394});
                      reg476 <= forvar405[(1'h1):(1'h0)];
                      reg477 <= forvar450;
                      reg478 <= $unsigned((forvar432[(3'h4):(1'h0)] ?
                          ((reg350 || reg385) ?
                              {reg373} : {forvar362}) : reg392));
                    end
                  else
                    begin
                      reg475 <= ((8'ha9) + $unsigned(((forvar463 >= reg387) ~^ forvar445[(1'h1):(1'h1)])));
                      reg476 <= (^$signed((-$signed(forvar395))));
                      reg477 <= $unsigned((&{$unsigned(reg447)}));
                    end
                end
              for (forvar479 = (1'h0); (forvar479 < (2'h3)); forvar479 = (forvar479 + (1'h1)))
                begin
                  for (forvar480 = (1'h0); (forvar480 < (2'h2)); forvar480 = (forvar480 + (1'h1)))
                    begin
                      reg481 <= ((!{$signed(forvar426)}) ?
                          ($signed((^~reg478)) ?
                              reg387[(4'hf):(4'hd)] : (((8'hb6) && reg436) ?
                                  (reg423 | reg389) : $unsigned(reg434))) : (8'ha8));
                      reg482 <= $signed(reg429[(4'hb):(1'h1)]);
                    end
                end
            end
          if ($unsigned(($unsigned($unsigned(reg422)) ?
              reg349[(3'h5):(3'h5)] : ($signed(reg376) <= (^(8'haa))))))
            begin
              reg483 <= $unsigned($unsigned((forvar385 ?
                  (~&reg414) : $unsigned(wire341))));
            end
          else
            begin
              if ($unsigned(reg462))
                begin
                  if ($unsigned($signed(({reg408} == forvar407))))
                    begin
                      reg483 <= (forvar389 ?
                          reg459[(4'ha):(1'h1)] : forvar393[(3'h7):(3'h5)]);
                      reg484 <= $unsigned((reg375[(1'h0):(1'h0)] ?
                          reg459 : reg350));
                      reg485 <= forvar346[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg483 <= (!$unsigned($signed((reg476 != reg477))));
                      reg484 <= $signed($unsigned($signed((~|reg414))));
                      reg485 <= $signed({$unsigned({(8'hb2)})});
                    end
                  if ($unsigned($signed(((forvar421 != (8'ha1)) + ((8'hb3) ^~ reg383)))))
                    begin
                      reg486 <= (~|(~|reg389[(2'h3):(1'h0)]));
                      reg487 <= ((!$signed(forvar393)) ?
                          (^~$unsigned({reg384})) : (({reg462} > $signed(reg449)) ?
                              $signed((reg433 ?
                                  forvar396 : reg422)) : $signed((forvar453 * reg387))));
                      reg488 <= reg370[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg486 <= reg406[(1'h1):(1'h1)];
                      reg487 <= ((&reg452[(4'h9):(3'h5)]) ?
                          (|((reg363 != forvar474) || (~&reg402))) : (forvar421[(3'h6):(1'h1)] ?
                              (^~(forvar344 ?
                                  forvar345 : forvar389)) : ((|(8'hb1)) <<< $signed((8'hb0)))));
                    end
                end
              else
                begin
                  if ((^~$signed($signed(forvar377[(2'h3):(1'h0)]))))
                    begin
                      reg483 <= $signed(($unsigned(reg452) <<< reg423));
                      reg484 <= reg389;
                    end
                  else
                    begin
                      reg483 <= $signed(($unsigned(reg406) ?
                          (forvar388 >>> wire341) : ((reg398 && reg360) ?
                              (forvar407 << forvar382) : reg430[(1'h1):(1'h0)])));
                    end
                  for (forvar485 = (1'h0); (forvar485 < (1'h1)); forvar485 = (forvar485 + (1'h1)))
                    begin
                      reg486 <= $signed($unsigned($signed(reg381[(2'h3):(1'h0)])));
                    end
                  for (forvar487 = (1'h0); (forvar487 < (2'h3)); forvar487 = (forvar487 + (1'h1)))
                    begin
                      reg488 <= ((+reg390[(3'h4):(2'h2)]) != reg389[(1'h0):(1'h0)]);
                      reg489 <= ((~|reg398) <<< (((reg392 ?
                          reg449 : (8'hac)) ^~ $signed((8'h9f))) == $signed(forvar404)));
                      reg490 <= reg484;
                      reg491 <= (&{($unsigned(reg379) ?
                              ((8'ha3) ^~ reg435) : (forvar344 ?
                                  reg357 : forvar413))});
                    end
                  if ((forvar453[(3'h6):(3'h6)] ?
                      ($signed({reg422}) << (reg397 >> $unsigned(forvar485))) : (~|forvar380[(3'h5):(2'h2)])))
                    begin
                      reg492 <= (($signed((~^(8'hb4))) ?
                              forvar485 : ($unsigned((8'hb5)) ?
                                  $signed(forvar348) : (forvar377 && reg374))) ?
                          ((~reg408[(1'h0):(1'h0)]) && $signed($unsigned(reg482))) : ({(forvar400 > reg458)} * ((reg409 | reg403) << (reg407 ?
                              reg379 : reg410))));
                      reg493 <= reg388[(3'h5):(1'h1)];
                      reg494 <= $signed($signed(($unsigned((8'ha8)) && reg451)));
                      reg495 <= forvar396;
                    end
                  else
                    begin
                      reg492 <= {$unsigned(((reg347 ?
                              forvar377 : (8'hb3)) && (reg417 >> reg462)))};
                    end
                end
              for (forvar496 = (1'h0); (forvar496 < (1'h1)); forvar496 = (forvar496 + (1'h1)))
                begin
                  for (forvar497 = (1'h0); (forvar497 < (1'h1)); forvar497 = (forvar497 + (1'h1)))
                    begin
                      reg498 <= $signed(forvar431[(3'h7):(3'h5)]);
                      reg499 <= ({(forvar463[(2'h3):(2'h3)] | reg451)} > $signed({$signed(reg403)}));
                    end
                  for (forvar500 = (1'h0); (forvar500 < (1'h0)); forvar500 = (forvar500 + (1'h1)))
                    begin
                      reg501 <= reg393[(2'h3):(1'h0)];
                    end
                end
              reg502 <= ((forvar487 ?
                      ({reg404} ?
                          forvar381[(2'h2):(1'h0)] : ((8'had) << reg350)) : ((~^forvar371) ?
                          $unsigned(reg373) : $signed(reg454))) ?
                  {(&(~^reg428))} : $unsigned(reg365[(1'h1):(1'h1)]));
            end
        end
      reg503 <= $unsigned(({(reg379 ? forvar453 : forvar348)} ?
          $signed((reg359 ? reg447 : reg411)) : {(reg358 ? reg423 : reg466)}));
    end
  assign wire504 = (~&(((reg449 | forvar396) >> (+(8'hb9))) ?
                       $unsigned((~|reg454)) : $signed(reg460)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module19
#( parameter param205 = (((((8'ha4) ? (8'hb2) : (8'hb9)) <<< ((8'ha0) ? (8'hba) : (8'had))) ? (((8'hb8) == (8'ha2)) && ((8'hb9) ? (8'had) : (8'ha6))) : (((8'hb4) & (8'hb4)) * ((8'ha6) ? (8'h9e) : (8'hb3)))) ? ((((8'hae) + (8'hb7)) == ((8'h9d) >>> (8'ha2))) > (((8'ha3) ? (8'h9f) : (8'h9c)) <<< ((8'ha0) ? (8'ha6) : (8'ha4)))) : ({((8'h9f) ? (8'haa) : (8'hb7))} ? (+(^~(8'ha3))) : ((-(8'ha5)) > ((8'ha2) ? (8'h9f) : (8'ha7))))) )
(y, clk, wire24, wire23, wire22, wire21, wire20);
  output wire [(32'h7bd):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire24;
  input wire signed [(3'h6):(1'h0)] wire23;
  input wire signed [(2'h2):(1'h0)] wire22;
  input wire [(4'hc):(1'h0)] wire21;
  input wire signed [(5'h10):(1'h0)] wire20;
  wire [(4'ha):(1'h0)] wire204;
  wire signed [(5'h10):(1'h0)] wire203;
  wire signed [(4'h9):(1'h0)] wire202;
  wire signed [(4'h9):(1'h0)] wire201;
  wire [(3'h7):(1'h0)] wire200;
  wire signed [(3'h7):(1'h0)] wire199;
  wire [(4'hd):(1'h0)] wire198;
  wire signed [(4'h9):(1'h0)] wire197;
  wire signed [(4'ha):(1'h0)] wire196;
  reg signed [(2'h2):(1'h0)] reg195 = (1'h0);
  reg [(5'h10):(1'h0)] reg194 = (1'h0);
  reg [(4'hf):(1'h0)] reg193 = (1'h0);
  reg [(3'h6):(1'h0)] reg192 = (1'h0);
  reg [(4'ha):(1'h0)] reg191 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg190 = (1'h0);
  reg [(4'h9):(1'h0)] forvar189 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg188 = (1'h0);
  reg [(2'h2):(1'h0)] forvar187 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar186 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg186 = (1'h0);
  reg [(2'h3):(1'h0)] reg185 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg184 = (1'h0);
  reg [(4'he):(1'h0)] reg183 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg182 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg180 = (1'h0);
  reg [(4'h9):(1'h0)] reg179 = (1'h0);
  reg [(4'h9):(1'h0)] reg178 = (1'h0);
  reg [(4'hd):(1'h0)] reg177 = (1'h0);
  reg [(3'h6):(1'h0)] forvar176 = (1'h0);
  reg [(4'hc):(1'h0)] forvar175 = (1'h0);
  reg [(4'hf):(1'h0)] forvar174 = (1'h0);
  reg [(2'h2):(1'h0)] forvar168 = (1'h0);
  reg [(3'h5):(1'h0)] forvar157 = (1'h0);
  reg [(4'hc):(1'h0)] reg171 = (1'h0);
  reg [(4'hd):(1'h0)] forvar170 = (1'h0);
  reg [(4'hb):(1'h0)] forvar166 = (1'h0);
  reg [(4'ha):(1'h0)] reg165 = (1'h0);
  reg [(3'h4):(1'h0)] forvar164 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg160 = (1'h0);
  reg [(2'h3):(1'h0)] forvar159 = (1'h0);
  reg [(4'hd):(1'h0)] reg154 = (1'h0);
  reg [(3'h5):(1'h0)] forvar150 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg143 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar142 = (1'h0);
  reg [(4'h8):(1'h0)] forvar139 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar138 = (1'h0);
  reg [(2'h2):(1'h0)] reg137 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar135 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg134 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar129 = (1'h0);
  reg [(4'hb):(1'h0)] reg128 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar127 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar117 = (1'h0);
  reg [(3'h7):(1'h0)] reg116 = (1'h0);
  reg [(3'h5):(1'h0)] forvar114 = (1'h0);
  reg [(3'h5):(1'h0)] forvar110 = (1'h0);
  reg signed [(4'he):(1'h0)] reg106 = (1'h0);
  reg [(4'he):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg175 = (1'h0);
  reg [(4'hf):(1'h0)] reg174 = (1'h0);
  reg [(3'h7):(1'h0)] reg173 = (1'h0);
  reg [(3'h6):(1'h0)] reg172 = (1'h0);
  reg [(2'h2):(1'h0)] forvar171 = (1'h0);
  reg [(3'h6):(1'h0)] reg170 = (1'h0);
  reg [(4'h8):(1'h0)] reg169 = (1'h0);
  reg [(4'ha):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg167 = (1'h0);
  reg [(4'hf):(1'h0)] reg166 = (1'h0);
  reg [(4'h8):(1'h0)] forvar165 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg164 = (1'h0);
  reg [(4'hd):(1'h0)] reg163 = (1'h0);
  reg [(5'h10):(1'h0)] reg162 = (1'h0);
  reg [(4'he):(1'h0)] reg161 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar160 = (1'h0);
  reg [(4'hd):(1'h0)] reg159 = (1'h0);
  reg [(4'he):(1'h0)] reg158 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg157 = (1'h0);
  reg [(4'ha):(1'h0)] reg156 = (1'h0);
  reg [(3'h6):(1'h0)] reg155 = (1'h0);
  reg [(4'ha):(1'h0)] forvar154 = (1'h0);
  reg [(4'hd):(1'h0)] reg153 = (1'h0);
  reg signed [(4'he):(1'h0)] reg152 = (1'h0);
  reg [(4'ha):(1'h0)] reg151 = (1'h0);
  reg [(3'h7):(1'h0)] reg150 = (1'h0);
  reg [(4'h8):(1'h0)] reg149 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg148 = (1'h0);
  reg [(4'hd):(1'h0)] reg147 = (1'h0);
  reg signed [(4'he):(1'h0)] reg146 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg145 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar144 = (1'h0);
  reg [(3'h5):(1'h0)] forvar143 = (1'h0);
  reg [(3'h6):(1'h0)] reg142 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg141 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg140 = (1'h0);
  reg [(4'he):(1'h0)] reg139 = (1'h0);
  reg [(4'hc):(1'h0)] reg138 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar137 = (1'h0);
  reg [(5'h10):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg135 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar134 = (1'h0);
  reg [(2'h3):(1'h0)] forvar133 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg132 = (1'h0);
  reg [(4'ha):(1'h0)] reg131 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg130 = (1'h0);
  reg [(4'h8):(1'h0)] reg129 = (1'h0);
  reg [(2'h3):(1'h0)] forvar128 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg127 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg126 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg125 = (1'h0);
  reg [(4'hc):(1'h0)] reg124 = (1'h0);
  reg [(3'h4):(1'h0)] reg123 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg122 = (1'h0);
  reg [(2'h2):(1'h0)] forvar121 = (1'h0);
  reg [(4'h9):(1'h0)] reg120 = (1'h0);
  reg [(2'h3):(1'h0)] reg119 = (1'h0);
  reg [(4'he):(1'h0)] forvar118 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg117 = (1'h0);
  reg [(3'h5):(1'h0)] forvar116 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg114 = (1'h0);
  reg [(3'h7):(1'h0)] reg113 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg112 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg111 = (1'h0);
  reg [(4'hd):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg108 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg107 = (1'h0);
  reg [(3'h7):(1'h0)] forvar106 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar105 = (1'h0);
  reg [(3'h4):(1'h0)] forvar99 = (1'h0);
  reg [(3'h4):(1'h0)] reg104 = (1'h0);
  reg [(2'h2):(1'h0)] reg103 = (1'h0);
  reg [(4'h9):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg101 = (1'h0);
  reg [(3'h6):(1'h0)] reg100 = (1'h0);
  reg [(2'h2):(1'h0)] reg99 = (1'h0);
  reg [(3'h7):(1'h0)] forvar98 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg83 = (1'h0);
  reg [(4'hc):(1'h0)] reg81 = (1'h0);
  reg [(2'h2):(1'h0)] forvar74 = (1'h0);
  reg [(3'h7):(1'h0)] forvar77 = (1'h0);
  reg [(4'hc):(1'h0)] reg76 = (1'h0);
  reg signed [(4'he):(1'h0)] reg72 = (1'h0);
  reg [(4'h9):(1'h0)] forvar64 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg97 = (1'h0);
  reg [(4'h8):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar95 = (1'h0);
  reg [(4'hb):(1'h0)] reg94 = (1'h0);
  reg [(2'h2):(1'h0)] reg93 = (1'h0);
  reg [(4'hf):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar91 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar90 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg89 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg88 = (1'h0);
  reg signed [(4'he):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg86 = (1'h0);
  reg [(4'h8):(1'h0)] reg85 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg84 = (1'h0);
  reg [(4'hc):(1'h0)] forvar83 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg82 = (1'h0);
  reg [(4'hd):(1'h0)] forvar81 = (1'h0);
  reg [(3'h7):(1'h0)] reg80 = (1'h0);
  reg [(3'h6):(1'h0)] reg79 = (1'h0);
  reg [(4'h9):(1'h0)] reg78 = (1'h0);
  reg [(4'ha):(1'h0)] reg77 = (1'h0);
  reg [(4'he):(1'h0)] forvar76 = (1'h0);
  reg [(3'h6):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg74 = (1'h0);
  reg [(4'ha):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar72 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg71 = (1'h0);
  reg [(4'ha):(1'h0)] reg70 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg69 = (1'h0);
  reg [(2'h2):(1'h0)] reg68 = (1'h0);
  reg [(4'hd):(1'h0)] reg67 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg65 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg64 = (1'h0);
  reg [(4'h9):(1'h0)] forvar63 = (1'h0);
  reg [(2'h2):(1'h0)] reg62 = (1'h0);
  reg signed [(4'he):(1'h0)] reg54 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg61 = (1'h0);
  reg [(4'h9):(1'h0)] reg60 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg59 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg58 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg57 = (1'h0);
  reg [(2'h3):(1'h0)] reg56 = (1'h0);
  reg [(4'hc):(1'h0)] reg55 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar54 = (1'h0);
  reg [(2'h3):(1'h0)] reg53 = (1'h0);
  reg [(4'hb):(1'h0)] reg52 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg51 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar50 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg49 = (1'h0);
  reg [(2'h2):(1'h0)] forvar48 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg42 = (1'h0);
  reg [(4'h8):(1'h0)] forvar41 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar39 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg44 = (1'h0);
  reg [(4'ha):(1'h0)] reg47 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg46 = (1'h0);
  reg [(4'h8):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar44 = (1'h0);
  reg [(2'h2):(1'h0)] reg43 = (1'h0);
  reg [(4'hf):(1'h0)] forvar42 = (1'h0);
  reg [(3'h5):(1'h0)] reg41 = (1'h0);
  reg [(2'h2):(1'h0)] reg40 = (1'h0);
  reg [(2'h3):(1'h0)] reg39 = (1'h0);
  reg [(2'h3):(1'h0)] reg38 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg37 = (1'h0);
  reg signed [(4'he):(1'h0)] reg36 = (1'h0);
  reg [(3'h6):(1'h0)] forvar35 = (1'h0);
  reg [(2'h3):(1'h0)] reg34 = (1'h0);
  reg [(2'h3):(1'h0)] reg33 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg32 = (1'h0);
  reg [(4'hd):(1'h0)] reg31 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg30 = (1'h0);
  reg [(3'h7):(1'h0)] reg29 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar27 = (1'h0);
  reg [(2'h3):(1'h0)] reg28 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg27 = (1'h0);
  reg [(4'hd):(1'h0)] forvar26 = (1'h0);
  reg [(4'h8):(1'h0)] reg25 = (1'h0);
  assign y = {wire204,
                 wire203,
                 wire202,
                 wire201,
                 wire200,
                 wire199,
                 wire198,
                 wire197,
                 wire196,
                 reg195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 forvar189,
                 reg188,
                 forvar187,
                 forvar186,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 forvar176,
                 forvar175,
                 forvar174,
                 forvar168,
                 forvar157,
                 reg171,
                 forvar170,
                 forvar166,
                 reg165,
                 forvar164,
                 reg160,
                 forvar159,
                 reg154,
                 forvar150,
                 reg144,
                 reg143,
                 forvar142,
                 forvar139,
                 forvar138,
                 reg137,
                 forvar135,
                 reg134,
                 reg133,
                 forvar129,
                 reg128,
                 forvar127,
                 reg118,
                 forvar117,
                 reg116,
                 forvar114,
                 forvar110,
                 reg106,
                 reg105,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 forvar171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 forvar165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 forvar160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 forvar154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 forvar144,
                 forvar143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 forvar137,
                 reg136,
                 reg135,
                 forvar134,
                 forvar133,
                 reg132,
                 reg131,
                 reg130,
                 reg129,
                 forvar128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 forvar121,
                 reg120,
                 reg119,
                 forvar118,
                 reg117,
                 forvar116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 forvar106,
                 forvar105,
                 forvar99,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 forvar98,
                 reg83,
                 reg81,
                 forvar74,
                 forvar77,
                 reg76,
                 reg72,
                 forvar64,
                 reg97,
                 reg96,
                 forvar95,
                 reg94,
                 reg93,
                 reg92,
                 forvar91,
                 forvar90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 forvar83,
                 reg82,
                 forvar81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 forvar76,
                 reg75,
                 reg74,
                 reg73,
                 forvar72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 forvar63,
                 reg62,
                 reg54,
                 reg61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 forvar54,
                 reg53,
                 reg52,
                 reg51,
                 forvar50,
                 reg49,
                 forvar48,
                 reg42,
                 forvar41,
                 forvar39,
                 reg44,
                 reg47,
                 reg46,
                 reg45,
                 forvar44,
                 reg43,
                 forvar42,
                 reg41,
                 reg40,
                 reg39,
                 reg38,
                 reg37,
                 reg36,
                 forvar35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 forvar27,
                 reg28,
                 reg27,
                 forvar26,
                 reg25,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg25 <= wire24;
      for (forvar26 = (1'h0); (forvar26 < (2'h2)); forvar26 = (forvar26 + (1'h1)))
        begin
          if ($signed(wire23))
            begin
              reg27 <= wire20[(2'h2):(1'h0)];
              reg28 <= (wire23 >>> ($unsigned(((8'h9f) ?
                  wire21 : (8'h9e))) > (~|$unsigned(reg25))));
            end
          else
            begin
              for (forvar27 = (1'h0); (forvar27 < (1'h0)); forvar27 = (forvar27 + (1'h1)))
                begin
                  if ($signed(wire22))
                    begin
                      reg28 <= $signed($signed(forvar27[(1'h1):(1'h0)]));
                      reg29 <= ((&((wire24 <<< forvar27) ?
                              (wire21 ?
                                  wire22 : wire20) : wire23[(3'h6):(3'h6)])) ?
                          (($unsigned(wire22) == (&reg28)) ?
                              ((reg25 >>> reg25) ?
                                  wire21 : (reg28 ^ reg25)) : wire21[(3'h4):(1'h0)]) : ($unsigned(((8'ha2) + wire22)) ^~ $unsigned(wire23[(1'h1):(1'h1)])));
                      reg30 <= forvar27[(2'h3):(2'h2)];
                      reg31 <= (!wire23);
                    end
                  else
                    begin
                      reg28 <= wire23[(2'h3):(2'h2)];
                    end
                  if ((forvar27 || ({$signed(reg29)} ?
                      $unsigned((wire24 ?
                          reg30 : wire23)) : ({forvar27} >= (reg28 - wire21)))))
                    begin
                      reg32 <= $signed($signed(($signed(wire23) ?
                          $signed(reg25) : (8'hb1))));
                      reg33 <= (((&reg29) < $unsigned((&wire22))) ^ $unsigned($unsigned(wire23)));
                      reg34 <= $unsigned($signed(($unsigned(reg27) ?
                          $signed((8'hae)) : {wire24})));
                    end
                  else
                    begin
                      reg32 <= (wire22 ?
                          ((8'haf) ?
                              (reg32 ?
                                  $unsigned(reg25) : reg27) : $unsigned((^~wire24))) : (|(~|reg31)));
                      reg33 <= (|(~&forvar27[(2'h2):(2'h2)]));
                    end
                end
              for (forvar35 = (1'h0); (forvar35 < (2'h3)); forvar35 = (forvar35 + (1'h1)))
                begin
                  reg36 <= $unsigned($unsigned((((8'ha3) || reg33) ?
                      $signed(wire23) : (wire22 || reg33))));
                end
              reg37 <= (reg31[(3'h6):(3'h5)] ?
                  $unsigned(($unsigned(reg28) != $signed(reg36))) : wire20[(4'hf):(3'h6)]);
              reg38 <= $unsigned(((!$unsigned(reg37)) <<< (reg27[(3'h4):(1'h1)] ?
                  (reg27 && reg29) : $signed(reg36))));
            end
          if (($signed(reg38[(2'h2):(1'h0)]) ? reg25 : $unsigned(reg29)))
            begin
              reg39 <= (+(~|reg25));
              reg40 <= ((((reg34 ? reg37 : (8'h9f)) <= wire24[(2'h3):(2'h2)]) ?
                  (~^reg27[(3'h4):(2'h2)]) : (reg36 ?
                      (wire21 && reg30) : (reg36 ?
                          forvar27 : forvar26))) >>> (reg33 <<< $signed((reg28 << reg27))));
              reg41 <= (8'hb6);
              if ((reg29 ?
                  $unsigned((wire20[(4'ha):(2'h3)] ?
                      ((8'hb4) <= reg28) : $signed((8'hac)))) : forvar26))
                begin
                  for (forvar42 = (1'h0); (forvar42 < (1'h1)); forvar42 = (forvar42 + (1'h1)))
                    begin
                      reg43 <= (~|(wire24[(2'h3):(1'h0)] * (-reg30)));
                    end
                  for (forvar44 = (1'h0); (forvar44 < (1'h0)); forvar44 = (forvar44 + (1'h1)))
                    begin
                      reg45 <= wire20[(1'h1):(1'h1)];
                    end
                  if ($signed(reg29[(2'h2):(2'h2)]))
                    begin
                      reg46 <= $signed({$signed(reg33)});
                    end
                  else
                    begin
                      reg46 <= $unsigned((!{$signed(reg29)}));
                      reg47 <= reg36[(4'he):(4'h9)];
                    end
                end
              else
                begin
                  for (forvar42 = (1'h0); (forvar42 < (2'h2)); forvar42 = (forvar42 + (1'h1)))
                    begin
                      reg43 <= $unsigned(wire24);
                      reg44 <= ($unsigned($signed((reg39 ?
                          (8'h9d) : wire20))) || (({reg27} * forvar44[(2'h3):(1'h1)]) ?
                          reg39 : ((!wire21) < $signed((8'hb7)))));
                      reg45 <= ((($signed(reg30) > (forvar42 || reg28)) >= wire24[(2'h3):(1'h0)]) ?
                          (!($unsigned(wire24) ?
                              (&forvar42) : $signed((8'ha3)))) : (!$unsigned($unsigned(forvar42))));
                    end
                  reg46 <= ($unsigned(reg38) - {(forvar42[(4'ha):(4'ha)] ?
                          (|reg25) : (reg44 && reg36))});
                end
            end
          else
            begin
              for (forvar39 = (1'h0); (forvar39 < (2'h2)); forvar39 = (forvar39 + (1'h1)))
                begin
                  reg40 <= ((+((!forvar26) + (reg25 ?
                      (8'h9f) : (8'ha6)))) >= ($unsigned((~&reg40)) ?
                      (wire24[(2'h2):(1'h0)] ?
                          {reg27} : $unsigned(wire21)) : forvar39));
                  for (forvar41 = (1'h0); (forvar41 < (2'h2)); forvar41 = (forvar41 + (1'h1)))
                    begin
                      reg42 <= {reg28[(2'h2):(2'h2)]};
                    end
                end
            end
          for (forvar48 = (1'h0); (forvar48 < (1'h0)); forvar48 = (forvar48 + (1'h1)))
            begin
              reg49 <= (forvar26[(3'h6):(2'h3)] ?
                  $signed((~reg28[(1'h1):(1'h0)])) : forvar42);
              for (forvar50 = (1'h0); (forvar50 < (1'h1)); forvar50 = (forvar50 + (1'h1)))
                begin
                  if ($unsigned({$unsigned($signed(reg39))}))
                    begin
                      reg51 <= $unsigned((~|{(forvar41 > (8'ha0))}));
                      reg52 <= $unsigned(reg36);
                      reg53 <= (reg27[(3'h6):(3'h6)] * $unsigned(($signed(reg44) + ((8'ha4) ?
                          (8'hb9) : reg51))));
                    end
                  else
                    begin
                      reg51 <= (reg47[(2'h2):(2'h2)] ?
                          $unsigned((!reg31)) : (~&reg52[(4'ha):(1'h1)]));
                    end
                end
              if ((~&($signed(reg31[(4'h8):(3'h4)]) > ((+forvar42) * (~reg31)))))
                begin
                  for (forvar54 = (1'h0); (forvar54 < (2'h3)); forvar54 = (forvar54 + (1'h1)))
                    begin
                      reg55 <= (^reg49);
                      reg56 <= wire22;
                      reg57 <= $unsigned($unsigned(($signed((8'hab)) << $signed(reg29))));
                    end
                  if ({(((~|forvar50) + $signed(forvar35)) == reg32[(1'h1):(1'h0)])})
                    begin
                      reg58 <= $unsigned((wire21[(4'h8):(1'h1)] ?
                          forvar27 : {(|reg28)}));
                    end
                  else
                    begin
                      reg58 <= ($signed(reg29) ?
                          ((reg47[(3'h4):(1'h0)] ?
                              $signed(reg56) : (~|reg44)) <= ($unsigned(reg58) ?
                              forvar42 : (^reg28))) : (forvar41[(3'h7):(1'h0)] ?
                              ($signed(reg34) ?
                                  (!forvar42) : (~^wire24)) : (-(reg49 | forvar26))));
                      reg59 <= $signed(reg29[(3'h6):(3'h4)]);
                      reg60 <= reg45[(4'h8):(2'h2)];
                      reg61 <= reg46[(3'h7):(3'h5)];
                    end
                end
              else
                begin
                  reg54 <= ({reg41} ?
                      ((~&$unsigned((8'had))) >>> $unsigned({reg60})) : $unsigned({(~&reg51)}));
                  if ((reg32[(2'h3):(2'h2)] || (^$signed((reg34 << reg41)))))
                    begin
                      reg55 <= (~|reg31[(4'ha):(1'h1)]);
                    end
                  else
                    begin
                      reg55 <= reg55;
                      reg56 <= (~|wire23);
                      reg57 <= $unsigned((reg33[(2'h2):(2'h2)] >= $signed($signed(reg46))));
                      reg58 <= (($unsigned({reg47}) ? reg53 : (^(~|reg42))) ?
                          reg42 : $signed(($unsigned(forvar41) >= (forvar39 ?
                              reg47 : (8'ha0)))));
                    end
                  if ($signed((forvar54 >= $signed($unsigned(reg49)))))
                    begin
                      reg59 <= reg37;
                      reg60 <= $signed($signed(((8'ha0) ?
                          (+reg59) : $signed(reg33))));
                    end
                  else
                    begin
                      reg59 <= (~&($signed((reg49 <<< reg29)) && $signed((forvar39 & reg31))));
                    end
                  reg61 <= reg37;
                end
              reg62 <= ($signed(reg45) == $signed({(8'h9f)}));
            end
          if ($unsigned($signed((!((8'hab) ? forvar27 : reg53)))))
            begin
              if ((($signed($signed(wire22)) ?
                  reg38[(2'h2):(1'h0)] : reg55) >> $unsigned((~|(reg54 ?
                  (8'h9f) : reg37)))))
                begin
                  for (forvar63 = (1'h0); (forvar63 < (1'h0)); forvar63 = (forvar63 + (1'h1)))
                    begin
                      reg64 <= reg34[(2'h3):(1'h1)];
                      reg65 <= ((+((!wire23) ~^ forvar48)) ?
                          forvar44 : ($unsigned($signed((8'ha7))) ?
                              {(reg25 >= (8'hb0))} : reg46));
                      reg66 <= forvar41;
                      reg67 <= (&(~&$signed({reg33})));
                    end
                  if ($signed((8'hb1)))
                    begin
                      reg68 <= {(^$signed(((8'ha9) ? reg37 : reg39)))};
                      reg69 <= (^~($unsigned((reg27 | forvar44)) >= $signed($unsigned(reg46))));
                      reg70 <= (reg68 ?
                          $signed($unsigned(reg46[(3'h6):(1'h1)])) : $unsigned($signed($signed(reg34))));
                    end
                  else
                    begin
                      reg68 <= (|$unsigned((-forvar39)));
                      reg69 <= $signed(((-reg37) ?
                          reg49[(1'h1):(1'h1)] : $unsigned((reg66 ?
                              reg65 : reg32))));
                      reg70 <= ($unsigned($unsigned((reg47 ?
                          reg51 : reg40))) || ($signed(reg65) ?
                          reg25[(1'h0):(1'h0)] : $unsigned((reg64 <<< forvar26))));
                      reg71 <= {(!forvar63)};
                    end
                end
              else
                begin
                  for (forvar63 = (1'h0); (forvar63 < (2'h2)); forvar63 = (forvar63 + (1'h1)))
                    begin
                      reg64 <= (|reg52);
                      reg65 <= (($unsigned((&reg61)) ?
                              reg27 : reg57[(3'h4):(3'h4)]) ?
                          (+(reg29 ^ $unsigned(reg71))) : reg61);
                      reg66 <= wire21[(4'h9):(3'h4)];
                    end
                  reg67 <= $signed(forvar42);
                  if (((^reg68[(1'h1):(1'h0)]) ? reg61 : reg66[(3'h4):(2'h2)]))
                    begin
                      reg68 <= wire20[(4'ha):(4'h9)];
                      reg69 <= (^~($signed({(8'hb0)}) ?
                          reg28[(1'h0):(1'h0)] : (~&(reg58 | reg47))));
                      reg70 <= $unsigned($unsigned(((forvar63 >>> forvar42) | reg42)));
                      reg71 <= $unsigned((|(8'hb5)));
                    end
                  else
                    begin
                      reg68 <= $unsigned((-((&reg43) <<< $signed(forvar44))));
                      reg69 <= (($signed((8'ha1)) ?
                              (~|(forvar39 & reg47)) : ($unsigned(reg29) ?
                                  forvar50 : $signed((8'hb4)))) ?
                          reg43[(1'h0):(1'h0)] : $unsigned(((reg59 ^ (8'hac)) * reg62[(1'h1):(1'h1)])));
                      reg70 <= forvar63;
                      reg71 <= (8'ha4);
                    end
                end
              for (forvar72 = (1'h0); (forvar72 < (2'h2)); forvar72 = (forvar72 + (1'h1)))
                begin
                  if ((&(({(8'hac)} ?
                      reg62[(1'h0):(1'h0)] : (forvar50 <= reg59)) && wire20)))
                    begin
                      reg73 <= reg27;
                      reg74 <= reg38[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg73 <= (-{reg71});
                      reg74 <= reg64;
                      reg75 <= wire20;
                    end
                  for (forvar76 = (1'h0); (forvar76 < (1'h0)); forvar76 = (forvar76 + (1'h1)))
                    begin
                      reg77 <= {$signed((8'hb9))};
                      reg78 <= $unsigned((-$signed(forvar39[(3'h5):(2'h3)])));
                      reg79 <= $signed(reg34[(2'h2):(2'h2)]);
                      reg80 <= $signed((+$unsigned($unsigned(wire20))));
                    end
                  for (forvar81 = (1'h0); (forvar81 < (2'h3)); forvar81 = (forvar81 + (1'h1)))
                    begin
                      reg82 <= (~|$unsigned({$signed(forvar35)}));
                    end
                end
              for (forvar83 = (1'h0); (forvar83 < (2'h3)); forvar83 = (forvar83 + (1'h1)))
                begin
                  reg84 <= reg82;
                  reg85 <= $signed($unsigned((reg77[(4'h8):(1'h1)] ?
                      reg53[(1'h1):(1'h0)] : wire20[(4'hb):(4'hb)])));
                  if (($unsigned((!$unsigned(reg60))) ?
                      ({reg34} ?
                          $unsigned($unsigned(forvar26)) : $signed($signed(reg64))) : (~($unsigned(reg62) ?
                          reg62[(1'h0):(1'h0)] : $signed(reg69)))))
                    begin
                      reg86 <= (reg85[(2'h2):(2'h2)] ?
                          wire24 : forvar44[(2'h3):(2'h2)]);
                      reg87 <= $signed((!$unsigned((forvar48 <= reg75))));
                      reg88 <= reg37[(1'h1):(1'h1)];
                      reg89 <= (forvar35[(1'h0):(1'h0)] << (~^reg55[(3'h7):(3'h7)]));
                    end
                  else
                    begin
                      reg86 <= $unsigned(((reg85 ?
                          (8'h9d) : $unsigned(forvar42)) << (-(reg84 ?
                          reg77 : reg87))));
                    end
                end
              for (forvar90 = (1'h0); (forvar90 < (2'h3)); forvar90 = (forvar90 + (1'h1)))
                begin
                  for (forvar91 = (1'h0); (forvar91 < (2'h2)); forvar91 = (forvar91 + (1'h1)))
                    begin
                      reg92 <= $signed({(|reg70[(1'h1):(1'h1)])});
                      reg93 <= $signed($signed((^~reg49)));
                      reg94 <= ($unsigned(reg79[(2'h2):(1'h1)]) & ($unsigned((forvar48 || reg25)) || {reg39[(1'h1):(1'h0)]}));
                    end
                  for (forvar95 = (1'h0); (forvar95 < (2'h3)); forvar95 = (forvar95 + (1'h1)))
                    begin
                      reg96 <= (~|$unsigned({$unsigned(reg69)}));
                      reg97 <= $unsigned($signed({$signed(reg45)}));
                    end
                end
            end
          else
            begin
              for (forvar63 = (1'h0); (forvar63 < (2'h2)); forvar63 = (forvar63 + (1'h1)))
                begin
                  for (forvar64 = (1'h0); (forvar64 < (2'h3)); forvar64 = (forvar64 + (1'h1)))
                    begin
                      reg65 <= (!($signed(reg61) ? (~|{(8'h9f)}) : wire21));
                      reg66 <= (forvar63 ?
                          (((8'ha7) ?
                                  $unsigned(forvar81) : $unsigned((8'h9d))) ?
                              forvar64[(2'h2):(1'h0)] : {$signed(reg38)}) : $unsigned(reg84[(2'h2):(1'h0)]));
                    end
                  if ($signed(((-$unsigned(forvar26)) <<< ({reg65} ^ (reg54 < forvar42)))))
                    begin
                      reg67 <= ({(-reg67[(3'h5):(2'h3)])} < reg58);
                      reg68 <= $unsigned({(reg74 - reg39)});
                      reg69 <= {{{(reg34 ? reg30 : reg73)}}};
                    end
                  else
                    begin
                      reg67 <= (^~reg43);
                      reg68 <= $signed($unsigned((-reg89)));
                      reg69 <= reg54;
                    end
                  reg70 <= reg25[(4'h8):(1'h0)];
                end
              reg71 <= reg66[(4'h9):(4'h8)];
              if ($unsigned($signed(forvar41[(3'h4):(2'h3)])))
                begin
                  if ((8'ha6))
                    begin
                      reg72 <= $unsigned($signed($unsigned(reg94)));
                      reg73 <= reg92[(3'h5):(3'h4)];
                      reg74 <= (8'ha2);
                      reg75 <= (reg64 || reg96[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg72 <= {(reg28[(1'h0):(1'h0)] ~^ $unsigned($unsigned(reg42)))};
                      reg73 <= reg80;
                    end
                  reg76 <= $signed(forvar95[(4'ha):(3'h7)]);
                  for (forvar77 = (1'h0); (forvar77 < (2'h2)); forvar77 = (forvar77 + (1'h1)))
                    begin
                      reg78 <= (!reg79);
                      reg79 <= ({($signed((8'h9e)) ^~ reg25)} == (-($unsigned(reg85) ?
                          {(8'ha7)} : (reg31 != reg70))));
                      reg80 <= $unsigned((8'hb1));
                    end
                end
              else
                begin
                  for (forvar72 = (1'h0); (forvar72 < (1'h0)); forvar72 = (forvar72 + (1'h1)))
                    begin
                      reg73 <= (((8'ha2) ? forvar64 : forvar77) ?
                          (reg31[(4'h8):(1'h0)] ~^ $signed({(8'ha0)})) : $unsigned({reg65[(2'h2):(1'h0)]}));
                    end
                  for (forvar74 = (1'h0); (forvar74 < (1'h0)); forvar74 = (forvar74 + (1'h1)))
                    begin
                      reg75 <= reg32;
                      reg76 <= (reg77 < (-$unsigned((reg42 >>> forvar76))));
                      reg77 <= $unsigned($unsigned((!((8'ha9) ?
                          (8'hac) : reg44))));
                    end
                  reg78 <= $signed(reg25);
                  if (reg54)
                    begin
                      reg79 <= reg28[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg79 <= ({(~&$unsigned(forvar27))} * reg88);
                      reg80 <= forvar95[(2'h2):(1'h1)];
                      reg81 <= ({$unsigned({reg36})} != reg61[(1'h1):(1'h0)]);
                      reg82 <= {reg27[(3'h6):(3'h6)]};
                    end
                end
              if ((reg92[(4'h8):(3'h6)] ? $signed((~^reg29)) : forvar81))
                begin
                  for (forvar83 = (1'h0); (forvar83 < (1'h0)); forvar83 = (forvar83 + (1'h1)))
                    begin
                      reg84 <= (forvar26 ? forvar74[(2'h2):(2'h2)] : reg27);
                      reg85 <= reg47;
                    end
                  reg86 <= (+reg93[(1'h0):(1'h0)]);
                  if ((~&{((-forvar76) ? $signed(reg25) : $signed((8'ha9)))}))
                    begin
                      reg87 <= (8'hb7);
                    end
                  else
                    begin
                      reg87 <= forvar77;
                      reg88 <= {$unsigned(((|reg46) | $signed((8'ha5))))};
                      reg89 <= $unsigned({($unsigned(reg33) > (^~reg40))});
                    end
                end
              else
                begin
                  if (((reg75 && ((reg73 << forvar74) ?
                      reg34 : reg40)) << (~|reg40[(1'h0):(1'h0)])))
                    begin
                      reg83 <= forvar76;
                      reg84 <= reg68[(2'h2):(2'h2)];
                      reg85 <= (&reg83[(1'h0):(1'h0)]);
                      reg86 <= reg34[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg83 <= ((reg86 ?
                          forvar95 : $signed(reg70[(4'h8):(1'h1)])) == forvar63[(4'h8):(2'h3)]);
                      reg84 <= $unsigned((forvar76[(4'ha):(1'h0)] >>> $signed($unsigned((8'h9e)))));
                    end
                end
            end
        end
      if ({reg59[(1'h0):(1'h0)]})
        begin
          for (forvar98 = (1'h0); (forvar98 < (1'h1)); forvar98 = (forvar98 + (1'h1)))
            begin
              if ((wire23 ?
                  {((reg42 - reg32) ?
                          (8'hb1) : ((8'ha2) - reg89))} : $signed(({reg36} ?
                      $signed(reg86) : reg49))))
                begin
                  if ((~$unsigned($unsigned(reg37))))
                    begin
                      reg99 <= forvar42[(4'hf):(3'h7)];
                      reg100 <= forvar90[(3'h6):(1'h1)];
                      reg101 <= $unsigned((8'ha4));
                    end
                  else
                    begin
                      reg99 <= reg32;
                      reg100 <= $unsigned(reg32[(3'h7):(1'h1)]);
                      reg101 <= (~^$unsigned($signed(reg68)));
                      reg102 <= {$signed($unsigned((+(8'haf))))};
                    end
                  if (($unsigned(((reg87 == reg33) || reg78)) >= ($unsigned($unsigned(reg66)) ?
                      (~|(^reg64)) : $unsigned((8'ha6)))))
                    begin
                      reg103 <= reg28;
                      reg104 <= $unsigned($signed(reg59[(3'h6):(1'h1)]));
                    end
                  else
                    begin
                      reg103 <= forvar64;
                    end
                end
              else
                begin
                  for (forvar99 = (1'h0); (forvar99 < (2'h3)); forvar99 = (forvar99 + (1'h1)))
                    begin
                      reg100 <= ($signed(({reg59} ?
                          (reg56 ?
                              forvar54 : wire21) : reg72[(4'h9):(3'h4)])) && $unsigned(reg75[(1'h1):(1'h0)]));
                    end
                end
              for (forvar105 = (1'h0); (forvar105 < (1'h0)); forvar105 = (forvar105 + (1'h1)))
                begin
                  for (forvar106 = (1'h0); (forvar106 < (2'h3)); forvar106 = (forvar106 + (1'h1)))
                    begin
                      reg107 <= (+reg47[(2'h3):(1'h0)]);
                      reg108 <= ((|forvar77[(1'h0):(1'h0)]) > reg38);
                      reg109 <= $signed((reg45[(4'h8):(3'h4)] ?
                          ((^(8'h9f)) >= (|reg65)) : reg61[(3'h4):(1'h1)]));
                      reg110 <= ({$signed(((8'ha3) & reg32))} >> $signed(reg34));
                    end
                  reg111 <= $unsigned((reg65 ?
                      $unsigned(reg81) : reg39[(1'h0):(1'h0)]));
                  if ((8'hb4))
                    begin
                      reg112 <= (&reg108);
                      reg113 <= forvar74;
                      reg114 <= reg45;
                      reg115 <= $unsigned((forvar64[(3'h7):(1'h1)] >> ((^reg53) ?
                          $signed(reg77) : {reg30})));
                    end
                  else
                    begin
                      reg112 <= {(~&reg73)};
                      reg113 <= reg85[(4'h8):(1'h1)];
                      reg114 <= $unsigned({(8'hba)});
                    end
                  for (forvar116 = (1'h0); (forvar116 < (2'h2)); forvar116 = (forvar116 + (1'h1)))
                    begin
                      reg117 <= (reg89[(3'h4):(3'h4)] <<< $unsigned({(^wire20)}));
                    end
                end
              for (forvar118 = (1'h0); (forvar118 < (1'h1)); forvar118 = (forvar118 + (1'h1)))
                begin
                  if ((~forvar74[(1'h1):(1'h1)]))
                    begin
                      reg119 <= reg51;
                      reg120 <= (((~reg110[(1'h0):(1'h0)]) ?
                          forvar26[(3'h6):(3'h5)] : ({reg77} && $signed(reg51))) + reg43);
                    end
                  else
                    begin
                      reg119 <= $unsigned(reg77[(4'h9):(3'h4)]);
                      reg120 <= $unsigned((reg65 ?
                          reg65[(2'h2):(1'h0)] : forvar42));
                    end
                  for (forvar121 = (1'h0); (forvar121 < (2'h2)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= (~^(^~((reg113 - reg93) ?
                          (!forvar26) : (reg115 == reg42))));
                      reg123 <= (8'ha3);
                      reg124 <= $unsigned((^((reg52 & reg68) > (reg34 ?
                          reg99 : reg86))));
                      reg125 <= reg64;
                    end
                  if ((^(^$unsigned((reg36 ~^ reg37)))))
                    begin
                      reg126 <= {reg82[(4'h8):(4'h8)]};
                      reg127 <= ((wire20[(3'h4):(3'h4)] >>> $signed($signed(forvar98))) ?
                          $signed((reg109 ?
                              (forvar106 ?
                                  reg65 : reg111) : $unsigned(reg124))) : reg117[(3'h6):(1'h1)]);
                    end
                  else
                    begin
                      reg126 <= (!$unsigned($unsigned((reg47 ?
                          reg102 : reg117))));
                      reg127 <= ($unsigned(($signed((8'hb0)) ^~ $unsigned(reg93))) ?
                          $unsigned(reg40) : reg42[(4'he):(4'h8)]);
                    end
                  for (forvar128 = (1'h0); (forvar128 < (2'h3)); forvar128 = (forvar128 + (1'h1)))
                    begin
                      reg129 <= ($unsigned($unsigned((-reg39))) ?
                          forvar39[(4'hb):(4'hb)] : ($signed($unsigned((8'ha8))) ?
                              $unsigned(reg92[(4'h9):(3'h6)]) : {$signed(reg30)}));
                      reg130 <= (|(^reg62[(2'h2):(1'h0)]));
                      reg131 <= (($unsigned(reg43) > (^~$unsigned(reg127))) ?
                          (~((+(8'ha5)) ^~ (reg110 ?
                              reg65 : forvar121))) : ({forvar63} >>> $unsigned($unsigned(reg73))));
                      reg132 <= $signed($unsigned({(-forvar41)}));
                    end
                end
            end
          for (forvar133 = (1'h0); (forvar133 < (1'h1)); forvar133 = (forvar133 + (1'h1)))
            begin
              for (forvar134 = (1'h0); (forvar134 < (2'h2)); forvar134 = (forvar134 + (1'h1)))
                begin
                  reg135 <= $signed(({reg97} <<< {(~reg130)}));
                  reg136 <= reg68;
                  for (forvar137 = (1'h0); (forvar137 < (1'h0)); forvar137 = (forvar137 + (1'h1)))
                    begin
                      reg138 <= (forvar137 ?
                          forvar27[(3'h6):(1'h0)] : (((reg122 ?
                                  reg125 : forvar128) < (reg67 & reg113)) ?
                              ((forvar81 ?
                                  reg47 : reg88) - (reg117 < wire21)) : (^$signed(reg100))));
                      reg139 <= $signed(((~&$unsigned(reg103)) >>> (-forvar77)));
                      reg140 <= $signed((((reg68 - forvar118) | $signed((8'ha2))) >>> reg82[(1'h0):(1'h0)]));
                    end
                  if (forvar74)
                    begin
                      reg141 <= (reg38 >> (^(reg83[(1'h1):(1'h1)] ?
                          $unsigned(reg125) : (reg136 ? reg74 : reg127))));
                      reg142 <= forvar81[(4'hd):(3'h4)];
                    end
                  else
                    begin
                      reg141 <= ($signed($unsigned($unsigned(reg107))) ?
                          ($unsigned((8'ha2)) - (&$signed((8'ha9)))) : {$signed((|reg44))});
                    end
                end
            end
          for (forvar143 = (1'h0); (forvar143 < (2'h3)); forvar143 = (forvar143 + (1'h1)))
            begin
              for (forvar144 = (1'h0); (forvar144 < (1'h1)); forvar144 = (forvar144 + (1'h1)))
                begin
                  if (forvar50[(3'h4):(2'h3)])
                    begin
                      reg145 <= (|$unsigned(($unsigned(reg61) ?
                          (-reg130) : ((8'ha9) <= reg131))));
                      reg146 <= (~&((forvar95 ^~ (8'ha8)) + (forvar74 <<< (reg25 ~^ reg77))));
                      reg147 <= (&($unsigned(forvar83) ?
                          forvar41 : (reg130 ?
                              ((8'hb1) & (8'ha6)) : $signed(forvar116))));
                      reg148 <= reg86;
                    end
                  else
                    begin
                      reg145 <= reg114[(4'hd):(3'h6)];
                      reg146 <= {$signed(wire20)};
                      reg147 <= (8'hb9);
                      reg148 <= (+$signed({(forvar64 + forvar121)}));
                    end
                  reg149 <= ($unsigned(({reg145} <<< (8'hb8))) ?
                      reg124[(3'h4):(1'h1)] : $signed(reg69[(1'h1):(1'h1)]));
                  if ((($unsigned((~|reg114)) ^~ (-$signed(reg47))) - reg54[(3'h7):(3'h4)]))
                    begin
                      reg150 <= ($unsigned(reg60) > {(&$signed(reg52))});
                      reg151 <= reg93;
                      reg152 <= $unsigned((|reg99[(1'h0):(1'h0)]));
                      reg153 <= $unsigned(((reg72 ? (!reg138) : reg127) ?
                          (reg61 * {reg47}) : (~(forvar83 == (8'hb1)))));
                    end
                  else
                    begin
                      reg150 <= ((-$unsigned($signed(forvar76))) ?
                          {$unsigned({forvar81})} : forvar76[(3'h7):(3'h6)]);
                      reg151 <= $signed({reg51[(4'h8):(3'h6)]});
                      reg152 <= reg25[(1'h0):(1'h0)];
                    end
                  for (forvar154 = (1'h0); (forvar154 < (2'h3)); forvar154 = (forvar154 + (1'h1)))
                    begin
                      reg155 <= reg83[(4'h9):(3'h5)];
                    end
                end
              if ((($signed($unsigned(reg59)) ?
                  $unsigned((~&reg27)) : reg117) < $unsigned(($unsigned(reg139) ?
                  reg34[(1'h0):(1'h0)] : $unsigned(reg53)))))
                begin
                  if (((-(reg146 ? (reg39 >= reg64) : $unsigned(reg37))) ?
                      {forvar81[(3'h7):(2'h3)]} : (!(^~(reg58 ?
                          (8'h9e) : (8'haf))))))
                    begin
                      reg156 <= $unsigned($signed($unsigned($unsigned(reg141))));
                      reg157 <= ({(~|(~reg61))} ?
                          reg34 : $signed(forvar121[(2'h2):(2'h2)]));
                      reg158 <= reg60;
                      reg159 <= (&$signed({$signed(reg94)}));
                    end
                  else
                    begin
                      reg156 <= reg96[(4'h8):(2'h3)];
                      reg157 <= reg140[(4'h8):(3'h6)];
                    end
                end
              else
                begin
                  reg156 <= (8'ha2);
                end
              if ((forvar76 ?
                  $signed($unsigned($unsigned(reg38))) : {$signed(reg140)}))
                begin
                  for (forvar160 = (1'h0); (forvar160 < (1'h0)); forvar160 = (forvar160 + (1'h1)))
                    begin
                      reg161 <= $unsigned((reg153[(4'hc):(3'h6)] ?
                          reg155 : $signed($signed(reg27))));
                      reg162 <= reg47[(2'h3):(1'h1)];
                      reg163 <= reg36;
                      reg164 <= (~|($signed(forvar134) ?
                          $unsigned($unsigned(reg52)) : $signed($signed(reg94))));
                    end
                end
              else
                begin
                  for (forvar160 = (1'h0); (forvar160 < (1'h1)); forvar160 = (forvar160 + (1'h1)))
                    begin
                      reg161 <= (|reg69[(2'h3):(2'h2)]);
                      reg162 <= $signed(forvar116[(2'h3):(1'h1)]);
                      reg163 <= (({reg104[(3'h4):(2'h3)]} ?
                          ((!reg75) ?
                              reg149 : ((8'hab) ?
                                  reg129 : reg83)) : (!$signed(forvar50))) ^ {forvar137[(3'h4):(1'h1)]});
                      reg164 <= (forvar90 >>> reg161[(3'h4):(1'h1)]);
                    end
                  for (forvar165 = (1'h0); (forvar165 < (2'h2)); forvar165 = (forvar165 + (1'h1)))
                    begin
                      reg166 <= $unsigned({$signed($signed(reg31))});
                    end
                  reg167 <= forvar72[(4'hd):(4'ha)];
                  if (reg129[(1'h0):(1'h0)])
                    begin
                      reg168 <= {$unsigned(($signed(reg103) ^ {reg76}))};
                      reg169 <= $unsigned(forvar99[(2'h2):(2'h2)]);
                      reg170 <= ($unsigned(reg25) ?
                          $signed($signed($signed(reg46))) : $unsigned(((-reg32) ?
                              $unsigned(reg32) : $signed(reg117))));
                    end
                  else
                    begin
                      reg168 <= reg114;
                      reg169 <= ($signed(forvar54) ?
                          $signed($signed(forvar42[(3'h4):(1'h0)])) : ($signed($unsigned(forvar105)) & reg51[(4'hd):(4'h9)]));
                      reg170 <= $unsigned((forvar98 ?
                          reg123 : (^(reg45 && reg73))));
                    end
                end
              for (forvar171 = (1'h0); (forvar171 < (1'h1)); forvar171 = (forvar171 + (1'h1)))
                begin
                  if ((($unsigned((reg41 ? reg79 : reg117)) != ((8'haa) ?
                      (reg146 ?
                          reg93 : reg166) : $unsigned(reg168))) || (-{(8'hb1)})))
                    begin
                      reg172 <= reg55[(1'h0):(1'h0)];
                      reg173 <= $signed($unsigned(($unsigned(reg83) + (reg82 || reg80))));
                      reg174 <= $signed({((forvar42 ? (8'hb9) : reg162) ?
                              $unsigned(forvar26) : forvar171[(1'h1):(1'h0)])});
                      reg175 <= $signed(((+(reg113 < (8'hb2))) != $unsigned($unsigned(reg152))));
                    end
                  else
                    begin
                      reg172 <= ($signed((^~$signed(reg30))) || $unsigned((~(~reg57))));
                      reg173 <= $unsigned($signed((~^$unsigned(reg130))));
                      reg174 <= ((wire24[(1'h1):(1'h0)] <= reg83[(4'h9):(2'h3)]) ?
                          $signed(($signed(reg94) != (reg101 ?
                              reg28 : reg163))) : reg93);
                    end
                end
            end
        end
      else
        begin
          for (forvar98 = (1'h0); (forvar98 < (1'h1)); forvar98 = (forvar98 + (1'h1)))
            begin
              for (forvar99 = (1'h0); (forvar99 < (2'h2)); forvar99 = (forvar99 + (1'h1)))
                begin
                  if ((forvar54[(3'h6):(3'h5)] ?
                      reg89 : ($unsigned($unsigned(reg89)) < ((forvar121 >>> reg167) ?
                          ((8'hb2) ?
                              forvar128 : forvar99) : (wire24 <= forvar50)))))
                    begin
                      reg100 <= ((($signed(reg153) >= (reg120 ?
                              reg119 : forvar64)) ?
                          (reg70[(2'h2):(2'h2)] > $signed(reg127)) : $signed(reg60[(3'h5):(1'h1)])) >= (^~(~&{forvar98})));
                      reg101 <= $signed((reg31 < $unsigned($signed(forvar121))));
                    end
                  else
                    begin
                      reg100 <= reg130[(3'h6):(3'h5)];
                      reg101 <= reg129[(2'h2):(2'h2)];
                      reg102 <= forvar165;
                      reg103 <= (($unsigned(reg161) >= (reg86[(3'h6):(3'h4)] & (reg108 - (8'hb5)))) ?
                          forvar116[(3'h5):(1'h0)] : reg112);
                    end
                  reg104 <= forvar95;
                  if ((|(reg30 ?
                      reg120[(3'h6):(2'h3)] : ($signed(reg81) * reg65[(2'h3):(1'h1)]))))
                    begin
                      reg105 <= $unsigned($unsigned((!{reg60})));
                    end
                  else
                    begin
                      reg105 <= forvar118;
                      reg106 <= (8'ha1);
                      reg107 <= forvar160[(1'h1):(1'h1)];
                      reg108 <= {$signed($signed($unsigned((8'hb4))))};
                    end
                end
              reg109 <= ($signed((~|(forvar121 >> forvar50))) && wire24[(4'h8):(3'h6)]);
              for (forvar110 = (1'h0); (forvar110 < (2'h2)); forvar110 = (forvar110 + (1'h1)))
                begin
                  if ((~|$unsigned((((8'haa) ? forvar72 : reg145) ?
                      {(8'hb4)} : (reg51 <<< reg96)))))
                    begin
                      reg111 <= (-{(reg150[(1'h1):(1'h1)] ?
                              $signed(wire23) : $signed(reg166))});
                      reg112 <= $signed(reg110[(2'h3):(1'h1)]);
                      reg113 <= ($unsigned((8'h9d)) ?
                          ({{reg25}} ?
                              $signed({(8'hb4)}) : (8'hae)) : ((^~reg105) ?
                              reg159 : (8'hba)));
                    end
                  else
                    begin
                      reg111 <= ((reg73 * (-reg82[(2'h3):(2'h3)])) || ($unsigned((8'hb1)) ?
                          {{reg173}} : {(~|reg84)}));
                    end
                  for (forvar114 = (1'h0); (forvar114 < (2'h2)); forvar114 = (forvar114 + (1'h1)))
                    begin
                      reg115 <= reg119;
                      reg116 <= $signed((~&{$signed(reg124)}));
                    end
                  for (forvar117 = (1'h0); (forvar117 < (1'h1)); forvar117 = (forvar117 + (1'h1)))
                    begin
                      reg118 <= (~&($unsigned($signed(forvar116)) + $unsigned((8'ha0))));
                      reg119 <= (forvar134 ?
                          {wire24} : $unsigned($signed((reg29 == forvar143))));
                      reg120 <= (forvar118 ~^ {forvar121});
                    end
                end
              if ({$unsigned({(forvar165 ? reg93 : reg161)})})
                begin
                  for (forvar121 = (1'h0); (forvar121 < (1'h1)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= forvar171;
                      reg123 <= ((^~forvar44) ?
                          reg109[(1'h0):(1'h0)] : reg132[(3'h6):(1'h0)]);
                      reg124 <= ((|$unsigned(reg97)) ?
                          $signed($unsigned(reg58)) : $signed((reg107 ?
                              ((8'h9d) ? reg53 : forvar72) : reg114)));
                      reg125 <= forvar54[(3'h6):(1'h1)];
                    end
                  reg126 <= forvar76;
                  for (forvar127 = (1'h0); (forvar127 < (1'h1)); forvar127 = (forvar127 + (1'h1)))
                    begin
                      reg128 <= ($unsigned($signed({reg68})) != {{$unsigned(reg42)}});
                    end
                end
              else
                begin
                  for (forvar121 = (1'h0); (forvar121 < (2'h2)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= forvar90;
                    end
                end
            end
          if ((((forvar90 ^~ (8'ha8)) > $unsigned((8'hb7))) ?
              {$signed((reg80 || reg97))} : $signed((&reg119[(2'h3):(1'h1)]))))
            begin
              if (reg80)
                begin
                  for (forvar129 = (1'h0); (forvar129 < (1'h0)); forvar129 = (forvar129 + (1'h1)))
                    begin
                      reg130 <= ($signed(forvar99) ~^ (forvar54 ^~ $signed(reg47)));
                      reg131 <= (forvar106 | {({(8'ha3)} ?
                              $unsigned(reg85) : $signed(reg99))});
                    end
                  if (forvar98)
                    begin
                      reg132 <= $unsigned($signed($unsigned(reg93[(2'h2):(2'h2)])));
                      reg133 <= (reg76[(4'h8):(3'h6)] ?
                          (($unsigned(reg57) || (reg147 ? reg79 : forvar95)) ?
                              $signed($unsigned(reg123)) : reg168[(3'h5):(3'h4)]) : reg123);
                      reg134 <= (~(({forvar26} ?
                          (reg88 | (8'ha3)) : reg173[(1'h0):(1'h0)]) < (~(&reg54))));
                    end
                  else
                    begin
                      reg132 <= (!{(reg31[(4'ha):(3'h6)] || reg122[(4'h8):(4'h8)])});
                      reg133 <= $signed($unsigned(reg93[(1'h1):(1'h0)]));
                    end
                  for (forvar135 = (1'h0); (forvar135 < (2'h3)); forvar135 = (forvar135 + (1'h1)))
                    begin
                      reg136 <= forvar117[(1'h1):(1'h0)];
                      reg137 <= ($unsigned({reg28}) >= $signed(((forvar160 >>> reg92) >> ((8'haa) << reg131))));
                    end
                end
              else
                begin
                  for (forvar129 = (1'h0); (forvar129 < (1'h1)); forvar129 = (forvar129 + (1'h1)))
                    begin
                      reg130 <= (+$unsigned((8'hb3)));
                    end
                  if (reg89)
                    begin
                      reg131 <= (8'ha6);
                    end
                  else
                    begin
                      reg131 <= ((+reg75[(2'h2):(1'h1)]) ?
                          (+(reg151[(3'h5):(3'h5)] ?
                              (reg148 | (8'ha1)) : $unsigned(reg169))) : reg105);
                      reg132 <= $unsigned($signed((&forvar54)));
                    end
                  for (forvar133 = (1'h0); (forvar133 < (1'h0)); forvar133 = (forvar133 + (1'h1)))
                    begin
                      reg134 <= ((($signed((8'ha9)) >>> (reg155 ?
                              reg33 : reg58)) ?
                          $signed(forvar26) : ((reg168 ?
                              reg96 : (8'h9c)) & (reg156 >>> reg32))) <<< (^~(reg89[(2'h2):(1'h1)] ?
                          (~&reg77) : $signed(reg106))));
                      reg135 <= (((forvar63 >> reg167[(5'h10):(4'hb)]) ?
                          reg32 : ({reg124} ?
                              (!reg40) : $unsigned(reg109))) <<< (((8'ha3) <= {reg88}) ^~ (reg138 ?
                          reg175 : reg172[(3'h6):(3'h4)])));
                    end
                end
              for (forvar138 = (1'h0); (forvar138 < (2'h3)); forvar138 = (forvar138 + (1'h1)))
                begin
                  for (forvar139 = (1'h0); (forvar139 < (1'h0)); forvar139 = (forvar139 + (1'h1)))
                    begin
                      reg140 <= $unsigned(reg36[(2'h3):(2'h2)]);
                    end
                end
              if (({$unsigned((8'hb1))} == (reg146 ?
                  (forvar116 ?
                      (reg28 > reg84) : $unsigned(forvar41)) : {(|reg137)})))
                begin
                  reg141 <= $unsigned(reg76[(4'hc):(3'h6)]);
                  for (forvar142 = (1'h0); (forvar142 < (1'h0)); forvar142 = (forvar142 + (1'h1)))
                    begin
                      reg143 <= ($unsigned($unsigned((forvar50 << reg106))) ?
                          (reg87[(1'h1):(1'h1)] ^ $unsigned($unsigned((8'hb2)))) : ((((8'ha3) < reg80) + (forvar144 ?
                              reg33 : reg92)) * (~^$unsigned(reg82))));
                    end
                  if (($signed($unsigned($unsigned(reg78))) ?
                      $unsigned((reg44 | $unsigned(forvar133))) : {($unsigned(forvar144) ?
                              (reg135 ^ reg92) : (reg56 >>> forvar72))}))
                    begin
                      reg144 <= $signed((((~&(8'ha2)) <<< (~^(8'hac))) + reg85[(3'h6):(2'h3)]));
                      reg145 <= (-$signed((8'ha8)));
                      reg146 <= ($signed($signed(reg27)) | $signed($unsigned((forvar127 < forvar127))));
                    end
                  else
                    begin
                      reg144 <= ((|reg173) ?
                          (~&reg147) : (^reg96[(3'h4):(2'h2)]));
                    end
                end
              else
                begin
                  if (reg89)
                    begin
                      reg141 <= reg112;
                      reg142 <= (reg71 ^ $unsigned($signed($unsigned(reg99))));
                      reg143 <= (&(!$unsigned((reg25 ? reg97 : reg138))));
                    end
                  else
                    begin
                      reg141 <= reg137;
                      reg142 <= reg119;
                      reg143 <= {(reg139 | (~&(reg69 <<< reg167)))};
                    end
                  for (forvar144 = (1'h0); (forvar144 < (1'h1)); forvar144 = (forvar144 + (1'h1)))
                    begin
                      reg145 <= reg97[(3'h5):(1'h0)];
                    end
                  if ($unsigned(({(reg62 || wire22)} | $unsigned((&reg67)))))
                    begin
                      reg146 <= (((^~reg97) >>> $unsigned(forvar50[(3'h7):(3'h7)])) || (forvar139[(1'h0):(1'h0)] ?
                          (8'hac) : $signed(forvar133)));
                      reg147 <= {(!reg29)};
                      reg148 <= reg34;
                      reg149 <= reg137[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg146 <= reg34;
                      reg147 <= (&$unsigned($signed((reg51 ~^ reg169))));
                    end
                end
            end
          else
            begin
              reg129 <= (|($signed((forvar44 ?
                  forvar105 : forvar77)) ~^ (^~(8'hba))));
            end
          if ($unsigned(reg99[(1'h0):(1'h0)]))
            begin
              for (forvar150 = (1'h0); (forvar150 < (1'h0)); forvar150 = (forvar150 + (1'h1)))
                begin
                  if (({{$unsigned(reg174)}} >>> $signed(reg57)))
                    begin
                      reg151 <= (reg38 ~^ $unsigned((((8'hb2) && reg58) ?
                          {reg56} : (~forvar137))));
                      reg152 <= reg166[(3'h6):(1'h0)];
                      reg153 <= wire22[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg151 <= reg175[(3'h4):(1'h1)];
                    end
                  reg154 <= $unsigned((~|reg68));
                  if ((-reg34[(1'h1):(1'h0)]))
                    begin
                      reg155 <= reg56;
                    end
                  else
                    begin
                      reg155 <= ($unsigned(reg71[(2'h3):(2'h2)]) ?
                          ($signed($signed((8'ha8))) ?
                              (^~$signed((8'ha5))) : $signed(reg79[(3'h6):(2'h3)])) : $unsigned($unsigned(forvar77[(3'h6):(2'h3)])));
                      reg156 <= forvar39;
                      reg157 <= (&((forvar121 | $signed(forvar118)) == ((wire21 ?
                              reg59 : reg69) ?
                          (forvar135 ? reg29 : (8'hb0)) : (forvar137 ?
                              reg28 : reg65))));
                      reg158 <= {(reg151[(2'h2):(1'h1)] ^ ($unsigned(reg64) << reg61))};
                    end
                end
              if ({reg120[(4'h9):(4'h8)]})
                begin
                  for (forvar159 = (1'h0); (forvar159 < (2'h2)); forvar159 = (forvar159 + (1'h1)))
                    begin
                      reg160 <= reg120[(4'h9):(3'h7)];
                      reg161 <= ($unsigned(($unsigned(forvar154) ?
                          $unsigned((8'hb9)) : ((8'haa) ?
                              reg104 : (8'haa)))) >>> $signed(reg135[(4'ha):(3'h7)]));
                      reg162 <= $signed(($signed((8'haf)) ^~ $unsigned(reg39)));
                      reg163 <= (($signed((|reg54)) ? reg37 : forvar83) ?
                          reg54[(4'h9):(3'h4)] : (($signed(reg169) ?
                                  {reg60} : $signed(reg49)) ?
                              $unsigned({reg102}) : reg29));
                    end
                  for (forvar164 = (1'h0); (forvar164 < (1'h0)); forvar164 = (forvar164 + (1'h1)))
                    begin
                      reg165 <= (reg119[(2'h3):(2'h3)] ^ reg61);
                    end
                  for (forvar166 = (1'h0); (forvar166 < (1'h1)); forvar166 = (forvar166 + (1'h1)))
                    begin
                      reg167 <= reg29;
                      reg168 <= reg131[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar159 = (1'h0); (forvar159 < (1'h0)); forvar159 = (forvar159 + (1'h1)))
                    begin
                      reg160 <= (reg140[(2'h3):(1'h0)] ?
                          $unsigned(forvar134) : {(~^forvar116[(3'h5):(3'h5)])});
                      reg161 <= (((~^{reg141}) ?
                          (~&(forvar159 ?
                              forvar133 : reg82)) : reg108[(2'h2):(1'h0)]) | $unsigned($unsigned($signed((8'ha8)))));
                      reg162 <= reg156;
                      reg163 <= (reg148 ?
                          $unsigned(((~reg119) ?
                              $unsigned(reg116) : (reg78 ?
                                  reg157 : reg46))) : (reg155[(3'h6):(3'h4)] && ((8'h9f) >= reg107[(2'h3):(1'h0)])));
                    end
                  reg164 <= reg27;
                  for (forvar165 = (1'h0); (forvar165 < (2'h2)); forvar165 = (forvar165 + (1'h1)))
                    begin
                      reg166 <= $signed(forvar166[(2'h3):(2'h3)]);
                      reg167 <= $signed($signed($unsigned(reg169[(4'h8):(1'h0)])));
                      reg168 <= reg30;
                      reg169 <= forvar54;
                    end
                  for (forvar170 = (1'h0); (forvar170 < (1'h1)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= $signed(forvar81[(3'h5):(3'h4)]);
                      reg172 <= reg162[(4'hc):(4'h9)];
                      reg173 <= reg170;
                    end
                end
            end
          else
            begin
              reg150 <= wire22;
              if (reg67[(3'h6):(1'h0)])
                begin
                  reg151 <= $signed($unsigned(reg171));
                  reg152 <= (!(8'ha4));
                  if ((~(|(8'h9d))))
                    begin
                      reg153 <= $signed($unsigned(reg62));
                      reg154 <= ((+(|$signed(reg122))) + $signed(($unsigned(reg164) * (!reg123))));
                    end
                  else
                    begin
                      reg153 <= {(reg112 ?
                              ($unsigned((8'h9d)) + ((8'h9e) == reg66)) : reg138[(4'h8):(1'h0)])};
                      reg154 <= ((8'h9d) << reg68);
                      reg155 <= $signed((8'ha1));
                      reg156 <= ((($signed(reg116) >> reg171[(2'h3):(1'h1)]) ?
                          $signed($signed(reg33)) : ((reg167 ~^ reg131) << (-reg69))) << forvar41);
                    end
                end
              else
                begin
                  if ($signed(((!(reg51 ?
                      reg126 : reg45)) < reg97[(2'h2):(1'h0)])))
                    begin
                      reg151 <= reg167[(4'hd):(4'h9)];
                      reg152 <= reg67;
                    end
                  else
                    begin
                      reg151 <= forvar160[(1'h1):(1'h1)];
                      reg152 <= (!($signed((reg126 << forvar81)) ?
                          reg136[(2'h2):(1'h1)] : reg122[(4'hf):(3'h5)]));
                      reg153 <= $unsigned((+$signed(((8'hb6) != reg103))));
                    end
                end
              if ((~reg102))
                begin
                  if ((-((reg119[(1'h1):(1'h0)] ?
                      forvar35 : (^~reg31)) <= reg138[(4'h8):(2'h2)])))
                    begin
                      reg157 <= (reg83 || ((-$unsigned(reg136)) & (reg148 ?
                          (wire21 ? wire20 : reg161) : $signed(forvar135))));
                      reg158 <= $signed($signed($signed($signed((8'hb5)))));
                      reg159 <= (-$unsigned($signed(reg76)));
                      reg160 <= $unsigned((reg160 ?
                          ($unsigned((8'ha5)) || $unsigned(reg34)) : reg49[(3'h4):(1'h0)]));
                    end
                  else
                    begin
                      reg157 <= $signed((($unsigned(reg61) ?
                              (~&reg166) : (reg92 != reg75)) ?
                          ((&forvar171) ?
                              $signed(reg40) : {(8'h9c)}) : ($signed(forvar129) ?
                              $unsigned(reg92) : reg115)));
                      reg158 <= (~|wire24);
                    end
                  if ((reg101 >= $unsigned(forvar98)))
                    begin
                      reg161 <= reg111;
                      reg162 <= forvar142;
                      reg163 <= {forvar165[(3'h4):(2'h2)]};
                      reg164 <= reg157;
                    end
                  else
                    begin
                      reg161 <= (~&(forvar116 * {reg40[(2'h2):(1'h0)]}));
                      reg162 <= (((&(reg47 ^ reg113)) ?
                          ($signed(reg151) ?
                              forvar164[(1'h0):(1'h0)] : (forvar98 ?
                                  reg83 : reg170)) : ((~|reg32) >>> (forvar26 ?
                              (8'ha7) : forvar116))) <<< ({$unsigned(reg75)} > (reg85[(3'h6):(3'h4)] ?
                          (reg153 ^ reg47) : (reg173 & reg163))));
                      reg163 <= {((+(^~reg88)) || (reg53 ?
                              wire22[(2'h2):(1'h1)] : $signed(reg150)))};
                    end
                  if ({$unsigned((~&(forvar110 ^~ reg68)))})
                    begin
                      reg165 <= forvar154[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg165 <= reg92;
                    end
                  if ((^forvar134))
                    begin
                      reg166 <= (8'ha6);
                      reg167 <= reg107;
                    end
                  else
                    begin
                      reg166 <= $signed(reg79[(3'h5):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar157 = (1'h0); (forvar157 < (2'h2)); forvar157 = (forvar157 + (1'h1)))
                    begin
                      reg158 <= (&forvar143[(1'h1):(1'h0)]);
                      reg159 <= (reg49[(3'h4):(1'h1)] & $signed({(!reg37)}));
                      reg160 <= ($unsigned((-$unsigned(reg105))) ?
                          (($signed(wire22) ?
                              (reg106 <= reg166) : $signed(forvar171)) || reg114[(4'ha):(4'ha)]) : ((~|wire22[(1'h0):(1'h0)]) && (+reg70[(4'ha):(3'h5)])));
                    end
                  reg161 <= (|{((^~(8'hb0)) ? (~&forvar137) : reg130)});
                  if ((~&(^~$signed({forvar166}))))
                    begin
                      reg162 <= reg143[(2'h3):(1'h1)];
                      reg163 <= (^~$unsigned(($signed((8'hb6)) ^~ $signed(forvar99))));
                      reg164 <= $signed((((~^reg53) ?
                              forvar129 : (reg37 ^~ forvar41)) ?
                          ($unsigned(reg119) <= $unsigned((8'hac))) : forvar91[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg162 <= {(((!reg107) ^ (+reg162)) ?
                              reg144[(1'h0):(1'h0)] : ((-reg65) | {forvar44}))};
                      reg163 <= $unsigned($signed(({forvar35} ^~ reg47[(3'h5):(2'h3)])));
                      reg164 <= $unsigned($unsigned(forvar134));
                    end
                end
              if ((~&reg71))
                begin
                  for (forvar168 = (1'h0); (forvar168 < (2'h3)); forvar168 = (forvar168 + (1'h1)))
                    begin
                      reg169 <= forvar121;
                    end
                  for (forvar170 = (1'h0); (forvar170 < (1'h1)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= (!$unsigned($signed((reg141 <<< reg126))));
                      reg172 <= reg78[(1'h0):(1'h0)];
                      reg173 <= $signed((^~forvar133));
                    end
                end
              else
                begin
                  for (forvar168 = (1'h0); (forvar168 < (1'h1)); forvar168 = (forvar168 + (1'h1)))
                    begin
                      reg169 <= $signed(reg108);
                    end
                  for (forvar170 = (1'h0); (forvar170 < (1'h0)); forvar170 = (forvar170 + (1'h1)))
                    begin
                      reg171 <= (($signed((reg149 == forvar133)) > {(reg40 || forvar81)}) >>> forvar26);
                      reg172 <= reg36[(2'h3):(2'h3)];
                    end
                end
            end
          for (forvar174 = (1'h0); (forvar174 < (1'h0)); forvar174 = (forvar174 + (1'h1)))
            begin
              for (forvar175 = (1'h0); (forvar175 < (2'h2)); forvar175 = (forvar175 + (1'h1)))
                begin
                  for (forvar176 = (1'h0); (forvar176 < (2'h3)); forvar176 = (forvar176 + (1'h1)))
                    begin
                      reg177 <= (reg61 ?
                          $signed($unsigned($signed(reg40))) : $signed({$unsigned(reg53)}));
                    end
                  if ($unsigned(reg111))
                    begin
                      reg178 <= (($signed($unsigned(reg81)) && $unsigned((~|reg46))) < $signed(($signed(forvar133) & (reg147 != forvar83))));
                    end
                  else
                    begin
                      reg178 <= $unsigned(reg172);
                      reg179 <= (((~^(~^reg167)) ^ (forvar76 ?
                              reg133 : $unsigned((8'ha8)))) ?
                          ($unsigned({reg39}) >> {reg32}) : $unsigned($unsigned(((8'ha2) && reg87))));
                      reg180 <= $unsigned({forvar63[(1'h0):(1'h0)]});
                    end
                  reg181 <= (8'ha1);
                  if ($unsigned($unsigned($signed((|forvar166)))))
                    begin
                      reg182 <= ($unsigned(($unsigned(reg94) ?
                          (~^reg156) : (-reg94))) << ($unsigned({reg46}) < reg150));
                    end
                  else
                    begin
                      reg182 <= (reg46 ?
                          $signed($signed($unsigned(reg112))) : $unsigned({{reg99}}));
                      reg183 <= $unsigned(reg163[(4'h9):(3'h5)]);
                      reg184 <= (^~(8'hb1));
                      reg185 <= $signed((^{$signed(reg134)}));
                    end
                end
            end
        end
      if ($unsigned(($signed((reg38 ? reg80 : (8'had))) ?
          $signed($signed(reg166)) : $unsigned(forvar157[(2'h3):(2'h2)]))))
        begin
          reg186 <= ($unsigned($signed($unsigned(reg49))) * (!reg73[(4'h8):(3'h6)]));
        end
      else
        begin
          for (forvar186 = (1'h0); (forvar186 < (2'h3)); forvar186 = (forvar186 + (1'h1)))
            begin
              for (forvar187 = (1'h0); (forvar187 < (1'h1)); forvar187 = (forvar187 + (1'h1)))
                begin
                  reg188 <= {((8'hb1) == reg47[(2'h3):(1'h0)])};
                  for (forvar189 = (1'h0); (forvar189 < (2'h3)); forvar189 = (forvar189 + (1'h1)))
                    begin
                      reg190 <= (reg163[(4'h9):(4'h9)] & (((8'hb4) ?
                              $unsigned(reg151) : $signed(reg120)) ?
                          ({reg105} < reg92[(4'h8):(3'h5)]) : (^~(reg84 ?
                              reg34 : (8'had)))));
                      reg191 <= forvar154;
                      reg192 <= ($signed((8'h9e)) && (reg123 ?
                          ($unsigned(reg180) | $unsigned(reg190)) : forvar164[(2'h2):(1'h0)]));
                      reg193 <= (((&wire20) ?
                              {(wire21 ~^ forvar171)} : {(reg161 ?
                                      reg32 : reg131)}) ?
                          (8'h9c) : $signed($unsigned((&forvar144))));
                    end
                end
              reg194 <= ({$unsigned((forvar41 == (8'hb2)))} <<< ((reg148[(1'h0):(1'h0)] ?
                  reg53 : (forvar186 ?
                      (8'hb1) : reg93)) >= $signed(reg135[(3'h7):(3'h6)])));
              reg195 <= $signed(reg104[(3'h4):(1'h0)]);
            end
        end
    end
  assign wire196 = reg146[(1'h1):(1'h1)];
  assign wire197 = ($unsigned(((reg195 ? reg109 : reg47) ?
                       $signed(reg94) : $signed(forvar121))) < {reg126});
  assign wire198 = ($unsigned((~&$signed(reg154))) ?
                       (^~reg169[(2'h2):(2'h2)]) : (~|$signed((~&reg120))));
  assign wire199 = $unsigned((!(|reg104[(1'h0):(1'h0)])));
  assign wire200 = (|$signed(((reg47 << reg185) ?
                       reg83[(3'h5):(3'h4)] : reg74)));
  assign wire201 = {((8'ha8) ?
                           ((~|forvar137) - (reg29 ^~ reg62)) : (-(~&reg67)))};
  assign wire202 = {$signed(reg116)};
  assign wire203 = $unsigned(reg192[(3'h4):(3'h4)]);
  assign wire204 = (8'hb5);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module675
#(parameter param7426 = (^~(~|((&(8'hba)) ? (^(8'hae)) : {(8'ha0)}))))
(y, clk, wire676, wire677, wire678, wire679);
  output wire [(32'h13ff):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire676;
  input wire signed [(3'h7):(1'h0)] wire677;
  input wire [(3'h7):(1'h0)] wire678;
  input wire [(4'he):(1'h0)] wire679;
  wire [(4'h8):(1'h0)] wire7425;
  wire [(2'h3):(1'h0)] wire7424;
  reg signed [(2'h2):(1'h0)] reg7420 = (1'h0);
  reg [(5'h10):(1'h0)] reg7416 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7423 = (1'h0);
  reg [(3'h7):(1'h0)] reg7422 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7421 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7420 = (1'h0);
  reg [(3'h7):(1'h0)] reg7419 = (1'h0);
  reg [(4'hb):(1'h0)] reg7418 = (1'h0);
  reg [(3'h6):(1'h0)] reg7417 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7416 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7415 = (1'h0);
  reg [(3'h5):(1'h0)] reg7414 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7413 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7412 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7411 = (1'h0);
  reg [(5'h10):(1'h0)] reg7410 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7409 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7408 = (1'h0);
  reg [(2'h2):(1'h0)] reg7407 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7406 = (1'h0);
  reg [(2'h2):(1'h0)] forvar7405 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7404 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7403 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7398 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7402 = (1'h0);
  reg [(4'hb):(1'h0)] reg7401 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7400 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7399 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7398 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7397 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7396 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7395 = (1'h0);
  reg [(3'h6):(1'h0)] reg7394 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7393 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7392 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7391 = (1'h0);
  reg [(4'ha):(1'h0)] reg7390 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7389 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7388 = (1'h0);
  reg [(4'hb):(1'h0)] reg7387 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7386 = (1'h0);
  reg [(4'he):(1'h0)] reg7385 = (1'h0);
  reg [(4'hc):(1'h0)] reg7384 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7383 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7382 = (1'h0);
  reg [(2'h3):(1'h0)] reg7381 = (1'h0);
  reg [(3'h6):(1'h0)] reg7380 = (1'h0);
  reg [(4'h9):(1'h0)] reg7379 = (1'h0);
  reg [(5'h10):(1'h0)] forvar7378 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7368 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7367 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7377 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7376 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7375 = (1'h0);
  reg [(5'h10):(1'h0)] reg7374 = (1'h0);
  reg [(2'h3):(1'h0)] reg7373 = (1'h0);
  reg [(3'h6):(1'h0)] reg7372 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7371 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7370 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7369 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7368 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar7367 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7366 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar7365 = (1'h0);
  reg [(4'hb):(1'h0)] reg7364 = (1'h0);
  wire [(5'h10):(1'h0)] wire7363;
  wire signed [(3'h7):(1'h0)] wire7362;
  reg [(4'hd):(1'h0)] reg7361 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7355 = (1'h0);
  reg [(2'h3):(1'h0)] reg7354 = (1'h0);
  reg [(3'h5):(1'h0)] reg7360 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7359 = (1'h0);
  reg [(3'h7):(1'h0)] reg7358 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7357 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7356 = (1'h0);
  reg [(3'h7):(1'h0)] reg7355 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7354 = (1'h0);
  reg [(4'hf):(1'h0)] reg7353 = (1'h0);
  reg [(4'ha):(1'h0)] reg7352 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7351 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7350 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7349 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7348 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7347 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7346 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7345 = (1'h0);
  reg [(4'h8):(1'h0)] reg7344 = (1'h0);
  reg [(4'hf):(1'h0)] reg7343 = (1'h0);
  reg [(4'he):(1'h0)] reg7342 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7341 = (1'h0);
  reg [(3'h5):(1'h0)] reg7340 = (1'h0);
  reg [(4'ha):(1'h0)] forvar7339 = (1'h0);
  reg [(2'h2):(1'h0)] reg7338 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7337 = (1'h0);
  reg [(3'h4):(1'h0)] reg7336 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar7335 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7334 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7333 = (1'h0);
  wire [(5'h10):(1'h0)] wire7331;
  wire signed [(4'h8):(1'h0)] wire4336;
  wire signed [(4'hc):(1'h0)] wire4335;
  reg signed [(3'h7):(1'h0)] reg4334 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4333 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4332 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4331 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4330 = (1'h0);
  reg [(3'h6):(1'h0)] reg4329 = (1'h0);
  reg [(4'he):(1'h0)] reg4328 = (1'h0);
  reg [(3'h5):(1'h0)] reg4327 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4324 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4316 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4311 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4308 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4307 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4296 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4326 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4322 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4321 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4320 = (1'h0);
  reg [(4'hb):(1'h0)] reg4318 = (1'h0);
  reg [(3'h6):(1'h0)] reg4325 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4324 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4323 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4322 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4321 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4320 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4319 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4318 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4317 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4316 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4315 = (1'h0);
  reg [(4'hb):(1'h0)] reg4305 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4304 = (1'h0);
  reg [(4'h9):(1'h0)] reg4299 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4298 = (1'h0);
  reg [(4'h8):(1'h0)] reg4295 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4314 = (1'h0);
  reg [(3'h6):(1'h0)] reg4313 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4312 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4311 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4310 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4309 = (1'h0);
  reg [(3'h4):(1'h0)] reg4308 = (1'h0);
  reg [(4'ha):(1'h0)] reg4307 = (1'h0);
  reg [(4'ha):(1'h0)] reg4306 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4305 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4304 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4303 = (1'h0);
  reg [(4'he):(1'h0)] reg4302 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4301 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4300 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4299 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4298 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4297 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4296 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4295 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4294 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4293 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4286 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4282 = (1'h0);
  reg [(4'ha):(1'h0)] reg4292 = (1'h0);
  reg [(4'h9):(1'h0)] reg4291 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4290 = (1'h0);
  reg [(5'h10):(1'h0)] reg4289 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4288 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4287 = (1'h0);
  reg [(4'ha):(1'h0)] reg4286 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4285 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4284 = (1'h0);
  reg [(4'he):(1'h0)] reg4283 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4282 = (1'h0);
  reg [(2'h2):(1'h0)] reg4281 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4280 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4279 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4278 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4277 = (1'h0);
  reg [(3'h5):(1'h0)] reg4276 = (1'h0);
  reg [(4'hf):(1'h0)] reg4275 = (1'h0);
  reg [(4'he):(1'h0)] reg4274 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4273 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4272 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4262 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4271 = (1'h0);
  reg [(4'hc):(1'h0)] reg4270 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4269 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4268 = (1'h0);
  reg [(4'ha):(1'h0)] reg4267 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4266 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4265 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4264 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4263 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4262 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4261 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4252 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4247 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4245 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4237 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4235 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4233 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4230 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4260 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4259 = (1'h0);
  reg [(5'h10):(1'h0)] reg4258 = (1'h0);
  reg [(2'h2):(1'h0)] reg4257 = (1'h0);
  reg [(3'h7):(1'h0)] reg4256 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4255 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4254 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4253 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4252 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4251 = (1'h0);
  reg [(2'h2):(1'h0)] reg4244 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4250 = (1'h0);
  reg [(4'hd):(1'h0)] reg4249 = (1'h0);
  reg [(3'h6):(1'h0)] reg4248 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4247 = (1'h0);
  reg [(4'hf):(1'h0)] reg4246 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4245 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4244 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4243 = (1'h0);
  reg [(3'h5):(1'h0)] reg4242 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4241 = (1'h0);
  reg [(4'h9):(1'h0)] reg4240 = (1'h0);
  reg [(3'h4):(1'h0)] reg4239 = (1'h0);
  reg [(4'hd):(1'h0)] reg4238 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4237 = (1'h0);
  reg [(5'h10):(1'h0)] reg4236 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4235 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4234 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4233 = (1'h0);
  reg [(4'hd):(1'h0)] reg4232 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4231 = (1'h0);
  reg [(3'h5):(1'h0)] reg4230 = (1'h0);
  reg [(4'he):(1'h0)] reg4229 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4228 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4227 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4226 = (1'h0);
  reg [(3'h5):(1'h0)] reg4183 = (1'h0);
  reg [(4'hc):(1'h0)] reg4216 = (1'h0);
  reg [(4'he):(1'h0)] reg4214 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4212 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4211 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4208 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4209 = (1'h0);
  reg [(4'h8):(1'h0)] reg4205 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4204 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4202 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4200 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4195 = (1'h0);
  reg [(4'he):(1'h0)] reg4191 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4187 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4172 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4225 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4224 = (1'h0);
  reg [(4'he):(1'h0)] reg4223 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4222 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4221 = (1'h0);
  reg [(2'h3):(1'h0)] reg4220 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4219 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4218 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4217 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4216 = (1'h0);
  reg [(5'h10):(1'h0)] reg4215 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4214 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4198 = (1'h0);
  reg [(2'h3):(1'h0)] reg4213 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4212 = (1'h0);
  reg [(4'he):(1'h0)] reg4211 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4210 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4209 = (1'h0);
  reg [(3'h7):(1'h0)] reg4208 = (1'h0);
  reg [(4'ha):(1'h0)] reg4207 = (1'h0);
  reg [(4'hf):(1'h0)] reg4206 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4205 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4204 = (1'h0);
  reg [(5'h10):(1'h0)] reg4203 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4202 = (1'h0);
  reg [(4'h9):(1'h0)] reg4201 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4200 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4199 = (1'h0);
  reg [(3'h6):(1'h0)] reg4198 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4197 = (1'h0);
  reg [(3'h4):(1'h0)] reg4196 = (1'h0);
  reg [(3'h6):(1'h0)] reg4195 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4192 = (1'h0);
  reg [(4'hd):(1'h0)] reg4194 = (1'h0);
  reg [(2'h2):(1'h0)] reg4193 = (1'h0);
  reg [(5'h10):(1'h0)] reg4192 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4191 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4190 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4189 = (1'h0);
  reg [(4'h9):(1'h0)] reg4188 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4187 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4186 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4185 = (1'h0);
  reg [(4'hc):(1'h0)] reg4184 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4183 = (1'h0);
  reg [(4'h8):(1'h0)] reg4182 = (1'h0);
  reg [(4'he):(1'h0)] forvar4181 = (1'h0);
  reg [(4'hc):(1'h0)] reg4174 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4180 = (1'h0);
  reg [(4'he):(1'h0)] reg4179 = (1'h0);
  reg [(4'h8):(1'h0)] reg4178 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4177 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4176 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4175 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4174 = (1'h0);
  reg [(4'hc):(1'h0)] reg4173 = (1'h0);
  reg [(4'hd):(1'h0)] reg4172 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4171 = (1'h0);
  reg [(4'ha):(1'h0)] forvar680 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar681 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar682 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg683 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg684 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg685 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg686 = (1'h0);
  reg [(3'h4):(1'h0)] forvar687 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar688 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar689 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg690 = (1'h0);
  reg [(3'h7):(1'h0)] reg691 = (1'h0);
  reg [(4'hb):(1'h0)] reg692 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg693 = (1'h0);
  reg [(4'he):(1'h0)] reg694 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg695 = (1'h0);
  reg [(3'h4):(1'h0)] reg696 = (1'h0);
  reg [(2'h2):(1'h0)] reg697 = (1'h0);
  reg [(3'h7):(1'h0)] reg698 = (1'h0);
  reg [(3'h6):(1'h0)] reg699 = (1'h0);
  reg [(4'h8):(1'h0)] reg700 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg701 = (1'h0);
  reg [(3'h5):(1'h0)] forvar702 = (1'h0);
  reg [(5'h10):(1'h0)] reg703 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg704 = (1'h0);
  reg [(3'h5):(1'h0)] reg705 = (1'h0);
  reg [(4'hc):(1'h0)] reg702 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar706 = (1'h0);
  reg [(3'h4):(1'h0)] reg707 = (1'h0);
  reg signed [(4'he):(1'h0)] reg708 = (1'h0);
  reg [(4'hf):(1'h0)] reg709 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar710 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg711 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg712 = (1'h0);
  reg [(4'h9):(1'h0)] reg713 = (1'h0);
  reg [(4'h9):(1'h0)] reg714 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg715 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg716 = (1'h0);
  reg [(3'h7):(1'h0)] reg717 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg718 = (1'h0);
  reg [(3'h4):(1'h0)] reg719 = (1'h0);
  reg [(4'hf):(1'h0)] reg720 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg721 = (1'h0);
  reg [(4'hc):(1'h0)] reg722 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg723 = (1'h0);
  reg [(3'h4):(1'h0)] reg724 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg725 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar719 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar724 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg726 = (1'h0);
  reg [(4'hf):(1'h0)] reg727 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg728 = (1'h0);
  reg [(5'h10):(1'h0)] reg729 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar730 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg731 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg732 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg733 = (1'h0);
  reg [(4'hc):(1'h0)] reg734 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar734 = (1'h0);
  reg [(2'h3):(1'h0)] reg735 = (1'h0);
  reg [(4'hf):(1'h0)] reg736 = (1'h0);
  reg [(3'h7):(1'h0)] reg737 = (1'h0);
  reg [(4'hd):(1'h0)] forvar707 = (1'h0);
  reg [(4'ha):(1'h0)] forvar709 = (1'h0);
  reg [(3'h7):(1'h0)] reg710 = (1'h0);
  reg [(4'hf):(1'h0)] forvar711 = (1'h0);
  reg [(4'hf):(1'h0)] forvar712 = (1'h0);
  reg [(3'h6):(1'h0)] forvar718 = (1'h0);
  reg [(2'h3):(1'h0)] forvar726 = (1'h0);
  reg [(4'hd):(1'h0)] reg730 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar715 = (1'h0);
  reg [(4'hc):(1'h0)] forvar716 = (1'h0);
  reg [(3'h6):(1'h0)] forvar729 = (1'h0);
  reg [(3'h7):(1'h0)] forvar731 = (1'h0);
  reg [(2'h2):(1'h0)] forvar733 = (1'h0);
  reg [(4'hb):(1'h0)] reg738 = (1'h0);
  reg [(3'h5):(1'h0)] reg739 = (1'h0);
  reg [(3'h6):(1'h0)] reg740 = (1'h0);
  reg [(4'he):(1'h0)] reg741 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg742 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg743 = (1'h0);
  reg [(4'hb):(1'h0)] forvar735 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg744 = (1'h0);
  reg [(4'h8):(1'h0)] reg745 = (1'h0);
  reg [(3'h5):(1'h0)] reg746 = (1'h0);
  reg [(4'ha):(1'h0)] reg747 = (1'h0);
  reg [(4'hc):(1'h0)] reg748 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar749 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg750 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg751 = (1'h0);
  reg [(2'h2):(1'h0)] reg752 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg753 = (1'h0);
  reg [(2'h2):(1'h0)] forvar754 = (1'h0);
  reg [(4'hf):(1'h0)] reg755 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg756 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg757 = (1'h0);
  reg [(2'h2):(1'h0)] reg758 = (1'h0);
  reg [(4'h8):(1'h0)] reg759 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg760 = (1'h0);
  reg [(4'h9):(1'h0)] reg761 = (1'h0);
  reg [(3'h4):(1'h0)] reg762 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar763 = (1'h0);
  reg [(3'h4):(1'h0)] forvar764 = (1'h0);
  reg [(3'h5):(1'h0)] reg765 = (1'h0);
  reg [(4'he):(1'h0)] reg766 = (1'h0);
  reg [(4'hd):(1'h0)] reg767 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg768 = (1'h0);
  reg [(3'h5):(1'h0)] reg769 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar770 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg771 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg772 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar773 = (1'h0);
  reg [(2'h2):(1'h0)] reg774 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg775 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg776 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg777 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar767 = (1'h0);
  reg [(2'h2):(1'h0)] reg770 = (1'h0);
  reg [(3'h6):(1'h0)] reg773 = (1'h0);
  reg [(4'h9):(1'h0)] forvar778 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar779 = (1'h0);
  reg [(3'h6):(1'h0)] forvar780 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg781 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar782 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg783 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg784 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg785 = (1'h0);
  reg [(4'h9):(1'h0)] reg786 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg787 = (1'h0);
  reg [(3'h7):(1'h0)] reg788 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar789 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar790 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg791 = (1'h0);
  reg [(4'he):(1'h0)] forvar792 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg793 = (1'h0);
  reg [(3'h5):(1'h0)] reg794 = (1'h0);
  reg signed [(4'he):(1'h0)] reg795 = (1'h0);
  reg [(3'h4):(1'h0)] reg796 = (1'h0);
  reg signed [(4'he):(1'h0)] reg790 = (1'h0);
  reg [(4'he):(1'h0)] forvar797 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg798 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar799 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg800 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg801 = (1'h0);
  reg [(4'hf):(1'h0)] reg802 = (1'h0);
  reg [(4'hb):(1'h0)] forvar803 = (1'h0);
  reg [(2'h2):(1'h0)] reg804 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg805 = (1'h0);
  reg [(4'ha):(1'h0)] reg806 = (1'h0);
  reg [(4'he):(1'h0)] reg807 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg799 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar802 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg803 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar808 = (1'h0);
  reg [(3'h4):(1'h0)] forvar809 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg810 = (1'h0);
  reg [(4'ha):(1'h0)] reg811 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg812 = (1'h0);
  reg [(4'he):(1'h0)] reg813 = (1'h0);
  reg [(4'ha):(1'h0)] forvar814 = (1'h0);
  reg [(5'h10):(1'h0)] reg815 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg816 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg817 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg818 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg820 = (1'h0);
  reg [(2'h3):(1'h0)] reg821 = (1'h0);
  reg [(3'h5):(1'h0)] forvar822 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg823 = (1'h0);
  reg [(4'hd):(1'h0)] reg824 = (1'h0);
  reg [(3'h6):(1'h0)] reg825 = (1'h0);
  reg signed [(4'he):(1'h0)] reg826 = (1'h0);
  reg [(4'h8):(1'h0)] reg827 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg828 = (1'h0);
  reg [(2'h2):(1'h0)] forvar791 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg792 = (1'h0);
  reg [(5'h10):(1'h0)] reg797 = (1'h0);
  reg [(4'he):(1'h0)] forvar804 = (1'h0);
  reg [(3'h6):(1'h0)] reg808 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg809 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar812 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg814 = (1'h0);
  reg [(4'hd):(1'h0)] reg829 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar830 = (1'h0);
  reg [(4'ha):(1'h0)] reg831 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg832 = (1'h0);
  reg [(5'h10):(1'h0)] forvar829 = (1'h0);
  reg [(5'h10):(1'h0)] reg830 = (1'h0);
  reg [(4'hd):(1'h0)] forvar832 = (1'h0);
  reg [(4'hc):(1'h0)] reg833 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg834 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg835 = (1'h0);
  reg [(4'ha):(1'h0)] reg836 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar837 = (1'h0);
  reg [(2'h2):(1'h0)] forvar838 = (1'h0);
  reg [(4'hf):(1'h0)] reg839 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg840 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg841 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg842 = (1'h0);
  reg [(4'ha):(1'h0)] reg843 = (1'h0);
  reg [(3'h5):(1'h0)] reg844 = (1'h0);
  reg [(3'h6):(1'h0)] reg845 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg846 = (1'h0);
  reg [(4'hc):(1'h0)] forvar847 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg848 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar831 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg837 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg838 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar842 = (1'h0);
  reg [(4'h9):(1'h0)] forvar844 = (1'h0);
  reg [(4'he):(1'h0)] reg847 = (1'h0);
  reg [(2'h3):(1'h0)] forvar848 = (1'h0);
  reg [(4'hc):(1'h0)] reg849 = (1'h0);
  reg [(4'hf):(1'h0)] reg850 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg851 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg852 = (1'h0);
  reg [(4'hb):(1'h0)] reg853 = (1'h0);
  reg signed [(4'he):(1'h0)] reg854 = (1'h0);
  reg [(4'hf):(1'h0)] reg855 = (1'h0);
  reg [(3'h6):(1'h0)] reg856 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar852 = (1'h0);
  reg [(3'h4):(1'h0)] reg857 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg858 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar859 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar860 = (1'h0);
  reg [(3'h6):(1'h0)] reg861 = (1'h0);
  reg [(4'he):(1'h0)] reg862 = (1'h0);
  reg [(4'he):(1'h0)] reg863 = (1'h0);
  reg [(4'hc):(1'h0)] reg864 = (1'h0);
  reg [(3'h7):(1'h0)] reg865 = (1'h0);
  reg [(3'h7):(1'h0)] forvar866 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg867 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar868 = (1'h0);
  reg [(4'hf):(1'h0)] reg869 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar870 = (1'h0);
  reg [(2'h2):(1'h0)] reg871 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg872 = (1'h0);
  reg [(4'hd):(1'h0)] reg873 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar874 = (1'h0);
  reg [(3'h5):(1'h0)] forvar875 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg876 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg877 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg878 = (1'h0);
  reg [(3'h5):(1'h0)] forvar879 = (1'h0);
  reg [(4'h9):(1'h0)] reg880 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg881 = (1'h0);
  reg [(4'ha):(1'h0)] reg882 = (1'h0);
  reg [(4'hc):(1'h0)] reg883 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg884 = (1'h0);
  reg [(4'h9):(1'h0)] reg885 = (1'h0);
  reg [(4'h9):(1'h0)] reg886 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg887 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire4169;
  assign y = {wire7425,
                 wire7424,
                 reg7420,
                 reg7416,
                 reg7423,
                 reg7422,
                 reg7421,
                 forvar7420,
                 reg7419,
                 reg7418,
                 reg7417,
                 forvar7416,
                 reg7415,
                 reg7414,
                 reg7413,
                 reg7412,
                 reg7411,
                 reg7410,
                 reg7409,
                 forvar7408,
                 reg7407,
                 reg7406,
                 forvar7405,
                 forvar7404,
                 forvar7403,
                 reg7398,
                 reg7402,
                 reg7401,
                 reg7400,
                 reg7399,
                 forvar7398,
                 reg7397,
                 reg7396,
                 reg7395,
                 reg7394,
                 reg7393,
                 reg7392,
                 forvar7391,
                 reg7390,
                 reg7389,
                 reg7388,
                 reg7387,
                 forvar7386,
                 reg7385,
                 reg7384,
                 forvar7383,
                 reg7382,
                 reg7381,
                 reg7380,
                 reg7379,
                 forvar7378,
                 forvar7368,
                 reg7367,
                 reg7377,
                 reg7376,
                 reg7375,
                 reg7374,
                 reg7373,
                 reg7372,
                 forvar7371,
                 reg7370,
                 reg7369,
                 reg7368,
                 forvar7367,
                 forvar7366,
                 forvar7365,
                 reg7364,
                 wire7363,
                 wire7362,
                 reg7361,
                 forvar7355,
                 reg7354,
                 reg7360,
                 forvar7359,
                 reg7358,
                 reg7357,
                 reg7356,
                 reg7355,
                 forvar7354,
                 reg7353,
                 reg7352,
                 reg7351,
                 reg7350,
                 reg7349,
                 reg7348,
                 reg7347,
                 reg7346,
                 forvar7345,
                 reg7344,
                 reg7343,
                 reg7342,
                 forvar7341,
                 reg7340,
                 forvar7339,
                 reg7338,
                 reg7337,
                 reg7336,
                 forvar7335,
                 forvar7334,
                 forvar7333,
                 wire7331,
                 wire4336,
                 wire4335,
                 reg4334,
                 reg4333,
                 reg4332,
                 reg4331,
                 forvar4330,
                 reg4329,
                 reg4328,
                 reg4327,
                 forvar4324,
                 reg4316,
                 forvar4311,
                 forvar4308,
                 forvar4307,
                 forvar4296,
                 reg4326,
                 forvar4322,
                 forvar4321,
                 reg4320,
                 reg4318,
                 reg4325,
                 reg4324,
                 reg4323,
                 reg4322,
                 reg4321,
                 forvar4320,
                 reg4319,
                 forvar4318,
                 reg4317,
                 forvar4316,
                 forvar4315,
                 reg4305,
                 forvar4304,
                 reg4299,
                 reg4298,
                 reg4295,
                 reg4314,
                 reg4313,
                 reg4312,
                 reg4311,
                 reg4310,
                 forvar4309,
                 reg4308,
                 reg4307,
                 reg4306,
                 forvar4305,
                 reg4304,
                 reg4303,
                 reg4302,
                 reg4301,
                 reg4300,
                 forvar4299,
                 forvar4298,
                 reg4297,
                 reg4296,
                 forvar4295,
                 reg4294,
                 forvar4293,
                 forvar4286,
                 reg4285,
                 reg4282,
                 reg4292,
                 reg4291,
                 reg4290,
                 reg4289,
                 reg4288,
                 reg4287,
                 reg4286,
                 forvar4285,
                 reg4284,
                 reg4283,
                 forvar4282,
                 reg4281,
                 reg4280,
                 forvar4279,
                 reg4278,
                 forvar4277,
                 reg4276,
                 reg4275,
                 reg4274,
                 reg4273,
                 forvar4272,
                 forvar4262,
                 reg4271,
                 reg4270,
                 reg4269,
                 forvar4268,
                 reg4267,
                 forvar4266,
                 reg4265,
                 reg4264,
                 reg4263,
                 reg4262,
                 forvar4261,
                 reg4252,
                 forvar4247,
                 forvar4245,
                 forvar4237,
                 forvar4235,
                 reg4233,
                 forvar4230,
                 reg4260,
                 reg4259,
                 reg4258,
                 reg4257,
                 reg4256,
                 reg4255,
                 reg4254,
                 reg4253,
                 forvar4252,
                 reg4251,
                 reg4244,
                 reg4250,
                 reg4249,
                 reg4248,
                 reg4247,
                 reg4246,
                 reg4245,
                 forvar4244,
                 reg4243,
                 reg4242,
                 reg4241,
                 reg4240,
                 reg4239,
                 reg4238,
                 reg4237,
                 reg4236,
                 reg4235,
                 reg4234,
                 forvar4233,
                 reg4232,
                 reg4231,
                 reg4230,
                 reg4229,
                 forvar4228,
                 forvar4227,
                 forvar4226,
                 reg4183,
                 reg4216,
                 reg4214,
                 forvar4212,
                 forvar4211,
                 forvar4208,
                 reg4209,
                 reg4205,
                 reg4204,
                 reg4202,
                 forvar4200,
                 forvar4195,
                 reg4191,
                 forvar4187,
                 forvar4172,
                 reg4225,
                 reg4224,
                 reg4223,
                 reg4222,
                 reg4221,
                 reg4220,
                 reg4219,
                 reg4218,
                 reg4217,
                 forvar4216,
                 reg4215,
                 forvar4214,
                 forvar4198,
                 reg4213,
                 reg4212,
                 reg4211,
                 reg4210,
                 forvar4209,
                 reg4208,
                 reg4207,
                 reg4206,
                 forvar4205,
                 forvar4204,
                 reg4203,
                 forvar4202,
                 reg4201,
                 reg4200,
                 reg4199,
                 reg4198,
                 reg4197,
                 reg4196,
                 reg4195,
                 forvar4192,
                 reg4194,
                 reg4193,
                 reg4192,
                 forvar4191,
                 reg4190,
                 reg4189,
                 reg4188,
                 reg4187,
                 reg4186,
                 reg4185,
                 reg4184,
                 forvar4183,
                 reg4182,
                 forvar4181,
                 reg4174,
                 reg4180,
                 reg4179,
                 reg4178,
                 reg4177,
                 reg4176,
                 reg4175,
                 forvar4174,
                 reg4173,
                 reg4172,
                 forvar4171,
                 forvar680,
                 forvar681,
                 forvar682,
                 reg683,
                 reg684,
                 reg685,
                 reg686,
                 forvar687,
                 forvar688,
                 forvar689,
                 reg690,
                 reg691,
                 reg692,
                 reg693,
                 reg694,
                 reg695,
                 reg696,
                 reg697,
                 reg698,
                 reg699,
                 reg700,
                 reg701,
                 forvar702,
                 reg703,
                 reg704,
                 reg705,
                 reg702,
                 forvar706,
                 reg707,
                 reg708,
                 reg709,
                 forvar710,
                 reg711,
                 reg712,
                 reg713,
                 reg714,
                 reg715,
                 reg716,
                 reg717,
                 reg718,
                 reg719,
                 reg720,
                 reg721,
                 reg722,
                 reg723,
                 reg724,
                 reg725,
                 forvar719,
                 forvar724,
                 reg726,
                 reg727,
                 reg728,
                 reg729,
                 forvar730,
                 reg731,
                 reg732,
                 reg733,
                 reg734,
                 forvar734,
                 reg735,
                 reg736,
                 reg737,
                 forvar707,
                 forvar709,
                 reg710,
                 forvar711,
                 forvar712,
                 forvar718,
                 forvar726,
                 reg730,
                 forvar715,
                 forvar716,
                 forvar729,
                 forvar731,
                 forvar733,
                 reg738,
                 reg739,
                 reg740,
                 reg741,
                 reg742,
                 reg743,
                 forvar735,
                 reg744,
                 reg745,
                 reg746,
                 reg747,
                 reg748,
                 forvar749,
                 reg750,
                 reg751,
                 reg752,
                 reg753,
                 forvar754,
                 reg755,
                 reg756,
                 reg757,
                 reg758,
                 reg759,
                 reg760,
                 reg761,
                 reg762,
                 forvar763,
                 forvar764,
                 reg765,
                 reg766,
                 reg767,
                 reg768,
                 reg769,
                 forvar770,
                 reg771,
                 reg772,
                 forvar773,
                 reg774,
                 reg775,
                 reg776,
                 reg777,
                 forvar767,
                 reg770,
                 reg773,
                 forvar778,
                 forvar779,
                 forvar780,
                 reg781,
                 forvar782,
                 reg783,
                 reg784,
                 reg785,
                 reg786,
                 reg787,
                 reg788,
                 forvar789,
                 forvar790,
                 reg791,
                 forvar792,
                 reg793,
                 reg794,
                 reg795,
                 reg796,
                 reg790,
                 forvar797,
                 reg798,
                 forvar799,
                 reg800,
                 reg801,
                 reg802,
                 forvar803,
                 reg804,
                 reg805,
                 reg806,
                 reg807,
                 reg799,
                 forvar802,
                 reg803,
                 forvar808,
                 forvar809,
                 reg810,
                 reg811,
                 reg812,
                 reg813,
                 forvar814,
                 reg815,
                 reg816,
                 reg817,
                 reg818,
                 reg819,
                 reg820,
                 reg821,
                 forvar822,
                 reg823,
                 reg824,
                 reg825,
                 reg826,
                 reg827,
                 reg828,
                 forvar791,
                 reg792,
                 reg797,
                 forvar804,
                 reg808,
                 reg809,
                 forvar812,
                 reg814,
                 reg829,
                 forvar830,
                 reg831,
                 reg832,
                 forvar829,
                 reg830,
                 forvar832,
                 reg833,
                 reg834,
                 reg835,
                 reg836,
                 forvar837,
                 forvar838,
                 reg839,
                 reg840,
                 reg841,
                 reg842,
                 reg843,
                 reg844,
                 reg845,
                 reg846,
                 forvar847,
                 reg848,
                 forvar831,
                 reg837,
                 reg838,
                 forvar842,
                 forvar844,
                 reg847,
                 forvar848,
                 reg849,
                 reg850,
                 reg851,
                 reg852,
                 reg853,
                 reg854,
                 reg855,
                 reg856,
                 forvar852,
                 reg857,
                 reg858,
                 forvar859,
                 forvar860,
                 reg861,
                 reg862,
                 reg863,
                 reg864,
                 reg865,
                 forvar866,
                 reg867,
                 forvar868,
                 reg869,
                 forvar870,
                 reg871,
                 reg872,
                 reg873,
                 forvar874,
                 forvar875,
                 reg876,
                 reg877,
                 reg878,
                 forvar879,
                 reg880,
                 reg881,
                 reg882,
                 reg883,
                 reg884,
                 reg885,
                 reg886,
                 reg887,
                 wire4169,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar680 = (1'h0); (forvar680 < (2'h2)); forvar680 = (forvar680 + (1'h1)))
        begin
          for (forvar681 = (1'h0); (forvar681 < (2'h3)); forvar681 = (forvar681 + (1'h1)))
            begin
              if (wire679)
                begin
                  for (forvar682 = (1'h0); (forvar682 < (1'h0)); forvar682 = (forvar682 + (1'h1)))
                    begin
                      reg683 <= (+wire678);
                      reg684 <= $unsigned(wire678);
                    end
                end
              else
                begin
                  for (forvar682 = (1'h0); (forvar682 < (1'h0)); forvar682 = (forvar682 + (1'h1)))
                    begin
                      reg683 <= forvar681;
                      reg684 <= forvar680;
                    end
                  reg685 <= forvar680[(4'ha):(4'ha)];
                  if (($unsigned(reg684[(1'h1):(1'h0)]) < (^~wire676)))
                    begin
                      reg686 <= $unsigned({(forvar680 && wire678)});
                    end
                  else
                    begin
                      reg686 <= forvar681[(3'h6):(2'h2)];
                    end
                end
            end
          for (forvar687 = (1'h0); (forvar687 < (2'h3)); forvar687 = (forvar687 + (1'h1)))
            begin
              for (forvar688 = (1'h0); (forvar688 < (1'h1)); forvar688 = (forvar688 + (1'h1)))
                begin
                  for (forvar689 = (1'h0); (forvar689 < (2'h2)); forvar689 = (forvar689 + (1'h1)))
                    begin
                      reg690 <= {(reg683 ^~ ($unsigned(forvar688) ?
                              $signed(forvar680) : $signed((8'ha0))))};
                      reg691 <= $unsigned({(~|$unsigned(reg685))});
                      reg692 <= $signed(((forvar689[(2'h2):(1'h0)] ~^ (reg690 ?
                              forvar681 : wire677)) ?
                          $unsigned({reg686}) : {wire679[(4'hd):(3'h6)]}));
                      reg693 <= reg692[(4'ha):(2'h3)];
                    end
                  if (forvar680)
                    begin
                      reg694 <= reg693;
                    end
                  else
                    begin
                      reg694 <= {(((forvar687 ? reg692 : reg685) ?
                              $signed(reg692) : (~|wire678)) ^~ $unsigned(forvar688))};
                      reg695 <= (forvar689 ?
                          $unsigned(((reg693 <<< forvar680) ?
                              (reg685 < reg684) : (8'h9c))) : ((|(reg686 >= reg683)) < {$signed(wire678)}));
                    end
                  if (reg693[(3'h5):(1'h0)])
                    begin
                      reg696 <= forvar687;
                      reg697 <= (^~(&(wire676[(3'h7):(1'h1)] ?
                          $unsigned(reg686) : (forvar689 ? reg695 : reg684))));
                      reg698 <= ($signed((8'hba)) == $unsigned($signed({reg694})));
                    end
                  else
                    begin
                      reg696 <= ($signed((~|(forvar680 ^~ reg690))) ?
                          reg692 : $unsigned(($signed(reg685) ?
                              wire679 : {reg696})));
                      reg697 <= $unsigned((~$unsigned((reg694 >> (8'hb6)))));
                    end
                  if ((((&wire678) || $unsigned((forvar682 ~^ reg684))) ^~ (!reg696)))
                    begin
                      reg699 <= $signed((wire676[(3'h6):(1'h1)] ?
                          $signed((reg691 ? reg697 : (8'ha9))) : forvar681));
                      reg700 <= $signed({$signed((&forvar688))});
                    end
                  else
                    begin
                      reg699 <= ({(8'hb8)} || $unsigned(reg694));
                      reg700 <= reg691[(3'h5):(1'h1)];
                      reg701 <= (reg685 - ($unsigned(reg696) & $signed(reg683)));
                    end
                end
              if ($signed(wire677[(1'h1):(1'h1)]))
                begin
                  for (forvar702 = (1'h0); (forvar702 < (2'h2)); forvar702 = (forvar702 + (1'h1)))
                    begin
                      reg703 <= reg699[(3'h4):(1'h1)];
                      reg704 <= reg693[(4'ha):(2'h2)];
                    end
                  reg705 <= wire678[(1'h0):(1'h0)];
                end
              else
                begin
                  reg702 <= (({$unsigned(reg704)} ?
                      ($unsigned(wire678) >> $signed(reg685)) : $signed((^~reg698))) & (~|reg695[(3'h5):(3'h4)]));
                  if (((~^(((8'hac) ?
                      (8'hb8) : reg694) < (forvar681 >> reg686))) > $unsigned(((-(8'h9e)) ?
                      forvar680[(3'h6):(2'h2)] : wire676))))
                    begin
                      reg703 <= $signed(forvar681);
                      reg704 <= {(|$signed((reg704 ? reg695 : reg685)))};
                    end
                  else
                    begin
                      reg703 <= (wire679 ?
                          forvar702[(2'h2):(1'h1)] : $signed(reg685));
                    end
                end
            end
        end
      if (reg702[(3'h5):(1'h1)])
        begin
          if (reg696[(1'h1):(1'h1)])
            begin
              for (forvar706 = (1'h0); (forvar706 < (1'h1)); forvar706 = (forvar706 + (1'h1)))
                begin
                  if ($unsigned(({(~&reg686)} ?
                      forvar682 : (~|(reg701 | reg702)))))
                    begin
                      reg707 <= ($signed(((forvar688 && reg698) + (reg691 ~^ wire678))) < forvar680[(3'h7):(3'h5)]);
                      reg708 <= $signed(reg698[(1'h0):(1'h0)]);
                      reg709 <= wire679[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg707 <= wire679[(1'h1):(1'h1)];
                      reg708 <= $unsigned(($unsigned((wire677 ?
                              wire677 : reg701)) ?
                          (reg697[(1'h0):(1'h0)] != {reg693}) : {(+wire678)}));
                      reg709 <= forvar682[(1'h0):(1'h0)];
                    end
                  for (forvar710 = (1'h0); (forvar710 < (2'h3)); forvar710 = (forvar710 + (1'h1)))
                    begin
                      reg711 <= $unsigned(($unsigned((reg697 ?
                          forvar687 : reg693)) << ((8'ha3) ?
                          ((8'hb7) ?
                              (8'ha6) : reg686) : forvar706[(2'h3):(1'h1)])));
                      reg712 <= $unsigned($unsigned($signed((forvar681 ^ (8'hab)))));
                      reg713 <= reg683;
                      reg714 <= $signed($unsigned($signed(reg704)));
                    end
                  if (reg697[(1'h1):(1'h1)])
                    begin
                      reg715 <= (!$unsigned(($unsigned(reg693) ?
                          $unsigned((8'ha8)) : $signed(forvar688))));
                      reg716 <= $signed(reg686[(2'h2):(1'h0)]);
                      reg717 <= $unsigned(reg711);
                      reg718 <= {((!(&wire677)) ? (8'hb6) : reg699)};
                    end
                  else
                    begin
                      reg715 <= $unsigned($signed($unsigned(forvar702)));
                      reg716 <= $signed(reg707[(1'h0):(1'h0)]);
                    end
                end
              if (reg684)
                begin
                  if (forvar702)
                    begin
                      reg719 <= $unsigned(($unsigned((~&reg711)) || (reg703[(4'hd):(4'hd)] ?
                          reg713 : (reg691 & wire679))));
                      reg720 <= ((reg700[(3'h4):(3'h4)] ?
                              ((reg704 ? reg719 : (8'hb4)) ?
                                  reg714 : forvar688) : (8'hae)) ?
                          $unsigned((~^$signed(wire676))) : reg716);
                      reg721 <= reg700;
                      reg722 <= (^~(((reg711 ? (8'hae) : reg721) ?
                              (~reg705) : {reg683}) ?
                          reg715[(4'h8):(3'h4)] : reg717));
                    end
                  else
                    begin
                      reg719 <= {reg696};
                    end
                  if ((~^{$signed($signed((8'ha8)))}))
                    begin
                      reg723 <= reg708;
                      reg724 <= $unsigned({(reg683[(3'h6):(3'h5)] && (~&reg699))});
                    end
                  else
                    begin
                      reg723 <= ({((reg692 < reg683) ?
                                  (reg685 ?
                                      reg695 : reg711) : reg693[(4'ha):(3'h5)])} ?
                          $signed($signed(((8'hb2) ?
                              reg691 : wire678))) : $unsigned(reg708[(2'h3):(2'h3)]));
                    end
                  reg725 <= (~(($unsigned(reg702) ?
                      forvar687[(1'h0):(1'h0)] : $signed(reg718)) - (~^(reg686 ?
                      reg684 : wire677))));
                end
              else
                begin
                  for (forvar719 = (1'h0); (forvar719 < (2'h2)); forvar719 = (forvar719 + (1'h1)))
                    begin
                      reg720 <= $signed((~&reg698[(1'h1):(1'h0)]));
                      reg721 <= $unsigned((reg697 < forvar688));
                      reg722 <= wire678[(2'h3):(2'h3)];
                      reg723 <= (|$unsigned((^~(forvar689 - (8'ha1)))));
                    end
                  for (forvar724 = (1'h0); (forvar724 < (2'h3)); forvar724 = (forvar724 + (1'h1)))
                    begin
                      reg725 <= $signed(($signed((reg698 || reg719)) ?
                          ($unsigned(reg708) ?
                              {reg704} : reg705[(1'h0):(1'h0)]) : ((+(8'ha5)) - (reg714 ?
                              forvar719 : reg722))));
                      reg726 <= ((^~((reg720 - reg717) ?
                          $unsigned((8'hb5)) : reg690[(4'h8):(2'h2)])) != reg698);
                      reg727 <= (8'ha1);
                      reg728 <= $signed(reg690[(3'h4):(2'h3)]);
                    end
                  reg729 <= $unsigned((({(8'ha4)} ?
                      (8'hb6) : $unsigned((8'hab))) * reg701));
                  for (forvar730 = (1'h0); (forvar730 < (1'h0)); forvar730 = (forvar730 + (1'h1)))
                    begin
                      reg731 <= ((8'ha9) ? reg715 : (+reg707));
                      reg732 <= forvar719;
                    end
                end
              reg733 <= ((~&$unsigned((-reg719))) * (~^(forvar689[(2'h3):(2'h3)] || $unsigned(reg697))));
              if ($unsigned(($signed(reg728) ?
                  ((reg683 + (8'ha1)) ?
                      (reg728 ?
                          reg700 : wire676) : $unsigned(reg708)) : forvar706[(1'h0):(1'h0)])))
                begin
                  if (reg709)
                    begin
                      reg734 <= (^~(~&$unsigned(reg699[(3'h5):(3'h4)])));
                    end
                  else
                    begin
                      reg734 <= ($unsigned(reg684[(1'h1):(1'h0)]) ?
                          reg723[(3'h5):(3'h5)] : $unsigned($signed(reg684[(2'h3):(2'h2)])));
                    end
                end
              else
                begin
                  for (forvar734 = (1'h0); (forvar734 < (2'h2)); forvar734 = (forvar734 + (1'h1)))
                    begin
                      reg735 <= $unsigned((^~$signed((forvar687 & reg712))));
                      reg736 <= (reg709 << forvar680);
                      reg737 <= $signed($unsigned($signed((&(8'ha3)))));
                    end
                end
            end
          else
            begin
              for (forvar706 = (1'h0); (forvar706 < (1'h0)); forvar706 = (forvar706 + (1'h1)))
                begin
                  for (forvar707 = (1'h0); (forvar707 < (1'h1)); forvar707 = (forvar707 + (1'h1)))
                    begin
                      reg708 <= forvar706;
                    end
                  for (forvar709 = (1'h0); (forvar709 < (2'h3)); forvar709 = (forvar709 + (1'h1)))
                    begin
                      reg710 <= $unsigned(($unsigned((-reg694)) ?
                          (forvar724 <= forvar680) : reg711));
                    end
                end
              for (forvar711 = (1'h0); (forvar711 < (2'h3)); forvar711 = (forvar711 + (1'h1)))
                begin
                  for (forvar712 = (1'h0); (forvar712 < (2'h2)); forvar712 = (forvar712 + (1'h1)))
                    begin
                      reg713 <= (&forvar687);
                      reg714 <= $unsigned(((((8'haa) ?
                          forvar687 : reg726) << {reg733}) & ({reg708} ?
                          (reg692 && reg715) : (forvar709 + (8'hb2)))));
                      reg715 <= reg705;
                      reg716 <= $signed($unsigned(($unsigned(forvar724) >>> (reg686 ?
                          forvar724 : reg700))));
                    end
                  reg717 <= {{$signed((forvar710 ? forvar702 : (8'h9c)))}};
                end
              for (forvar718 = (1'h0); (forvar718 < (1'h1)); forvar718 = (forvar718 + (1'h1)))
                begin
                  for (forvar719 = (1'h0); (forvar719 < (1'h1)); forvar719 = (forvar719 + (1'h1)))
                    begin
                      reg720 <= reg712[(1'h0):(1'h0)];
                      reg721 <= (&reg709);
                    end
                  if ((+{$unsigned($unsigned((8'hb7)))}))
                    begin
                      reg722 <= (8'ha1);
                      reg723 <= ($signed(($signed(wire677) && $unsigned(reg733))) ?
                          (8'had) : reg690[(2'h2):(1'h1)]);
                      reg724 <= (8'had);
                      reg725 <= (reg717 != ($signed(reg709[(4'hc):(3'h4)]) ?
                          (8'hb9) : (+(forvar681 ? reg694 : reg690))));
                    end
                  else
                    begin
                      reg722 <= reg720[(3'h5):(2'h3)];
                      reg723 <= {((!(^reg733)) >= forvar718)};
                    end
                  for (forvar726 = (1'h0); (forvar726 < (2'h2)); forvar726 = (forvar726 + (1'h1)))
                    begin
                      reg727 <= (-reg732[(3'h5):(3'h5)]);
                      reg728 <= (((~&(reg727 <= forvar734)) && (~^$unsigned(reg726))) ~^ (((reg698 == forvar718) < $unsigned(forvar682)) | ($signed(reg725) & reg700[(3'h5):(1'h0)])));
                      reg729 <= $signed($signed(reg704));
                      reg730 <= $unsigned((!{{reg714}}));
                    end
                  if ({($signed(reg712[(1'h0):(1'h0)]) ?
                          {(forvar726 ^ (8'ha8))} : ((reg717 | forvar712) || (reg716 - reg728)))})
                    begin
                      reg731 <= ($unsigned(forvar730) ?
                          $signed(forvar719) : ($unsigned($signed(reg724)) ?
                              $unsigned(((8'ha9) ?
                                  forvar734 : reg718)) : ((reg686 ?
                                      reg730 : (8'hb5)) ?
                                  (~^reg703) : reg723[(1'h0):(1'h0)])));
                      reg732 <= (($signed($unsigned(forvar702)) ~^ ($signed(forvar718) && $signed(reg735))) + (((8'hb4) ?
                              (~&(8'ha3)) : (+reg726)) ?
                          (~(~^reg728)) : forvar724));
                    end
                  else
                    begin
                      reg731 <= ($signed(reg726[(1'h1):(1'h0)]) ^~ forvar724);
                    end
                end
            end
        end
      else
        begin
          if ((^~$unsigned($signed((wire677 ? reg691 : wire676)))))
            begin
              for (forvar706 = (1'h0); (forvar706 < (1'h1)); forvar706 = (forvar706 + (1'h1)))
                begin
                  for (forvar707 = (1'h0); (forvar707 < (1'h0)); forvar707 = (forvar707 + (1'h1)))
                    begin
                      reg708 <= $unsigned($unsigned(((!(8'ha6)) && $unsigned((8'ha3)))));
                      reg709 <= $signed(({reg705} - $signed(reg696)));
                    end
                  if ($unsigned(reg703))
                    begin
                      reg710 <= $unsigned((|(&forvar709[(4'h9):(4'h9)])));
                      reg711 <= (~|$signed(reg722));
                      reg712 <= $signed((((+reg728) ~^ (forvar718 <= forvar730)) ?
                          (forvar718 ?
                              $signed((8'h9d)) : (reg724 ?
                                  forvar710 : (8'hac))) : reg730[(4'h8):(3'h5)]));
                      reg713 <= (reg698 ^~ (reg723 ?
                          {$unsigned(forvar682)} : (8'ha4)));
                    end
                  else
                    begin
                      reg710 <= $unsigned({(^~(reg683 ? forvar711 : (8'hb0)))});
                      reg711 <= reg713;
                      reg712 <= {$unsigned($unsigned($unsigned(forvar711)))};
                      reg713 <= {forvar706};
                    end
                end
              reg714 <= reg698;
              for (forvar715 = (1'h0); (forvar715 < (1'h1)); forvar715 = (forvar715 + (1'h1)))
                begin
                  reg716 <= ((-reg735[(2'h2):(2'h2)]) && wire677);
                  if (forvar682)
                    begin
                      reg717 <= $signed((wire676[(2'h3):(2'h2)] ?
                          ({(8'had)} ?
                              (reg720 ? forvar709 : (8'ha1)) : (forvar712 ?
                                  reg725 : (8'ha3))) : $unsigned((+reg737))));
                    end
                  else
                    begin
                      reg717 <= (^~((forvar687[(2'h3):(1'h1)] - {(8'hab)}) ?
                          ((reg719 ?
                              (8'h9d) : reg718) && (reg686 && reg718)) : {(reg730 & reg707)}));
                      reg718 <= ({((^~(8'hb8)) << (forvar680 + (8'ha2)))} ?
                          (($signed(wire678) ^ {reg718}) ?
                              ((8'hb5) & (reg730 ^ reg712)) : wire679[(4'h8):(1'h0)]) : forvar724[(4'ha):(1'h1)]);
                    end
                  if ((^forvar718))
                    begin
                      reg719 <= {{reg692}};
                      reg720 <= (+$signed($signed((8'h9d))));
                      reg721 <= {reg737};
                      reg722 <= reg735;
                    end
                  else
                    begin
                      reg719 <= ((~^(^(reg725 ? reg729 : reg697))) ?
                          $unsigned(wire676[(1'h0):(1'h0)]) : $unsigned(({reg724} << ((8'h9e) ?
                              reg726 : forvar730))));
                      reg720 <= (reg735[(1'h0):(1'h0)] ?
                          reg684 : ($signed((reg710 ? reg715 : reg709)) ?
                              forvar734[(1'h1):(1'h0)] : forvar689[(2'h3):(1'h1)]));
                      reg721 <= (!reg724);
                      reg722 <= ($unsigned(((-forvar730) ~^ forvar702[(2'h2):(1'h0)])) <<< reg685);
                    end
                end
            end
          else
            begin
              for (forvar706 = (1'h0); (forvar706 < (2'h3)); forvar706 = (forvar706 + (1'h1)))
                begin
                  for (forvar707 = (1'h0); (forvar707 < (2'h2)); forvar707 = (forvar707 + (1'h1)))
                    begin
                      reg708 <= (~&forvar726[(2'h2):(1'h0)]);
                    end
                  if (reg716)
                    begin
                      reg709 <= $unsigned(((~&{reg710}) ?
                          ($signed((8'hb1)) & $signed(reg726)) : reg734));
                      reg710 <= $unsigned((({reg696} >= $signed(forvar709)) ?
                          $signed(reg691) : $signed($signed(reg722))));
                    end
                  else
                    begin
                      reg709 <= (~|{$unsigned(reg719)});
                      reg710 <= $signed((-((wire677 > reg719) ?
                          (forvar707 - forvar687) : $unsigned(reg690))));
                      reg711 <= ($unsigned($unsigned(reg712[(3'h4):(2'h2)])) || forvar724);
                    end
                  for (forvar712 = (1'h0); (forvar712 < (1'h1)); forvar712 = (forvar712 + (1'h1)))
                    begin
                      reg713 <= (|(^$signed((forvar712 ? wire676 : reg690))));
                      reg714 <= {(~|$signed($unsigned(reg733)))};
                      reg715 <= (~reg726[(1'h1):(1'h0)]);
                    end
                end
              for (forvar716 = (1'h0); (forvar716 < (2'h2)); forvar716 = (forvar716 + (1'h1)))
                begin
                  if ($unsigned((((reg703 ? (8'ha4) : (8'hb8)) ?
                          $unsigned(reg718) : (forvar718 ? reg719 : reg709)) ?
                      (((8'ha4) ? reg696 : (8'hb7)) ?
                          forvar711 : (reg719 ?
                              forvar709 : reg722)) : {(reg724 != reg708)})))
                    begin
                      reg717 <= (((&reg702) ?
                              reg714 : (reg735 ?
                                  reg702[(4'h9):(1'h1)] : reg732)) ?
                          $unsigned((reg711[(2'h2):(1'h1)] | (reg692 ?
                              reg691 : forvar702))) : (reg684[(1'h0):(1'h0)] + forvar730));
                      reg718 <= ({reg722[(4'h9):(3'h6)]} ? reg737 : (8'h9f));
                      reg719 <= (~&reg711);
                      reg720 <= (8'hae);
                    end
                  else
                    begin
                      reg717 <= reg684;
                      reg718 <= (forvar711 || reg734[(4'hb):(4'h9)]);
                      reg719 <= forvar689;
                      reg720 <= forvar707;
                    end
                  if (($unsigned(forvar724[(4'hb):(4'h8)]) ?
                      $signed($signed((forvar710 ?
                          reg726 : (8'hba)))) : forvar688))
                    begin
                      reg721 <= (~^$unsigned($unsigned($signed(reg735))));
                      reg722 <= reg701[(3'h4):(2'h3)];
                      reg723 <= $signed((({forvar716} ^ reg731[(4'ha):(4'h8)]) ?
                          reg701 : forvar719));
                    end
                  else
                    begin
                      reg721 <= (-((~$unsigned(forvar689)) << (-$unsigned(reg705))));
                      reg722 <= {(^~wire679[(2'h3):(1'h1)])};
                      reg723 <= reg692[(2'h2):(2'h2)];
                    end
                  for (forvar724 = (1'h0); (forvar724 < (2'h2)); forvar724 = (forvar724 + (1'h1)))
                    begin
                      reg725 <= {reg696};
                    end
                end
              if ($signed(reg702[(4'h9):(4'h8)]))
                begin
                  if ($signed($signed((^reg736[(4'h8):(2'h3)]))))
                    begin
                      reg726 <= $unsigned({(-wire677)});
                      reg727 <= ($unsigned((^reg731[(1'h1):(1'h1)])) <<< $signed(reg696));
                      reg728 <= reg737;
                    end
                  else
                    begin
                      reg726 <= ($unsigned((|$unsigned(reg710))) ?
                          reg735[(1'h1):(1'h1)] : $unsigned($signed(reg710)));
                      reg727 <= {$signed({(reg722 - (8'hae))})};
                    end
                  for (forvar729 = (1'h0); (forvar729 < (1'h1)); forvar729 = (forvar729 + (1'h1)))
                    begin
                      reg730 <= (8'ha5);
                    end
                end
              else
                begin
                  if (({(&forvar711[(3'h7):(3'h4)])} < reg730))
                    begin
                      reg726 <= forvar710[(4'h8):(3'h7)];
                    end
                  else
                    begin
                      reg726 <= (~|$signed(reg690));
                      reg727 <= $signed(reg728);
                    end
                  if ((($unsigned(forvar719[(3'h6):(3'h4)]) + reg729[(4'hf):(3'h6)]) ?
                      (!reg716[(2'h3):(1'h0)]) : (|{$unsigned(reg728)})))
                    begin
                      reg728 <= $signed($unsigned($unsigned({reg708})));
                      reg729 <= (|reg737[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg728 <= ((^~$signed(reg708[(4'h8):(4'h8)])) != ({reg731[(2'h2):(2'h2)]} ?
                          (^$unsigned(wire679)) : forvar712[(3'h7):(3'h6)]));
                      reg729 <= $unsigned(($unsigned(reg728[(1'h1):(1'h0)]) & $signed({reg727})));
                      reg730 <= (reg707[(2'h3):(1'h0)] < reg700[(3'h6):(3'h5)]);
                    end
                  for (forvar731 = (1'h0); (forvar731 < (2'h2)); forvar731 = (forvar731 + (1'h1)))
                    begin
                      reg732 <= $signed((reg723[(3'h5):(3'h5)] + forvar706[(1'h1):(1'h0)]));
                    end
                  for (forvar733 = (1'h0); (forvar733 < (2'h2)); forvar733 = (forvar733 + (1'h1)))
                    begin
                      reg734 <= (reg721 && {reg724});
                    end
                end
              if (reg736[(4'ha):(1'h0)])
                begin
                  if ($signed($signed((-(forvar712 > reg718)))))
                    begin
                      reg735 <= reg724[(2'h3):(2'h2)];
                      reg736 <= $unsigned((forvar733[(1'h0):(1'h0)] ?
                          ($unsigned((8'hab)) - $signed(forvar718)) : (8'haf)));
                      reg737 <= (^{(8'haf)});
                      reg738 <= ((+(8'ha3)) >>> (((forvar682 ?
                              wire678 : forvar707) <= (8'hb6)) ?
                          (((8'h9e) < forvar706) <= (~reg720)) : (~(reg717 ?
                              (8'h9d) : reg695))));
                    end
                  else
                    begin
                      reg735 <= (|{$unsigned(reg696[(3'h4):(2'h3)])});
                      reg736 <= forvar734;
                    end
                  if ((reg705[(3'h5):(3'h5)] + $signed({$unsigned((8'haf))})))
                    begin
                      reg739 <= (((|$unsigned(reg738)) ?
                          (-$unsigned((8'hb0))) : reg683) && wire676[(2'h2):(2'h2)]);
                      reg740 <= reg693[(4'hb):(4'hb)];
                    end
                  else
                    begin
                      reg739 <= (8'ha2);
                      reg740 <= reg731;
                      reg741 <= {reg709[(2'h2):(1'h0)]};
                    end
                  reg742 <= $signed((8'ha8));
                  reg743 <= $signed({($signed(forvar710) << reg742)});
                end
              else
                begin
                  for (forvar735 = (1'h0); (forvar735 < (1'h1)); forvar735 = (forvar735 + (1'h1)))
                    begin
                      reg736 <= ((($signed(reg690) > (-forvar711)) ?
                          reg713[(4'h9):(1'h0)] : $signed(((8'hba) - wire677))) - ((reg705[(1'h1):(1'h0)] ?
                          forvar702[(3'h5):(2'h3)] : (~&reg690)) & ((~reg724) ?
                          (!(8'hb3)) : (reg701 ? forvar681 : reg724))));
                      reg737 <= forvar707[(3'h6):(2'h3)];
                      reg738 <= (((|$unsigned(forvar731)) ?
                          wire677 : (~|$signed(forvar712))) < $unsigned((^~(+reg694))));
                      reg739 <= forvar687[(1'h1):(1'h1)];
                    end
                  if ({(-(&(reg736 & forvar735)))})
                    begin
                      reg740 <= forvar709[(3'h5):(2'h2)];
                      reg741 <= (~&($signed($unsigned((8'hb9))) ?
                          forvar734 : ((forvar681 << forvar735) <= (~reg690))));
                      reg742 <= reg710;
                      reg743 <= (|$signed((!wire678[(2'h3):(1'h1)])));
                    end
                  else
                    begin
                      reg740 <= $unsigned(reg696);
                    end
                  if ($signed(((((8'hae) | (8'hb2)) ?
                          $unsigned((8'haf)) : (reg738 ?
                              forvar682 : forvar689)) ?
                      {$signed((8'ha2))} : reg685)))
                    begin
                      reg744 <= $signed(forvar716[(3'h7):(3'h5)]);
                      reg745 <= (+reg729);
                      reg746 <= (reg686[(1'h0):(1'h0)] ?
                          reg694 : {$signed((-forvar724))});
                      reg747 <= $unsigned($signed($signed(reg730)));
                    end
                  else
                    begin
                      reg744 <= (+(^($signed((8'h9c)) ? reg737 : (|reg708))));
                      reg745 <= (^~(($signed(reg696) + (reg732 <<< (8'ha8))) ^ (8'hb9)));
                    end
                end
            end
          reg748 <= {(((-reg684) << {forvar715}) ^ $unsigned(forvar707))};
          for (forvar749 = (1'h0); (forvar749 < (1'h1)); forvar749 = (forvar749 + (1'h1)))
            begin
              if (wire677[(1'h1):(1'h1)])
                begin
                  if ({({(^~reg743)} ?
                          {{reg720}} : ((reg732 & reg685) ?
                              $unsigned(reg727) : (reg685 >>> reg703)))})
                    begin
                      reg750 <= forvar730;
                      reg751 <= $unsigned($unsigned(forvar716[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg750 <= ($signed((reg743 < forvar680[(3'h4):(2'h3)])) ?
                          $signed(reg746) : (8'had));
                      reg751 <= {({(reg723 ? reg710 : forvar689)} ?
                              forvar733 : ({reg700} ?
                                  (+(8'hb8)) : $unsigned(reg698)))};
                      reg752 <= $signed($signed({$signed(reg737)}));
                      reg753 <= {((reg716[(2'h2):(1'h0)] ?
                              $unsigned(reg709) : (8'hb8)) ^~ reg705)};
                    end
                  for (forvar754 = (1'h0); (forvar754 < (1'h0)); forvar754 = (forvar754 + (1'h1)))
                    begin
                      reg755 <= ((8'hae) <<< (((~forvar681) ?
                              (forvar681 < reg726) : reg752[(2'h2):(1'h1)]) ?
                          $signed($signed(reg727)) : reg734[(4'h9):(1'h0)]));
                      reg756 <= $signed((!$signed($signed(forvar710))));
                      reg757 <= ({wire676} ?
                          ($signed((reg741 & reg694)) >= $unsigned($unsigned(reg724))) : (({reg756} < reg730[(4'hd):(3'h4)]) ?
                              (|$unsigned((8'hae))) : reg726));
                    end
                  if ((8'hb6))
                    begin
                      reg758 <= {reg737[(3'h5):(3'h5)]};
                      reg759 <= {reg700};
                      reg760 <= $unsigned(reg753[(4'h9):(3'h6)]);
                    end
                  else
                    begin
                      reg758 <= (forvar689[(2'h2):(1'h0)] > (forvar735[(1'h0):(1'h0)] ?
                          $unsigned((!(8'haf))) : ({reg732} ?
                              forvar712[(1'h1):(1'h1)] : $signed(reg750))));
                      reg759 <= (({wire677} & forvar689) ?
                          $signed(forvar715) : $signed((8'ha2)));
                    end
                  reg761 <= $unsigned(reg685);
                end
              else
                begin
                  if (reg700[(3'h6):(1'h0)])
                    begin
                      reg750 <= {reg714[(2'h2):(1'h0)]};
                      reg751 <= {reg725[(3'h4):(3'h4)]};
                    end
                  else
                    begin
                      reg750 <= forvar707;
                      reg751 <= (8'ha5);
                      reg752 <= reg713[(1'h0):(1'h0)];
                      reg753 <= ($unsigned((8'hb5)) ?
                          ($unsigned($signed(forvar709)) ~^ (wire677[(1'h1):(1'h0)] ?
                              $unsigned(reg690) : reg747[(4'ha):(2'h2)])) : (($unsigned(reg745) ?
                                  forvar719[(3'h4):(1'h0)] : $signed(forvar688)) ?
                              $signed({reg721}) : (8'hb9)));
                    end
                  for (forvar754 = (1'h0); (forvar754 < (2'h2)); forvar754 = (forvar754 + (1'h1)))
                    begin
                      reg755 <= ($unsigned(((reg735 ?
                          wire678 : reg684) ^~ $signed(reg710))) && $unsigned(($unsigned(reg695) ?
                          (reg697 ~^ (8'ha4)) : reg709)));
                      reg756 <= ((reg711 ? (8'ha3) : (^(^reg704))) ?
                          ((~{forvar730}) > {((8'h9e) ^ forvar709)}) : reg748);
                      reg757 <= $unsigned({reg757});
                    end
                end
              reg762 <= (forvar689[(1'h1):(1'h0)] ?
                  ((8'ha0) ^ {reg761[(3'h6):(3'h4)]}) : ((reg702 ?
                          (reg719 <<< reg748) : (forvar716 ?
                              (8'hb7) : forvar754)) ?
                      (reg699[(1'h0):(1'h0)] && reg709[(4'hb):(3'h4)]) : reg721));
              for (forvar763 = (1'h0); (forvar763 < (2'h3)); forvar763 = (forvar763 + (1'h1)))
                begin
                  for (forvar764 = (1'h0); (forvar764 < (1'h0)); forvar764 = (forvar764 + (1'h1)))
                    begin
                      reg765 <= reg710[(3'h4):(1'h1)];
                    end
                  reg766 <= $unsigned($unsigned(reg750));
                end
              if (reg719[(1'h0):(1'h0)])
                begin
                  if (reg708[(4'h8):(4'h8)])
                    begin
                      reg767 <= $unsigned(((reg755 || reg709[(3'h7):(1'h1)]) ?
                          reg735 : reg694));
                      reg768 <= $unsigned({{$unsigned((8'h9e))}});
                    end
                  else
                    begin
                      reg767 <= (^~$signed({(reg756 * reg742)}));
                      reg768 <= reg766[(4'hb):(1'h0)];
                      reg769 <= (&forvar726);
                    end
                  for (forvar770 = (1'h0); (forvar770 < (2'h3)); forvar770 = (forvar770 + (1'h1)))
                    begin
                      reg771 <= $signed($signed((8'hb4)));
                      reg772 <= $unsigned({(reg691 ?
                              $unsigned(wire679) : (reg709 >> (8'h9f)))});
                    end
                  for (forvar773 = (1'h0); (forvar773 < (1'h0)); forvar773 = (forvar773 + (1'h1)))
                    begin
                      reg774 <= forvar749;
                      reg775 <= ((-reg690) >>> forvar707);
                      reg776 <= ((($unsigned((8'hb6)) != forvar724) || (|forvar707[(1'h1):(1'h0)])) ?
                          forvar702 : (~|reg762[(1'h1):(1'h1)]));
                      reg777 <= reg697[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar767 = (1'h0); (forvar767 < (2'h2)); forvar767 = (forvar767 + (1'h1)))
                    begin
                      reg768 <= reg777[(2'h2):(2'h2)];
                      reg769 <= reg691[(3'h7):(3'h7)];
                      reg770 <= forvar711;
                      reg771 <= (reg693 ?
                          $unsigned(reg735) : $unsigned((-$signed(reg720))));
                    end
                  if (reg751[(4'h8):(1'h1)])
                    begin
                      reg772 <= (forvar702 & ((&(forvar773 ?
                              wire676 : reg761)) ?
                          $signed($signed(forvar734)) : (8'haa)));
                      reg773 <= ($signed(forvar731[(3'h5):(3'h4)]) ^~ ((&forvar735[(2'h3):(2'h3)]) ^ {forvar726}));
                      reg774 <= (+reg736[(1'h1):(1'h1)]);
                      reg775 <= reg726[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg772 <= $unsigned($unsigned(($signed(reg716) ?
                          $signed(reg692) : (reg714 ? reg747 : reg685))));
                      reg773 <= $unsigned(((!$unsigned((8'ha9))) < reg771[(3'h4):(2'h2)]));
                    end
                end
            end
          for (forvar778 = (1'h0); (forvar778 < (2'h2)); forvar778 = (forvar778 + (1'h1)))
            begin
              for (forvar779 = (1'h0); (forvar779 < (1'h0)); forvar779 = (forvar779 + (1'h1)))
                begin
                  for (forvar780 = (1'h0); (forvar780 < (2'h3)); forvar780 = (forvar780 + (1'h1)))
                    begin
                      reg781 <= $unsigned(((reg741[(3'h4):(1'h0)] ?
                              forvar778 : ((8'hb6) >> reg765)) ?
                          reg699 : ($signed(reg697) >>> reg718[(3'h4):(1'h1)])));
                    end
                  for (forvar782 = (1'h0); (forvar782 < (2'h3)); forvar782 = (forvar782 + (1'h1)))
                    begin
                      reg783 <= $unsigned((!reg736));
                      reg784 <= forvar767;
                      reg785 <= wire676;
                      reg786 <= (forvar709 || reg710[(1'h1):(1'h0)]);
                    end
                  reg787 <= (8'h9c);
                  reg788 <= reg750[(2'h3):(1'h1)];
                end
            end
        end
      for (forvar789 = (1'h0); (forvar789 < (1'h1)); forvar789 = (forvar789 + (1'h1)))
        begin
          if (forvar719[(1'h0):(1'h0)])
            begin
              if ($unsigned((forvar719[(2'h3):(2'h3)] ^ $signed(forvar719[(1'h1):(1'h1)]))))
                begin
                  for (forvar790 = (1'h0); (forvar790 < (1'h0)); forvar790 = (forvar790 + (1'h1)))
                    begin
                      reg791 <= reg733;
                    end
                  for (forvar792 = (1'h0); (forvar792 < (1'h0)); forvar792 = (forvar792 + (1'h1)))
                    begin
                      reg793 <= reg775;
                      reg794 <= $signed(($signed((reg738 | (8'hb3))) ?
                          reg684 : $signed(reg718[(1'h1):(1'h0)])));
                      reg795 <= (((~|forvar754[(1'h0):(1'h0)]) ^ (&(reg753 * reg724))) ?
                          (forvar689 >= $unsigned((-reg701))) : {wire678});
                      reg796 <= ({reg751[(3'h5):(3'h4)]} & $unsigned((forvar719 <= (forvar689 ?
                          reg795 : reg786))));
                    end
                end
              else
                begin
                  reg790 <= ($unsigned((8'ha7)) ^~ forvar767[(1'h0):(1'h0)]);
                end
              if ($signed(($unsigned($signed(reg708)) > reg788)))
                begin
                  for (forvar797 = (1'h0); (forvar797 < (2'h2)); forvar797 = (forvar797 + (1'h1)))
                    begin
                      reg798 <= reg697;
                    end
                  for (forvar799 = (1'h0); (forvar799 < (2'h2)); forvar799 = (forvar799 + (1'h1)))
                    begin
                      reg800 <= {(|((|reg726) * $unsigned((8'hae))))};
                      reg801 <= forvar729[(1'h0):(1'h0)];
                      reg802 <= ({$signed($unsigned(reg776))} && (~&$unsigned($signed((8'ha7)))));
                    end
                  for (forvar803 = (1'h0); (forvar803 < (1'h0)); forvar803 = (forvar803 + (1'h1)))
                    begin
                      reg804 <= {(reg693[(3'h7):(2'h2)] == {$unsigned(reg755)})};
                      reg805 <= reg712[(1'h0):(1'h0)];
                      reg806 <= $unsigned({$unsigned((reg709 | forvar773))});
                      reg807 <= reg728;
                    end
                end
              else
                begin
                  for (forvar797 = (1'h0); (forvar797 < (2'h3)); forvar797 = (forvar797 + (1'h1)))
                    begin
                      reg798 <= ($signed($unsigned($unsigned((8'ha7)))) ?
                          (~^{$signed(reg760)}) : $unsigned((forvar780 ?
                              $signed(reg758) : ((8'ha7) ? reg729 : reg690))));
                    end
                  if ($signed((~^$unsigned((reg709 == reg683)))))
                    begin
                      reg799 <= ($signed(forvar789[(2'h2):(1'h1)]) >>> $unsigned(((~^reg771) << reg691)));
                      reg800 <= (({$unsigned(forvar734)} - {{(8'ha9)}}) ?
                          (^~(-(~&(8'hb9)))) : $unsigned(reg743));
                      reg801 <= (forvar729 ?
                          ($unsigned(((8'ha1) | (8'h9e))) ?
                              forvar790[(3'h4):(2'h2)] : (-$unsigned(forvar763))) : {reg805[(1'h1):(1'h1)]});
                    end
                  else
                    begin
                      reg799 <= forvar706;
                    end
                  for (forvar802 = (1'h0); (forvar802 < (2'h2)); forvar802 = (forvar802 + (1'h1)))
                    begin
                      reg803 <= (forvar802[(4'hc):(4'h8)] ?
                          $unsigned(reg728) : $signed($unsigned($signed(reg769))));
                      reg804 <= ((|(|(forvar687 | reg729))) <<< reg686);
                    end
                end
              for (forvar808 = (1'h0); (forvar808 < (1'h1)); forvar808 = (forvar808 + (1'h1)))
                begin
                  for (forvar809 = (1'h0); (forvar809 < (2'h2)); forvar809 = (forvar809 + (1'h1)))
                    begin
                      reg810 <= (-(~^forvar778[(2'h3):(2'h2)]));
                      reg811 <= (wire678 + $unsigned((+$unsigned((8'haf)))));
                      reg812 <= ((8'hb8) << forvar764);
                      reg813 <= (8'hae);
                    end
                end
              if ($signed({reg786[(4'h9):(3'h5)]}))
                begin
                  for (forvar814 = (1'h0); (forvar814 < (1'h1)); forvar814 = (forvar814 + (1'h1)))
                    begin
                      reg815 <= (reg722 ? reg811 : {$unsigned((-reg799))});
                      reg816 <= (-reg701);
                    end
                end
              else
                begin
                  for (forvar814 = (1'h0); (forvar814 < (2'h3)); forvar814 = (forvar814 + (1'h1)))
                    begin
                      reg815 <= (reg765[(1'h0):(1'h0)] ?
                          ($signed((reg753 ?
                              reg693 : forvar715)) ^~ $signed(forvar778)) : $signed({(~&(8'ha9))}));
                      reg816 <= reg700[(1'h1):(1'h1)];
                      reg817 <= ($signed((!$unsigned(reg804))) ?
                          {forvar731} : reg745);
                    end
                  if (reg714[(3'h4):(1'h0)])
                    begin
                      reg818 <= (8'hb4);
                      reg819 <= ($unsigned($unsigned((reg746 ?
                          reg697 : reg728))) ^ $unsigned((~|{forvar767})));
                      reg820 <= $signed(((|(~reg734)) ?
                          reg707 : $signed((reg807 << reg755))));
                      reg821 <= reg756[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg818 <= {$unsigned(((reg694 < reg769) <= (reg762 ~^ reg815)))};
                      reg819 <= (reg787[(1'h1):(1'h0)] | $unsigned({reg771}));
                      reg820 <= (((forvar799 <= reg727[(2'h2):(2'h2)]) ~^ ($unsigned(reg791) <= $signed(reg730))) <<< forvar782);
                      reg821 <= ($unsigned({forvar716[(1'h0):(1'h0)]}) ?
                          $unsigned((|$signed(forvar767))) : (~($unsigned((8'h9c)) ?
                              (8'hb3) : $unsigned(reg752))));
                    end
                  for (forvar822 = (1'h0); (forvar822 < (2'h3)); forvar822 = (forvar822 + (1'h1)))
                    begin
                      reg823 <= ($unsigned({(reg698 == reg772)}) ?
                          (forvar808 ?
                              (reg810 ?
                                  forvar706[(3'h5):(1'h0)] : $unsigned((8'h9f))) : (reg777 ?
                                  {(8'hb3)} : $unsigned(reg710))) : {$unsigned({(8'hae)})});
                      reg824 <= forvar702;
                      reg825 <= {(($signed(forvar735) == (reg729 ?
                              reg802 : (8'ha4))) == reg805[(1'h1):(1'h0)])};
                      reg826 <= $signed(({reg686} ?
                          $signed($signed(forvar809)) : $signed(reg708)));
                    end
                  if (reg825[(1'h1):(1'h0)])
                    begin
                      reg827 <= ((reg750 * reg695[(3'h5):(2'h2)]) ?
                          ($signed((|reg700)) <= (|$unsigned(reg725))) : reg815);
                    end
                  else
                    begin
                      reg827 <= ((~^reg715) ?
                          (!$signed((reg722 & (8'hb2)))) : reg774[(1'h0):(1'h0)]);
                      reg828 <= reg775[(4'hc):(4'ha)];
                    end
                end
            end
          else
            begin
              for (forvar790 = (1'h0); (forvar790 < (2'h2)); forvar790 = (forvar790 + (1'h1)))
                begin
                  for (forvar791 = (1'h0); (forvar791 < (1'h0)); forvar791 = (forvar791 + (1'h1)))
                    begin
                      reg792 <= ($signed(((!forvar688) || reg760)) ?
                          (~(reg800[(3'h4):(2'h3)] ?
                              $signed(reg694) : $unsigned(reg786))) : (8'h9f));
                      reg793 <= $unsigned($unsigned(reg696[(2'h2):(2'h2)]));
                      reg794 <= reg714[(1'h1):(1'h0)];
                      reg795 <= ((~$unsigned($unsigned(reg698))) ?
                          reg775 : $unsigned(({forvar754} + $signed(forvar716))));
                    end
                  if ((~reg700))
                    begin
                      reg796 <= $unsigned(reg777);
                    end
                  else
                    begin
                      reg796 <= (((!$signed(forvar718)) ?
                              $unsigned(((8'h9c) ~^ reg802)) : reg743[(1'h0):(1'h0)]) ?
                          {(^reg813[(3'h7):(3'h5)])} : $unsigned($signed((^~reg737))));
                      reg797 <= ((reg776[(2'h3):(1'h0)] ?
                          ($signed(reg729) && reg719[(3'h4):(2'h3)]) : ($unsigned(forvar782) - {reg773})) ^ (^~((^forvar689) ?
                          (forvar780 & wire677) : reg788[(2'h2):(2'h2)])));
                      reg798 <= $unsigned($unsigned($unsigned(reg730[(4'hb):(3'h4)])));
                    end
                end
              for (forvar799 = (1'h0); (forvar799 < (1'h0)); forvar799 = (forvar799 + (1'h1)))
                begin
                  if (reg733)
                    begin
                      reg800 <= reg810[(1'h1):(1'h0)];
                      reg801 <= $unsigned(forvar716[(3'h5):(2'h3)]);
                      reg802 <= (((reg739 ?
                              $unsigned(forvar749) : $unsigned(reg794)) ?
                          (^$unsigned(reg798)) : $unsigned(reg686)) ^~ reg745);
                      reg803 <= $signed(reg790[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg800 <= ((8'ha1) ?
                          $signed(($unsigned(reg698) ?
                              {reg790} : (reg790 ?
                                  (8'ha7) : reg691))) : (8'ha9));
                      reg801 <= reg690;
                      reg802 <= (reg760 ?
                          reg710[(3'h5):(3'h4)] : ({forvar802[(3'h6):(3'h6)]} && $signed(reg759)));
                    end
                  for (forvar804 = (1'h0); (forvar804 < (1'h1)); forvar804 = (forvar804 + (1'h1)))
                    begin
                      reg805 <= reg816[(4'ha):(4'h8)];
                    end
                  reg806 <= {((reg772[(3'h7):(3'h6)] ?
                              (+forvar802) : forvar803) ?
                          (!(!reg793)) : $signed(reg699))};
                end
              if ((~&$unsigned(reg759)))
                begin
                  if (forvar707[(3'h4):(1'h1)])
                    begin
                      reg807 <= ({$signed($unsigned(reg719))} && $signed($unsigned((wire677 ?
                          forvar706 : reg737))));
                    end
                  else
                    begin
                      reg807 <= $unsigned((+$unsigned((reg724 || reg775))));
                      reg808 <= (reg719[(1'h0):(1'h0)] ^ ($signed((wire676 * reg737)) ?
                          reg803[(4'hb):(1'h1)] : (8'h9f)));
                      reg809 <= (reg744 ?
                          reg800[(3'h4):(2'h3)] : $signed($signed((reg707 != forvar822))));
                    end
                  if ((+$signed(reg714[(3'h5):(3'h5)])))
                    begin
                      reg810 <= (~|{$unsigned((reg700 < (8'hac)))});
                      reg811 <= $unsigned(reg802);
                    end
                  else
                    begin
                      reg810 <= (reg695 ?
                          $signed(forvar688[(1'h1):(1'h0)]) : reg815);
                      reg811 <= $unsigned((~|(8'ha2)));
                    end
                  for (forvar812 = (1'h0); (forvar812 < (1'h1)); forvar812 = (forvar812 + (1'h1)))
                    begin
                      reg813 <= (+forvar724[(3'h5):(1'h0)]);
                      reg814 <= $unsigned(reg762[(3'h4):(1'h1)]);
                    end
                end
              else
                begin
                  if (reg759[(1'h1):(1'h1)])
                    begin
                      reg807 <= $unsigned($signed(((reg787 ?
                          reg684 : forvar763) > reg701[(3'h5):(1'h1)])));
                      reg808 <= (^reg769);
                      reg809 <= (reg774 ?
                          reg759[(3'h4):(1'h1)] : $signed(((^reg707) ?
                              (!reg784) : (reg709 ? forvar808 : (8'ha1)))));
                    end
                  else
                    begin
                      reg807 <= reg698;
                    end
                  if (reg770[(1'h0):(1'h0)])
                    begin
                      reg810 <= $unsigned({($signed(reg765) ?
                              forvar782[(1'h1):(1'h0)] : $unsigned(reg810))});
                      reg811 <= $unsigned(((forvar680[(3'h4):(1'h0)] >= $unsigned(reg693)) ?
                          ((reg824 && forvar681) ?
                              $signed(forvar803) : (reg805 ?
                                  (8'had) : reg691)) : reg752[(1'h1):(1'h0)]));
                      reg812 <= (~|($signed((~^reg802)) ~^ (8'haa)));
                      reg813 <= reg791;
                    end
                  else
                    begin
                      reg810 <= reg685[(3'h4):(1'h1)];
                      reg811 <= reg752[(1'h1):(1'h0)];
                    end
                end
            end
          if (reg692)
            begin
              if (((+(reg708 ?
                  reg767[(4'hd):(4'hc)] : forvar791)) > reg768[(2'h2):(2'h2)]))
                begin
                  reg829 <= reg788;
                  for (forvar830 = (1'h0); (forvar830 < (1'h1)); forvar830 = (forvar830 + (1'h1)))
                    begin
                      reg831 <= reg785;
                      reg832 <= $unsigned($unsigned($unsigned(forvar719[(2'h2):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar829 = (1'h0); (forvar829 < (2'h3)); forvar829 = (forvar829 + (1'h1)))
                    begin
                      reg830 <= $signed(reg711[(3'h4):(1'h0)]);
                      reg831 <= $unsigned($unsigned(($signed(forvar710) ?
                          (forvar729 ? reg797 : reg771) : $signed(reg736))));
                    end
                  for (forvar832 = (1'h0); (forvar832 < (1'h0)); forvar832 = (forvar832 + (1'h1)))
                    begin
                      reg833 <= (8'ha2);
                      reg834 <= (-$unsigned(reg725[(2'h2):(1'h0)]));
                      reg835 <= forvar804[(1'h0):(1'h0)];
                    end
                  reg836 <= $signed(forvar770);
                end
              for (forvar837 = (1'h0); (forvar837 < (1'h1)); forvar837 = (forvar837 + (1'h1)))
                begin
                  for (forvar838 = (1'h0); (forvar838 < (1'h1)); forvar838 = (forvar838 + (1'h1)))
                    begin
                      reg839 <= (-(^reg759[(4'h8):(1'h1)]));
                      reg840 <= $signed({reg836});
                      reg841 <= ((+(reg801 ?
                          (~&reg704) : reg744)) >> reg714[(1'h1):(1'h1)]);
                      reg842 <= (reg807 ~^ reg762);
                    end
                  if ((+(reg815 ?
                      reg727[(1'h1):(1'h1)] : (~reg747[(1'h0):(1'h0)]))))
                    begin
                      reg843 <= reg755[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg843 <= (reg836 ?
                          $unsigned(((8'had) ^ $unsigned(forvar779))) : reg750[(2'h3):(2'h2)]);
                      reg844 <= forvar733[(1'h1):(1'h1)];
                      reg845 <= $unsigned(reg788[(1'h1):(1'h1)]);
                    end
                end
              reg846 <= $signed(forvar718[(1'h0):(1'h0)]);
              for (forvar847 = (1'h0); (forvar847 < (2'h2)); forvar847 = (forvar847 + (1'h1)))
                begin
                  reg848 <= (~|((~(reg701 <<< reg785)) ?
                      (((8'h9e) && reg736) | $unsigned(reg747)) : ($signed(reg759) ?
                          reg815 : (~&reg727))));
                end
            end
          else
            begin
              reg829 <= ($unsigned(reg685[(3'h4):(2'h3)]) ?
                  (reg696 && {reg752}) : $signed($signed($signed(reg752))));
              for (forvar830 = (1'h0); (forvar830 < (1'h1)); forvar830 = (forvar830 + (1'h1)))
                begin
                  for (forvar831 = (1'h0); (forvar831 < (2'h2)); forvar831 = (forvar831 + (1'h1)))
                    begin
                      reg832 <= (~reg738[(1'h0):(1'h0)]);
                      reg833 <= $signed(($signed(forvar792[(4'h9):(3'h4)]) >= ($signed(reg785) >> $signed(reg783))));
                    end
                  if ({(reg693 <= ($signed(reg825) ?
                          (forvar779 ?
                              reg714 : wire679) : forvar688[(4'ha):(2'h2)]))})
                    begin
                      reg834 <= ((^~{reg771}) ?
                          ((8'hb3) ?
                              reg844[(3'h5):(3'h5)] : forvar706) : reg818);
                      reg835 <= ($unsigned($signed({reg839})) ?
                          (8'ha1) : (reg787[(2'h2):(1'h0)] ?
                              (|(~^(8'haf))) : $signed({reg745})));
                      reg836 <= $signed($unsigned(reg800));
                      reg837 <= {((~|(|forvar710)) != ($unsigned(forvar764) ?
                              $signed(forvar808) : (8'ha8)))};
                    end
                  else
                    begin
                      reg834 <= wire679;
                    end
                  if (forvar792[(3'h4):(3'h4)])
                    begin
                      reg838 <= {{({reg819} ?
                                  (forvar719 ^~ reg699) : $signed(reg788))}};
                      reg839 <= ({reg723} >> $unsigned({(forvar790 ?
                              reg816 : reg807)}));
                      reg840 <= $signed($signed((reg844[(3'h5):(3'h4)] | $unsigned((8'hb4)))));
                      reg841 <= (!(($signed(reg745) ~^ (reg720 ?
                              reg698 : (8'ha3))) ?
                          {reg760} : reg692));
                    end
                  else
                    begin
                      reg838 <= {reg761};
                    end
                end
              for (forvar842 = (1'h0); (forvar842 < (1'h0)); forvar842 = (forvar842 + (1'h1)))
                begin
                  reg843 <= {($signed($unsigned((8'hb3))) * reg824)};
                  for (forvar844 = (1'h0); (forvar844 < (2'h2)); forvar844 = (forvar844 + (1'h1)))
                    begin
                      reg845 <= {(forvar831 >= {forvar797[(3'h5):(2'h2)]})};
                      reg846 <= $unsigned({(8'had)});
                      reg847 <= ($signed((((8'ha0) >> forvar733) < (&(8'ha2)))) ?
                          ((reg685[(1'h0):(1'h0)] ?
                              $signed(reg715) : reg783) - (~|(reg845 ?
                              (8'ha6) : forvar803))) : $signed({$unsigned(reg831)}));
                    end
                  for (forvar848 = (1'h0); (forvar848 < (2'h3)); forvar848 = (forvar848 + (1'h1)))
                    begin
                      reg849 <= $signed(reg746);
                      reg850 <= (8'hba);
                      reg851 <= (reg748 > reg777);
                    end
                end
              if ($unsigned(forvar688[(3'h4):(1'h1)]))
                begin
                  if (reg743[(1'h1):(1'h0)])
                    begin
                      reg852 <= (^reg825);
                    end
                  else
                    begin
                      reg852 <= ($signed((|reg755)) ?
                          ($signed((|reg761)) ?
                              $unsigned((reg771 ? reg692 : reg831)) : {(reg852 ?
                                      reg790 : reg824)}) : {forvar702});
                      reg853 <= forvar754[(1'h1):(1'h0)];
                      reg854 <= $signed(((!reg723[(3'h6):(3'h5)]) ?
                          $unsigned(forvar716[(3'h6):(1'h1)]) : $unsigned(reg760)));
                      reg855 <= reg811[(3'h7):(1'h1)];
                    end
                  reg856 <= reg849[(1'h0):(1'h0)];
                end
              else
                begin
                  for (forvar852 = (1'h0); (forvar852 < (2'h2)); forvar852 = (forvar852 + (1'h1)))
                    begin
                      reg853 <= (~&(+((~^(8'had)) < (&reg836))));
                    end
                  reg854 <= $signed(forvar724[(4'hd):(3'h5)]);
                  if (((((~reg720) ?
                      reg787[(2'h3):(2'h3)] : {forvar718}) && (reg856 ?
                      (8'ha6) : (reg832 ~^ forvar812))) ^~ $unsigned({(reg809 ^ reg726)})))
                    begin
                      reg855 <= ((8'hb2) ?
                          $signed($unsigned(reg817)) : $signed($signed(forvar687[(1'h0):(1'h0)])));
                      reg856 <= reg705[(3'h5):(1'h1)];
                      reg857 <= reg758;
                      reg858 <= ({$signed((&(8'haa)))} ?
                          (8'hac) : (~|{(reg850 >> forvar767)}));
                    end
                  else
                    begin
                      reg855 <= (-reg757[(1'h0):(1'h0)]);
                      reg856 <= reg776;
                      reg857 <= reg753[(2'h2):(1'h1)];
                      reg858 <= (~^$unsigned(($signed(reg857) & reg829)));
                    end
                end
            end
          for (forvar859 = (1'h0); (forvar859 < (2'h2)); forvar859 = (forvar859 + (1'h1)))
            begin
              if ($unsigned($signed(reg761[(4'h8):(2'h3)])))
                begin
                  for (forvar860 = (1'h0); (forvar860 < (2'h2)); forvar860 = (forvar860 + (1'h1)))
                    begin
                      reg861 <= $signed({$signed((reg714 ? reg770 : reg834))});
                      reg862 <= ($signed((reg774[(1'h1):(1'h1)] ?
                              forvar688[(5'h10):(4'hc)] : $signed(reg848))) ?
                          forvar829[(4'ha):(4'h9)] : forvar734[(1'h1):(1'h1)]);
                    end
                  if ((8'ha6))
                    begin
                      reg863 <= {reg710[(3'h5):(1'h0)]};
                      reg864 <= reg709[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg863 <= forvar710[(4'hc):(2'h2)];
                      reg864 <= {($signed({reg816}) ?
                              $signed(reg739[(2'h3):(2'h3)]) : $signed($signed(reg709)))};
                      reg865 <= reg802[(3'h6):(2'h3)];
                    end
                end
              else
                begin
                  for (forvar860 = (1'h0); (forvar860 < (2'h2)); forvar860 = (forvar860 + (1'h1)))
                    begin
                      reg861 <= ((($signed(reg702) <= $unsigned(forvar719)) ?
                          $signed({(8'haa)}) : reg852) < reg711);
                      reg862 <= $signed((8'ha4));
                    end
                  reg863 <= forvar729;
                end
              for (forvar866 = (1'h0); (forvar866 < (1'h1)); forvar866 = (forvar866 + (1'h1)))
                begin
                  reg867 <= (!$signed((~&$unsigned(reg832))));
                  for (forvar868 = (1'h0); (forvar868 < (1'h1)); forvar868 = (forvar868 + (1'h1)))
                    begin
                      reg869 <= $signed((8'ha9));
                    end
                  for (forvar870 = (1'h0); (forvar870 < (2'h2)); forvar870 = (forvar870 + (1'h1)))
                    begin
                      reg871 <= (8'hb8);
                      reg872 <= (~(&$signed({reg745})));
                      reg873 <= (reg720[(2'h2):(2'h2)] ?
                          $signed(reg842[(1'h1):(1'h1)]) : reg806);
                    end
                end
              for (forvar874 = (1'h0); (forvar874 < (1'h0)); forvar874 = (forvar874 + (1'h1)))
                begin
                  for (forvar875 = (1'h0); (forvar875 < (2'h2)); forvar875 = (forvar875 + (1'h1)))
                    begin
                      reg876 <= {reg808};
                      reg877 <= (((!reg746) > (~&$unsigned(forvar763))) ?
                          ($signed(reg783[(4'hc):(4'hb)]) < (8'hb9)) : (reg783 ?
                              $unsigned((forvar831 || reg862)) : $signed($signed(reg823))));
                      reg878 <= reg736[(3'h7):(2'h2)];
                    end
                  for (forvar879 = (1'h0); (forvar879 < (2'h3)); forvar879 = (forvar879 + (1'h1)))
                    begin
                      reg880 <= $signed(reg736[(2'h3):(1'h1)]);
                      reg881 <= $unsigned($unsigned(($unsigned(forvar688) ?
                          reg762[(1'h1):(1'h1)] : $signed(reg821))));
                      reg882 <= {(-({reg775} < reg816))};
                      reg883 <= $unsigned(forvar838);
                    end
                  if (forvar804)
                    begin
                      reg884 <= ($signed(((8'hba) - (8'hab))) & (~^reg810));
                      reg885 <= (-forvar831);
                      reg886 <= $signed(forvar682[(1'h0):(1'h0)]);
                      reg887 <= (8'haf);
                    end
                  else
                    begin
                      reg884 <= ({(|reg837[(4'h8):(3'h7)])} ?
                          ($signed($signed(reg777)) ?
                              $unsigned((^~reg750)) : reg871[(1'h0):(1'h0)]) : $unsigned(forvar712[(2'h3):(2'h2)]));
                    end
                end
            end
        end
    end
  module888 modinst4170 (.wire889(wire678), .clk(clk), .y(wire4169), .wire890(reg887), .wire891(reg861), .wire892(forvar724), .wire893(forvar799));
  always
    @(posedge clk) begin
      if ((8'hae))
        begin
          for (forvar4171 = (1'h0); (forvar4171 < (1'h1)); forvar4171 = (forvar4171 + (1'h1)))
            begin
              reg4172 <= $unsigned($unsigned((~forvar719)));
              reg4173 <= (~|$signed(($signed((8'hb3)) ?
                  (8'hb0) : (!forvar848))));
              if (((+$signed($signed(forvar706))) | $signed(((reg718 <= (8'h9f)) || reg877))))
                begin
                  for (forvar4174 = (1'h0); (forvar4174 < (2'h2)); forvar4174 = (forvar4174 + (1'h1)))
                    begin
                      reg4175 <= {({{reg811}} ? {(^~forvar842)} : {(8'ha9)})};
                      reg4176 <= ($signed({(&reg776)}) ?
                          (-((forvar710 <<< reg844) * (^~reg852))) : (($signed(wire676) ?
                              (reg740 ?
                                  reg725 : reg720) : reg794) >>> (reg762[(3'h4):(2'h3)] * $unsigned(reg705))));
                    end
                  if ((~^(+reg831[(2'h3):(1'h0)])))
                    begin
                      reg4177 <= {(!(^~forvar749[(3'h5):(2'h3)]))};
                      reg4178 <= $signed(reg745);
                      reg4179 <= (($unsigned((+(8'h9f))) ?
                              $signed((reg848 << reg774)) : $unsigned((forvar767 ^~ reg760))) ?
                          ($signed($signed(reg816)) - reg759) : $signed(reg697));
                      reg4180 <= (forvar767[(4'hb):(1'h0)] ~^ $signed((~|$unsigned(reg696))));
                    end
                  else
                    begin
                      reg4177 <= $signed(forvar778);
                      reg4178 <= reg793;
                      reg4179 <= reg722;
                      reg4180 <= (+((((8'ha2) >= reg785) ?
                          reg837 : $unsigned(reg720)) >> (8'hac)));
                    end
                end
              else
                begin
                  if ({(&((forvar790 ? reg713 : reg776) << $unsigned(reg805)))})
                    begin
                      reg4174 <= ($signed((~forvar731)) ?
                          (reg821 ^~ {reg791[(1'h1):(1'h0)]}) : ((&(!reg770)) == (~&(~|(8'hb8)))));
                      reg4175 <= forvar715;
                      reg4176 <= (reg805[(3'h4):(2'h3)] > forvar734[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4174 <= (8'h9c);
                      reg4175 <= $signed($unsigned(((reg731 ?
                              reg824 : forvar734) ?
                          $signed(reg719) : ((8'h9d) > reg824))));
                    end
                  reg4177 <= $signed(($unsigned((reg774 ? reg4174 : (8'hb5))) ?
                      {(reg846 ?
                              reg752 : forvar719)} : ($signed(reg711) != $unsigned(forvar791))));
                end
              for (forvar4181 = (1'h0); (forvar4181 < (1'h1)); forvar4181 = (forvar4181 + (1'h1)))
                begin
                  reg4182 <= ({$unsigned(forvar715[(1'h1):(1'h1)])} > (-reg704[(1'h0):(1'h0)]));
                  for (forvar4183 = (1'h0); (forvar4183 < (1'h1)); forvar4183 = (forvar4183 + (1'h1)))
                    begin
                      reg4184 <= ((-$signed((forvar731 != forvar709))) != (8'hb1));
                      reg4185 <= $signed(((+reg746[(3'h4):(3'h4)]) != reg854));
                    end
                  reg4186 <= $signed((-(~^$unsigned(reg4177))));
                  if (reg808)
                    begin
                      reg4187 <= (wire676 < reg722);
                      reg4188 <= forvar868[(3'h5):(3'h4)];
                      reg4189 <= ({((forvar814 >= reg4175) != reg684)} >>> $unsigned((-(reg756 ?
                          reg686 : reg684))));
                      reg4190 <= ((((8'h9f) ?
                          {forvar688} : reg730) >= $signed((~^reg813))) >>> ((reg850[(3'h6):(3'h5)] ?
                              ((8'hb3) || reg707) : {reg730}) ?
                          reg742[(2'h2):(1'h1)] : {reg853[(3'h4):(2'h3)]}));
                    end
                  else
                    begin
                      reg4187 <= ($unsigned($unsigned($signed(reg854))) ?
                          reg753 : $signed(reg817[(3'h4):(2'h2)]));
                      reg4188 <= (&$unsigned((-(forvar879 ?
                          (8'had) : (8'hac)))));
                      reg4189 <= forvar773;
                    end
                end
            end
          for (forvar4191 = (1'h0); (forvar4191 < (1'h1)); forvar4191 = (forvar4191 + (1'h1)))
            begin
              if (reg685[(2'h3):(2'h3)])
                begin
                  if (reg769[(1'h0):(1'h0)])
                    begin
                      reg4192 <= reg788[(2'h2):(1'h1)];
                      reg4193 <= reg4174;
                    end
                  else
                    begin
                      reg4192 <= ({$signed({reg801})} <= $signed({(reg837 < reg721)}));
                    end
                  reg4194 <= reg705[(1'h1):(1'h0)];
                end
              else
                begin
                  for (forvar4192 = (1'h0); (forvar4192 < (1'h1)); forvar4192 = (forvar4192 + (1'h1)))
                    begin
                      reg4193 <= (reg855 ?
                          (8'hb6) : (((forvar689 ?
                                  reg719 : reg832) ^ $unsigned(reg717)) ?
                              $unsigned($signed(reg733)) : ($unsigned(reg684) + $unsigned((8'ha8)))));
                    end
                end
            end
          if ($signed(reg697))
            begin
              if (forvar789[(1'h0):(1'h0)])
                begin
                  if ({(~|(8'ha4))})
                    begin
                      reg4195 <= (!$signed((reg751 ?
                          reg692[(4'hb):(4'h9)] : (~^(8'hb8)))));
                      reg4196 <= reg4177;
                    end
                  else
                    begin
                      reg4195 <= (($unsigned((reg848 ?
                          reg4184 : forvar790)) != $signed(reg697[(1'h0):(1'h0)])) <= reg852[(1'h1):(1'h0)]);
                      reg4196 <= (^~(^~reg742[(1'h0):(1'h0)]));
                      reg4197 <= $unsigned(reg799[(4'ha):(2'h2)]);
                    end
                end
              else
                begin
                  if (reg768[(3'h6):(3'h5)])
                    begin
                      reg4195 <= $unsigned((($unsigned(forvar689) ?
                          ((8'ha3) != (8'ha7)) : forvar868) != $unsigned(forvar780[(3'h5):(3'h5)])));
                      reg4196 <= ((8'haf) ?
                          reg777[(2'h2):(1'h0)] : $signed((^~((8'hb4) && reg770))));
                      reg4197 <= ($unsigned(reg817[(2'h3):(1'h1)]) | reg774[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg4195 <= ((~^({forvar749} > ((8'ha8) ?
                              reg806 : forvar779))) ?
                          forvar687[(3'h4):(1'h1)] : (~(&(reg837 & reg4195))));
                      reg4196 <= ($unsigned(forvar715) ?
                          (~^forvar782) : (|$unsigned((forvar803 ?
                              reg751 : (8'hb7)))));
                    end
                  if (forvar4171)
                    begin
                      reg4198 <= (^(&(8'hb5)));
                    end
                  else
                    begin
                      reg4198 <= ((~&({forvar767} <= forvar716[(3'h4):(1'h0)])) ^ (!$signed($unsigned(reg714))));
                      reg4199 <= ({reg842[(3'h5):(1'h0)]} != {$unsigned($unsigned(forvar847))});
                      reg4200 <= (reg878[(3'h5):(1'h1)] ?
                          reg816[(3'h7):(2'h2)] : reg705);
                    end
                  reg4201 <= forvar767;
                  for (forvar4202 = (1'h0); (forvar4202 < (1'h0)); forvar4202 = (forvar4202 + (1'h1)))
                    begin
                      reg4203 <= reg719[(2'h3):(2'h3)];
                    end
                end
              for (forvar4204 = (1'h0); (forvar4204 < (1'h0)); forvar4204 = (forvar4204 + (1'h1)))
                begin
                  for (forvar4205 = (1'h0); (forvar4205 < (2'h2)); forvar4205 = (forvar4205 + (1'h1)))
                    begin
                      reg4206 <= {($unsigned((reg738 ? reg797 : (8'hb8))) ?
                              {((8'hb2) ?
                                      (8'ha5) : reg4186)} : $unsigned((reg4172 ?
                                  reg864 : forvar868)))};
                      reg4207 <= {(~^(~^(+reg883)))};
                      reg4208 <= {({(reg745 ^ forvar724)} != reg768)};
                    end
                  for (forvar4209 = (1'h0); (forvar4209 < (2'h2)); forvar4209 = (forvar4209 + (1'h1)))
                    begin
                      reg4210 <= reg828[(3'h6):(2'h2)];
                      reg4211 <= $unsigned((((forvar852 ? (8'hb8) : reg811) ?
                          reg708[(2'h3):(1'h0)] : reg845[(2'h2):(1'h1)]) || reg781));
                      reg4212 <= $signed($unsigned(forvar687[(2'h3):(2'h2)]));
                      reg4213 <= $signed(forvar832[(4'h9):(1'h1)]);
                    end
                end
            end
          else
            begin
              if (reg4174)
                begin
                  reg4195 <= reg843;
                  if ($unsigned(((forvar868 ?
                          (wire679 ^ forvar681) : $signed(forvar681)) ?
                      ($unsigned(reg784) ~^ (wire678 ?
                          reg817 : forvar804)) : forvar711)))
                    begin
                      reg4196 <= (~|$unsigned(($signed(reg750) ?
                          (reg4182 <<< reg705) : reg873)));
                    end
                  else
                    begin
                      reg4196 <= (reg685 ?
                          (reg802[(4'hb):(1'h1)] & (|$signed(reg4174))) : (({reg693} ?
                                  (^(8'hb3)) : forvar718[(3'h5):(2'h3)]) ?
                              (8'ha9) : forvar4209));
                      reg4197 <= (+{{reg771[(3'h6):(3'h6)]}});
                      reg4198 <= {reg831};
                    end
                end
              else
                begin
                  if (((&(8'hb5)) ?
                      reg774[(2'h2):(2'h2)] : (reg716[(2'h2):(1'h0)] || ($signed(reg729) ?
                          (reg743 ? reg770 : reg792) : $unsigned(reg704)))))
                    begin
                      reg4195 <= (reg773[(1'h1):(1'h0)] ~^ $unsigned($unsigned((~|reg4194))));
                      reg4196 <= (&(~|{(reg4178 ? reg734 : reg831)}));
                    end
                  else
                    begin
                      reg4195 <= (8'h9e);
                      reg4196 <= ((^~reg4197) >= (^(-reg843)));
                    end
                  reg4197 <= $signed({$unsigned((reg832 ? (8'hb1) : reg708))});
                  for (forvar4198 = (1'h0); (forvar4198 < (1'h1)); forvar4198 = (forvar4198 + (1'h1)))
                    begin
                      reg4199 <= reg762;
                    end
                  reg4200 <= reg819;
                end
              reg4201 <= reg4210[(1'h0):(1'h0)];
            end
          for (forvar4214 = (1'h0); (forvar4214 < (1'h1)); forvar4214 = (forvar4214 + (1'h1)))
            begin
              reg4215 <= $unsigned((((reg776 ? (8'hba) : reg721) ?
                      $unsigned((8'hac)) : reg733[(2'h3):(2'h2)]) ?
                  reg727[(4'h8):(3'h7)] : reg849[(4'hb):(3'h4)]));
              if (((($signed(reg745) < {reg769}) ?
                  reg840 : (reg4211 + $unsigned(reg828))) || (((&reg717) + (forvar4204 >= (8'ha7))) + (((8'hb6) ^~ reg884) >>> (|forvar837)))))
                begin
                  for (forvar4216 = (1'h0); (forvar4216 < (1'h0)); forvar4216 = (forvar4216 + (1'h1)))
                    begin
                      reg4217 <= {reg795[(3'h4):(2'h2)]};
                      reg4218 <= $unsigned(reg880);
                      reg4219 <= (+(forvar735[(1'h0):(1'h0)] ?
                          reg871 : $signed({reg832})));
                    end
                end
              else
                begin
                  for (forvar4216 = (1'h0); (forvar4216 < (1'h1)); forvar4216 = (forvar4216 + (1'h1)))
                    begin
                      reg4217 <= (reg758[(2'h2):(2'h2)] <= (^((reg4174 ?
                              reg846 : reg733) ?
                          reg790[(4'hc):(2'h3)] : (|reg848))));
                    end
                  if (($signed(reg711[(2'h2):(2'h2)]) ^ (8'ha1)))
                    begin
                      reg4218 <= $signed(((~(reg4210 ?
                          reg836 : forvar870)) != ($signed(reg767) || $unsigned(forvar4198))));
                      reg4219 <= ((((reg807 << reg834) ?
                              reg849 : reg4194[(3'h6):(2'h3)]) ?
                          $signed(forvar870[(2'h3):(2'h2)]) : $unsigned(reg4211)) & $unsigned(({reg774} ?
                          reg767[(1'h0):(1'h0)] : $signed(forvar4209))));
                      reg4220 <= (($unsigned((reg721 || (8'hb7))) ?
                              $unsigned(reg798[(1'h0):(1'h0)]) : $unsigned((reg766 ?
                                  forvar838 : reg798))) ?
                          $signed($unsigned((forvar688 < forvar733))) : ({$signed(reg4190)} != (reg871 ?
                              forvar790[(4'hc):(4'hc)] : forvar754)));
                      reg4221 <= $signed(reg801);
                    end
                  else
                    begin
                      reg4218 <= $signed(((~^(reg690 << wire676)) >>> ((8'ha2) ?
                          (^reg882) : $signed(reg821))));
                    end
                  if (($unsigned(forvar689) >>> (reg4174 ?
                      reg850[(2'h3):(2'h2)] : ((&forvar875) ?
                          $unsigned(reg785) : (^~reg4218)))))
                    begin
                      reg4222 <= (reg717[(1'h1):(1'h0)] ?
                          {{(forvar724 ?
                                      reg708 : forvar707)}} : (-(~^reg719[(1'h1):(1'h0)])));
                      reg4223 <= ((+(+$signed(reg711))) ?
                          $unsigned($signed($unsigned(forvar847))) : reg4200[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg4222 <= reg4182[(2'h3):(2'h2)];
                      reg4223 <= {(~&{{forvar809}})};
                      reg4224 <= ($signed(($unsigned(reg4218) - (-reg692))) ^~ reg730[(3'h4):(3'h4)]);
                      reg4225 <= $unsigned({{reg862}});
                    end
                end
            end
        end
      else
        begin
          for (forvar4171 = (1'h0); (forvar4171 < (2'h3)); forvar4171 = (forvar4171 + (1'h1)))
            begin
              for (forvar4172 = (1'h0); (forvar4172 < (2'h3)); forvar4172 = (forvar4172 + (1'h1)))
                begin
                  reg4173 <= ((forvar735[(3'h5):(1'h0)] ?
                          (reg703[(4'hb):(3'h5)] ?
                              $unsigned(reg747) : reg854[(4'hd):(4'ha)]) : $unsigned(((8'hb5) ?
                              reg728 : reg4210))) ?
                      $unsigned(($unsigned(reg705) ?
                          {(8'hb4)} : forvar735[(4'ha):(2'h2)])) : $unsigned(reg4197));
                  for (forvar4174 = (1'h0); (forvar4174 < (1'h1)); forvar4174 = (forvar4174 + (1'h1)))
                    begin
                      reg4175 <= reg845[(3'h5):(2'h2)];
                      reg4176 <= forvar681;
                    end
                  if ($unsigned($unsigned(($signed(reg802) ?
                      {forvar4209} : reg759[(3'h4):(1'h1)]))))
                    begin
                      reg4177 <= (reg690[(1'h1):(1'h0)] ^ (($signed(reg698) ?
                          (8'hb2) : (reg821 ? forvar716 : reg766)) >= (8'hb5)));
                    end
                  else
                    begin
                      reg4177 <= $signed((&reg4211[(4'hb):(3'h7)]));
                      reg4178 <= reg801[(4'hd):(3'h4)];
                      reg4179 <= $signed(forvar790[(3'h5):(2'h3)]);
                    end
                  reg4180 <= reg4192[(2'h2):(2'h2)];
                end
            end
          if ((reg808 ?
              $unsigned(({reg4218} ~^ (forvar791 | reg829))) : reg716))
            begin
              for (forvar4181 = (1'h0); (forvar4181 < (2'h2)); forvar4181 = (forvar4181 + (1'h1)))
                begin
                  reg4182 <= forvar715;
                  for (forvar4183 = (1'h0); (forvar4183 < (1'h1)); forvar4183 = (forvar4183 + (1'h1)))
                    begin
                      reg4184 <= forvar790[(3'h6):(3'h5)];
                      reg4185 <= reg827;
                      reg4186 <= $signed($unsigned((wire677[(3'h6):(1'h0)] + $signed(reg869))));
                    end
                  for (forvar4187 = (1'h0); (forvar4187 < (2'h3)); forvar4187 = (forvar4187 + (1'h1)))
                    begin
                      reg4188 <= forvar808;
                      reg4189 <= {reg750[(3'h5):(1'h0)]};
                      reg4190 <= forvar860[(1'h0):(1'h0)];
                    end
                  if (({(forvar4198 ?
                          $unsigned(reg4223) : forvar726)} * $unsigned(reg728[(3'h4):(3'h4)])))
                    begin
                      reg4191 <= $signed((~|forvar868[(2'h3):(1'h1)]));
                      reg4192 <= $unsigned(forvar681);
                      reg4193 <= ({$signed(reg4187[(4'h8):(3'h7)])} <<< (^~(^reg869[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg4191 <= reg784;
                      reg4192 <= (!$signed((8'ha0)));
                      reg4193 <= reg685[(1'h1):(1'h1)];
                      reg4194 <= (~|{$unsigned(reg4194[(3'h7):(3'h5)])});
                    end
                end
              for (forvar4195 = (1'h0); (forvar4195 < (1'h0)); forvar4195 = (forvar4195 + (1'h1)))
                begin
                  if (forvar773)
                    begin
                      reg4196 <= ($unsigned(reg695[(4'h8):(3'h4)]) * $signed($unsigned(reg740)));
                      reg4197 <= reg758;
                      reg4198 <= (-$unsigned(forvar719));
                      reg4199 <= {({forvar791} ~^ forvar799[(3'h6):(3'h4)])};
                    end
                  else
                    begin
                      reg4196 <= $unsigned($signed((^reg845[(1'h1):(1'h1)])));
                      reg4197 <= $signed($signed((!forvar4172[(3'h5):(2'h3)])));
                      reg4198 <= $signed($unsigned((!$signed(reg4200))));
                    end
                  for (forvar4200 = (1'h0); (forvar4200 < (1'h0)); forvar4200 = (forvar4200 + (1'h1)))
                    begin
                      reg4201 <= (reg717[(3'h7):(3'h6)] ?
                          ((~|(~reg711)) > forvar814) : (({reg4187} <= {forvar4187}) ?
                              ($signed(forvar799) ?
                                  $signed(forvar780) : ((8'ha9) ?
                                      reg711 : (8'ha2))) : $unsigned(((8'ha5) ^ forvar680))));
                      reg4202 <= reg800[(2'h2):(2'h2)];
                      reg4203 <= ((($signed(reg796) && (forvar860 <<< forvar859)) ?
                          reg819[(3'h6):(3'h6)] : $signed(((8'hb2) >>> forvar868))) != reg887);
                    end
                end
              if ({(~^(!(~|reg4206)))})
                begin
                  if (($signed($signed(reg4208[(3'h6):(2'h3)])) * (~&($signed(reg804) ?
                      reg733[(3'h6):(3'h6)] : $unsigned(reg799)))))
                    begin
                      reg4204 <= $signed((forvar844 ? reg4173 : (~^{reg758})));
                      reg4205 <= {(8'hac)};
                      reg4206 <= $unsigned({reg759[(1'h0):(1'h0)]});
                    end
                  else
                    begin
                      reg4204 <= $unsigned(reg867[(3'h6):(3'h4)]);
                    end
                  if ($signed($unsigned((~$unsigned(forvar4209)))))
                    begin
                      reg4207 <= reg817[(3'h4):(1'h0)];
                      reg4208 <= (($unsigned(forvar4191) - (reg4220 ?
                              reg4212[(4'h8):(1'h1)] : (forvar799 <<< (8'hb7)))) ?
                          $unsigned($unsigned((&reg801))) : $unsigned($signed($signed(reg776))));
                      reg4209 <= $signed($signed($signed(reg714[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg4207 <= reg760;
                      reg4208 <= (($unsigned(reg810[(2'h2):(1'h1)]) ?
                              $unsigned((forvar681 >> (8'hb3))) : ((&reg710) <= (&reg738))) ?
                          (-reg785) : $unsigned($signed(forvar735[(3'h4):(1'h0)])));
                      reg4209 <= (((8'ha2) > (^reg746)) >>> forvar831);
                      reg4210 <= (($signed((&reg4221)) << reg817[(1'h1):(1'h1)]) << $signed(reg877));
                    end
                end
              else
                begin
                  for (forvar4204 = (1'h0); (forvar4204 < (1'h1)); forvar4204 = (forvar4204 + (1'h1)))
                    begin
                      reg4205 <= reg878[(2'h3):(1'h0)];
                      reg4206 <= (+(({reg803} ?
                              $unsigned(reg4194) : (wire677 <= reg775)) ?
                          $signed((reg769 >>> reg733)) : reg820));
                      reg4207 <= $unsigned(reg769[(1'h1):(1'h1)]);
                    end
                  for (forvar4208 = (1'h0); (forvar4208 < (2'h2)); forvar4208 = (forvar4208 + (1'h1)))
                    begin
                      reg4209 <= reg728[(2'h2):(1'h0)];
                      reg4210 <= $unsigned((reg4207[(2'h2):(1'h0)] ^ reg4217[(2'h2):(1'h1)]));
                    end
                end
              for (forvar4211 = (1'h0); (forvar4211 < (1'h1)); forvar4211 = (forvar4211 + (1'h1)))
                begin
                  for (forvar4212 = (1'h0); (forvar4212 < (2'h2)); forvar4212 = (forvar4212 + (1'h1)))
                    begin
                      reg4213 <= $unsigned(reg869[(2'h2):(1'h1)]);
                      reg4214 <= reg755[(4'hf):(4'ha)];
                      reg4215 <= $signed((8'hb4));
                      reg4216 <= $signed(((~|((8'hb7) ? reg842 : reg885)) ?
                          forvar804[(4'h9):(4'h9)] : {$unsigned((8'hae))}));
                    end
                end
            end
          else
            begin
              if ($unsigned((($unsigned(reg741) ?
                      forvar681 : (reg755 ? reg871 : forvar4192)) ?
                  $signed($signed(forvar4171)) : $signed(forvar779))))
                begin
                  for (forvar4181 = (1'h0); (forvar4181 < (2'h3)); forvar4181 = (forvar4181 + (1'h1)))
                    begin
                      reg4182 <= $signed((~|(~|$unsigned(reg862))));
                      reg4183 <= reg4208[(3'h5):(2'h2)];
                    end
                  if (reg816[(1'h0):(1'h0)])
                    begin
                      reg4184 <= forvar4198;
                      reg4185 <= (^~$signed((8'hb8)));
                      reg4186 <= {(~^forvar710[(4'hb):(1'h1)])};
                    end
                  else
                    begin
                      reg4184 <= ((reg883 ?
                          (((8'hb9) ?
                              reg4204 : forvar682) || forvar4209) : (forvar874 && $unsigned(reg4200))) || (reg878[(2'h3):(2'h2)] <<< (|{reg766})));
                      reg4185 <= reg4222[(1'h0):(1'h0)];
                      reg4186 <= reg806;
                    end
                  if ((reg4201 ?
                      {$unsigned(((8'hb7) ?
                              (8'hba) : forvar4211))} : ($unsigned(reg828[(2'h2):(2'h2)]) ^~ $signed($signed(reg844)))))
                    begin
                      reg4187 <= $signed((reg776[(2'h2):(1'h0)] ?
                          (reg4224[(2'h3):(2'h3)] & (reg738 >>> reg745)) : $unsigned(reg750)));
                    end
                  else
                    begin
                      reg4187 <= (~(&$unsigned($signed(reg803))));
                      reg4188 <= (^~$signed((((8'ha3) << reg852) ?
                          $unsigned(reg736) : (forvar687 <<< reg742))));
                      reg4189 <= reg714;
                      reg4190 <= ((8'hb5) ?
                          (~$unsigned((reg702 <= forvar842))) : ($unsigned(reg861[(3'h6):(1'h0)]) == (|$signed(reg833))));
                    end
                end
              else
                begin
                  for (forvar4181 = (1'h0); (forvar4181 < (2'h3)); forvar4181 = (forvar4181 + (1'h1)))
                    begin
                      reg4182 <= reg4211;
                      reg4183 <= $unsigned($signed($signed((reg713 ?
                          reg737 : (8'hae)))));
                      reg4184 <= ($unsigned({$signed(reg4193)}) * (~|{reg810[(1'h1):(1'h0)]}));
                      reg4185 <= (^~forvar749);
                    end
                  reg4186 <= ((&(!$unsigned(reg839))) ? (8'ha5) : reg4220);
                  for (forvar4187 = (1'h0); (forvar4187 < (2'h2)); forvar4187 = (forvar4187 + (1'h1)))
                    begin
                      reg4188 <= $signed(forvar682[(1'h0):(1'h0)]);
                      reg4189 <= ((~^reg821[(1'h0):(1'h0)]) >>> reg855[(4'hf):(4'hd)]);
                      reg4190 <= (&$unsigned($unsigned((forvar689 ?
                          (8'h9e) : reg4209))));
                      reg4191 <= reg806;
                    end
                  for (forvar4192 = (1'h0); (forvar4192 < (2'h3)); forvar4192 = (forvar4192 + (1'h1)))
                    begin
                      reg4193 <= forvar682;
                      reg4194 <= forvar874[(3'h6):(3'h6)];
                      reg4195 <= (reg827[(4'h8):(3'h7)] >= $unsigned({(~&reg746)}));
                      reg4196 <= {({(reg4220 + wire676)} ?
                              (reg762[(1'h0):(1'h0)] ?
                                  (~^reg4197) : (&(8'ha9))) : (~&(reg801 != forvar838)))};
                    end
                end
              reg4197 <= $unsigned(($signed((^~reg4203)) > ((reg4217 ?
                      reg774 : reg700) ?
                  (-forvar4208) : $unsigned(forvar735))));
            end
        end
      for (forvar4226 = (1'h0); (forvar4226 < (2'h3)); forvar4226 = (forvar4226 + (1'h1)))
        begin
          if ((reg765 ?
              $unsigned(({forvar680} ?
                  forvar702 : (reg777 ?
                      reg761 : reg719))) : ($unsigned((reg717 ?
                      reg712 : (8'hb8))) ?
                  reg758 : (~(reg700 == reg856)))))
            begin
              for (forvar4227 = (1'h0); (forvar4227 < (2'h3)); forvar4227 = (forvar4227 + (1'h1)))
                begin
                  for (forvar4228 = (1'h0); (forvar4228 < (1'h0)); forvar4228 = (forvar4228 + (1'h1)))
                    begin
                      reg4229 <= ((reg774 ?
                          ((forvar837 ? reg862 : forvar706) ?
                              $unsigned(reg796) : reg826) : reg724) < $signed($unsigned(reg836[(4'h8):(3'h5)])));
                      reg4230 <= reg4209;
                      reg4231 <= $unsigned({(~&(^~reg4172))});
                      reg4232 <= forvar782;
                    end
                  for (forvar4233 = (1'h0); (forvar4233 < (2'h3)); forvar4233 = (forvar4233 + (1'h1)))
                    begin
                      reg4234 <= reg828[(3'h4):(2'h3)];
                      reg4235 <= $unsigned(reg714);
                      reg4236 <= $unsigned($signed(($signed(reg798) > (reg740 ?
                          reg746 : forvar778))));
                      reg4237 <= $unsigned((((wire678 <= (8'ha3)) ?
                          {reg820} : reg818) <= (!reg730[(4'hc):(3'h5)])));
                    end
                  if ((!reg865[(3'h6):(3'h5)]))
                    begin
                      reg4238 <= (($unsigned((reg698 <= reg766)) <<< (|$signed(reg730))) ?
                          $unsigned((((8'hab) ?
                              forvar860 : reg730) >> $unsigned(reg731))) : reg4205);
                    end
                  else
                    begin
                      reg4238 <= ($unsigned(forvar789) ?
                          ((reg849[(1'h0):(1'h0)] ?
                                  (forvar847 ?
                                      (8'hb2) : (8'hb9)) : $signed(reg770)) ?
                              $unsigned($unsigned(forvar716)) : (reg4185[(4'h8):(3'h6)] ~^ $signed(reg742))) : (({(8'ha7)} ?
                                  reg772[(3'h7):(3'h7)] : forvar4187) ?
                              {(&reg737)} : $unsigned($signed(reg805))));
                      reg4239 <= $unsigned(reg802);
                      reg4240 <= $signed(reg845);
                      reg4241 <= reg881[(1'h1):(1'h0)];
                    end
                end
              reg4242 <= reg857;
              reg4243 <= {reg684};
              if (reg721[(3'h5):(1'h1)])
                begin
                  for (forvar4244 = (1'h0); (forvar4244 < (2'h2)); forvar4244 = (forvar4244 + (1'h1)))
                    begin
                      reg4245 <= $unsigned(forvar809[(2'h3):(2'h2)]);
                      reg4246 <= ($signed(forvar734) || (&$signed(reg864[(4'hb):(4'ha)])));
                      reg4247 <= reg707;
                      reg4248 <= reg867[(1'h0):(1'h0)];
                    end
                  if ((reg4234[(1'h0):(1'h0)] ?
                      (((+reg4232) >= (reg728 != forvar4227)) - (^~{(8'ha8)})) : reg772[(1'h0):(1'h0)]))
                    begin
                      reg4249 <= $unsigned(forvar848[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg4249 <= ($signed($unsigned(wire677[(3'h7):(2'h3)])) <<< (8'hb0));
                      reg4250 <= $unsigned(((reg761 > (~|forvar844)) & {reg4239}));
                    end
                end
              else
                begin
                  if ((-$signed($unsigned(reg707))))
                    begin
                      reg4244 <= forvar832[(3'h7):(1'h0)];
                      reg4245 <= (~|forvar842[(4'h9):(3'h6)]);
                    end
                  else
                    begin
                      reg4244 <= $unsigned((reg839[(4'h8):(1'h1)] ?
                          forvar709[(4'h8):(2'h3)] : (reg784 ?
                              $signed(forvar689) : reg841)));
                      reg4245 <= reg4213[(1'h1):(1'h1)];
                      reg4246 <= ($signed($signed($signed(reg824))) ?
                          reg723 : (~$unsigned($signed(reg771))));
                      reg4247 <= ($unsigned($unsigned((forvar4216 + reg759))) ^ $signed(reg709[(1'h1):(1'h0)]));
                    end
                  if (forvar4244)
                    begin
                      reg4248 <= ((((forvar711 ?
                          reg796 : forvar4209) > (~reg727)) ^~ reg842) + reg744[(4'hc):(4'hb)]);
                      reg4249 <= (reg4192 || ((reg751[(3'h4):(3'h4)] ?
                          $unsigned(forvar4226) : $signed(reg837)) <<< $signed((reg769 ?
                          reg4250 : (8'haa)))));
                      reg4250 <= (-((8'h9e) >>> (~(forvar4228 | reg710))));
                      reg4251 <= ((reg4221 == (8'hb6)) * {($unsigned((8'had)) || ((8'hba) ^~ reg725))});
                    end
                  else
                    begin
                      reg4248 <= ($signed(reg751[(3'h7):(2'h3)]) <= ((|$signed((8'hb6))) <= (forvar829 ?
                          (|(8'hb5)) : (reg711 ? reg726 : reg747))));
                      reg4249 <= ((reg4194 ?
                              ({forvar718} ?
                                  reg4244 : reg884[(2'h3):(1'h1)]) : ((~|reg840) ?
                                  {(8'ha7)} : ((8'had) ? reg855 : reg4212))) ?
                          ((^~$signed(forvar842)) >= {$signed(reg4220)}) : {$unsigned($unsigned(forvar702))});
                    end
                  for (forvar4252 = (1'h0); (forvar4252 < (2'h2)); forvar4252 = (forvar4252 + (1'h1)))
                    begin
                      reg4253 <= $signed(forvar866[(1'h1):(1'h0)]);
                      reg4254 <= $unsigned($unsigned(($signed(forvar764) ?
                          {reg720} : (forvar682 ? forvar4252 : reg703))));
                      reg4255 <= $unsigned((wire677 ?
                          reg797 : ($signed(reg766) == (reg4180 ?
                              reg790 : reg4198))));
                      reg4256 <= $signed($signed($signed(forvar702[(3'h5):(2'h3)])));
                    end
                  if (wire678[(3'h6):(3'h5)])
                    begin
                      reg4257 <= {$unsigned($unsigned((reg806 ?
                              reg4202 : reg851)))};
                      reg4258 <= (forvar4233 && ((8'had) * ($signed(reg729) * reg4232)));
                      reg4259 <= {reg4208};
                      reg4260 <= reg883;
                    end
                  else
                    begin
                      reg4257 <= $signed($signed(reg848[(1'h0):(1'h0)]));
                    end
                end
            end
          else
            begin
              for (forvar4227 = (1'h0); (forvar4227 < (2'h3)); forvar4227 = (forvar4227 + (1'h1)))
                begin
                  for (forvar4228 = (1'h0); (forvar4228 < (2'h3)); forvar4228 = (forvar4228 + (1'h1)))
                    begin
                      reg4229 <= (reg767[(4'hd):(2'h3)] ?
                          $unsigned(reg4254) : {(+forvar809[(3'h4):(2'h3)])});
                    end
                  for (forvar4230 = (1'h0); (forvar4230 < (1'h1)); forvar4230 = (forvar4230 + (1'h1)))
                    begin
                      reg4231 <= {(^~$signed((!forvar859)))};
                      reg4232 <= $signed((forvar831 << {(^~(8'hb8))}));
                      reg4233 <= reg723[(1'h1):(1'h1)];
                      reg4234 <= ((((forvar803 == reg4244) <= (reg4256 ?
                              forvar4174 : forvar731)) >> (~|(reg702 ?
                              (8'ha0) : reg872))) ?
                          reg800 : forvar837[(1'h0):(1'h0)]);
                    end
                  for (forvar4235 = (1'h0); (forvar4235 < (1'h0)); forvar4235 = (forvar4235 + (1'h1)))
                    begin
                      reg4236 <= $unsigned(forvar4226[(3'h6):(1'h0)]);
                    end
                end
              for (forvar4237 = (1'h0); (forvar4237 < (1'h0)); forvar4237 = (forvar4237 + (1'h1)))
                begin
                  if (reg717)
                    begin
                      reg4238 <= ((((reg4235 != reg690) >> {(8'had)}) ?
                          {$unsigned(reg721)} : (8'hba)) <<< (reg722 ?
                          reg832[(2'h2):(2'h2)] : (~|reg884)));
                      reg4239 <= $unsigned(({$unsigned((8'hb6))} || $signed($unsigned(forvar837))));
                      reg4240 <= reg4175;
                      reg4241 <= (~|(reg806 ^ (reg4200 ~^ reg813[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg4238 <= $unsigned($unsigned((~&((8'ha8) >= reg710))));
                      reg4239 <= ((forvar829 > (-(reg737 * reg850))) | forvar4192);
                    end
                  reg4242 <= (^reg4255);
                  if (($unsigned($signed(reg716[(2'h2):(2'h2)])) ?
                      $signed((|{reg4247})) : (-$unsigned(reg4250[(3'h5):(1'h0)]))))
                    begin
                      reg4243 <= (reg722 << forvar875[(3'h5):(2'h3)]);
                      reg4244 <= $signed({$unsigned((reg851 ?
                              forvar808 : reg777))});
                    end
                  else
                    begin
                      reg4243 <= forvar4208[(3'h6):(3'h4)];
                    end
                  for (forvar4245 = (1'h0); (forvar4245 < (2'h3)); forvar4245 = (forvar4245 + (1'h1)))
                    begin
                      reg4246 <= $signed((reg716 >= $signed((reg760 ?
                          reg787 : reg4173))));
                    end
                end
              if (((forvar726 ?
                      ((|reg683) ?
                          reg835[(4'hf):(4'he)] : reg757) : $unsigned((~reg729))) ?
                  (!reg708[(3'h4):(1'h0)]) : $signed({{forvar715}})))
                begin
                  if ($signed($unsigned({(reg708 ? reg4248 : forvar832)})))
                    begin
                      reg4247 <= $signed(reg862[(4'h8):(3'h7)]);
                    end
                  else
                    begin
                      reg4247 <= forvar829[(4'he):(2'h2)];
                    end
                  if ($signed(reg4178))
                    begin
                      reg4248 <= forvar680[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg4248 <= ((reg876 ?
                          (!$signed(forvar875)) : forvar789) || forvar4214[(2'h3):(2'h2)]);
                      reg4249 <= $signed($signed(((reg4256 ?
                          forvar792 : forvar733) >= {forvar837})));
                    end
                end
              else
                begin
                  for (forvar4247 = (1'h0); (forvar4247 < (2'h2)); forvar4247 = (forvar4247 + (1'h1)))
                    begin
                      reg4248 <= $unsigned({reg820});
                    end
                  reg4249 <= {reg843};
                  if ((~((reg4194[(4'hc):(2'h2)] ?
                          (reg726 ? reg692 : forvar4174) : $unsigned(reg849)) ?
                      (!reg883[(3'h7):(2'h3)]) : (reg814 <= ((8'ha4) ^ forvar711)))))
                    begin
                      reg4250 <= ({$unsigned(reg696)} != reg4244);
                      reg4251 <= (reg761[(3'h5):(2'h3)] ?
                          (reg4237 << reg4242[(1'h1):(1'h1)]) : (^~(reg722[(4'hb):(2'h3)] <<< $unsigned(reg743))));
                      reg4252 <= ((+forvar830[(3'h7):(3'h4)]) ?
                          $unsigned(($unsigned(reg871) <<< $unsigned((8'ha1)))) : forvar729[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg4250 <= $signed(((reg871 ?
                          $unsigned((8'hb6)) : (forvar715 >>> reg819)) != $signed($signed(reg843))));
                      reg4251 <= ((|(forvar729 | $unsigned((8'h9e)))) <<< (((forvar4226 != reg4233) - (reg877 * reg843)) >= $unsigned($unsigned(reg4238))));
                    end
                end
              reg4253 <= (~reg4250);
            end
          for (forvar4261 = (1'h0); (forvar4261 < (1'h1)); forvar4261 = (forvar4261 + (1'h1)))
            begin
              if ($unsigned(reg4186))
                begin
                  if (forvar4244[(1'h0):(1'h0)])
                    begin
                      reg4262 <= (((~&forvar4174[(4'he):(1'h0)]) + (reg769 >> {(8'ha3)})) << ((~&(^(8'had))) ?
                          forvar4214 : $unsigned((reg716 ~^ reg4205))));
                    end
                  else
                    begin
                      reg4262 <= (reg719 ^~ $unsigned({$unsigned((8'ha1))}));
                    end
                  if ($unsigned($unsigned($signed((reg788 ?
                      forvar782 : reg769)))))
                    begin
                      reg4263 <= (~|$signed(((forvar4230 != reg737) ?
                          (reg848 << reg786) : {reg840})));
                      reg4264 <= reg4208[(2'h2):(1'h0)];
                      reg4265 <= (!reg717);
                    end
                  else
                    begin
                      reg4263 <= $unsigned($unsigned((^~(forvar710 ?
                          reg4230 : forvar844))));
                    end
                  for (forvar4266 = (1'h0); (forvar4266 < (2'h2)); forvar4266 = (forvar4266 + (1'h1)))
                    begin
                      reg4267 <= (reg4172[(3'h6):(1'h0)] ?
                          $unsigned(reg765) : $signed((forvar4191[(4'ha):(3'h4)] ?
                              forvar729[(3'h4):(3'h4)] : ((8'haa) ?
                                  (8'ha4) : reg873))));
                    end
                  for (forvar4268 = (1'h0); (forvar4268 < (2'h3)); forvar4268 = (forvar4268 + (1'h1)))
                    begin
                      reg4269 <= ((^~reg872) == $unsigned(reg750[(3'h4):(2'h3)]));
                      reg4270 <= (-(($unsigned(reg696) ?
                          (|(8'hb1)) : $signed(forvar4181)) ^ ((reg698 ^ reg887) ?
                          (~|forvar709) : forvar847)));
                      reg4271 <= $unsigned($signed($unsigned((forvar4202 <<< reg4210))));
                    end
                end
              else
                begin
                  for (forvar4262 = (1'h0); (forvar4262 < (2'h2)); forvar4262 = (forvar4262 + (1'h1)))
                    begin
                      reg4263 <= $unsigned((((~^reg721) ?
                              reg759 : $signed(forvar804)) ?
                          forvar852 : (8'h9f)));
                      reg4264 <= reg809[(3'h6):(3'h5)];
                      reg4265 <= (reg796 ?
                          $signed(($signed(reg4197) ?
                              reg773 : (&reg760))) : {reg766});
                    end
                end
              for (forvar4272 = (1'h0); (forvar4272 < (2'h2)); forvar4272 = (forvar4272 + (1'h1)))
                begin
                  if (reg4244)
                    begin
                      reg4273 <= $signed(reg697);
                      reg4274 <= $unsigned((-(^reg813)));
                    end
                  else
                    begin
                      reg4273 <= reg806;
                      reg4274 <= forvar870[(4'hf):(1'h0)];
                      reg4275 <= reg4199;
                      reg4276 <= reg717;
                    end
                end
              for (forvar4277 = (1'h0); (forvar4277 < (1'h1)); forvar4277 = (forvar4277 + (1'h1)))
                begin
                  reg4278 <= ((8'ha9) <<< (((8'h9c) != forvar792[(4'h9):(3'h4)]) ?
                      ((^reg698) ^~ (!(8'ha4))) : (~|(|reg831))));
                  for (forvar4279 = (1'h0); (forvar4279 < (1'h0)); forvar4279 = (forvar4279 + (1'h1)))
                    begin
                      reg4280 <= reg802;
                      reg4281 <= (~{($signed(reg869) <<< (reg4200 ?
                              (8'hb9) : (8'haf)))});
                    end
                end
              if (reg884)
                begin
                  for (forvar4282 = (1'h0); (forvar4282 < (2'h3)); forvar4282 = (forvar4282 + (1'h1)))
                    begin
                      reg4283 <= reg4253[(1'h1):(1'h0)];
                      reg4284 <= reg4252[(1'h1):(1'h0)];
                    end
                  for (forvar4285 = (1'h0); (forvar4285 < (2'h3)); forvar4285 = (forvar4285 + (1'h1)))
                    begin
                      reg4286 <= forvar822[(3'h5):(2'h2)];
                      reg4287 <= ((reg4252[(3'h4):(2'h2)] * ($signed(reg781) ?
                              (reg4221 ?
                                  reg4172 : forvar790) : $signed(reg828))) ?
                          ((^{reg796}) ?
                              $unsigned(forvar709[(3'h5):(1'h0)]) : (&$signed(reg830))) : $unsigned(reg770));
                      reg4288 <= {$unsigned(reg4213[(2'h2):(2'h2)])};
                      reg4289 <= $signed(reg4204);
                    end
                  if ($signed($signed((~$unsigned(forvar4261)))))
                    begin
                      reg4290 <= forvar773;
                    end
                  else
                    begin
                      reg4290 <= $unsigned(wire677[(3'h4):(2'h2)]);
                      reg4291 <= reg853;
                    end
                  reg4292 <= ($signed({(reg777 ?
                          (8'h9e) : forvar837)}) || forvar831[(1'h0):(1'h0)]);
                end
              else
                begin
                  if (($signed(reg4175) ?
                      reg4225 : $signed((~(reg883 - forvar754)))))
                    begin
                      reg4282 <= (($signed($signed(forvar842)) ?
                              ((forvar681 ? reg4204 : reg4197) ?
                                  $signed(reg4242) : (reg739 >>> reg4252)) : {(!reg4208)}) ?
                          reg709 : $unsigned($signed(((8'had) ?
                              forvar4262 : forvar778))));
                    end
                  else
                    begin
                      reg4282 <= $unsigned(reg4236);
                      reg4283 <= reg746;
                      reg4284 <= forvar719;
                    end
                  reg4285 <= forvar763;
                  for (forvar4286 = (1'h0); (forvar4286 < (1'h0)); forvar4286 = (forvar4286 + (1'h1)))
                    begin
                      reg4287 <= (^{$signed((|reg4206))});
                      reg4288 <= (reg857[(1'h1):(1'h1)] ?
                          ($unsigned(reg815) ?
                              (8'hb3) : ((&reg830) ^ $signed(forvar792))) : reg4241);
                      reg4289 <= $unsigned($unsigned(((~&reg4255) ?
                          {reg826} : reg695)));
                      reg4290 <= $signed({forvar4198[(1'h0):(1'h0)]});
                    end
                end
            end
        end
      if ($signed((((|(8'haf)) ?
              (reg742 || forvar724) : (reg4215 << forvar754)) ?
          forvar680[(3'h6):(1'h1)] : ((^reg4284) ? reg4263 : (+reg716)))))
        begin
          if (forvar709[(2'h2):(1'h1)])
            begin
              for (forvar4293 = (1'h0); (forvar4293 < (1'h1)); forvar4293 = (forvar4293 + (1'h1)))
                begin
                  reg4294 <= ((+(~$unsigned(reg4238))) ?
                      (^$unsigned($signed(reg762))) : (forvar4192 < reg846[(3'h7):(2'h3)]));
                  for (forvar4295 = (1'h0); (forvar4295 < (1'h0)); forvar4295 = (forvar4295 + (1'h1)))
                    begin
                      reg4296 <= forvar814;
                    end
                end
              reg4297 <= $unsigned((reg4263 | forvar879));
              for (forvar4298 = (1'h0); (forvar4298 < (2'h2)); forvar4298 = (forvar4298 + (1'h1)))
                begin
                  for (forvar4299 = (1'h0); (forvar4299 < (2'h2)); forvar4299 = (forvar4299 + (1'h1)))
                    begin
                      reg4300 <= forvar4209;
                      reg4301 <= reg878[(4'h9):(4'h9)];
                      reg4302 <= reg699;
                    end
                  if ((|(reg4287 && (~$unsigned((8'hb2))))))
                    begin
                      reg4303 <= reg4292;
                      reg4304 <= $unsigned((reg705 ?
                          ({reg4217} + forvar4262[(1'h0):(1'h0)]) : $signed($signed((8'ha4)))));
                    end
                  else
                    begin
                      reg4303 <= ($signed((^reg685)) ~^ $signed((((8'had) ?
                          forvar822 : reg848) && (reg4194 ?
                          (8'ha9) : (8'hb7)))));
                      reg4304 <= $signed(forvar4237);
                    end
                  for (forvar4305 = (1'h0); (forvar4305 < (1'h1)); forvar4305 = (forvar4305 + (1'h1)))
                    begin
                      reg4306 <= (~&reg4285[(3'h4):(2'h2)]);
                      reg4307 <= reg4255[(4'hd):(1'h0)];
                      reg4308 <= $unsigned($signed(($signed(forvar688) ?
                          reg685[(2'h2):(1'h0)] : (reg798 > reg4217))));
                    end
                  for (forvar4309 = (1'h0); (forvar4309 < (2'h3)); forvar4309 = (forvar4309 + (1'h1)))
                    begin
                      reg4310 <= ({$signed((reg4201 ?
                              reg833 : reg819))} || (~|((+reg4206) <<< (^forvar4295))));
                      reg4311 <= $signed((forvar4277[(3'h5):(1'h0)] | $signed($signed(reg787))));
                      reg4312 <= ($unsigned($signed($signed(forvar4230))) != $unsigned(({reg693} < forvar847[(2'h3):(2'h2)])));
                      reg4313 <= $unsigned($signed($unsigned(reg807)));
                    end
                end
              reg4314 <= {$unsigned({$unsigned(reg4297)})};
            end
          else
            begin
              for (forvar4293 = (1'h0); (forvar4293 < (2'h2)); forvar4293 = (forvar4293 + (1'h1)))
                begin
                  if ({((^$signed(forvar726)) || wire676)})
                    begin
                      reg4294 <= (($signed($signed(reg769)) << (~(8'h9c))) != (($unsigned(reg4291) ?
                              reg781[(4'hc):(4'h8)] : (forvar4174 ~^ reg851)) ?
                          ($signed(forvar874) ~^ $unsigned(forvar4279)) : (-reg4313)));
                      reg4295 <= reg4213[(1'h1):(1'h0)];
                      reg4296 <= ((reg814[(1'h0):(1'h0)] ?
                              (reg833[(2'h3):(1'h1)] >>> $unsigned(forvar809)) : reg4187[(4'h8):(3'h5)]) ?
                          {$signed((+(8'ha0)))} : (~|reg710));
                    end
                  else
                    begin
                      reg4294 <= ($signed($unsigned($unsigned(reg4195))) ?
                          (^$unsigned(reg810)) : reg4252[(1'h0):(1'h0)]);
                      reg4295 <= (8'hb0);
                    end
                  if ((|({(forvar789 ?
                          reg4201 : (8'ha2))} & (((8'hb7) != reg4215) != (reg4285 || reg744)))))
                    begin
                      reg4297 <= $signed({$signed(reg4249)});
                      reg4298 <= reg4243;
                      reg4299 <= $signed((^((forvar4192 ? reg845 : forvar829) ?
                          (!forvar4295) : $signed(reg873))));
                      reg4300 <= $signed({reg4306});
                    end
                  else
                    begin
                      reg4297 <= reg803[(4'h8):(2'h2)];
                    end
                  reg4301 <= (|$unsigned($signed(reg729[(1'h0):(1'h0)])));
                  if ((8'ha0))
                    begin
                      reg4302 <= ($signed((+(~^reg692))) ?
                          (reg803 - (~^$unsigned(reg705))) : $signed(({reg4220} ?
                              $unsigned((8'hb9)) : $signed(reg4271))));
                    end
                  else
                    begin
                      reg4302 <= {$unsigned({reg4282})};
                      reg4303 <= forvar852;
                    end
                end
              for (forvar4304 = (1'h0); (forvar4304 < (2'h3)); forvar4304 = (forvar4304 + (1'h1)))
                begin
                  reg4305 <= (8'ha0);
                  reg4306 <= $signed((~|((8'hb2) ?
                      (reg753 ? reg691 : reg756) : $signed(forvar4298))));
                end
            end
          if ($signed(({reg4230} >> reg4310[(1'h1):(1'h1)])))
            begin
              for (forvar4315 = (1'h0); (forvar4315 < (2'h2)); forvar4315 = (forvar4315 + (1'h1)))
                begin
                  for (forvar4316 = (1'h0); (forvar4316 < (2'h3)); forvar4316 = (forvar4316 + (1'h1)))
                    begin
                      reg4317 <= $unsigned((|{(forvar4171 ? reg819 : reg821)}));
                    end
                end
              for (forvar4318 = (1'h0); (forvar4318 < (2'h2)); forvar4318 = (forvar4318 + (1'h1)))
                begin
                  reg4319 <= reg873[(1'h1):(1'h0)];
                  for (forvar4320 = (1'h0); (forvar4320 < (1'h0)); forvar4320 = (forvar4320 + (1'h1)))
                    begin
                      reg4321 <= (reg767 ^~ (^$signed((reg783 ?
                          reg4210 : (8'ha3)))));
                      reg4322 <= $signed({$signed($signed(reg733))});
                      reg4323 <= ($signed(reg4215[(3'h7):(1'h0)]) ?
                          reg725 : (8'hae));
                    end
                  reg4324 <= (~(-forvar4212));
                  reg4325 <= $signed(((reg797[(3'h4):(3'h4)] ^ (reg848 - reg885)) >>> ($unsigned(reg4260) + $signed((8'hac)))));
                end
            end
          else
            begin
              for (forvar4315 = (1'h0); (forvar4315 < (1'h1)); forvar4315 = (forvar4315 + (1'h1)))
                begin
                  for (forvar4316 = (1'h0); (forvar4316 < (1'h1)); forvar4316 = (forvar4316 + (1'h1)))
                    begin
                      reg4317 <= {$signed((~|(reg691 ? reg766 : forvar4181)))};
                      reg4318 <= $unsigned((reg4213[(2'h2):(1'h1)] ?
                          reg705[(3'h4):(1'h0)] : reg826));
                      reg4319 <= forvar733;
                    end
                  reg4320 <= (8'ha9);
                end
              for (forvar4321 = (1'h0); (forvar4321 < (1'h1)); forvar4321 = (forvar4321 + (1'h1)))
                begin
                  for (forvar4322 = (1'h0); (forvar4322 < (2'h3)); forvar4322 = (forvar4322 + (1'h1)))
                    begin
                      reg4323 <= (reg4178 ?
                          forvar875[(1'h1):(1'h1)] : (~&(8'ha7)));
                    end
                end
            end
          reg4326 <= {$unsigned(forvar687)};
        end
      else
        begin
          for (forvar4293 = (1'h0); (forvar4293 < (1'h1)); forvar4293 = (forvar4293 + (1'h1)))
            begin
              reg4294 <= reg4218;
              for (forvar4295 = (1'h0); (forvar4295 < (2'h3)); forvar4295 = (forvar4295 + (1'h1)))
                begin
                  for (forvar4296 = (1'h0); (forvar4296 < (1'h1)); forvar4296 = (forvar4296 + (1'h1)))
                    begin
                      reg4297 <= reg4255[(1'h1):(1'h0)];
                      reg4298 <= forvar4272[(1'h0):(1'h0)];
                    end
                  for (forvar4299 = (1'h0); (forvar4299 < (1'h1)); forvar4299 = (forvar4299 + (1'h1)))
                    begin
                      reg4300 <= reg4317;
                      reg4301 <= (((forvar4198 + reg685) ?
                              {{reg736}} : forvar868) ?
                          (forvar724[(4'h9):(3'h7)] ?
                              (-reg4264[(3'h4):(1'h0)]) : (reg4185[(3'h6):(2'h3)] != reg800)) : (^reg800));
                      reg4302 <= ($unsigned({(reg700 ?
                              reg759 : (8'hac))}) == (|$unsigned(forvar838)));
                      reg4303 <= $signed({($signed(reg824) ?
                              $signed(reg853) : forvar837)});
                    end
                  for (forvar4304 = (1'h0); (forvar4304 < (1'h1)); forvar4304 = (forvar4304 + (1'h1)))
                    begin
                      reg4305 <= $unsigned(forvar814[(3'h5):(2'h3)]);
                    end
                  reg4306 <= reg702[(1'h1):(1'h0)];
                end
            end
          for (forvar4307 = (1'h0); (forvar4307 < (1'h1)); forvar4307 = (forvar4307 + (1'h1)))
            begin
              for (forvar4308 = (1'h0); (forvar4308 < (1'h1)); forvar4308 = (forvar4308 + (1'h1)))
                begin
                  for (forvar4309 = (1'h0); (forvar4309 < (1'h0)); forvar4309 = (forvar4309 + (1'h1)))
                    begin
                      reg4310 <= forvar709;
                    end
                end
              if ((((~^(&forvar875)) ?
                  (-$unsigned(forvar879)) : forvar733) && $signed($unsigned((reg699 ?
                  reg4306 : forvar4172)))))
                begin
                  for (forvar4311 = (1'h0); (forvar4311 < (1'h0)); forvar4311 = (forvar4311 + (1'h1)))
                    begin
                      reg4312 <= ((^{forvar842[(4'h9):(4'h8)]}) ?
                          forvar773 : $unsigned((8'hb6)));
                      reg4313 <= $unsigned($unsigned((((8'hb7) - forvar763) * ((8'h9e) ^~ forvar4209))));
                      reg4314 <= (+$unsigned(reg748));
                    end
                end
              else
                begin
                  reg4311 <= (~^reg740[(3'h5):(2'h2)]);
                end
              for (forvar4315 = (1'h0); (forvar4315 < (1'h1)); forvar4315 = (forvar4315 + (1'h1)))
                begin
                  if ((^~{$unsigned($signed(reg4253))}))
                    begin
                      reg4316 <= {(((reg4296 * reg698) ?
                              (reg852 ?
                                  reg797 : (8'h9c)) : (forvar4205 ~^ forvar4235)) * ((~reg867) || $unsigned(reg758)))};
                    end
                  else
                    begin
                      reg4316 <= reg4229[(4'h8):(2'h3)];
                      reg4317 <= (~|({reg786[(3'h4):(2'h3)]} ?
                          $unsigned((reg863 ^~ reg4284)) : ((reg774 >> reg853) ?
                              (~^reg4260) : $unsigned(forvar707))));
                      reg4318 <= $unsigned((~|(+$unsigned(forvar4171))));
                      reg4319 <= ({(~|$unsigned(reg4300))} <<< {$signed((!reg878))});
                    end
                  for (forvar4320 = (1'h0); (forvar4320 < (1'h1)); forvar4320 = (forvar4320 + (1'h1)))
                    begin
                      reg4321 <= reg849;
                      reg4322 <= ($unsigned(($signed(reg4294) ?
                              reg695[(3'h7):(2'h2)] : (reg4245 | forvar754))) ?
                          (($unsigned(forvar724) ?
                                  $signed(reg775) : $signed((8'hb0))) ?
                              (8'ha6) : reg876) : $signed({(reg4199 ?
                                  reg739 : wire676)}));
                      reg4323 <= reg692;
                    end
                end
              for (forvar4324 = (1'h0); (forvar4324 < (2'h3)); forvar4324 = (forvar4324 + (1'h1)))
                begin
                  if ((reg4281 ~^ (reg4175 ^ reg723)))
                    begin
                      reg4325 <= $signed(wire677[(2'h3):(2'h2)]);
                      reg4326 <= (reg4235[(1'h1):(1'h1)] < ($signed((~^reg783)) >>> $unsigned({forvar797})));
                      reg4327 <= (^(~|(reg4244[(1'h0):(1'h0)] ^ $unsigned(reg4205))));
                      reg4328 <= reg4219[(3'h6):(3'h6)];
                    end
                  else
                    begin
                      reg4325 <= reg693;
                      reg4326 <= $unsigned(reg4251[(3'h5):(1'h0)]);
                      reg4327 <= forvar803[(1'h0):(1'h0)];
                    end
                  reg4329 <= (~forvar782);
                  for (forvar4330 = (1'h0); (forvar4330 < (1'h1)); forvar4330 = (forvar4330 + (1'h1)))
                    begin
                      reg4331 <= reg850;
                      reg4332 <= (reg770 ?
                          (&$unsigned((reg709 ?
                              (8'hb1) : forvar4262))) : $signed(forvar804));
                      reg4333 <= $signed((forvar779[(1'h1):(1'h0)] >>> ((!(8'had)) << (~|forvar681))));
                      reg4334 <= $signed({((+reg4270) ~^ forvar831)});
                    end
                end
            end
        end
    end
  assign wire4335 = (~{((|forvar4299) <<< forvar782)});
  assign wire4336 = (((reg4175 ?
                        (forvar4307 << (8'ha3)) : reg772) >>> {(+reg4199)}) <<< reg727[(4'hc):(4'hb)]);
  module4337 modinst7332 (.y(wire7331), .wire4338(reg4197), .wire4339(forvar4315), .wire4340(reg882), .wire4341(reg873), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar7333 = (1'h0); (forvar7333 < (2'h2)); forvar7333 = (forvar7333 + (1'h1)))
        begin
          for (forvar7334 = (1'h0); (forvar7334 < (2'h3)); forvar7334 = (forvar7334 + (1'h1)))
            begin
              for (forvar7335 = (1'h0); (forvar7335 < (1'h1)); forvar7335 = (forvar7335 + (1'h1)))
                begin
                  if (forvar4285[(2'h3):(1'h1)])
                    begin
                      reg7336 <= ($signed($unsigned($signed(reg730))) ?
                          forvar724[(2'h2):(1'h1)] : (+(forvar4202 ?
                              $unsigned(forvar814) : (reg880 ?
                                  (8'hb1) : (8'hb0)))));
                      reg7337 <= {reg855};
                      reg7338 <= $signed($signed({(reg709 - forvar4252)}));
                    end
                  else
                    begin
                      reg7336 <= forvar4268[(1'h1):(1'h1)];
                      reg7337 <= $unsigned({$signed((+forvar4315))});
                      reg7338 <= $signed(((-(forvar4293 ^~ reg819)) ?
                          ((forvar4311 << (8'ha4)) ?
                              reg746[(3'h4):(3'h4)] : reg4250[(1'h0):(1'h0)]) : $unsigned((reg4229 ?
                              (8'ha4) : reg741))));
                    end
                end
              for (forvar7339 = (1'h0); (forvar7339 < (2'h2)); forvar7339 = (forvar7339 + (1'h1)))
                begin
                  reg7340 <= reg738;
                  for (forvar7341 = (1'h0); (forvar7341 < (2'h2)); forvar7341 = (forvar7341 + (1'h1)))
                    begin
                      reg7342 <= ((reg801[(4'hc):(4'h8)] | forvar729) == reg842[(1'h0):(1'h0)]);
                      reg7343 <= (reg7340 ?
                          {(8'ha6)} : (^~reg760[(2'h3):(2'h3)]));
                      reg7344 <= (~^reg710[(1'h1):(1'h1)]);
                    end
                  for (forvar7345 = (1'h0); (forvar7345 < (1'h0)); forvar7345 = (forvar7345 + (1'h1)))
                    begin
                      reg7346 <= $unsigned((forvar879[(3'h5):(2'h2)] && $signed((|reg727))));
                    end
                  if ($signed(reg4244))
                    begin
                      reg7347 <= ($signed(reg721[(4'h9):(3'h5)]) ^~ $unsigned($unsigned($signed(reg4191))));
                    end
                  else
                    begin
                      reg7347 <= reg4259[(1'h1):(1'h0)];
                      reg7348 <= reg817[(2'h3):(1'h0)];
                      reg7349 <= forvar715[(3'h5):(3'h5)];
                    end
                end
              if (($signed($signed((8'hb1))) ?
                  forvar682[(2'h2):(2'h2)] : ($signed({reg800}) == reg4329[(1'h0):(1'h0)])))
                begin
                  if (forvar4268[(3'h7):(3'h4)])
                    begin
                      reg7350 <= ($unsigned(reg858[(3'h7):(3'h4)]) ^~ (forvar767 ^ ((reg4280 && (8'hac)) ?
                          $unsigned(reg697) : (8'hb2))));
                      reg7351 <= ((^~((reg4248 ? reg865 : forvar790) ?
                              (reg4275 + reg807) : (reg886 ?
                                  reg877 : reg4175))) ?
                          reg871 : reg747[(1'h0):(1'h0)]);
                      reg7352 <= $unsigned($unsigned((^~(reg4221 >>> reg685))));
                      reg7353 <= (($signed(forvar4320[(2'h2):(2'h2)]) ?
                              forvar4216 : forvar734) ?
                          (~(&$signed(reg800))) : $unsigned(reg4301[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg7350 <= forvar4295[(4'hb):(1'h1)];
                      reg7351 <= $unsigned($signed($signed(((8'hb4) ?
                          reg827 : reg867))));
                      reg7352 <= $signed((-$unsigned($unsigned(reg752))));
                    end
                  for (forvar7354 = (1'h0); (forvar7354 < (2'h2)); forvar7354 = (forvar7354 + (1'h1)))
                    begin
                      reg7355 <= $unsigned(($unsigned(forvar830) ^~ ((reg773 >= reg738) & $signed(reg4300))));
                      reg7356 <= ((($unsigned(forvar7341) > reg4276) ?
                              (~&(^reg867)) : ({reg4184} == $signed(reg4260))) ?
                          reg4190 : (forvar4192[(1'h0):(1'h0)] ?
                              forvar4286[(4'h8):(2'h3)] : {(~reg715)}));
                      reg7357 <= (&((reg4281 >>> reg4318[(4'ha):(4'ha)]) ?
                          ((forvar702 - forvar797) ?
                              (reg4200 ?
                                  reg845 : (8'h9e)) : wire4336[(1'h1):(1'h0)]) : reg4283[(2'h3):(1'h0)]));
                      reg7358 <= wire7331;
                    end
                  for (forvar7359 = (1'h0); (forvar7359 < (2'h3)); forvar7359 = (forvar7359 + (1'h1)))
                    begin
                      reg7360 <= reg4219[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if (($unsigned(((reg795 || reg4174) ?
                      ((8'hb4) ? reg4205 : (8'ha5)) : ((8'ha8) ?
                          reg4255 : reg4187))) - wire678))
                    begin
                      reg7350 <= {(|reg7346)};
                    end
                  else
                    begin
                      reg7350 <= (~&{forvar7359[(3'h4):(3'h4)]});
                      reg7351 <= {$signed(forvar4174)};
                      reg7352 <= (^~reg4321[(1'h1):(1'h1)]);
                      reg7353 <= ((~&$unsigned(reg708)) ? reg4287 : reg685);
                    end
                  reg7354 <= (($signed((reg7360 | (8'ha3))) == forvar749) ?
                      (^~$signed((~reg693))) : (^~$unsigned($unsigned((8'ha1)))));
                  for (forvar7355 = (1'h0); (forvar7355 < (1'h0)); forvar7355 = (forvar7355 + (1'h1)))
                    begin
                      reg7356 <= $signed($signed((8'h9e)));
                      reg7357 <= ((&((|reg709) ?
                          forvar718[(1'h1):(1'h0)] : (reg4289 ?
                              reg695 : reg4212))) * forvar4244);
                    end
                end
            end
        end
      reg7361 <= reg4179;
    end
  assign wire7362 = $signed((^~($signed(forvar4321) >> {reg4255})));
  assign wire7363 = {reg737[(3'h7):(1'h0)]};
  always
    @(posedge clk) begin
      reg7364 <= ((reg695[(3'h4):(1'h1)] >> $signed($signed(reg834))) ?
          reg7351 : forvar7333[(3'h7):(2'h3)]);
      for (forvar7365 = (1'h0); (forvar7365 < (2'h3)); forvar7365 = (forvar7365 + (1'h1)))
        begin
          for (forvar7366 = (1'h0); (forvar7366 < (2'h2)); forvar7366 = (forvar7366 + (1'h1)))
            begin
              if ((|($signed(forvar848) ?
                  ((8'hb6) - (!reg716)) : $signed(reg4302[(2'h2):(1'h0)]))))
                begin
                  for (forvar7367 = (1'h0); (forvar7367 < (1'h1)); forvar7367 = (forvar7367 + (1'h1)))
                    begin
                      reg7368 <= {(~$signed((+(8'hb5))))};
                      reg7369 <= $unsigned((-({reg4291} || (reg721 >= reg851))));
                      reg7370 <= {{$signed(reg4290[(2'h2):(1'h1)])}};
                    end
                  for (forvar7371 = (1'h0); (forvar7371 < (1'h1)); forvar7371 = (forvar7371 + (1'h1)))
                    begin
                      reg7372 <= reg4175[(3'h5):(3'h5)];
                      reg7373 <= $signed((~&reg4183[(1'h1):(1'h1)]));
                      reg7374 <= (forvar799 ?
                          (^~$unsigned($signed(reg850))) : $signed($unsigned(reg696)));
                      reg7375 <= $signed({$signed(((8'ha2) ?
                              (8'h9d) : reg729))});
                    end
                  reg7376 <= $unsigned((($signed((8'ha8)) || forvar4216) ?
                      (!(^~reg858)) : $signed(forvar4279[(3'h5):(3'h5)])));
                  reg7377 <= {reg853[(4'ha):(3'h5)]};
                end
              else
                begin
                  reg7367 <= (-reg4245);
                  for (forvar7368 = (1'h0); (forvar7368 < (2'h3)); forvar7368 = (forvar7368 + (1'h1)))
                    begin
                      reg7369 <= $signed(((^~reg4313[(3'h6):(2'h2)]) ?
                          {$unsigned(forvar4181)} : (|(reg7374 ?
                              reg4248 : reg4327))));
                      reg7370 <= (((8'haf) ^~ (-(^~reg4299))) ~^ reg696);
                    end
                end
              for (forvar7378 = (1'h0); (forvar7378 < (2'h3)); forvar7378 = (forvar7378 + (1'h1)))
                begin
                  if (((^~(+(reg711 * (8'ha0)))) ?
                      (((+wire4336) - reg4259) > reg799[(3'h5):(2'h3)]) : (~$signed(((8'hb3) ?
                          reg726 : reg4326)))))
                    begin
                      reg7379 <= $unsigned(forvar790);
                      reg7380 <= ($signed(forvar735) & {((reg723 ?
                              reg4327 : reg4198) != (forvar870 >= forvar4226))});
                      reg7381 <= ($signed((&(+reg7374))) ?
                          reg4260 : $unsigned(($unsigned(forvar879) + $signed(reg712))));
                      reg7382 <= $signed(((~(reg4265 ? forvar4192 : reg4220)) ?
                          (~|(!reg4172)) : reg4229[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg7379 <= reg7350;
                      reg7380 <= $signed($unsigned(($signed(reg841) << forvar852[(4'hd):(1'h0)])));
                      reg7381 <= reg4273[(4'h8):(1'h0)];
                    end
                  for (forvar7383 = (1'h0); (forvar7383 < (1'h0)); forvar7383 = (forvar7383 + (1'h1)))
                    begin
                      reg7384 <= (~&($unsigned((+reg767)) >> $signed($signed(reg4290))));
                      reg7385 <= reg4326[(2'h3):(2'h2)];
                    end
                  for (forvar7386 = (1'h0); (forvar7386 < (1'h1)); forvar7386 = (forvar7386 + (1'h1)))
                    begin
                      reg7387 <= (~|(({reg810} * (+(8'ha2))) ?
                          reg775[(4'he):(4'h8)] : (reg4196[(2'h2):(1'h1)] ?
                              (reg7381 > (8'hb5)) : forvar4308[(4'h8):(3'h4)])));
                      reg7388 <= $unsigned($signed({$unsigned(reg693)}));
                      reg7389 <= reg7349[(2'h2):(2'h2)];
                    end
                  reg7390 <= (+$signed($unsigned((~^(8'hb5)))));
                end
              for (forvar7391 = (1'h0); (forvar7391 < (2'h3)); forvar7391 = (forvar7391 + (1'h1)))
                begin
                  if (((~|(8'had)) < reg830))
                    begin
                      reg7392 <= {reg759};
                    end
                  else
                    begin
                      reg7392 <= (&forvar4216);
                      reg7393 <= {((~|(|reg885)) ^ ((forvar780 + reg4173) && $signed(reg4231)))};
                      reg7394 <= (reg4305 >> reg4262[(1'h1):(1'h0)]);
                      reg7395 <= ((^~(~|((8'h9d) ?
                          reg7392 : reg4307))) ^ $signed($signed((reg843 ?
                          forvar4324 : forvar681))));
                    end
                  if (($signed(forvar4204[(1'h0):(1'h0)]) ?
                      (reg7364[(4'h8):(1'h0)] * $unsigned({reg4184})) : reg833))
                    begin
                      reg7396 <= $unsigned($signed(($unsigned(reg4231) * (reg7376 ?
                          reg4306 : forvar4268))));
                      reg7397 <= $signed($signed(forvar711));
                    end
                  else
                    begin
                      reg7396 <= ($signed(((reg4233 == reg857) ?
                          (!reg691) : forvar726[(1'h0):(1'h0)])) & reg784[(4'h8):(1'h0)]);
                      reg7397 <= $unsigned((((^~reg820) & $signed(forvar4268)) ?
                          reg4178[(1'h1):(1'h1)] : forvar4181[(4'h9):(4'h8)]));
                    end
                end
              if ((~{{reg4247[(2'h2):(1'h1)]}}))
                begin
                  for (forvar7398 = (1'h0); (forvar7398 < (1'h0)); forvar7398 = (forvar7398 + (1'h1)))
                    begin
                      reg7399 <= reg7356;
                      reg7400 <= (reg4177[(4'ha):(2'h3)] ?
                          $signed((reg4193[(1'h1):(1'h1)] ?
                              $signed(forvar4307) : forvar719[(3'h4):(1'h1)])) : ((((8'hb7) ?
                                  forvar875 : (8'h9e)) <= (reg4262 ?
                                  reg849 : wire677)) ?
                              forvar707 : (&reg4328)));
                      reg7401 <= (8'ha7);
                      reg7402 <= forvar4195;
                    end
                end
              else
                begin
                  reg7398 <= (-({(forvar4214 >>> reg726)} ~^ reg865));
                end
            end
          for (forvar7403 = (1'h0); (forvar7403 < (1'h0)); forvar7403 = (forvar7403 + (1'h1)))
            begin
              for (forvar7404 = (1'h0); (forvar7404 < (2'h2)); forvar7404 = (forvar7404 + (1'h1)))
                begin
                  for (forvar7405 = (1'h0); (forvar7405 < (1'h0)); forvar7405 = (forvar7405 + (1'h1)))
                    begin
                      reg7406 <= ({$unsigned($unsigned(forvar4293))} | (|((8'hb0) <= forvar4172[(3'h6):(2'h2)])));
                      reg7407 <= (~^$unsigned(reg694));
                    end
                  for (forvar7408 = (1'h0); (forvar7408 < (1'h1)); forvar7408 = (forvar7408 + (1'h1)))
                    begin
                      reg7409 <= $signed((-reg768));
                      reg7410 <= (^reg823[(4'ha):(3'h4)]);
                      reg7411 <= reg4230;
                      reg7412 <= (^$unsigned(forvar4226));
                    end
                  reg7413 <= $signed($signed(forvar718));
                end
              if (($unsigned(reg7357) ?
                  reg869 : (((8'hba) <= reg718) ?
                      reg871[(1'h0):(1'h0)] : ((reg683 ?
                          reg785 : (8'hba)) & forvar879))))
                begin
                  if ((~|{reg7352}))
                    begin
                      reg7414 <= ((((-(8'ha8)) ?
                          reg4190[(2'h2):(1'h0)] : (-reg819)) <<< $unsigned(forvar789)) != (forvar7371[(3'h5):(2'h2)] ?
                          $signed((reg684 == forvar4320)) : (&forvar866)));
                      reg7415 <= $signed(reg805);
                    end
                  else
                    begin
                      reg7414 <= ($unsigned($signed($signed(reg738))) ?
                          (~&{$unsigned(reg772)}) : forvar779[(2'h2):(1'h1)]);
                    end
                  for (forvar7416 = (1'h0); (forvar7416 < (1'h1)); forvar7416 = (forvar7416 + (1'h1)))
                    begin
                      reg7417 <= $unsigned(((~^$signed((8'hb7))) ?
                          reg4237 : (reg4326 ?
                              (reg701 ? reg4253 : reg702) : (forvar4316 ?
                                  reg4243 : reg777))));
                      reg7418 <= (~^reg785);
                      reg7419 <= ((reg4317 ?
                          (&$signed(reg840)) : (8'ha5)) <<< forvar4205);
                    end
                  for (forvar7420 = (1'h0); (forvar7420 < (1'h1)); forvar7420 = (forvar7420 + (1'h1)))
                    begin
                      reg7421 <= $unsigned({{forvar4330[(3'h4):(2'h2)]}});
                      reg7422 <= reg7415;
                      reg7423 <= (~forvar7341);
                    end
                end
              else
                begin
                  if (reg4280)
                    begin
                      reg7414 <= (8'h9d);
                      reg7415 <= (!$unsigned($signed((reg776 ?
                          forvar832 : reg4291))));
                      reg7416 <= $unsigned($unsigned((^~((8'had) ~^ (8'hab)))));
                    end
                  else
                    begin
                      reg7414 <= (reg4313[(1'h1):(1'h0)] ?
                          reg4265[(4'h8):(2'h2)] : (($unsigned((8'ha2)) ?
                              $signed(forvar4192) : forvar682) | $signed($signed(reg7384))));
                    end
                  if (reg748[(2'h2):(2'h2)])
                    begin
                      reg7417 <= (|$unsigned(reg713[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg7417 <= $unsigned(((~|(reg774 ?
                          reg691 : reg4321)) > $signed((^~reg844))));
                      reg7418 <= forvar4252;
                      reg7419 <= forvar7391[(1'h1):(1'h1)];
                      reg7420 <= $signed(reg7396[(2'h2):(1'h1)]);
                    end
                end
            end
        end
    end
  assign wire7424 = $unsigned(reg4321[(1'h1):(1'h1)]);
  assign wire7425 = $unsigned($unsigned(forvar7368));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4337
#(parameter param7330 = (~^(+((~&(8'h9f)) >= (&(8'hac))))))
(y, clk, wire4341, wire4340, wire4339, wire4338);
  output wire [(32'h1795):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire4341;
  input wire [(4'ha):(1'h0)] wire4340;
  input wire [(3'h5):(1'h0)] wire4339;
  input wire [(3'h7):(1'h0)] wire4338;
  reg signed [(3'h4):(1'h0)] reg7329 = (1'h0);
  reg [(4'h9):(1'h0)] reg7328 = (1'h0);
  reg [(4'h8):(1'h0)] reg7327 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7326 = (1'h0);
  reg [(4'hf):(1'h0)] reg7325 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7324 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7323 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7322 = (1'h0);
  reg [(4'hc):(1'h0)] reg7321 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7320 = (1'h0);
  reg [(2'h3):(1'h0)] reg7319 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7318 = (1'h0);
  reg [(4'hf):(1'h0)] reg7317 = (1'h0);
  reg [(5'h10):(1'h0)] reg7316 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7315 = (1'h0);
  reg [(3'h7):(1'h0)] reg7314 = (1'h0);
  reg [(4'hc):(1'h0)] reg7313 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7312 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7311 = (1'h0);
  reg [(3'h6):(1'h0)] reg7310 = (1'h0);
  reg [(4'hd):(1'h0)] reg7309 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7308 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7307 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7306 = (1'h0);
  reg [(3'h6):(1'h0)] reg7302 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7300 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7299 = (1'h0);
  reg [(4'h8):(1'h0)] reg7305 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7304 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7303 = (1'h0);
  reg [(3'h6):(1'h0)] forvar7302 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7301 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7300 = (1'h0);
  reg [(3'h7):(1'h0)] reg7299 = (1'h0);
  reg [(2'h2):(1'h0)] reg7298 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7297 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7296 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7295 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7293 = (1'h0);
  reg [(4'h9):(1'h0)] reg7287 = (1'h0);
  reg [(4'he):(1'h0)] reg7294 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7293 = (1'h0);
  reg [(4'hb):(1'h0)] reg7292 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7291 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7290 = (1'h0);
  reg [(4'hd):(1'h0)] reg7289 = (1'h0);
  reg [(5'h10):(1'h0)] reg7288 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar7287 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7286 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7285 = (1'h0);
  reg [(3'h6):(1'h0)] reg7284 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7283 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7282 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7281 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7280 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7279 = (1'h0);
  reg [(4'ha):(1'h0)] reg7278 = (1'h0);
  reg [(3'h4):(1'h0)] reg7277 = (1'h0);
  reg [(3'h5):(1'h0)] reg7276 = (1'h0);
  reg [(2'h3):(1'h0)] reg7275 = (1'h0);
  reg [(4'he):(1'h0)] reg7274 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7273 = (1'h0);
  reg [(4'he):(1'h0)] reg7272 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7271 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7270 = (1'h0);
  reg [(4'hb):(1'h0)] reg7269 = (1'h0);
  reg [(4'hf):(1'h0)] reg7268 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7267 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7266 = (1'h0);
  reg [(4'ha):(1'h0)] reg7265 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7264 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7263 = (1'h0);
  reg [(3'h4):(1'h0)] reg7262 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7261 = (1'h0);
  reg [(3'h7):(1'h0)] forvar7260 = (1'h0);
  reg [(4'h8):(1'h0)] reg7259 = (1'h0);
  reg [(2'h3):(1'h0)] reg7258 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7257 = (1'h0);
  reg [(3'h4):(1'h0)] reg7254 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7253 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7257 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7256 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7255 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7254 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7253 = (1'h0);
  reg [(4'ha):(1'h0)] reg7249 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7245 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7242 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7252 = (1'h0);
  reg [(2'h3):(1'h0)] reg7251 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7250 = (1'h0);
  reg [(4'hd):(1'h0)] forvar7249 = (1'h0);
  reg [(4'h8):(1'h0)] reg7248 = (1'h0);
  reg [(2'h3):(1'h0)] reg7247 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7246 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7245 = (1'h0);
  reg [(4'h8):(1'h0)] reg7244 = (1'h0);
  reg [(4'ha):(1'h0)] reg7243 = (1'h0);
  reg [(4'hc):(1'h0)] reg7242 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar7241 = (1'h0);
  reg [(4'h8):(1'h0)] reg7240 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7239 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7238 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7237 = (1'h0);
  reg [(5'h10):(1'h0)] reg7236 = (1'h0);
  reg [(4'hb):(1'h0)] reg7235 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7234 = (1'h0);
  reg [(4'hd):(1'h0)] reg7233 = (1'h0);
  reg [(4'hb):(1'h0)] reg7232 = (1'h0);
  reg [(4'hb):(1'h0)] reg7231 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7230 = (1'h0);
  reg [(5'h10):(1'h0)] reg7229 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7228 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7227 = (1'h0);
  reg [(3'h6):(1'h0)] reg7226 = (1'h0);
  reg [(4'he):(1'h0)] reg7225 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7224 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7223 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7222 = (1'h0);
  reg [(4'hd):(1'h0)] reg7221 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7220 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7219 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7218 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7217 = (1'h0);
  reg [(4'he):(1'h0)] reg7216 = (1'h0);
  reg [(4'ha):(1'h0)] reg7215 = (1'h0);
  reg [(3'h5):(1'h0)] forvar7214 = (1'h0);
  reg [(2'h2):(1'h0)] forvar7213 = (1'h0);
  reg [(3'h7):(1'h0)] reg7212 = (1'h0);
  reg [(3'h5):(1'h0)] reg7211 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7210 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7209 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7208 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7207 = (1'h0);
  reg [(4'hb):(1'h0)] reg7206 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7205 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7201 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7205 = (1'h0);
  reg [(3'h5):(1'h0)] reg7204 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7203 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7202 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7201 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7200 = (1'h0);
  reg [(4'hb):(1'h0)] reg7199 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7196 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7193 = (1'h0);
  reg [(3'h4):(1'h0)] reg7198 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7197 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7196 = (1'h0);
  reg [(4'h8):(1'h0)] reg7195 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7194 = (1'h0);
  reg [(4'he):(1'h0)] reg7193 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7192 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7191 = (1'h0);
  reg [(4'hb):(1'h0)] reg7170 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7190 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7189 = (1'h0);
  reg [(5'h10):(1'h0)] reg7188 = (1'h0);
  reg [(4'ha):(1'h0)] reg7187 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7186 = (1'h0);
  reg [(4'hc):(1'h0)] reg7185 = (1'h0);
  reg [(4'he):(1'h0)] reg7184 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7183 = (1'h0);
  reg [(4'h8):(1'h0)] reg7182 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7181 = (1'h0);
  reg [(4'he):(1'h0)] reg7180 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7179 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7178 = (1'h0);
  reg [(3'h6):(1'h0)] reg7177 = (1'h0);
  reg [(4'h8):(1'h0)] reg7176 = (1'h0);
  reg [(5'h10):(1'h0)] reg7175 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7174 = (1'h0);
  reg [(4'hf):(1'h0)] reg7173 = (1'h0);
  reg [(3'h7):(1'h0)] reg7172 = (1'h0);
  reg [(2'h2):(1'h0)] reg7171 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar7170 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7169 = (1'h0);
  reg [(4'h8):(1'h0)] reg7168 = (1'h0);
  reg [(4'he):(1'h0)] reg7167 = (1'h0);
  reg [(4'he):(1'h0)] reg7166 = (1'h0);
  reg [(4'hc):(1'h0)] reg7165 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7164 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7163 = (1'h0);
  reg [(4'ha):(1'h0)] reg7162 = (1'h0);
  reg [(4'he):(1'h0)] reg7161 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7160 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7159 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7158 = (1'h0);
  reg [(4'hd):(1'h0)] reg7157 = (1'h0);
  reg [(4'he):(1'h0)] forvar7154 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7153 = (1'h0);
  reg [(4'hf):(1'h0)] reg7152 = (1'h0);
  reg [(5'h10):(1'h0)] forvar7150 = (1'h0);
  reg [(2'h3):(1'h0)] reg7149 = (1'h0);
  reg [(3'h4):(1'h0)] reg7156 = (1'h0);
  reg [(4'hf):(1'h0)] reg7155 = (1'h0);
  reg [(3'h7):(1'h0)] reg7154 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7153 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7152 = (1'h0);
  reg [(4'he):(1'h0)] reg7151 = (1'h0);
  reg [(3'h6):(1'h0)] reg7150 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7149 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7148 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7147 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7142 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7141 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar7134 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7132 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar7129 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar7125 = (1'h0);
  reg [(4'h9):(1'h0)] forvar7116 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7118 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7115 = (1'h0);
  reg [(3'h6):(1'h0)] forvar7114 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar7103 = (1'h0);
  reg [(2'h2):(1'h0)] forvar7099 = (1'h0);
  reg [(4'hb):(1'h0)] forvar7098 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7093 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7094 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7090 = (1'h0);
  reg [(4'hd):(1'h0)] reg7089 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7086 = (1'h0);
  reg [(3'h7):(1'h0)] reg7146 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar7139 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7145 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7143 = (1'h0);
  reg [(3'h6):(1'h0)] reg7140 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar7138 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar7136 = (1'h0);
  reg [(3'h4):(1'h0)] reg7135 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar7131 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7130 = (1'h0);
  reg [(4'hb):(1'h0)] reg7126 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar7123 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7120 = (1'h0);
  reg [(4'h9):(1'h0)] forvar7112 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7111 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar7106 = (1'h0);
  reg [(4'he):(1'h0)] reg7144 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7143 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7142 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7141 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7140 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7139 = (1'h0);
  reg [(2'h3):(1'h0)] reg7138 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7137 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7136 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7135 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7134 = (1'h0);
  reg [(3'h6):(1'h0)] reg7133 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7132 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg7131 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar7130 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7129 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7128 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7127 = (1'h0);
  reg [(3'h4):(1'h0)] forvar7126 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7125 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7124 = (1'h0);
  reg [(4'h9):(1'h0)] reg7123 = (1'h0);
  reg [(4'hf):(1'h0)] reg7122 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7121 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7120 = (1'h0);
  reg [(2'h2):(1'h0)] reg7119 = (1'h0);
  reg [(4'hd):(1'h0)] reg7118 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7117 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7116 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7115 = (1'h0);
  reg [(3'h5):(1'h0)] reg7114 = (1'h0);
  reg [(4'hb):(1'h0)] reg7113 = (1'h0);
  reg [(4'he):(1'h0)] reg7112 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7111 = (1'h0);
  reg [(4'h9):(1'h0)] reg7110 = (1'h0);
  reg [(4'hb):(1'h0)] reg7109 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7108 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7107 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7106 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg7105 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7104 = (1'h0);
  reg [(3'h5):(1'h0)] reg7088 = (1'h0);
  reg [(3'h6):(1'h0)] forvar7087 = (1'h0);
  reg [(4'ha):(1'h0)] reg7103 = (1'h0);
  reg [(4'he):(1'h0)] reg7102 = (1'h0);
  reg [(4'ha):(1'h0)] reg7101 = (1'h0);
  reg [(2'h2):(1'h0)] reg7100 = (1'h0);
  reg [(4'hf):(1'h0)] reg7099 = (1'h0);
  reg [(3'h7):(1'h0)] reg7098 = (1'h0);
  reg [(4'h8):(1'h0)] reg7097 = (1'h0);
  reg [(4'h9):(1'h0)] reg7096 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7095 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar7094 = (1'h0);
  reg [(5'h10):(1'h0)] reg7093 = (1'h0);
  reg [(3'h7):(1'h0)] reg7092 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7091 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7090 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7089 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7088 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7087 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7086 = (1'h0);
  reg [(4'hd):(1'h0)] reg7085 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7084 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7083 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7082 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7081 = (1'h0);
  reg [(2'h3):(1'h0)] reg7080 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7079 = (1'h0);
  reg [(4'hc):(1'h0)] reg7078 = (1'h0);
  reg [(5'h10):(1'h0)] reg7077 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7076 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7075 = (1'h0);
  reg [(4'h9):(1'h0)] reg7074 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7071 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7073 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7072 = (1'h0);
  reg [(4'he):(1'h0)] reg7071 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7070 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7069 = (1'h0);
  reg [(4'h9):(1'h0)] forvar7068 = (1'h0);
  reg [(4'hf):(1'h0)] reg7067 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7066 = (1'h0);
  reg [(2'h2):(1'h0)] reg7065 = (1'h0);
  reg [(3'h4):(1'h0)] reg7064 = (1'h0);
  reg [(2'h3):(1'h0)] forvar7063 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg7062 = (1'h0);
  reg [(3'h7):(1'h0)] reg7061 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7060 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7059 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg7058 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7057 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7056 = (1'h0);
  reg [(4'he):(1'h0)] reg7055 = (1'h0);
  reg [(2'h2):(1'h0)] forvar7054 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7053 = (1'h0);
  reg [(4'hd):(1'h0)] reg7052 = (1'h0);
  reg [(4'ha):(1'h0)] reg7051 = (1'h0);
  reg [(3'h5):(1'h0)] reg7050 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7049 = (1'h0);
  reg [(4'hf):(1'h0)] forvar7048 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar7047 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7044 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar7040 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7046 = (1'h0);
  reg [(4'hd):(1'h0)] reg7045 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg7044 = (1'h0);
  reg [(4'h8):(1'h0)] reg7043 = (1'h0);
  reg [(4'hc):(1'h0)] reg7042 = (1'h0);
  reg [(5'h10):(1'h0)] reg7041 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg7040 = (1'h0);
  reg [(2'h2):(1'h0)] reg7039 = (1'h0);
  reg [(4'h9):(1'h0)] reg7038 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar7037 = (1'h0);
  reg [(3'h5):(1'h0)] forvar7033 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7030 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg7036 = (1'h0);
  reg [(4'he):(1'h0)] reg7035 = (1'h0);
  reg [(5'h10):(1'h0)] reg7034 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7033 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7032 = (1'h0);
  reg [(2'h3):(1'h0)] reg7031 = (1'h0);
  reg [(5'h10):(1'h0)] forvar7030 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg7029 = (1'h0);
  reg [(2'h3):(1'h0)] reg7028 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg7027 = (1'h0);
  reg [(2'h2):(1'h0)] reg7026 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg7025 = (1'h0);
  reg [(2'h2):(1'h0)] reg7024 = (1'h0);
  reg [(4'h9):(1'h0)] forvar7023 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg7022 = (1'h0);
  reg [(4'hb):(1'h0)] reg7021 = (1'h0);
  reg [(4'hd):(1'h0)] reg7020 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg7019 = (1'h0);
  reg [(4'he):(1'h0)] reg7018 = (1'h0);
  reg signed [(4'he):(1'h0)] reg7017 = (1'h0);
  reg [(4'hb):(1'h0)] reg7016 = (1'h0);
  reg [(4'h8):(1'h0)] reg7015 = (1'h0);
  reg [(2'h2):(1'h0)] reg7014 = (1'h0);
  reg [(2'h2):(1'h0)] reg7013 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar7012 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7011 = (1'h0);
  reg [(4'h8):(1'h0)] forvar7010 = (1'h0);
  wire [(2'h3):(1'h0)] wire7009;
  wire signed [(3'h4):(1'h0)] wire7008;
  wire signed [(4'h8):(1'h0)] wire7006;
  wire [(4'hc):(1'h0)] wire4571;
  reg [(3'h5):(1'h0)] reg4570 = (1'h0);
  reg [(4'hb):(1'h0)] reg4569 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4568 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4567 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4566 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4565 = (1'h0);
  reg [(4'hc):(1'h0)] reg4564 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4563 = (1'h0);
  reg [(4'ha):(1'h0)] reg4562 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4561 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4560 = (1'h0);
  reg [(4'h8):(1'h0)] reg4559 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4558 = (1'h0);
  reg [(4'hb):(1'h0)] reg4557 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4556 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4555 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4554 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4553 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4552 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4551 = (1'h0);
  reg [(4'hd):(1'h0)] reg4550 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4549 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4548 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4547 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4546 = (1'h0);
  reg [(4'h9):(1'h0)] reg4545 = (1'h0);
  reg [(4'h9):(1'h0)] reg4544 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4543 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4542 = (1'h0);
  reg [(5'h10):(1'h0)] reg4538 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4537 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4542 = (1'h0);
  reg [(4'hc):(1'h0)] reg4541 = (1'h0);
  reg [(4'h8):(1'h0)] reg4540 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4539 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4538 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4537 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4536 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4535 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4522 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4520 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4534 = (1'h0);
  reg [(3'h4):(1'h0)] reg4533 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4532 = (1'h0);
  reg [(3'h5):(1'h0)] reg4531 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4530 = (1'h0);
  reg [(3'h4):(1'h0)] reg4529 = (1'h0);
  reg [(4'hf):(1'h0)] reg4528 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4527 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4526 = (1'h0);
  reg [(3'h7):(1'h0)] reg4525 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4524 = (1'h0);
  reg [(4'hf):(1'h0)] reg4523 = (1'h0);
  reg [(5'h10):(1'h0)] reg4522 = (1'h0);
  reg [(4'hb):(1'h0)] reg4521 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4520 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4519 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4518 = (1'h0);
  reg [(4'hd):(1'h0)] reg4517 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4510 = (1'h0);
  reg [(4'he):(1'h0)] forvar4509 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4506 = (1'h0);
  reg [(4'hc):(1'h0)] reg4516 = (1'h0);
  reg [(3'h7):(1'h0)] reg4515 = (1'h0);
  reg [(3'h6):(1'h0)] reg4514 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4513 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4512 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4511 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4510 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4509 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4508 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4503 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4496 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4490 = (1'h0);
  reg [(2'h2):(1'h0)] reg4489 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4487 = (1'h0);
  reg [(4'ha):(1'h0)] reg4486 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4485 = (1'h0);
  reg [(4'hf):(1'h0)] reg4482 = (1'h0);
  reg [(3'h7):(1'h0)] reg4507 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4504 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4501 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4500 = (1'h0);
  reg [(4'hd):(1'h0)] reg4506 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4505 = (1'h0);
  reg [(4'hc):(1'h0)] reg4504 = (1'h0);
  reg [(5'h10):(1'h0)] reg4503 = (1'h0);
  reg [(2'h2):(1'h0)] reg4502 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4501 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4500 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4499 = (1'h0);
  reg [(2'h2):(1'h0)] reg4498 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4497 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4496 = (1'h0);
  reg [(4'hf):(1'h0)] reg4495 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4494 = (1'h0);
  reg [(4'h9):(1'h0)] reg4493 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4492 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4491 = (1'h0);
  reg [(4'ha):(1'h0)] reg4490 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4489 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4488 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4487 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4486 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4485 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4484 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4483 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4481 = (1'h0);
  reg [(5'h10):(1'h0)] reg4480 = (1'h0);
  reg [(4'hf):(1'h0)] reg4479 = (1'h0);
  reg [(4'hb):(1'h0)] reg4478 = (1'h0);
  reg [(5'h10):(1'h0)] reg4477 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4476 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4475 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4474 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4473 = (1'h0);
  reg [(4'h8):(1'h0)] reg4472 = (1'h0);
  reg [(2'h2):(1'h0)] reg4471 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4470 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4469 = (1'h0);
  reg [(4'ha):(1'h0)] reg4468 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4467 = (1'h0);
  reg [(4'hb):(1'h0)] reg4466 = (1'h0);
  reg [(3'h4):(1'h0)] reg4465 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4464 = (1'h0);
  reg [(4'h8):(1'h0)] reg4463 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4462 = (1'h0);
  reg [(2'h2):(1'h0)] reg4461 = (1'h0);
  reg [(3'h6):(1'h0)] reg4459 = (1'h0);
  reg [(4'hb):(1'h0)] reg4457 = (1'h0);
  reg [(4'hb):(1'h0)] reg4460 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4459 = (1'h0);
  reg [(3'h4):(1'h0)] reg4458 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4457 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4456 = (1'h0);
  reg [(2'h2):(1'h0)] reg4455 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4454 = (1'h0);
  reg [(2'h3):(1'h0)] reg4453 = (1'h0);
  reg [(4'hf):(1'h0)] reg4452 = (1'h0);
  reg [(4'hb):(1'h0)] reg4451 = (1'h0);
  reg [(4'h9):(1'h0)] reg4450 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4449 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4448 = (1'h0);
  reg [(4'h8):(1'h0)] reg4447 = (1'h0);
  reg [(4'hd):(1'h0)] reg4446 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4445 = (1'h0);
  reg [(4'hd):(1'h0)] reg4444 = (1'h0);
  reg [(4'hf):(1'h0)] reg4443 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4442 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4441 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4440 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4439 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4438 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4437 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4436 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4435 = (1'h0);
  reg [(4'hc):(1'h0)] reg4434 = (1'h0);
  reg [(4'h9):(1'h0)] reg4433 = (1'h0);
  reg [(4'h9):(1'h0)] reg4432 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4427 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4424 = (1'h0);
  reg [(2'h3):(1'h0)] reg4423 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4422 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4414 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4412 = (1'h0);
  reg [(4'hb):(1'h0)] reg4431 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4430 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4429 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4428 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4427 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4426 = (1'h0);
  reg [(3'h6):(1'h0)] reg4425 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4424 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4423 = (1'h0);
  reg [(4'he):(1'h0)] reg4422 = (1'h0);
  reg [(4'hb):(1'h0)] reg4418 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4413 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4421 = (1'h0);
  reg [(4'h9):(1'h0)] reg4420 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4419 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4418 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4417 = (1'h0);
  reg [(4'ha):(1'h0)] reg4416 = (1'h0);
  reg [(3'h7):(1'h0)] reg4415 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4414 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4413 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4411 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4410 = (1'h0);
  reg [(3'h6):(1'h0)] reg4409 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4408 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4407 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4406 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4405 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4404 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4403 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4402 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4401 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4400 = (1'h0);
  reg [(4'ha):(1'h0)] reg4391 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4386 = (1'h0);
  reg [(4'ha):(1'h0)] reg4399 = (1'h0);
  reg [(3'h6):(1'h0)] reg4398 = (1'h0);
  reg [(3'h4):(1'h0)] reg4397 = (1'h0);
  reg [(5'h10):(1'h0)] reg4396 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4395 = (1'h0);
  reg [(4'h8):(1'h0)] reg4394 = (1'h0);
  reg [(4'ha):(1'h0)] reg4393 = (1'h0);
  reg [(3'h7):(1'h0)] reg4392 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4391 = (1'h0);
  reg [(5'h10):(1'h0)] reg4390 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4389 = (1'h0);
  reg [(4'he):(1'h0)] reg4388 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4387 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4386 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4385 = (1'h0);
  reg [(3'h4):(1'h0)] reg4384 = (1'h0);
  reg [(3'h5):(1'h0)] reg4383 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4382 = (1'h0);
  reg [(4'ha):(1'h0)] reg4381 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4380 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4379 = (1'h0);
  reg [(4'hf):(1'h0)] reg4378 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4377 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4375 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4372 = (1'h0);
  reg [(2'h2):(1'h0)] reg4369 = (1'h0);
  reg [(4'he):(1'h0)] reg4376 = (1'h0);
  reg [(5'h10):(1'h0)] reg4375 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4374 = (1'h0);
  reg [(4'h9):(1'h0)] reg4373 = (1'h0);
  reg [(4'hb):(1'h0)] reg4372 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4371 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4370 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4369 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4368 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4367 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4366 = (1'h0);
  reg [(4'hd):(1'h0)] reg4365 = (1'h0);
  reg [(4'he):(1'h0)] forvar4364 = (1'h0);
  reg [(4'h8):(1'h0)] reg4359 = (1'h0);
  reg [(4'h8):(1'h0)] reg4363 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4362 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4361 = (1'h0);
  reg [(4'ha):(1'h0)] reg4360 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4359 = (1'h0);
  reg [(4'hf):(1'h0)] reg4356 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4353 = (1'h0);
  reg [(4'he):(1'h0)] reg4352 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4350 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4347 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4345 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4358 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4357 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4356 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4355 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4354 = (1'h0);
  reg [(4'ha):(1'h0)] reg4353 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4352 = (1'h0);
  reg [(2'h3):(1'h0)] reg4351 = (1'h0);
  reg [(2'h2):(1'h0)] reg4350 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4349 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4348 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4347 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4346 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4345 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4344 = (1'h0);
  wire [(4'hb):(1'h0)] wire4343;
  wire signed [(4'hf):(1'h0)] wire4342;
  assign y = {reg7329,
                 reg7328,
                 reg7327,
                 reg7326,
                 reg7325,
                 reg7324,
                 reg7323,
                 reg7322,
                 reg7321,
                 forvar7320,
                 reg7319,
                 reg7318,
                 reg7317,
                 reg7316,
                 forvar7315,
                 reg7314,
                 reg7313,
                 reg7312,
                 forvar7311,
                 reg7310,
                 reg7309,
                 reg7308,
                 forvar7307,
                 forvar7306,
                 reg7302,
                 reg7300,
                 forvar7299,
                 reg7305,
                 reg7304,
                 reg7303,
                 forvar7302,
                 reg7301,
                 forvar7300,
                 reg7299,
                 reg7298,
                 forvar7297,
                 reg7296,
                 forvar7295,
                 forvar7293,
                 reg7287,
                 reg7294,
                 reg7293,
                 reg7292,
                 reg7291,
                 forvar7290,
                 reg7289,
                 reg7288,
                 forvar7287,
                 reg7286,
                 forvar7285,
                 reg7284,
                 reg7283,
                 reg7282,
                 forvar7281,
                 forvar7280,
                 forvar7279,
                 reg7278,
                 reg7277,
                 reg7276,
                 reg7275,
                 reg7274,
                 forvar7273,
                 reg7272,
                 reg7271,
                 reg7270,
                 reg7269,
                 reg7268,
                 reg7267,
                 reg7266,
                 reg7265,
                 reg7264,
                 reg7263,
                 reg7262,
                 forvar7261,
                 forvar7260,
                 reg7259,
                 reg7258,
                 forvar7257,
                 reg7254,
                 reg7253,
                 reg7257,
                 reg7256,
                 reg7255,
                 forvar7254,
                 forvar7253,
                 reg7249,
                 reg7245,
                 forvar7242,
                 reg7252,
                 reg7251,
                 reg7250,
                 forvar7249,
                 reg7248,
                 reg7247,
                 reg7246,
                 forvar7245,
                 reg7244,
                 reg7243,
                 reg7242,
                 forvar7241,
                 reg7240,
                 reg7239,
                 forvar7238,
                 forvar7237,
                 reg7236,
                 reg7235,
                 reg7234,
                 reg7233,
                 reg7232,
                 reg7231,
                 reg7230,
                 reg7229,
                 forvar7228,
                 forvar7227,
                 reg7226,
                 reg7225,
                 reg7224,
                 reg7223,
                 reg7222,
                 reg7221,
                 reg7220,
                 forvar7219,
                 reg7218,
                 reg7217,
                 reg7216,
                 reg7215,
                 forvar7214,
                 forvar7213,
                 reg7212,
                 reg7211,
                 reg7210,
                 reg7209,
                 reg7208,
                 forvar7207,
                 reg7206,
                 forvar7205,
                 forvar7201,
                 reg7205,
                 reg7204,
                 reg7203,
                 reg7202,
                 reg7201,
                 reg7200,
                 reg7199,
                 reg7196,
                 forvar7193,
                 reg7198,
                 reg7197,
                 forvar7196,
                 reg7195,
                 reg7194,
                 reg7193,
                 reg7192,
                 forvar7191,
                 reg7170,
                 reg7190,
                 reg7189,
                 reg7188,
                 reg7187,
                 reg7186,
                 reg7185,
                 reg7184,
                 forvar7183,
                 reg7182,
                 forvar7181,
                 reg7180,
                 reg7179,
                 reg7178,
                 reg7177,
                 reg7176,
                 reg7175,
                 reg7174,
                 reg7173,
                 reg7172,
                 reg7171,
                 forvar7170,
                 forvar7169,
                 reg7168,
                 reg7167,
                 reg7166,
                 reg7165,
                 reg7164,
                 reg7163,
                 reg7162,
                 reg7161,
                 forvar7160,
                 forvar7159,
                 reg7158,
                 reg7157,
                 forvar7154,
                 forvar7153,
                 reg7152,
                 forvar7150,
                 reg7149,
                 reg7156,
                 reg7155,
                 reg7154,
                 reg7153,
                 forvar7152,
                 reg7151,
                 reg7150,
                 forvar7149,
                 forvar7148,
                 reg7147,
                 forvar7142,
                 forvar7141,
                 forvar7134,
                 forvar7132,
                 forvar7129,
                 forvar7125,
                 forvar7116,
                 forvar7118,
                 forvar7115,
                 forvar7114,
                 forvar7103,
                 forvar7099,
                 forvar7098,
                 forvar7093,
                 reg7094,
                 forvar7090,
                 reg7089,
                 forvar7086,
                 reg7146,
                 forvar7139,
                 reg7145,
                 forvar7143,
                 reg7140,
                 forvar7138,
                 forvar7136,
                 reg7135,
                 forvar7131,
                 reg7130,
                 reg7126,
                 forvar7123,
                 forvar7121,
                 reg7120,
                 forvar7112,
                 forvar7111,
                 forvar7106,
                 reg7144,
                 reg7143,
                 reg7142,
                 reg7141,
                 forvar7140,
                 reg7139,
                 reg7138,
                 reg7137,
                 reg7136,
                 forvar7135,
                 reg7134,
                 reg7133,
                 reg7132,
                 reg7131,
                 forvar7130,
                 reg7129,
                 reg7128,
                 reg7127,
                 forvar7126,
                 reg7125,
                 reg7124,
                 reg7123,
                 reg7122,
                 reg7121,
                 forvar7120,
                 reg7119,
                 reg7118,
                 reg7117,
                 reg7116,
                 reg7115,
                 reg7114,
                 reg7113,
                 reg7112,
                 reg7111,
                 reg7110,
                 reg7109,
                 reg7108,
                 reg7107,
                 reg7106,
                 reg7105,
                 forvar7104,
                 reg7088,
                 forvar7087,
                 reg7103,
                 reg7102,
                 reg7101,
                 reg7100,
                 reg7099,
                 reg7098,
                 reg7097,
                 reg7096,
                 reg7095,
                 forvar7094,
                 reg7093,
                 reg7092,
                 reg7091,
                 reg7090,
                 forvar7089,
                 forvar7088,
                 reg7087,
                 reg7086,
                 reg7085,
                 reg7084,
                 reg7083,
                 reg7082,
                 reg7081,
                 reg7080,
                 forvar7079,
                 reg7078,
                 reg7077,
                 reg7076,
                 reg7075,
                 reg7074,
                 forvar7071,
                 reg7073,
                 reg7072,
                 reg7071,
                 reg7070,
                 forvar7069,
                 forvar7068,
                 reg7067,
                 reg7066,
                 reg7065,
                 reg7064,
                 forvar7063,
                 reg7062,
                 reg7061,
                 reg7060,
                 reg7059,
                 reg7058,
                 reg7057,
                 reg7056,
                 reg7055,
                 forvar7054,
                 reg7053,
                 reg7052,
                 reg7051,
                 reg7050,
                 forvar7049,
                 forvar7048,
                 forvar7047,
                 forvar7044,
                 forvar7040,
                 reg7046,
                 reg7045,
                 reg7044,
                 reg7043,
                 reg7042,
                 reg7041,
                 reg7040,
                 reg7039,
                 reg7038,
                 forvar7037,
                 forvar7033,
                 reg7030,
                 reg7036,
                 reg7035,
                 reg7034,
                 reg7033,
                 reg7032,
                 reg7031,
                 forvar7030,
                 reg7029,
                 reg7028,
                 reg7027,
                 reg7026,
                 reg7025,
                 reg7024,
                 forvar7023,
                 reg7022,
                 reg7021,
                 reg7020,
                 reg7019,
                 reg7018,
                 reg7017,
                 reg7016,
                 reg7015,
                 reg7014,
                 reg7013,
                 forvar7012,
                 forvar7011,
                 forvar7010,
                 wire7009,
                 wire7008,
                 wire7006,
                 wire4571,
                 reg4570,
                 reg4569,
                 forvar4568,
                 forvar4567,
                 reg4566,
                 reg4565,
                 reg4564,
                 reg4563,
                 reg4562,
                 forvar4561,
                 reg4560,
                 reg4559,
                 forvar4558,
                 reg4557,
                 forvar4556,
                 reg4555,
                 forvar4554,
                 forvar4553,
                 reg4552,
                 reg4551,
                 reg4550,
                 reg4549,
                 reg4548,
                 forvar4547,
                 forvar4546,
                 reg4545,
                 reg4544,
                 reg4543,
                 forvar4542,
                 reg4538,
                 forvar4537,
                 reg4542,
                 reg4541,
                 reg4540,
                 reg4539,
                 forvar4538,
                 reg4537,
                 reg4536,
                 forvar4535,
                 forvar4522,
                 reg4520,
                 reg4534,
                 reg4533,
                 reg4532,
                 reg4531,
                 forvar4530,
                 reg4529,
                 reg4528,
                 forvar4527,
                 reg4526,
                 reg4525,
                 reg4524,
                 reg4523,
                 reg4522,
                 reg4521,
                 forvar4520,
                 reg4519,
                 forvar4518,
                 reg4517,
                 reg4510,
                 forvar4509,
                 forvar4506,
                 reg4516,
                 reg4515,
                 reg4514,
                 reg4513,
                 reg4512,
                 reg4511,
                 forvar4510,
                 reg4509,
                 reg4508,
                 forvar4503,
                 reg4496,
                 forvar4490,
                 reg4489,
                 reg4487,
                 reg4486,
                 forvar4485,
                 reg4482,
                 reg4507,
                 forvar4504,
                 forvar4501,
                 reg4500,
                 reg4506,
                 reg4505,
                 reg4504,
                 reg4503,
                 reg4502,
                 reg4501,
                 forvar4500,
                 reg4499,
                 reg4498,
                 reg4497,
                 forvar4496,
                 reg4495,
                 reg4494,
                 reg4493,
                 reg4492,
                 reg4491,
                 reg4490,
                 forvar4489,
                 reg4488,
                 forvar4487,
                 forvar4486,
                 reg4485,
                 reg4484,
                 reg4483,
                 forvar4482,
                 reg4481,
                 reg4480,
                 reg4479,
                 reg4478,
                 reg4477,
                 forvar4476,
                 forvar4475,
                 reg4474,
                 reg4473,
                 reg4472,
                 reg4471,
                 reg4470,
                 reg4469,
                 reg4468,
                 forvar4467,
                 reg4466,
                 reg4465,
                 forvar4464,
                 reg4463,
                 reg4462,
                 reg4461,
                 reg4459,
                 reg4457,
                 reg4460,
                 forvar4459,
                 reg4458,
                 forvar4457,
                 forvar4456,
                 reg4455,
                 forvar4454,
                 reg4453,
                 reg4452,
                 reg4451,
                 reg4450,
                 forvar4449,
                 reg4448,
                 reg4447,
                 reg4446,
                 reg4445,
                 reg4444,
                 reg4443,
                 reg4442,
                 reg4441,
                 forvar4440,
                 reg4439,
                 reg4438,
                 forvar4437,
                 forvar4436,
                 reg4435,
                 reg4434,
                 reg4433,
                 reg4432,
                 forvar4427,
                 reg4424,
                 reg4423,
                 forvar4422,
                 forvar4414,
                 forvar4412,
                 reg4431,
                 reg4430,
                 reg4429,
                 reg4428,
                 reg4427,
                 reg4426,
                 reg4425,
                 forvar4424,
                 forvar4423,
                 reg4422,
                 reg4418,
                 forvar4413,
                 reg4421,
                 reg4420,
                 reg4419,
                 forvar4418,
                 reg4417,
                 reg4416,
                 reg4415,
                 reg4414,
                 reg4413,
                 reg4412,
                 reg4411,
                 reg4410,
                 reg4409,
                 forvar4408,
                 reg4407,
                 reg4406,
                 reg4405,
                 reg4404,
                 forvar4403,
                 reg4402,
                 forvar4401,
                 reg4400,
                 reg4391,
                 forvar4386,
                 reg4399,
                 reg4398,
                 reg4397,
                 reg4396,
                 reg4395,
                 reg4394,
                 reg4393,
                 reg4392,
                 forvar4391,
                 reg4390,
                 forvar4389,
                 reg4388,
                 reg4387,
                 reg4386,
                 reg4385,
                 reg4384,
                 reg4383,
                 reg4382,
                 reg4381,
                 reg4380,
                 reg4379,
                 reg4378,
                 reg4377,
                 forvar4375,
                 forvar4372,
                 reg4369,
                 reg4376,
                 reg4375,
                 forvar4374,
                 reg4373,
                 reg4372,
                 reg4371,
                 reg4370,
                 forvar4369,
                 forvar4368,
                 reg4367,
                 reg4366,
                 reg4365,
                 forvar4364,
                 reg4359,
                 reg4363,
                 reg4362,
                 reg4361,
                 reg4360,
                 forvar4359,
                 reg4356,
                 forvar4353,
                 reg4352,
                 forvar4350,
                 reg4347,
                 forvar4345,
                 reg4358,
                 reg4357,
                 forvar4356,
                 reg4355,
                 reg4354,
                 reg4353,
                 forvar4352,
                 reg4351,
                 reg4350,
                 reg4349,
                 reg4348,
                 forvar4347,
                 forvar4346,
                 reg4345,
                 forvar4344,
                 wire4343,
                 wire4342,
                 (1'h0)};
  assign wire4342 = wire4338;
  assign wire4343 = wire4342[(1'h1):(1'h1)];
  always
    @(posedge clk) begin
      if (wire4341)
        begin
          for (forvar4344 = (1'h0); (forvar4344 < (2'h3)); forvar4344 = (forvar4344 + (1'h1)))
            begin
              reg4345 <= ({wire4343[(2'h3):(1'h0)]} ?
                  wire4338 : $unsigned(wire4339[(2'h3):(1'h0)]));
              for (forvar4346 = (1'h0); (forvar4346 < (2'h3)); forvar4346 = (forvar4346 + (1'h1)))
                begin
                  for (forvar4347 = (1'h0); (forvar4347 < (2'h3)); forvar4347 = (forvar4347 + (1'h1)))
                    begin
                      reg4348 <= (forvar4344[(4'h8):(1'h0)] ?
                          $unsigned(wire4343[(4'h9):(3'h7)]) : $signed(($signed(forvar4344) ?
                              forvar4346[(4'ha):(1'h1)] : {forvar4344})));
                      reg4349 <= (^~$signed(($unsigned(forvar4347) ?
                          (8'ha4) : ((8'ha1) || wire4341))));
                      reg4350 <= $signed($signed($signed(wire4339[(1'h1):(1'h0)])));
                    end
                end
              reg4351 <= ($unsigned((-$unsigned(wire4340))) <= $signed(wire4342));
              for (forvar4352 = (1'h0); (forvar4352 < (1'h0)); forvar4352 = (forvar4352 + (1'h1)))
                begin
                  if ((^($signed((forvar4352 || wire4341)) ^ $signed({forvar4347}))))
                    begin
                      reg4353 <= ($unsigned((-{wire4342})) ?
                          wire4340[(2'h3):(2'h2)] : $signed((((8'hba) ?
                              wire4338 : (8'ha2)) < $unsigned(wire4343))));
                    end
                  else
                    begin
                      reg4353 <= (+forvar4344);
                      reg4354 <= forvar4346[(2'h3):(2'h3)];
                    end
                end
            end
          reg4355 <= (~&(((~^forvar4352) + (~|reg4349)) ?
              (((8'ha3) ? reg4345 : wire4338) < (+reg4348)) : (8'had)));
          for (forvar4356 = (1'h0); (forvar4356 < (1'h1)); forvar4356 = (forvar4356 + (1'h1)))
            begin
              reg4357 <= (reg4345 ?
                  ($unsigned($unsigned(wire4342)) == (forvar4356[(3'h6):(3'h4)] ?
                      forvar4346[(2'h3):(1'h1)] : (reg4354 ?
                          forvar4344 : (8'haf)))) : $signed($signed((forvar4356 ?
                      reg4353 : reg4345))));
              reg4358 <= (^~(($signed(reg4355) ?
                  $signed(wire4340) : reg4345) < $signed((~|reg4349))));
            end
        end
      else
        begin
          for (forvar4344 = (1'h0); (forvar4344 < (1'h0)); forvar4344 = (forvar4344 + (1'h1)))
            begin
              for (forvar4345 = (1'h0); (forvar4345 < (2'h3)); forvar4345 = (forvar4345 + (1'h1)))
                begin
                  for (forvar4346 = (1'h0); (forvar4346 < (1'h0)); forvar4346 = (forvar4346 + (1'h1)))
                    begin
                      reg4347 <= (8'hb0);
                      reg4348 <= $unsigned((forvar4344 >>> {{forvar4352}}));
                      reg4349 <= ({((forvar4347 <= forvar4347) != reg4354)} ?
                          (8'haf) : (~&$unsigned($unsigned(wire4339))));
                    end
                  for (forvar4350 = (1'h0); (forvar4350 < (2'h3)); forvar4350 = (forvar4350 + (1'h1)))
                    begin
                      reg4351 <= ($signed(reg4345[(3'h7):(3'h7)]) ?
                          forvar4346[(1'h0):(1'h0)] : (!((reg4357 || wire4338) != forvar4356[(2'h2):(1'h0)])));
                      reg4352 <= {(wire4340 ?
                              forvar4356[(3'h4):(2'h2)] : (|(reg4357 - forvar4356)))};
                    end
                end
              for (forvar4353 = (1'h0); (forvar4353 < (1'h1)); forvar4353 = (forvar4353 + (1'h1)))
                begin
                  if ((^~($signed(forvar4345) > (8'ha6))))
                    begin
                      reg4354 <= $signed((~^(^~(reg4358 ? reg4350 : reg4348))));
                      reg4355 <= wire4343;
                      reg4356 <= (~(8'ha6));
                    end
                  else
                    begin
                      reg4354 <= (~forvar4344);
                      reg4355 <= reg4351[(1'h1):(1'h0)];
                      reg4356 <= (-forvar4350[(1'h0):(1'h0)]);
                      reg4357 <= ((($signed(reg4351) >> (|reg4355)) >= {(^reg4345)}) ?
                          $unsigned((reg4357[(1'h1):(1'h1)] ?
                              $unsigned((8'ha1)) : {forvar4347})) : (+forvar4356));
                    end
                end
              if ({$signed(reg4358)})
                begin
                  reg4358 <= wire4339[(3'h5):(2'h2)];
                  for (forvar4359 = (1'h0); (forvar4359 < (1'h1)); forvar4359 = (forvar4359 + (1'h1)))
                    begin
                      reg4360 <= wire4339;
                    end
                  if (wire4343)
                    begin
                      reg4361 <= reg4354;
                      reg4362 <= ($signed((-(8'hb8))) ^~ {$signed($signed(forvar4359))});
                    end
                  else
                    begin
                      reg4361 <= forvar4347;
                      reg4362 <= forvar4346;
                      reg4363 <= {forvar4359};
                    end
                end
              else
                begin
                  if (($unsigned(((wire4339 - forvar4346) & $signed(wire4340))) ~^ $unsigned($signed(reg4347))))
                    begin
                      reg4358 <= forvar4359;
                      reg4359 <= $unsigned(((reg4349 ^~ $signed(reg4347)) ?
                          ((wire4342 ? wire4342 : reg4348) ?
                              $signed(reg4361) : (reg4347 >> (8'ha8))) : (reg4354[(3'h6):(1'h0)] ?
                              {reg4357} : wire4338)));
                      reg4360 <= ($signed({$unsigned(reg4354)}) ?
                          (((forvar4350 && forvar4344) ?
                                  (wire4342 ?
                                      reg4349 : reg4345) : (reg4354 << reg4360)) ?
                              (&(forvar4344 >>> reg4352)) : $signed($unsigned((8'ha7)))) : reg4356);
                      reg4361 <= {$signed($unsigned($signed(forvar4344)))};
                    end
                  else
                    begin
                      reg4358 <= ($signed($unsigned((reg4352 ~^ forvar4345))) ?
                          $signed($unsigned($signed(reg4348))) : $unsigned((((8'ha1) ?
                                  forvar4346 : wire4342) ?
                              (forvar4356 != forvar4344) : wire4341)));
                      reg4359 <= forvar4345;
                      reg4360 <= $unsigned((({reg4345} * {wire4342}) != {$signed(forvar4359)}));
                    end
                  reg4362 <= $unsigned((reg4351[(1'h0):(1'h0)] ?
                      {wire4343[(3'h4):(2'h3)]} : forvar4346[(4'h9):(3'h5)]));
                  reg4363 <= reg4355;
                end
              for (forvar4364 = (1'h0); (forvar4364 < (2'h3)); forvar4364 = (forvar4364 + (1'h1)))
                begin
                  if (((8'ha4) << {($unsigned(reg4363) * {wire4341})}))
                    begin
                      reg4365 <= ((({(8'hb7)} <= (^~(8'had))) ?
                              reg4352 : $signed($signed(reg4363))) ?
                          (((reg4347 <<< reg4349) ?
                                  wire4342[(3'h4):(2'h2)] : (~&forvar4364)) ?
                              forvar4359[(1'h1):(1'h1)] : reg4350[(1'h0):(1'h0)]) : ($unsigned({forvar4347}) && (^~reg4359[(2'h3):(2'h2)])));
                      reg4366 <= (reg4362[(1'h0):(1'h0)] || (&(-(reg4351 > wire4341))));
                    end
                  else
                    begin
                      reg4365 <= ($unsigned($signed((~|reg4347))) ?
                          $signed({(reg4349 ?
                                  forvar4350 : reg4350)}) : $signed(forvar4346));
                      reg4366 <= ((reg4353[(4'ha):(2'h2)] ?
                              (((8'hb6) ? forvar4364 : forvar4364) ?
                                  $unsigned(reg4350) : $unsigned(forvar4352)) : ((reg4349 ?
                                      forvar4346 : wire4340) ?
                                  (reg4359 ?
                                      forvar4346 : reg4365) : (wire4343 >>> forvar4347))) ?
                          reg4360 : reg4352[(1'h1):(1'h1)]);
                      reg4367 <= ((reg4358[(1'h1):(1'h1)] ?
                              (((8'ha8) ? reg4352 : reg4357) ?
                                  wire4341 : forvar4364[(1'h0):(1'h0)]) : (&$unsigned(reg4355))) ?
                          wire4339[(2'h2):(1'h1)] : (((reg4354 <= reg4357) ?
                              (-reg4352) : $unsigned(reg4354)) == (-(forvar4345 ?
                              reg4345 : forvar4353))));
                    end
                end
            end
        end
      for (forvar4368 = (1'h0); (forvar4368 < (2'h2)); forvar4368 = (forvar4368 + (1'h1)))
        begin
          if ($signed((($signed(wire4339) >= $unsigned(reg4352)) ^ (reg4365 ?
              (!forvar4353) : $signed(forvar4353)))))
            begin
              for (forvar4369 = (1'h0); (forvar4369 < (1'h0)); forvar4369 = (forvar4369 + (1'h1)))
                begin
                  if ($signed($signed(forvar4346[(4'he):(4'hc)])))
                    begin
                      reg4370 <= wire4338;
                      reg4371 <= ($signed($signed(reg4363)) < $unsigned((8'hb6)));
                      reg4372 <= $signed(reg4356[(4'hd):(3'h5)]);
                    end
                  else
                    begin
                      reg4370 <= wire4343;
                      reg4371 <= reg4348[(4'h9):(1'h1)];
                      reg4372 <= {(forvar4364 - ($signed(wire4338) >= (~reg4349)))};
                      reg4373 <= ($unsigned(forvar4347[(2'h3):(1'h1)]) ?
                          (reg4371 << {reg4358[(3'h7):(3'h5)]}) : reg4355[(3'h6):(1'h0)]);
                    end
                end
              for (forvar4374 = (1'h0); (forvar4374 < (2'h2)); forvar4374 = (forvar4374 + (1'h1)))
                begin
                  reg4375 <= (forvar4356[(4'h9):(4'h8)] >= $unsigned($signed((^~forvar4369))));
                  reg4376 <= reg4355[(3'h5):(3'h5)];
                end
            end
          else
            begin
              if ((8'h9e))
                begin
                  if ($signed((reg4376 ? reg4359 : $unsigned((~|(8'ha4))))))
                    begin
                      reg4369 <= (forvar4352[(1'h1):(1'h0)] ?
                          ($unsigned(reg4359[(3'h6):(3'h5)]) ?
                              forvar4374[(1'h1):(1'h0)] : (reg4352[(4'hb):(1'h0)] ?
                                  (reg4365 ? (8'hb7) : reg4347) : (reg4359 ?
                                      reg4375 : wire4338))) : reg4376);
                      reg4370 <= (reg4348[(1'h0):(1'h0)] && reg4351);
                      reg4371 <= $signed(forvar4350);
                    end
                  else
                    begin
                      reg4369 <= reg4356;
                      reg4370 <= ((~|$signed($signed(forvar4347))) | {(((8'hae) >> reg4352) ^~ {wire4342})});
                    end
                  for (forvar4372 = (1'h0); (forvar4372 < (1'h1)); forvar4372 = (forvar4372 + (1'h1)))
                    begin
                      reg4373 <= reg4350[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  if ({(+(+wire4339[(3'h5):(1'h0)]))})
                    begin
                      reg4369 <= (-reg4359);
                      reg4370 <= (reg4347 + ((-(^~(8'ha4))) + wire4340));
                      reg4371 <= {(~|(~$unsigned(reg4356)))};
                    end
                  else
                    begin
                      reg4369 <= reg4354[(3'h6):(3'h5)];
                      reg4370 <= (reg4372[(1'h0):(1'h0)] != $unsigned($signed(reg4360[(2'h3):(1'h0)])));
                      reg4371 <= reg4360[(3'h6):(3'h6)];
                    end
                  reg4372 <= $signed($unsigned(((reg4375 * reg4373) && (8'ha9))));
                end
              for (forvar4374 = (1'h0); (forvar4374 < (2'h3)); forvar4374 = (forvar4374 + (1'h1)))
                begin
                  for (forvar4375 = (1'h0); (forvar4375 < (1'h0)); forvar4375 = (forvar4375 + (1'h1)))
                    begin
                      reg4376 <= $signed({(^(~&reg4348))});
                    end
                  reg4377 <= $unsigned(($unsigned(forvar4353) >>> (forvar4352 >= $unsigned(wire4339))));
                  if (reg4353[(4'ha):(3'h5)])
                    begin
                      reg4378 <= $unsigned($signed($signed((reg4352 ?
                          reg4367 : reg4348))));
                      reg4379 <= ($signed($signed((forvar4356 ?
                              reg4371 : (8'hb6)))) ?
                          (reg4357[(1'h0):(1'h0)] ?
                              ($signed(reg4349) ?
                                  (~reg4366) : $signed(forvar4347)) : (~(wire4341 >> forvar4375))) : (($signed(reg4355) ?
                                  reg4355 : (forvar4344 ^~ reg4366)) ?
                              {(~reg4350)} : {$signed(reg4365)}));
                      reg4380 <= (&{$unsigned((reg4353 ? reg4350 : reg4376))});
                      reg4381 <= reg4378[(4'hd):(3'h5)];
                    end
                  else
                    begin
                      reg4378 <= reg4362[(1'h1):(1'h1)];
                      reg4379 <= reg4353;
                    end
                  if ((8'hb1))
                    begin
                      reg4382 <= (^(~&reg4375));
                      reg4383 <= (~((~|$unsigned(forvar4368)) ?
                          (reg4354[(3'h7):(2'h3)] ?
                              $signed((8'hb3)) : $unsigned(reg4352)) : (|(forvar4353 >>> reg4373))));
                      reg4384 <= (~($signed({reg4350}) | (+(~^forvar4353))));
                    end
                  else
                    begin
                      reg4382 <= (reg4383[(3'h5):(1'h0)] || $signed(($unsigned((8'ha0)) ?
                          reg4379 : (wire4340 || (8'hab)))));
                      reg4383 <= forvar4368;
                      reg4384 <= (~|$unsigned($unsigned(reg4362[(3'h7):(3'h5)])));
                      reg4385 <= wire4342;
                    end
                end
            end
          if ((&$signed({wire4338})))
            begin
              reg4386 <= reg4369;
            end
          else
            begin
              if ($unsigned(forvar4372[(1'h1):(1'h0)]))
                begin
                  if ($unsigned((-(reg4366[(3'h7):(3'h7)] ?
                      (^reg4360) : reg4383))))
                    begin
                      reg4386 <= (~^($signed($signed(forvar4346)) ?
                          reg4351[(1'h0):(1'h0)] : wire4343[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg4386 <= $signed(wire4339[(3'h5):(3'h5)]);
                      reg4387 <= forvar4364;
                      reg4388 <= (~&$signed(wire4341[(4'h9):(4'h9)]));
                    end
                  for (forvar4389 = (1'h0); (forvar4389 < (2'h3)); forvar4389 = (forvar4389 + (1'h1)))
                    begin
                      reg4390 <= (^$signed($signed($unsigned(reg4353))));
                    end
                  for (forvar4391 = (1'h0); (forvar4391 < (1'h0)); forvar4391 = (forvar4391 + (1'h1)))
                    begin
                      reg4392 <= ($unsigned(((~^wire4341) ?
                          (8'hab) : $unsigned(reg4365))) ^~ (($signed(reg4363) == (forvar4391 ?
                              reg4357 : reg4365)) ?
                          reg4386 : reg4387[(4'he):(3'h5)]));
                      reg4393 <= $signed($signed((forvar4369 ?
                          reg4359 : reg4347)));
                      reg4394 <= ($signed((!reg4365[(3'h5):(2'h2)])) ?
                          ($signed($unsigned(forvar4353)) ~^ ((forvar4364 <<< forvar4346) ^ (forvar4359 ?
                              forvar4374 : reg4345))) : ({(~reg4348)} ?
                              (~reg4376) : (|{reg4379})));
                      reg4395 <= $signed(((8'hba) ?
                          forvar4352 : ({reg4388} ?
                              $signed(reg4380) : (forvar4389 == (8'hb2)))));
                    end
                  if (forvar4347)
                    begin
                      reg4396 <= reg4380[(4'h9):(3'h4)];
                      reg4397 <= reg4347[(4'hb):(3'h4)];
                    end
                  else
                    begin
                      reg4396 <= $signed(($unsigned(reg4347[(1'h1):(1'h0)]) + (8'h9f)));
                      reg4397 <= $unsigned(reg4387);
                      reg4398 <= reg4395;
                      reg4399 <= (~$unsigned($signed({forvar4368})));
                    end
                end
              else
                begin
                  for (forvar4386 = (1'h0); (forvar4386 < (2'h3)); forvar4386 = (forvar4386 + (1'h1)))
                    begin
                      reg4387 <= (reg4349 ? reg4348 : $unsigned(reg4379));
                    end
                  reg4388 <= (+reg4365);
                  for (forvar4389 = (1'h0); (forvar4389 < (2'h2)); forvar4389 = (forvar4389 + (1'h1)))
                    begin
                      reg4390 <= wire4339;
                      reg4391 <= (wire4342[(4'hc):(4'hc)] ?
                          $signed($unsigned($signed(reg4373))) : forvar4369[(3'h5):(3'h4)]);
                      reg4392 <= $signed($signed($signed($signed(forvar4372))));
                      reg4393 <= ($signed($unsigned((reg4362 <= (8'hac)))) ?
                          ($signed($unsigned((8'ha6))) ?
                              ($unsigned(reg4393) ~^ $signed(forvar4386)) : $unsigned($signed((8'ha9)))) : $signed($signed(reg4371)));
                    end
                  if (reg4345)
                    begin
                      reg4394 <= ((forvar4352[(1'h1):(1'h0)] ?
                              reg4352 : (forvar4359[(1'h1):(1'h1)] < reg4350[(1'h0):(1'h0)])) ?
                          forvar4372 : (~^$unsigned($unsigned(forvar4359))));
                    end
                  else
                    begin
                      reg4394 <= $unsigned((reg4348[(3'h5):(1'h1)] ?
                          (-{forvar4347}) : $signed({reg4385})));
                      reg4395 <= reg4388;
                      reg4396 <= $signed((reg4373 >= forvar4345));
                    end
                end
              if ($signed($unsigned($signed(forvar4359))))
                begin
                  reg4400 <= {$signed((&(~reg4376)))};
                end
              else
                begin
                  reg4400 <= ((reg4399[(3'h7):(2'h2)] > (-forvar4350[(4'h9):(4'h8)])) ?
                      $unsigned(($unsigned(forvar4375) >= reg4360)) : (8'had));
                end
              for (forvar4401 = (1'h0); (forvar4401 < (1'h1)); forvar4401 = (forvar4401 + (1'h1)))
                begin
                  reg4402 <= (reg4350[(2'h2):(1'h1)] ?
                      reg4397[(2'h2):(1'h0)] : $unsigned((8'hb0)));
                  for (forvar4403 = (1'h0); (forvar4403 < (1'h0)); forvar4403 = (forvar4403 + (1'h1)))
                    begin
                      reg4404 <= {(((-(8'ha2)) <<< $unsigned(reg4375)) ?
                              $unsigned(reg4394) : reg4396)};
                      reg4405 <= ((8'hae) ?
                          ({{reg4370}} == ((forvar4374 ? reg4392 : forvar4386) ?
                              (reg4384 ?
                                  forvar4369 : forvar4368) : (^~reg4371))) : wire4339);
                      reg4406 <= (~^($signed($unsigned(reg4365)) < ((|(8'hb3)) <= reg4378)));
                      reg4407 <= $signed($signed(forvar4352));
                    end
                  for (forvar4408 = (1'h0); (forvar4408 < (2'h2)); forvar4408 = (forvar4408 + (1'h1)))
                    begin
                      reg4409 <= ((^~$unsigned($signed(reg4366))) ?
                          forvar4350[(3'h6):(3'h5)] : $unsigned((((8'ha5) << reg4355) ?
                              $signed(wire4340) : reg4393)));
                      reg4410 <= {({reg4400} ?
                              $signed((reg4406 ^~ reg4379)) : $unsigned($signed(forvar4345)))};
                    end
                  reg4411 <= reg4404;
                end
            end
          if ($signed(reg4394))
            begin
              reg4412 <= $signed({forvar4368[(2'h3):(1'h1)]});
              if (reg4400[(3'h5):(1'h0)])
                begin
                  if (reg4400)
                    begin
                      reg4413 <= reg4412[(1'h1):(1'h0)];
                      reg4414 <= $signed((8'hac));
                    end
                  else
                    begin
                      reg4413 <= wire4339;
                      reg4414 <= ((~^(^~(wire4341 && wire4342))) >= reg4407);
                    end
                  reg4415 <= $signed($signed($unsigned(reg4363[(3'h4):(3'h4)])));
                  if ($unsigned((reg4405[(3'h6):(2'h2)] ?
                      $signed((&reg4383)) : $signed({reg4363}))))
                    begin
                      reg4416 <= $signed((((wire4339 ?
                              reg4395 : reg4366) && reg4397) ?
                          ((8'hb3) | $unsigned(forvar4372)) : reg4388[(4'hb):(2'h3)]));
                    end
                  else
                    begin
                      reg4416 <= $signed((reg4355 != (~|(|(8'h9c)))));
                      reg4417 <= (&(8'hab));
                    end
                  for (forvar4418 = (1'h0); (forvar4418 < (1'h0)); forvar4418 = (forvar4418 + (1'h1)))
                    begin
                      reg4419 <= ((!(8'ha5)) >>> ((wire4343[(2'h3):(2'h2)] ?
                          ((8'h9d) ?
                              reg4359 : forvar4345) : reg4409) - ((~^reg4398) <<< (reg4354 * (8'hb8)))));
                      reg4420 <= (~|(~&$unsigned((reg4376 != forvar4391))));
                      reg4421 <= (reg4377[(1'h1):(1'h0)] ?
                          ({reg4378[(4'he):(2'h2)]} ?
                              $signed((~^wire4339)) : (~&(8'h9d))) : reg4356[(3'h4):(3'h4)]);
                    end
                end
              else
                begin
                  for (forvar4413 = (1'h0); (forvar4413 < (2'h3)); forvar4413 = (forvar4413 + (1'h1)))
                    begin
                      reg4414 <= reg4361[(4'h8):(2'h2)];
                    end
                  if ($unsigned($unsigned((reg4372 ? {reg4385} : forvar4386))))
                    begin
                      reg4415 <= reg4370;
                    end
                  else
                    begin
                      reg4415 <= {reg4367};
                      reg4416 <= wire4338;
                      reg4417 <= $signed((forvar4391[(3'h6):(1'h1)] ?
                          $unsigned($signed((8'hb0))) : (&reg4369[(2'h2):(1'h1)])));
                      reg4418 <= forvar4403[(3'h7):(2'h2)];
                    end
                  if (($unsigned(reg4421) ?
                      ((~^(reg4385 ?
                          reg4418 : reg4361)) | reg4369[(1'h1):(1'h1)]) : $signed(((reg4413 ?
                          reg4347 : reg4395) | (forvar4372 >>> forvar4403)))))
                    begin
                      reg4419 <= (&reg4412);
                      reg4420 <= $signed($unsigned(reg4351[(2'h3):(2'h3)]));
                      reg4421 <= ($signed((!(^reg4378))) << $unsigned($signed((reg4375 > reg4376))));
                      reg4422 <= reg4354;
                    end
                  else
                    begin
                      reg4419 <= reg4412;
                      reg4420 <= ((-$signed((reg4417 || reg4410))) ?
                          {(reg4417[(3'h6):(2'h3)] ~^ $unsigned((8'ha0)))} : ((!{(8'ha7)}) ?
                              reg4352[(3'h5):(3'h5)] : ((reg4359 ?
                                  forvar4375 : reg4394) ~^ reg4390)));
                    end
                end
              for (forvar4423 = (1'h0); (forvar4423 < (2'h2)); forvar4423 = (forvar4423 + (1'h1)))
                begin
                  for (forvar4424 = (1'h0); (forvar4424 < (1'h0)); forvar4424 = (forvar4424 + (1'h1)))
                    begin
                      reg4425 <= reg4351[(2'h2):(1'h1)];
                      reg4426 <= $signed((|$signed($signed(reg4407))));
                      reg4427 <= forvar4408[(1'h1):(1'h1)];
                    end
                  if (reg4391)
                    begin
                      reg4428 <= ($unsigned(($unsigned(reg4426) ^~ $signed(reg4394))) ?
                          wire4343[(2'h3):(1'h0)] : ({(reg4421 * (8'haf))} << $unsigned(reg4406[(1'h1):(1'h1)])));
                      reg4429 <= reg4416[(4'ha):(4'h8)];
                      reg4430 <= (|reg4414[(1'h1):(1'h1)]);
                      reg4431 <= ($unsigned((^reg4365[(3'h5):(1'h0)])) <= {$unsigned(reg4357[(2'h2):(1'h0)])});
                    end
                  else
                    begin
                      reg4428 <= (reg4347 ^ $unsigned(reg4370));
                      reg4429 <= forvar4418[(4'h9):(3'h7)];
                      reg4430 <= (((^forvar4408) ^ $unsigned((wire4339 ?
                              (8'h9c) : reg4412))) ?
                          ((|$unsigned((8'ha2))) > forvar4369) : (reg4365[(4'h9):(4'h8)] <<< ($signed(reg4391) ?
                              forvar4423[(4'h8):(1'h0)] : (reg4384 ?
                                  forvar4359 : forvar4389))));
                    end
                end
            end
          else
            begin
              if ($signed(reg4421))
                begin
                  for (forvar4412 = (1'h0); (forvar4412 < (1'h1)); forvar4412 = (forvar4412 + (1'h1)))
                    begin
                      reg4413 <= {((reg4379[(4'h8):(3'h6)] - (reg4422 ?
                                  reg4398 : forvar4369)) ?
                              (-(reg4426 < reg4360)) : $unsigned($unsigned(reg4376)))};
                    end
                  for (forvar4414 = (1'h0); (forvar4414 < (1'h1)); forvar4414 = (forvar4414 + (1'h1)))
                    begin
                      reg4415 <= $unsigned((~|$unsigned({forvar4424})));
                      reg4416 <= $signed((reg4415[(1'h0):(1'h0)] - reg4381[(3'h6):(1'h0)]));
                      reg4417 <= {{forvar4413[(2'h2):(2'h2)]}};
                    end
                  for (forvar4418 = (1'h0); (forvar4418 < (2'h2)); forvar4418 = (forvar4418 + (1'h1)))
                    begin
                      reg4419 <= (reg4384[(3'h4):(1'h1)] & reg4385);
                      reg4420 <= (!reg4394[(1'h0):(1'h0)]);
                      reg4421 <= {wire4342};
                    end
                  for (forvar4422 = (1'h0); (forvar4422 < (1'h1)); forvar4422 = (forvar4422 + (1'h1)))
                    begin
                      reg4423 <= (+((reg4351 || $signed((8'hb3))) ?
                          ($unsigned(reg4372) ?
                              (reg4405 ? reg4404 : forvar4347) : (reg4394 ?
                                  (8'h9f) : reg4358)) : $signed($signed(reg4411))));
                      reg4424 <= reg4390;
                      reg4425 <= $signed({reg4355});
                      reg4426 <= reg4420[(4'h9):(1'h1)];
                    end
                end
              else
                begin
                  if ($signed((reg4430[(3'h7):(2'h3)] ?
                      reg4423 : ({reg4427} | (forvar4346 ~^ reg4349)))))
                    begin
                      reg4412 <= $unsigned((8'haf));
                      reg4413 <= reg4402[(1'h1):(1'h0)];
                      reg4414 <= reg4371;
                      reg4415 <= $unsigned((reg4422 ?
                          reg4398 : (reg4369 ?
                              ((8'ha8) ?
                                  (8'ha3) : reg4392) : (wire4338 * (8'hac)))));
                    end
                  else
                    begin
                      reg4412 <= (reg4418[(3'h7):(3'h5)] <= reg4428[(1'h1):(1'h1)]);
                      reg4413 <= (!$unsigned($unsigned((8'ha8))));
                      reg4414 <= ($unsigned($unsigned((forvar4347 ?
                          forvar4391 : reg4413))) * {(~(reg4404 ^ (8'hb4)))});
                    end
                end
              if (reg4349[(4'hb):(4'h8)])
                begin
                  for (forvar4427 = (1'h0); (forvar4427 < (2'h2)); forvar4427 = (forvar4427 + (1'h1)))
                    begin
                      reg4428 <= reg4423[(2'h2):(1'h0)];
                    end
                  if ({(|(^~(reg4357 ? (8'had) : wire4340)))})
                    begin
                      reg4429 <= ($signed($unsigned((8'hab))) ?
                          $signed($signed((|reg4355))) : ((8'hb1) ^ forvar4372[(2'h3):(2'h2)]));
                      reg4430 <= forvar4353[(3'h6):(1'h0)];
                      reg4431 <= reg4366[(3'h4):(2'h2)];
                      reg4432 <= $unsigned($unsigned({$unsigned(reg4404)}));
                    end
                  else
                    begin
                      reg4429 <= $signed($unsigned((|(reg4432 ?
                          reg4400 : reg4421))));
                      reg4430 <= ($signed((reg4415 & $signed(reg4412))) - (|reg4399[(4'h9):(4'h8)]));
                      reg4431 <= {reg4409};
                      reg4432 <= reg4409;
                    end
                  if (forvar4422)
                    begin
                      reg4433 <= forvar4346;
                    end
                  else
                    begin
                      reg4433 <= ($unsigned(wire4342[(4'hf):(3'h7)]) ?
                          reg4428 : $signed(($signed(forvar4412) ?
                              (8'ha6) : wire4342[(3'h4):(1'h1)])));
                      reg4434 <= $unsigned(forvar4389[(2'h3):(1'h1)]);
                    end
                  reg4435 <= ((-reg4423[(1'h0):(1'h0)]) ?
                      ($unsigned((8'hb3)) ?
                          $unsigned($unsigned(reg4350)) : ($signed(reg4404) ?
                              reg4394[(1'h0):(1'h0)] : forvar4364)) : $signed((~^$unsigned(reg4399))));
                end
              else
                begin
                  reg4427 <= {(reg4409[(1'h0):(1'h0)] ?
                          reg4426[(3'h4):(2'h3)] : ((reg4393 || reg4347) ?
                              $unsigned((8'haf)) : $unsigned(reg4371)))};
                  reg4428 <= $unsigned($signed($signed(reg4377)));
                  if ((~|reg4433[(3'h6):(2'h3)]))
                    begin
                      reg4429 <= $unsigned($signed(forvar4427));
                      reg4430 <= $unsigned(((~$unsigned(forvar4347)) | (~$signed(reg4397))));
                      reg4431 <= reg4429[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4429 <= $signed(($unsigned(reg4365) ?
                          ((reg4429 ^~ (8'ha1)) ?
                              ((8'hb6) ?
                                  reg4431 : reg4353) : $unsigned(reg4350)) : $signed($unsigned(reg4357))));
                    end
                end
              for (forvar4436 = (1'h0); (forvar4436 < (1'h0)); forvar4436 = (forvar4436 + (1'h1)))
                begin
                  for (forvar4437 = (1'h0); (forvar4437 < (1'h1)); forvar4437 = (forvar4437 + (1'h1)))
                    begin
                      reg4438 <= $signed(forvar4437[(3'h5):(2'h3)]);
                      reg4439 <= reg4427;
                    end
                  for (forvar4440 = (1'h0); (forvar4440 < (1'h0)); forvar4440 = (forvar4440 + (1'h1)))
                    begin
                      reg4441 <= $signed(wire4339);
                      reg4442 <= ($signed($unsigned({forvar4424})) + {((!forvar4413) <= reg4417)});
                      reg4443 <= $unsigned((|{$unsigned(reg4359)}));
                    end
                  reg4444 <= reg4391[(4'h9):(3'h5)];
                  reg4445 <= ($unsigned(reg4410[(1'h0):(1'h0)]) <= wire4342[(3'h4):(2'h2)]);
                end
              if (forvar4368)
                begin
                  if (wire4338)
                    begin
                      reg4446 <= $unsigned($signed($unsigned((reg4439 && (8'ha3)))));
                      reg4447 <= reg4419;
                      reg4448 <= (8'ha1);
                    end
                  else
                    begin
                      reg4446 <= forvar4364;
                      reg4447 <= (reg4369[(1'h0):(1'h0)] ~^ ($unsigned($unsigned((8'ha8))) < (!(~(8'hb4)))));
                      reg4448 <= $signed($signed(($unsigned(reg4433) >> (&forvar4440))));
                    end
                  for (forvar4449 = (1'h0); (forvar4449 < (2'h2)); forvar4449 = (forvar4449 + (1'h1)))
                    begin
                      reg4450 <= forvar4427[(2'h2):(1'h0)];
                      reg4451 <= (forvar4359[(3'h4):(2'h2)] - reg4356[(4'he):(2'h2)]);
                      reg4452 <= $signed($unsigned($signed(reg4419)));
                      reg4453 <= $unsigned((~|((reg4432 <= (8'hb6)) > (8'ha1))));
                    end
                  for (forvar4454 = (1'h0); (forvar4454 < (1'h1)); forvar4454 = (forvar4454 + (1'h1)))
                    begin
                      reg4455 <= $signed($signed(($unsigned(reg4438) <= reg4356)));
                    end
                end
              else
                begin
                  if (reg4359[(1'h0):(1'h0)])
                    begin
                      reg4446 <= (reg4413[(2'h2):(1'h0)] <<< reg4410[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg4446 <= reg4423;
                    end
                  if ($unsigned((~$unsigned((-(8'hb2))))))
                    begin
                      reg4447 <= ((((^reg4432) ^~ forvar4408) > ((-reg4446) ?
                          reg4381 : reg4433)) + (wire4340 ^~ reg4425));
                      reg4448 <= reg4427;
                    end
                  else
                    begin
                      reg4447 <= ($signed($unsigned($signed(reg4439))) ?
                          forvar4344[(3'h4):(2'h2)] : $signed((reg4432[(3'h4):(2'h2)] > $unsigned(forvar4350))));
                      reg4448 <= (!reg4433[(1'h0):(1'h0)]);
                    end
                  for (forvar4449 = (1'h0); (forvar4449 < (2'h2)); forvar4449 = (forvar4449 + (1'h1)))
                    begin
                      reg4450 <= (^forvar4440);
                      reg4451 <= ($signed($unsigned((|wire4342))) != {$unsigned(reg4371)});
                      reg4452 <= (^~(|({(8'h9e)} - $signed(reg4345))));
                    end
                end
            end
          for (forvar4456 = (1'h0); (forvar4456 < (1'h0)); forvar4456 = (forvar4456 + (1'h1)))
            begin
              if ((~|{reg4375[(3'h6):(3'h4)]}))
                begin
                  for (forvar4457 = (1'h0); (forvar4457 < (2'h2)); forvar4457 = (forvar4457 + (1'h1)))
                    begin
                      reg4458 <= ($unsigned((-(!forvar4389))) ?
                          ((forvar4389 ?
                              reg4345 : $signed(forvar4391)) == ({(8'hb7)} <= (reg4358 != wire4339))) : reg4352);
                    end
                  for (forvar4459 = (1'h0); (forvar4459 < (2'h2)); forvar4459 = (forvar4459 + (1'h1)))
                    begin
                      reg4460 <= reg4387;
                    end
                end
              else
                begin
                  if (forvar4350[(3'h6):(3'h6)])
                    begin
                      reg4457 <= reg4417;
                      reg4458 <= {reg4360};
                      reg4459 <= ($unsigned(((forvar4427 >> forvar4356) ?
                              (8'haa) : reg4445)) ?
                          (8'h9f) : (reg4376 & reg4386[(4'h8):(4'h8)]));
                    end
                  else
                    begin
                      reg4457 <= (^$unsigned(reg4419));
                      reg4458 <= $signed(($unsigned((reg4444 ?
                              wire4338 : forvar4423)) ?
                          $unsigned(reg4446[(3'h6):(3'h4)]) : reg4385));
                      reg4459 <= $unsigned((~((forvar4353 ? (8'hae) : reg4434) ?
                          reg4361 : reg4416[(3'h4):(1'h1)])));
                      reg4460 <= reg4455[(1'h0):(1'h0)];
                    end
                end
              reg4461 <= (forvar4347 > reg4425[(2'h3):(1'h1)]);
              if ($unsigned(({{reg4352}} ?
                  {$signed((8'h9e))} : reg4370[(4'ha):(3'h6)])))
                begin
                  reg4462 <= forvar4374;
                  reg4463 <= (($signed((reg4356 ? reg4409 : reg4453)) ?
                          ((~forvar4423) <<< (reg4372 <<< (8'hab))) : (reg4375 ?
                              $unsigned(forvar4374) : $unsigned(reg4345))) ?
                      reg4399 : $unsigned(((reg4359 == wire4343) && $unsigned(reg4447))));
                  for (forvar4464 = (1'h0); (forvar4464 < (2'h2)); forvar4464 = (forvar4464 + (1'h1)))
                    begin
                      reg4465 <= $unsigned($unsigned(forvar4424));
                      reg4466 <= (&$signed((~^(!wire4340))));
                    end
                end
              else
                begin
                  if (reg4379)
                    begin
                      reg4462 <= ((^reg4407) ?
                          $signed($unsigned({forvar4369})) : forvar4368[(1'h1):(1'h0)]);
                      reg4463 <= reg4376[(4'h8):(3'h6)];
                    end
                  else
                    begin
                      reg4462 <= (reg4352[(3'h7):(3'h7)] ?
                          {reg4350} : $signed((^~reg4443)));
                    end
                end
              for (forvar4467 = (1'h0); (forvar4467 < (1'h1)); forvar4467 = (forvar4467 + (1'h1)))
                begin
                  if (((reg4423[(1'h1):(1'h1)] >>> (8'haf)) + {forvar4456}))
                    begin
                      reg4468 <= reg4453[(1'h0):(1'h0)];
                      reg4469 <= $signed({(^~(forvar4440 >>> reg4351))});
                      reg4470 <= reg4378[(4'h8):(3'h4)];
                    end
                  else
                    begin
                      reg4468 <= $unsigned($unsigned(($unsigned(reg4365) ?
                          ((8'hae) + reg4382) : $signed(reg4427))));
                      reg4469 <= (+(|reg4445));
                    end
                  if ((^~reg4369[(1'h0):(1'h0)]))
                    begin
                      reg4471 <= {(reg4442 != ((reg4413 ?
                                  reg4383 : forvar4456) ?
                              reg4410[(1'h0):(1'h0)] : (reg4416 ?
                                  reg4387 : reg4372)))};
                      reg4472 <= (|forvar4457[(4'h9):(3'h7)]);
                    end
                  else
                    begin
                      reg4471 <= (^~$unsigned(($signed(reg4391) & {(8'haf)})));
                      reg4472 <= (($signed(forvar4413) - reg4369) ^~ forvar4352);
                      reg4473 <= (reg4369 * {{(reg4372 && reg4417)}});
                      reg4474 <= (&reg4426);
                    end
                end
            end
        end
      if (($unsigned(((+reg4463) == reg4380[(3'h4):(3'h4)])) != ($signed((~&(8'hb2))) ?
          (~&(reg4390 >>> reg4404)) : reg4348[(1'h1):(1'h1)])))
        begin
          for (forvar4475 = (1'h0); (forvar4475 < (2'h2)); forvar4475 = (forvar4475 + (1'h1)))
            begin
              for (forvar4476 = (1'h0); (forvar4476 < (1'h1)); forvar4476 = (forvar4476 + (1'h1)))
                begin
                  if ($signed(($signed($unsigned(forvar4372)) << (|forvar4345))))
                    begin
                      reg4477 <= $unsigned((!$unsigned($unsigned(forvar4454))));
                      reg4478 <= ((!$signed(reg4418[(4'ha):(3'h5)])) ?
                          ($unsigned(((8'ha8) ? reg4426 : (8'ha1))) ?
                              (~forvar4440[(2'h3):(2'h2)]) : $signed((|(8'ha5)))) : reg4361);
                      reg4479 <= $signed(((^reg4370) >= ((~^forvar4422) ?
                          (^wire4339) : reg4433[(4'h8):(3'h7)])));
                      reg4480 <= ($unsigned($unsigned({reg4451})) ?
                          (reg4404[(2'h2):(1'h1)] ?
                              reg4375[(3'h7):(3'h6)] : reg4441[(4'he):(2'h3)]) : {forvar4374});
                    end
                  else
                    begin
                      reg4477 <= $unsigned(forvar4413[(2'h2):(2'h2)]);
                    end
                  reg4481 <= forvar4353;
                  for (forvar4482 = (1'h0); (forvar4482 < (1'h0)); forvar4482 = (forvar4482 + (1'h1)))
                    begin
                      reg4483 <= (reg4438[(2'h2):(1'h1)] ?
                          (($unsigned(forvar4424) <<< $signed(reg4443)) > $signed({(8'ha5)})) : (($signed(reg4479) ?
                                  reg4439[(3'h6):(1'h0)] : forvar4467) ?
                              reg4463[(2'h3):(1'h0)] : $unsigned(reg4441)));
                      reg4484 <= (forvar4352[(1'h1):(1'h0)] ?
                          reg4427[(1'h0):(1'h0)] : $signed((((8'haf) ?
                              reg4422 : reg4411) < $unsigned(forvar4346))));
                      reg4485 <= $unsigned($unsigned(reg4446));
                    end
                end
            end
          for (forvar4486 = (1'h0); (forvar4486 < (2'h2)); forvar4486 = (forvar4486 + (1'h1)))
            begin
              for (forvar4487 = (1'h0); (forvar4487 < (1'h0)); forvar4487 = (forvar4487 + (1'h1)))
                begin
                  reg4488 <= $signed($signed(((~^forvar4427) ?
                      $signed(forvar4427) : reg4386[(4'hf):(1'h0)])));
                end
              for (forvar4489 = (1'h0); (forvar4489 < (2'h3)); forvar4489 = (forvar4489 + (1'h1)))
                begin
                  if (forvar4422[(3'h7):(3'h6)])
                    begin
                      reg4490 <= (&(~|$unsigned($unsigned(reg4412))));
                      reg4491 <= (reg4359 ?
                          $signed(reg4466[(3'h7):(1'h1)]) : $unsigned((((8'hb6) & reg4427) ?
                              (-reg4478) : $signed(reg4435))));
                      reg4492 <= (|(reg4444 ? $unsigned((8'hb1)) : (8'hb4)));
                      reg4493 <= reg4386[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg4490 <= (!$signed((reg4352[(4'h9):(2'h2)] ~^ {reg4356})));
                      reg4491 <= $signed($unsigned($unsigned({reg4462})));
                    end
                  reg4494 <= forvar4344[(4'hc):(3'h7)];
                  if ({(reg4385[(3'h5):(1'h0)] ~^ $signed((forvar4412 ?
                          forvar4353 : wire4339)))})
                    begin
                      reg4495 <= reg4463;
                    end
                  else
                    begin
                      reg4495 <= $unsigned($signed((((8'hb5) ?
                              wire4340 : (8'had)) ?
                          wire4342[(3'h5):(1'h1)] : (^~(8'hb9)))));
                    end
                  for (forvar4496 = (1'h0); (forvar4496 < (2'h3)); forvar4496 = (forvar4496 + (1'h1)))
                    begin
                      reg4497 <= reg4425;
                      reg4498 <= ((reg4424[(2'h3):(2'h3)] ?
                              (8'hb8) : $unsigned((reg4360 + reg4443))) ?
                          $unsigned(forvar4350[(3'h7):(3'h4)]) : {((~^(8'hb5)) >= reg4369)});
                    end
                end
              reg4499 <= ((^$signed((reg4462 == reg4405))) ?
                  (!$unsigned((-reg4457))) : reg4419);
              if (forvar4440)
                begin
                  for (forvar4500 = (1'h0); (forvar4500 < (1'h1)); forvar4500 = (forvar4500 + (1'h1)))
                    begin
                      reg4501 <= {(reg4431 ?
                              ($unsigned((8'ha4)) == {forvar4350}) : $signed((~reg4423)))};
                      reg4502 <= $signed($signed({$unsigned(forvar4449)}));
                    end
                  if (((~$unsigned($unsigned((8'haa)))) - ({reg4455[(2'h2):(1'h0)]} ?
                      reg4395[(2'h2):(2'h2)] : {{reg4388}})))
                    begin
                      reg4503 <= {{({forvar4475} ~^ $signed(reg4502))}};
                      reg4504 <= {$signed(reg4411[(4'h8):(3'h6)])};
                      reg4505 <= $signed($signed((((8'ha0) ?
                              (8'h9e) : reg4390) ?
                          forvar4422[(2'h3):(1'h0)] : $unsigned(forvar4391))));
                    end
                  else
                    begin
                      reg4503 <= (((reg4413 || $unsigned(reg4370)) << reg4407[(3'h6):(3'h6)]) == $signed(reg4409[(2'h2):(1'h0)]));
                    end
                  reg4506 <= reg4499[(3'h4):(1'h1)];
                end
              else
                begin
                  reg4500 <= (($signed((~&reg4380)) ?
                      (8'h9c) : forvar4375[(1'h0):(1'h0)]) & forvar4359[(1'h0):(1'h0)]);
                  for (forvar4501 = (1'h0); (forvar4501 < (1'h1)); forvar4501 = (forvar4501 + (1'h1)))
                    begin
                      reg4502 <= $unsigned(((^~(reg4377 ? reg4473 : (8'hae))) ?
                          forvar4427[(3'h5):(3'h5)] : (+(reg4396 <<< reg4439))));
                      reg4503 <= $signed((~^((-forvar4353) | reg4405[(4'hb):(3'h5)])));
                    end
                  for (forvar4504 = (1'h0); (forvar4504 < (2'h2)); forvar4504 = (forvar4504 + (1'h1)))
                    begin
                      reg4505 <= (!reg4447[(3'h4):(1'h0)]);
                      reg4506 <= $signed($signed(reg4365[(3'h4):(2'h2)]));
                      reg4507 <= {(forvar4504 | (reg4412 <= reg4384))};
                    end
                end
            end
        end
      else
        begin
          for (forvar4475 = (1'h0); (forvar4475 < (2'h3)); forvar4475 = (forvar4475 + (1'h1)))
            begin
              for (forvar4476 = (1'h0); (forvar4476 < (2'h3)); forvar4476 = (forvar4476 + (1'h1)))
                begin
                  if ($unsigned(($signed($signed((8'ha0))) ?
                      (reg4362 ?
                          (forvar4386 ?
                              reg4393 : (8'hb2)) : reg4425) : {forvar4500[(3'h7):(2'h2)]})))
                    begin
                      reg4477 <= reg4388;
                      reg4478 <= (~reg4446);
                      reg4479 <= ({reg4465[(1'h0):(1'h0)]} >>> $unsigned((!(reg4396 ?
                          (8'haf) : reg4358))));
                      reg4480 <= (&($unsigned((!forvar4456)) << ($signed(forvar4368) ?
                          (8'hb0) : reg4379[(2'h3):(1'h1)])));
                    end
                  else
                    begin
                      reg4477 <= (+(^{$signed(reg4395)}));
                    end
                  if (($unsigned(reg4376[(3'h5):(2'h3)]) & $unsigned((&forvar4389[(1'h0):(1'h0)]))))
                    begin
                      reg4481 <= $signed($signed({{(8'hac)}}));
                      reg4482 <= ($signed((~|$signed(forvar4487))) >> forvar4464[(3'h4):(1'h1)]);
                      reg4483 <= ((~^$signed($unsigned((8'hba)))) >>> reg4498);
                    end
                  else
                    begin
                      reg4481 <= $unsigned((reg4481[(4'hd):(4'hb)] ?
                          reg4381 : reg4428[(3'h4):(2'h3)]));
                      reg4482 <= ($unsigned($signed(reg4366[(2'h2):(1'h1)])) ?
                          reg4444 : (forvar4413[(1'h0):(1'h0)] && (-(reg4348 < (8'ha7)))));
                      reg4483 <= $signed(($unsigned(((8'h9f) ~^ reg4493)) ?
                          reg4390 : reg4459[(2'h3):(1'h1)]));
                      reg4484 <= {(~&$unsigned((^~reg4506)))};
                    end
                  for (forvar4485 = (1'h0); (forvar4485 < (1'h0)); forvar4485 = (forvar4485 + (1'h1)))
                    begin
                      reg4486 <= forvar4414[(1'h1):(1'h0)];
                      reg4487 <= $signed((~|$unsigned((reg4348 ?
                          (8'haa) : reg4424))));
                      reg4488 <= {$signed(forvar4413)};
                      reg4489 <= reg4432[(2'h3):(1'h1)];
                    end
                end
              if (forvar4436)
                begin
                  for (forvar4490 = (1'h0); (forvar4490 < (1'h1)); forvar4490 = (forvar4490 + (1'h1)))
                    begin
                      reg4491 <= ($signed($signed($signed(reg4488))) | reg4350);
                    end
                  reg4492 <= $signed({{$signed(reg4486)}});
                end
              else
                begin
                  if (reg4503)
                    begin
                      reg4490 <= reg4433[(4'h8):(3'h7)];
                      reg4491 <= reg4489;
                    end
                  else
                    begin
                      reg4490 <= ((forvar4482[(3'h7):(3'h4)] & forvar4489) != $unsigned(reg4497));
                      reg4491 <= $signed(((reg4485[(1'h0):(1'h0)] ?
                              $signed(wire4338) : {reg4377}) ?
                          ((-reg4375) == reg4348) : reg4377[(4'h9):(1'h1)]));
                      reg4492 <= {reg4451[(3'h4):(2'h3)]};
                      reg4493 <= $unsigned($unsigned((forvar4501[(4'hb):(3'h5)] < (reg4490 >> reg4451))));
                    end
                  if ($signed($signed($unsigned((~|forvar4389)))))
                    begin
                      reg4494 <= ((|$unsigned(((8'hae) - reg4448))) ?
                          (+(forvar4403[(3'h4):(1'h0)] ?
                              $signed(reg4470) : reg4383[(1'h1):(1'h0)])) : reg4431);
                      reg4495 <= {reg4442};
                      reg4496 <= $unsigned((8'ha3));
                    end
                  else
                    begin
                      reg4494 <= $signed(forvar4364[(4'ha):(3'h5)]);
                      reg4495 <= (~|{(8'hb6)});
                      reg4496 <= reg4461;
                    end
                  if ((~|$signed((~|$unsigned(reg4379)))))
                    begin
                      reg4497 <= {(reg4429 <= (!((8'ha3) ?
                              reg4415 : reg4385)))};
                      reg4498 <= {$unsigned($signed(reg4442))};
                      reg4499 <= reg4430[(4'h8):(4'h8)];
                      reg4500 <= (wire4341[(4'hb):(3'h5)] ?
                          {(reg4377 ?
                                  (forvar4423 == (8'hb6)) : ((8'hb2) ^~ reg4406))} : forvar4437[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg4497 <= ((reg4457[(3'h4):(1'h0)] ?
                              $signed((reg4407 ^~ reg4377)) : $signed((~^(8'hae)))) ?
                          $signed($signed($signed(reg4494))) : ($unsigned(reg4485) > (8'ha2)));
                      reg4498 <= ((((forvar4423 <<< reg4472) ?
                          (|reg4452) : {reg4407}) << reg4469[(2'h2):(1'h0)]) <= {$unsigned(forvar4500[(2'h3):(2'h2)])});
                    end
                  if ($signed($signed($unsigned(forvar4449))))
                    begin
                      reg4501 <= $unsigned(reg4420);
                      reg4502 <= reg4447[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg4501 <= (8'hb0);
                    end
                end
              if ((reg4462[(2'h3):(1'h1)] > forvar4490))
                begin
                  for (forvar4503 = (1'h0); (forvar4503 < (1'h1)); forvar4503 = (forvar4503 + (1'h1)))
                    begin
                      reg4504 <= ($unsigned({reg4400}) >> (-{(-reg4386)}));
                      reg4505 <= $signed(reg4441[(5'h10):(2'h2)]);
                    end
                  if ((^~(($unsigned((8'hb6)) ? (^(8'hba)) : reg4452) ?
                      ((+reg4394) * (reg4350 ?
                          reg4402 : reg4383)) : (^~reg4496))))
                    begin
                      reg4506 <= (($unsigned((~&forvar4350)) ?
                          ({reg4473} >>> $signed(forvar4408)) : ((reg4371 ?
                                  reg4443 : reg4466) ?
                              $unsigned(reg4376) : {(8'hb5)})) << ($signed({forvar4346}) > ($unsigned(reg4410) ?
                          $unsigned(forvar4345) : forvar4386)));
                      reg4507 <= {(~|$signed($unsigned((8'hb7))))};
                      reg4508 <= reg4370[(4'hb):(3'h7)];
                      reg4509 <= $signed($signed(($signed(forvar4449) & reg4458)));
                    end
                  else
                    begin
                      reg4506 <= $signed($signed((+(reg4349 || forvar4467))));
                      reg4507 <= (~&(8'hb1));
                      reg4508 <= $unsigned($signed(($signed(reg4473) ?
                          reg4450[(1'h1):(1'h1)] : (8'ha2))));
                    end
                  for (forvar4510 = (1'h0); (forvar4510 < (2'h2)); forvar4510 = (forvar4510 + (1'h1)))
                    begin
                      reg4511 <= $unsigned((^~$signed(forvar4457[(3'h5):(2'h2)])));
                      reg4512 <= $unsigned(reg4409[(3'h4):(1'h0)]);
                    end
                  if ((reg4438[(2'h2):(1'h1)] ?
                      reg4459[(1'h0):(1'h0)] : $unsigned((reg4460[(2'h3):(1'h1)] | reg4402[(2'h3):(2'h2)]))))
                    begin
                      reg4513 <= $signed(forvar4500);
                      reg4514 <= reg4366;
                      reg4515 <= (reg4493[(4'h9):(1'h1)] * reg4503[(3'h7):(3'h5)]);
                      reg4516 <= (reg4350[(1'h1):(1'h0)] - $unsigned(reg4481[(2'h3):(1'h1)]));
                    end
                  else
                    begin
                      reg4513 <= $unsigned($unsigned($signed((reg4345 ?
                          reg4481 : (8'had)))));
                    end
                end
              else
                begin
                  for (forvar4503 = (1'h0); (forvar4503 < (2'h2)); forvar4503 = (forvar4503 + (1'h1)))
                    begin
                      reg4504 <= (~&(((reg4473 ?
                              reg4439 : forvar4347) << (8'hab)) ?
                          (reg4512 ?
                              (^~reg4470) : reg4381[(2'h3):(1'h0)]) : (8'ha3)));
                      reg4505 <= reg4395;
                    end
                  for (forvar4506 = (1'h0); (forvar4506 < (1'h1)); forvar4506 = (forvar4506 + (1'h1)))
                    begin
                      reg4507 <= (8'ha9);
                      reg4508 <= $signed(forvar4350[(1'h1):(1'h0)]);
                    end
                  for (forvar4509 = (1'h0); (forvar4509 < (1'h0)); forvar4509 = (forvar4509 + (1'h1)))
                    begin
                      reg4510 <= forvar4391;
                    end
                end
              reg4517 <= {$signed($unsigned($signed(reg4400)))};
            end
        end
      for (forvar4518 = (1'h0); (forvar4518 < (2'h2)); forvar4518 = (forvar4518 + (1'h1)))
        begin
          reg4519 <= {(!$signed(forvar4359))};
          if ({(({forvar4437} ? $signed(reg4393) : $unsigned(reg4463)) ?
                  (-$signed(reg4378)) : ((^reg4357) ^~ (^forvar4486)))})
            begin
              for (forvar4520 = (1'h0); (forvar4520 < (1'h0)); forvar4520 = (forvar4520 + (1'h1)))
                begin
                  reg4521 <= ($signed(({(8'hb5)} ^ (reg4357 <= reg4400))) | (reg4496[(2'h2):(1'h0)] != (~|{(8'hb7)})));
                end
              reg4522 <= {reg4406};
            end
          else
            begin
              if (reg4428)
                begin
                  for (forvar4520 = (1'h0); (forvar4520 < (1'h1)); forvar4520 = (forvar4520 + (1'h1)))
                    begin
                      reg4521 <= reg4371;
                      reg4522 <= (&reg4498);
                      reg4523 <= ($signed($signed($unsigned(wire4342))) == $signed(((reg4365 - forvar4386) ?
                          reg4347 : (reg4419 ? reg4480 : reg4479))));
                    end
                  if ($signed((~^(!((8'h9f) > reg4448)))))
                    begin
                      reg4524 <= (^~(-$unsigned($signed(reg4508))));
                      reg4525 <= reg4469;
                      reg4526 <= ((8'hb0) != ((~^$signed((8'h9e))) ?
                          $unsigned(reg4525) : ((reg4470 ?
                              reg4361 : reg4513) <= $unsigned(reg4447))));
                    end
                  else
                    begin
                      reg4524 <= (|{reg4392});
                      reg4525 <= ((~(-{reg4503})) <= reg4369[(2'h2):(1'h0)]);
                      reg4526 <= (|$unsigned(forvar4372[(1'h0):(1'h0)]));
                    end
                  for (forvar4527 = (1'h0); (forvar4527 < (2'h3)); forvar4527 = (forvar4527 + (1'h1)))
                    begin
                      reg4528 <= reg4498;
                      reg4529 <= {{$unsigned(reg4474[(3'h4):(3'h4)])}};
                    end
                  for (forvar4530 = (1'h0); (forvar4530 < (2'h2)); forvar4530 = (forvar4530 + (1'h1)))
                    begin
                      reg4531 <= $unsigned((reg4515 ?
                          forvar4530 : (reg4462[(3'h7):(2'h2)] >= {(8'ha5)})));
                      reg4532 <= reg4499;
                      reg4533 <= {reg4432};
                      reg4534 <= {$signed(forvar4414[(1'h0):(1'h0)])};
                    end
                end
              else
                begin
                  reg4520 <= (~{$unsigned((^~reg4379))});
                  reg4521 <= reg4384;
                  for (forvar4522 = (1'h0); (forvar4522 < (1'h1)); forvar4522 = (forvar4522 + (1'h1)))
                    begin
                      reg4523 <= {reg4451[(4'ha):(3'h5)]};
                      reg4524 <= reg4350[(1'h0):(1'h0)];
                      reg4525 <= (8'ha3);
                    end
                  reg4526 <= reg4388;
                end
              if ($unsigned((&((reg4520 | reg4490) >= forvar4401[(2'h2):(1'h0)]))))
                begin
                  for (forvar4535 = (1'h0); (forvar4535 < (2'h2)); forvar4535 = (forvar4535 + (1'h1)))
                    begin
                      reg4536 <= reg4459[(3'h6):(2'h2)];
                      reg4537 <= $signed(((reg4532 * reg4442) & ({forvar4436} || $unsigned((8'hb1)))));
                    end
                  for (forvar4538 = (1'h0); (forvar4538 < (2'h2)); forvar4538 = (forvar4538 + (1'h1)))
                    begin
                      reg4539 <= $signed(($signed((&reg4517)) * wire4341));
                      reg4540 <= (^~$signed((+reg4362)));
                      reg4541 <= $signed((forvar4476 >>> $unsigned(reg4406)));
                      reg4542 <= (^~{$unsigned(wire4339)});
                    end
                end
              else
                begin
                  for (forvar4535 = (1'h0); (forvar4535 < (2'h2)); forvar4535 = (forvar4535 + (1'h1)))
                    begin
                      reg4536 <= forvar4414[(1'h0):(1'h0)];
                    end
                  for (forvar4537 = (1'h0); (forvar4537 < (2'h3)); forvar4537 = (forvar4537 + (1'h1)))
                    begin
                      reg4538 <= forvar4375;
                      reg4539 <= $unsigned($unsigned((reg4502[(2'h2):(1'h0)] ?
                          (&(8'hb6)) : (|reg4386))));
                      reg4540 <= {reg4382[(1'h1):(1'h0)]};
                      reg4541 <= ((-(|(!reg4494))) ?
                          (~$unsigned(((8'hb3) <= forvar4506))) : $unsigned((+reg4379[(2'h3):(2'h3)])));
                    end
                  for (forvar4542 = (1'h0); (forvar4542 < (1'h1)); forvar4542 = (forvar4542 + (1'h1)))
                    begin
                      reg4543 <= forvar4487;
                      reg4544 <= reg4420;
                    end
                  reg4545 <= reg4515;
                end
              for (forvar4546 = (1'h0); (forvar4546 < (2'h2)); forvar4546 = (forvar4546 + (1'h1)))
                begin
                  for (forvar4547 = (1'h0); (forvar4547 < (2'h3)); forvar4547 = (forvar4547 + (1'h1)))
                    begin
                      reg4548 <= ((8'hae) + (8'hac));
                      reg4549 <= reg4373[(4'h8):(2'h3)];
                      reg4550 <= (~|((8'hae) & ({reg4413} * $unsigned(forvar4422))));
                      reg4551 <= ({$unsigned($unsigned(forvar4412))} & (~^(8'hb3)));
                    end
                  reg4552 <= (~&($unsigned(((8'ha1) ?
                      (8'h9e) : reg4434)) < ((+reg4524) ?
                      forvar4482[(4'hb):(3'h4)] : reg4470)));
                end
            end
          for (forvar4553 = (1'h0); (forvar4553 < (2'h2)); forvar4553 = (forvar4553 + (1'h1)))
            begin
              for (forvar4554 = (1'h0); (forvar4554 < (1'h0)); forvar4554 = (forvar4554 + (1'h1)))
                begin
                  reg4555 <= (^(|(wire4338[(3'h4):(2'h2)] ?
                      ((8'hb5) ^ reg4381) : (+forvar4401))));
                  for (forvar4556 = (1'h0); (forvar4556 < (2'h2)); forvar4556 = (forvar4556 + (1'h1)))
                    begin
                      reg4557 <= (forvar4427 * $unsigned(reg4480));
                    end
                end
              for (forvar4558 = (1'h0); (forvar4558 < (1'h0)); forvar4558 = (forvar4558 + (1'h1)))
                begin
                  if ((!$signed($signed((reg4505 ? forvar4530 : forvar4459)))))
                    begin
                      reg4559 <= (~&$unsigned(((~reg4412) << (reg4489 & reg4360))));
                      reg4560 <= reg4349[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg4559 <= (^~{($signed(wire4341) <= reg4461)});
                      reg4560 <= ((reg4497[(2'h2):(2'h2)] && $unsigned({(8'hac)})) * ((8'had) ?
                          ({wire4339} ?
                              (reg4365 ? reg4534 : (8'ha2)) : (reg4461 ?
                                  reg4416 : reg4482)) : $signed($unsigned(reg4517))));
                    end
                  for (forvar4561 = (1'h0); (forvar4561 < (2'h3)); forvar4561 = (forvar4561 + (1'h1)))
                    begin
                      reg4562 <= $unsigned({(-(reg4373 ? reg4496 : reg4509))});
                      reg4563 <= (($signed($unsigned((8'hab))) >>> forvar4372[(3'h4):(2'h2)]) ?
                          (reg4425[(1'h1):(1'h0)] ?
                              forvar4344[(4'h9):(1'h1)] : (8'ha1)) : (^~(8'ha6)));
                      reg4564 <= reg4537;
                    end
                  if ({($signed($signed(reg4488)) ^~ {{forvar4347}})})
                    begin
                      reg4565 <= (&(~$unsigned((8'hb9))));
                      reg4566 <= ($unsigned(($unsigned((8'ha3)) - (forvar4437 ?
                              forvar4364 : reg4540))) ?
                          (+$unsigned($signed(reg4458))) : (-$signed({forvar4500})));
                    end
                  else
                    begin
                      reg4565 <= (!forvar4347);
                      reg4566 <= $signed(forvar4535);
                    end
                end
              for (forvar4567 = (1'h0); (forvar4567 < (2'h3)); forvar4567 = (forvar4567 + (1'h1)))
                begin
                  for (forvar4568 = (1'h0); (forvar4568 < (2'h3)); forvar4568 = (forvar4568 + (1'h1)))
                    begin
                      reg4569 <= (reg4487[(4'hc):(4'h9)] <= $signed((forvar4359 | forvar4518[(2'h2):(2'h2)])));
                    end
                end
              reg4570 <= {(forvar4476[(1'h0):(1'h0)] && forvar4486[(3'h6):(1'h0)])};
            end
        end
    end
  assign wire4571 = (~|(|{reg4525[(1'h0):(1'h0)]}));
  module4572 modinst7007 (.wire4573(reg4378), .y(wire7006), .wire4575(reg4409), .clk(clk), .wire4576(reg4459), .wire4574(reg4379));
  assign wire7008 = forvar4374;
  assign wire7009 = $unsigned($unsigned($unsigned(forvar4506[(3'h5):(1'h1)])));
  always
    @(posedge clk) begin
      for (forvar7010 = (1'h0); (forvar7010 < (2'h2)); forvar7010 = (forvar7010 + (1'h1)))
        begin
          for (forvar7011 = (1'h0); (forvar7011 < (1'h0)); forvar7011 = (forvar7011 + (1'h1)))
            begin
              for (forvar7012 = (1'h0); (forvar7012 < (2'h3)); forvar7012 = (forvar7012 + (1'h1)))
                begin
                  if ({reg4380})
                    begin
                      reg7013 <= ((+(forvar4423 ~^ (reg4479 >> reg4382))) >= $unsigned($signed({reg4529})));
                      reg7014 <= $signed($unsigned((8'hb3)));
                    end
                  else
                    begin
                      reg7013 <= $signed({$signed((reg4525 ?
                              reg4514 : reg4545))});
                      reg7014 <= (forvar4464[(2'h2):(1'h1)] ?
                          (reg4455 ?
                              forvar4391 : ({reg4366} >>> {reg4444})) : ($signed((reg4365 ?
                              reg4489 : reg4363)) <= reg4423[(1'h1):(1'h1)]));
                      reg7015 <= $signed($signed($signed((~^reg4514))));
                    end
                  if (reg4516)
                    begin
                      reg7016 <= {{((~reg4541) ?
                                  {(8'hb9)} : reg4387[(4'hf):(4'he)])}};
                      reg7017 <= reg4483;
                      reg7018 <= $unsigned((^~(((8'hb4) >= reg4417) ?
                          {reg4353} : (reg4376 ^~ reg4545))));
                    end
                  else
                    begin
                      reg7016 <= ($signed($unsigned({wire4571})) | ({(~^reg4426)} ^ (reg4485[(4'h9):(3'h6)] <<< (reg4383 ?
                          reg4413 : reg4492))));
                      reg7017 <= ($unsigned({$signed(reg4544)}) ?
                          reg4570 : (($signed(forvar4518) ?
                              (reg4523 < forvar4464) : forvar4364) >= ($signed(wire7009) ?
                              (8'hb5) : $unsigned(reg7016))));
                      reg7018 <= (reg4367[(1'h0):(1'h0)] ?
                          reg4395[(1'h1):(1'h0)] : reg4399[(4'ha):(3'h6)]);
                    end
                  if (reg4386[(2'h2):(2'h2)])
                    begin
                      reg7019 <= $signed(forvar4352[(2'h2):(2'h2)]);
                      reg7020 <= (~|(forvar4347 & wire4340));
                    end
                  else
                    begin
                      reg7019 <= reg4512;
                      reg7020 <= $signed((reg4548[(2'h3):(1'h0)] >> reg4407[(3'h5):(3'h5)]));
                      reg7021 <= (-$signed((^(forvar4364 ?
                          forvar4489 : (8'ha4)))));
                      reg7022 <= (8'hb6);
                    end
                end
            end
        end
      for (forvar7023 = (1'h0); (forvar7023 < (2'h2)); forvar7023 = (forvar7023 + (1'h1)))
        begin
          if ({$signed((reg4448 ? $signed(reg4400) : $unsigned(reg4386)))})
            begin
              reg7024 <= $unsigned(wire4341[(3'h5):(2'h2)]);
              if ($unsigned($signed($unsigned(reg4383))))
                begin
                  if (reg4483[(1'h0):(1'h0)])
                    begin
                      reg7025 <= reg4525[(2'h2):(1'h1)];
                      reg7026 <= (8'hb3);
                      reg7027 <= reg7014[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg7025 <= (~|$unsigned($unsigned((~&forvar7023))));
                      reg7026 <= (reg4504[(3'h5):(2'h3)] ?
                          ((reg4370 ~^ $unsigned(reg4517)) ?
                              $signed($unsigned(reg4504)) : forvar4413) : ({(forvar4422 & reg4418)} < reg4426[(3'h4):(3'h4)]));
                      reg7027 <= forvar4422;
                      reg7028 <= $signed(($unsigned((reg4359 ?
                              forvar4482 : reg4474)) ?
                          $signed(forvar7011[(3'h5):(3'h4)]) : $signed($unsigned(forvar4490))));
                    end
                  reg7029 <= ($unsigned(reg4504[(3'h7):(3'h6)]) ~^ reg4462);
                  for (forvar7030 = (1'h0); (forvar7030 < (2'h3)); forvar7030 = (forvar7030 + (1'h1)))
                    begin
                      reg7031 <= $unsigned($unsigned($signed($unsigned(forvar4547))));
                      reg7032 <= reg4351[(1'h1):(1'h0)];
                      reg7033 <= (($signed((8'ha8)) ?
                              reg4354[(4'ha):(3'h7)] : ((forvar4485 ?
                                  reg4443 : forvar4418) >= reg7029)) ?
                          (8'hb0) : ({(-reg4536)} ^~ ((reg4425 || reg4367) ?
                              $signed(reg4500) : (reg4502 ?
                                  forvar4344 : (8'hb9)))));
                    end
                  if ((&{(8'ha7)}))
                    begin
                      reg7034 <= reg4416[(1'h0):(1'h0)];
                      reg7035 <= $signed($signed(($signed(reg7024) ^~ reg4367)));
                      reg7036 <= forvar7030;
                    end
                  else
                    begin
                      reg7034 <= ((8'hae) >>> (~reg4414[(2'h2):(2'h2)]));
                      reg7035 <= $signed((reg4529 - $unsigned({reg4359})));
                    end
                end
              else
                begin
                  if ({$signed($unsigned(reg4405))})
                    begin
                      reg7025 <= $signed(($unsigned((^~(8'haf))) ?
                          forvar4486[(3'h6):(2'h2)] : {wire4340[(4'ha):(3'h7)]}));
                      reg7026 <= reg4562[(4'h9):(2'h3)];
                    end
                  else
                    begin
                      reg7025 <= reg4441[(3'h4):(2'h3)];
                      reg7026 <= (($unsigned($unsigned(reg4526)) ?
                          wire7009 : forvar4487) <= (8'ha0));
                      reg7027 <= reg4514;
                    end
                  if (((((forvar4500 == (8'hb0)) ?
                          (reg4501 ~^ (8'ha2)) : (~forvar4356)) <<< $unsigned($signed(reg4461))) ?
                      forvar4567[(4'h8):(2'h2)] : forvar4537))
                    begin
                      reg7028 <= $signed((^($unsigned(forvar4369) ?
                          reg4565 : (8'ha3))));
                      reg7029 <= ($unsigned(forvar4506[(1'h0):(1'h0)]) ?
                          reg4345 : (reg7016[(4'h8):(3'h5)] ?
                              ((reg4384 + reg4495) ?
                                  reg4382[(1'h0):(1'h0)] : $unsigned(forvar4464)) : (^~reg4365[(3'h7):(3'h7)])));
                      reg7030 <= $unsigned(reg7035[(4'h9):(1'h0)]);
                      reg7031 <= ((^~{(^(8'hb7))}) < (reg4521 ?
                          $unsigned((^reg4388)) : $unsigned($unsigned(forvar4364))));
                    end
                  else
                    begin
                      reg7028 <= (forvar4464[(2'h2):(1'h1)] ?
                          reg4514 : reg4404[(2'h3):(2'h2)]);
                      reg7029 <= ((((reg4498 ?
                              forvar4386 : reg4563) * (~reg4387)) ?
                          (forvar4561[(3'h5):(2'h2)] & (reg4441 ?
                              reg4381 : forvar4368)) : wire4571[(3'h4):(2'h2)]) != $unsigned(forvar4344));
                    end
                  reg7032 <= $signed((|(!(reg4482 | reg4529))));
                  for (forvar7033 = (1'h0); (forvar7033 < (2'h2)); forvar7033 = (forvar7033 + (1'h1)))
                    begin
                      reg7034 <= (^(((wire7006 - reg7016) ?
                              (~&(8'h9c)) : $unsigned(forvar4456)) ?
                          {$signed(reg4361)} : $unsigned(reg4380)));
                    end
                end
              if ($unsigned($unsigned(reg4398)))
                begin
                  for (forvar7037 = (1'h0); (forvar7037 < (2'h2)); forvar7037 = (forvar7037 + (1'h1)))
                    begin
                      reg7038 <= (((^~(reg4439 ?
                              reg4501 : reg4450)) & $signed(forvar4424[(2'h3):(1'h0)])) ?
                          reg4537[(3'h4):(1'h0)] : ($unsigned((reg4505 > forvar4389)) ?
                              $unsigned($signed((8'hb7))) : reg4357));
                    end
                  if ((($unsigned((reg4363 * (8'ha7))) ?
                          reg7029[(1'h0):(1'h0)] : ((forvar4459 ?
                              (8'hac) : reg4498) <<< reg7029)) ?
                      (({reg7024} ^ ((8'hae) ? reg4396 : reg4551)) ?
                          ($signed(reg4371) && $unsigned(reg4426)) : (reg4438 ~^ $signed(reg4393))) : $signed(wire4338[(2'h2):(1'h1)])))
                    begin
                      reg7039 <= $signed(reg4384[(2'h3):(1'h1)]);
                      reg7040 <= $signed(forvar7023);
                      reg7041 <= (reg4532[(1'h1):(1'h1)] == reg4395[(2'h2):(2'h2)]);
                      reg7042 <= reg4509[(4'ha):(2'h3)];
                    end
                  else
                    begin
                      reg7039 <= (reg4541 << $unsigned((reg4349 ?
                          {forvar4352} : reg4533)));
                      reg7040 <= $unsigned((~^(forvar4556 < {forvar4386})));
                      reg7041 <= ($signed($unsigned((^~reg4404))) ?
                          ((~|{forvar4556}) == $unsigned((reg4397 > reg4549))) : ({(+reg4492)} ?
                              (8'hab) : $unsigned($signed(forvar4449))));
                      reg7042 <= {(~^{(reg4529 ? forvar4389 : reg4513)})};
                    end
                  if (forvar4558[(3'h6):(2'h3)])
                    begin
                      reg7043 <= $signed(reg4457);
                      reg7044 <= {$signed(($signed(reg4392) ?
                              (reg4566 ?
                                  forvar4553 : reg4492) : $unsigned(forvar7033)))};
                      reg7045 <= (-$signed((^~forvar4530[(2'h2):(2'h2)])));
                      reg7046 <= reg4512;
                    end
                  else
                    begin
                      reg7043 <= (8'ha3);
                    end
                end
              else
                begin
                  for (forvar7037 = (1'h0); (forvar7037 < (2'h3)); forvar7037 = (forvar7037 + (1'h1)))
                    begin
                      reg7038 <= {$unsigned(((forvar4487 ?
                                  forvar4527 : reg4444) ?
                              (~&(8'ha2)) : $signed(reg4523)))};
                      reg7039 <= $unsigned({{(8'hb9)}});
                    end
                  for (forvar7040 = (1'h0); (forvar7040 < (2'h2)); forvar7040 = (forvar7040 + (1'h1)))
                    begin
                      reg7041 <= (^reg7036[(4'he):(4'he)]);
                      reg7042 <= ($signed(((8'ha1) ?
                          (reg7019 ?
                              reg7045 : reg4543) : reg4542)) <= {reg7046[(2'h3):(2'h2)]});
                      reg7043 <= reg4540[(4'h8):(1'h1)];
                    end
                  for (forvar7044 = (1'h0); (forvar7044 < (2'h2)); forvar7044 = (forvar7044 + (1'h1)))
                    begin
                      reg7045 <= reg7035;
                    end
                end
            end
          else
            begin
              reg7024 <= $signed(($unsigned((reg7044 >>> reg4433)) ?
                  $unsigned((^~reg4538)) : $unsigned(reg4414)));
            end
          for (forvar7047 = (1'h0); (forvar7047 < (2'h3)); forvar7047 = (forvar7047 + (1'h1)))
            begin
              for (forvar7048 = (1'h0); (forvar7048 < (2'h2)); forvar7048 = (forvar7048 + (1'h1)))
                begin
                  for (forvar7049 = (1'h0); (forvar7049 < (2'h2)); forvar7049 = (forvar7049 + (1'h1)))
                    begin
                      reg7050 <= (({(~reg4353)} - forvar4440[(1'h0):(1'h0)]) < (~^((|reg4407) != (~&(8'h9c)))));
                      reg7051 <= (reg7027[(3'h5):(3'h4)] ?
                          (!$signed(reg7014[(2'h2):(2'h2)])) : $unsigned(((8'hb8) ^~ reg4534)));
                      reg7052 <= {(+$signed(reg4490[(1'h1):(1'h1)]))};
                    end
                  if (({(8'hb7)} ?
                      ((forvar7030[(1'h1):(1'h1)] | forvar4547[(2'h2):(1'h0)]) ~^ $signed(reg7018[(3'h5):(3'h4)])) : ($signed(reg4543[(1'h1):(1'h1)]) - (reg4425[(2'h2):(2'h2)] ?
                          (^reg7044) : $unsigned(forvar4386)))))
                    begin
                      reg7053 <= (!$signed(wire4343[(4'h9):(3'h5)]));
                    end
                  else
                    begin
                      reg7053 <= {reg4486[(2'h2):(1'h0)]};
                    end
                end
              for (forvar7054 = (1'h0); (forvar7054 < (2'h3)); forvar7054 = (forvar7054 + (1'h1)))
                begin
                  if ($unsigned($unsigned({forvar7011[(4'h8):(3'h4)]})))
                    begin
                      reg7055 <= $unsigned(reg4541[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg7055 <= (~$unsigned({$signed(reg4500)}));
                      reg7056 <= reg4420[(3'h7):(1'h0)];
                      reg7057 <= (8'h9f);
                      reg7058 <= $signed(reg4517);
                    end
                  if (forvar7010)
                    begin
                      reg7059 <= (&(({reg4465} && $unsigned(wire7009)) ?
                          (forvar7047 ^~ (^~reg4372)) : $unsigned($signed(reg4423))));
                    end
                  else
                    begin
                      reg7059 <= (!$signed({(+forvar4500)}));
                      reg7060 <= ($unsigned((~^(^~forvar4454))) || (reg4569 < ((reg4459 ?
                          wire4571 : forvar4464) && reg4382[(2'h2):(1'h0)])));
                      reg7061 <= $unsigned(forvar4542);
                      reg7062 <= (~^reg4366);
                    end
                  for (forvar7063 = (1'h0); (forvar7063 < (2'h3)); forvar7063 = (forvar7063 + (1'h1)))
                    begin
                      reg7064 <= (~^forvar4437[(1'h1):(1'h1)]);
                      reg7065 <= $unsigned((^~{$unsigned(reg4410)}));
                      reg7066 <= $unsigned(reg4358[(4'hd):(1'h1)]);
                      reg7067 <= reg4363[(2'h2):(1'h0)];
                    end
                end
            end
          for (forvar7068 = (1'h0); (forvar7068 < (1'h1)); forvar7068 = (forvar7068 + (1'h1)))
            begin
              if ((reg4493[(1'h1):(1'h0)] ^~ ($unsigned($signed(forvar4490)) <= $unsigned($signed(reg4413)))))
                begin
                  for (forvar7069 = (1'h0); (forvar7069 < (1'h0)); forvar7069 = (forvar7069 + (1'h1)))
                    begin
                      reg7070 <= reg4564[(4'hc):(1'h1)];
                      reg7071 <= reg7026[(1'h1):(1'h1)];
                      reg7072 <= reg4520[(1'h1):(1'h1)];
                      reg7073 <= {reg7062[(1'h1):(1'h0)]};
                    end
                end
              else
                begin
                  for (forvar7069 = (1'h0); (forvar7069 < (1'h0)); forvar7069 = (forvar7069 + (1'h1)))
                    begin
                      reg7070 <= reg4353;
                    end
                  for (forvar7071 = (1'h0); (forvar7071 < (1'h0)); forvar7071 = (forvar7071 + (1'h1)))
                    begin
                      reg7072 <= forvar4403[(4'ha):(3'h6)];
                      reg7073 <= {(($signed(reg4488) ?
                              (forvar4558 ?
                                  forvar4345 : reg4499) : {reg4495}) ~^ $unsigned($unsigned(forvar4538)))};
                      reg7074 <= reg4421[(4'he):(1'h0)];
                      reg7075 <= {reg4347[(4'ha):(4'h9)]};
                    end
                  if (({$unsigned($unsigned(reg4367))} >= reg4548[(2'h3):(2'h3)]))
                    begin
                      reg7076 <= ($unsigned($unsigned((&reg4432))) == reg7016[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg7076 <= reg4417;
                      reg7077 <= (^(reg4418[(3'h5):(2'h2)] ?
                          reg7044 : {(reg4543 ? reg4503 : forvar4504)}));
                      reg7078 <= (reg4361[(2'h3):(2'h3)] ?
                          forvar4496 : ({(~|reg4544)} <<< {(reg4508 ~^ forvar4414)}));
                    end
                  for (forvar7079 = (1'h0); (forvar7079 < (2'h3)); forvar7079 = (forvar7079 + (1'h1)))
                    begin
                      reg7080 <= ($unsigned(reg4484[(1'h1):(1'h0)]) ?
                          reg4427[(4'h8):(4'h8)] : (8'hb4));
                      reg7081 <= reg4400[(1'h1):(1'h0)];
                      reg7082 <= {reg4381};
                      reg7083 <= (|reg4473);
                    end
                end
            end
        end
      reg7084 <= $unsigned($signed($signed((forvar7010 ? (8'h9d) : reg4370))));
      reg7085 <= ((reg4528[(1'h1):(1'h1)] * reg4505) * ($signed(reg4570[(3'h4):(1'h1)]) ?
          {{reg4511}} : (+(reg4361 ? reg4560 : reg7032))));
    end
  always
    @(posedge clk) begin
      if (forvar7054)
        begin
          reg7086 <= (-forvar4356[(1'h1):(1'h0)]);
          if ($signed($unsigned(reg7043[(4'h8):(3'h5)])))
            begin
              reg7087 <= $unsigned((reg4404[(2'h2):(1'h1)] ?
                  (~$unsigned(reg7051)) : $signed({reg4356})));
              for (forvar7088 = (1'h0); (forvar7088 < (2'h2)); forvar7088 = (forvar7088 + (1'h1)))
                begin
                  for (forvar7089 = (1'h0); (forvar7089 < (1'h1)); forvar7089 = (forvar7089 + (1'h1)))
                    begin
                      reg7090 <= (reg4552[(2'h2):(2'h2)] ?
                          $unsigned(({reg4361} - $signed((8'ha4)))) : $signed(((8'ha7) <<< reg4510)));
                      reg7091 <= reg4415;
                      reg7092 <= $signed(reg4570[(2'h3):(2'h3)]);
                      reg7093 <= $signed((~^((reg4536 < reg4460) & (&reg7040))));
                    end
                  for (forvar7094 = (1'h0); (forvar7094 < (1'h1)); forvar7094 = (forvar7094 + (1'h1)))
                    begin
                      reg7095 <= reg4452[(3'h6):(2'h3)];
                      reg7096 <= $unsigned({reg4369[(2'h2):(2'h2)]});
                      reg7097 <= (forvar4476 ?
                          $unsigned(({reg4550} >= (forvar4522 ?
                              reg4483 : forvar4561))) : $signed(((+reg4423) <<< $signed(reg7080))));
                    end
                end
              if ($unsigned(((((8'ha2) ? reg4525 : reg4358) ?
                      $unsigned(reg4526) : ((8'hb6) ? reg7020 : reg4486)) ?
                  reg7026[(1'h1):(1'h1)] : $unsigned(reg4458))))
                begin
                  if (($signed(($signed(reg4506) > (~|reg7015))) ?
                      {(8'haa)} : ((reg4361[(3'h6):(2'h2)] * $signed((8'ha9))) ?
                          (^(forvar4476 >>> forvar4537)) : (reg7064[(1'h1):(1'h0)] ?
                              (-forvar7089) : (forvar4464 ~^ forvar7033)))))
                    begin
                      reg7098 <= forvar4538[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg7098 <= (!reg4468[(1'h1):(1'h0)]);
                    end
                  reg7099 <= ($unsigned($unsigned($signed(reg4444))) ?
                      $signed((-reg7061)) : $signed({{reg7058}}));
                  if ((((((8'haf) ? reg7030 : reg7044) ?
                              (reg4415 ? forvar4506 : reg7053) : reg4359) ?
                          (reg4482[(2'h3):(1'h0)] >= (reg4463 ?
                              forvar7094 : reg4565)) : reg4489) ?
                      reg4524[(4'h8):(2'h3)] : reg4468))
                    begin
                      reg7100 <= $unsigned(reg7027[(3'h4):(1'h1)]);
                      reg7101 <= forvar4456[(3'h5):(1'h0)];
                    end
                  else
                    begin
                      reg7100 <= reg4541;
                      reg7101 <= $unsigned({($unsigned((8'hb3)) && $unsigned(reg4520))});
                      reg7102 <= (~^reg4524);
                      reg7103 <= {$signed(reg7062)};
                    end
                end
              else
                begin
                  if ((~(reg4398[(2'h3):(1'h0)] ?
                      forvar4456 : forvar4553[(1'h1):(1'h1)])))
                    begin
                      reg7098 <= (~forvar7010[(4'h8):(3'h4)]);
                    end
                  else
                    begin
                      reg7098 <= ({$unsigned((forvar4364 << reg4472))} ?
                          reg4570 : (^{{reg4529}}));
                    end
                  if (reg7071[(4'h8):(3'h6)])
                    begin
                      reg7099 <= forvar4558[(3'h5):(2'h2)];
                      reg7100 <= reg4406;
                      reg7101 <= ($unsigned(((reg7100 ^ reg4545) >= (8'haf))) ?
                          {$unsigned((&reg7090))} : $unsigned({(&reg7086)}));
                      reg7102 <= ($signed((^forvar4535)) ?
                          reg7070 : (((reg4416 ? reg4413 : reg4544) ?
                                  reg4487[(2'h2):(1'h1)] : (reg4472 ?
                                      reg4390 : reg4533)) ?
                              (^$signed(forvar4364)) : $unsigned(((8'hae) ?
                                  forvar4408 : forvar4542))));
                    end
                  else
                    begin
                      reg7099 <= {forvar4542[(1'h1):(1'h1)]};
                      reg7100 <= ($unsigned({(+reg7099)}) ~^ $unsigned(reg4423[(2'h3):(1'h0)]));
                      reg7101 <= ($signed((^~$unsigned((8'haf)))) ?
                          (reg7041 ?
                              $signed($unsigned(reg4360)) : forvar4391[(3'h5):(2'h3)]) : $signed(($signed(forvar7088) ?
                              (forvar4537 > reg4461) : (forvar4554 ?
                                  reg4400 : forvar4522))));
                    end
                end
            end
          else
            begin
              for (forvar7087 = (1'h0); (forvar7087 < (2'h2)); forvar7087 = (forvar7087 + (1'h1)))
                begin
                  reg7088 <= (forvar4372[(3'h5):(1'h0)] ?
                      (-reg4405) : $signed((forvar4486 ?
                          reg4468[(4'ha):(3'h6)] : reg4550[(3'h7):(1'h0)])));
                end
            end
          if ($signed(forvar7094))
            begin
              if ((|(^$unsigned(forvar4509[(1'h1):(1'h0)]))))
                begin
                  for (forvar7104 = (1'h0); (forvar7104 < (1'h0)); forvar7104 = (forvar7104 + (1'h1)))
                    begin
                      reg7105 <= (^~reg4451[(4'ha):(3'h6)]);
                      reg7106 <= {$unsigned(reg7062)};
                      reg7107 <= (+(((reg4452 >> (8'ha4)) ?
                          reg7073 : {reg4433}) || $unsigned((!reg4523))));
                    end
                  if (($signed({$signed(reg4488)}) + ($signed({reg4376}) ?
                      $unsigned({reg4380}) : {(8'hae)})))
                    begin
                      reg7108 <= (({{(8'ha0)}} ?
                              reg7085[(4'ha):(3'h6)] : forvar4558) ?
                          (reg4470[(1'h1):(1'h1)] == $unsigned({(8'ha2)})) : (($signed((8'hb6)) ?
                              (reg4503 > (8'ha7)) : (+reg4387)) ^~ (reg7088[(1'h1):(1'h0)] ?
                              $signed(reg4539) : (^reg4502))));
                      reg7109 <= reg7056[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg7108 <= $unsigned($signed(reg4407));
                      reg7109 <= reg4492;
                      reg7110 <= $unsigned($unsigned(($signed(forvar4427) & (reg4481 ?
                          reg4407 : reg7040))));
                    end
                  if (((|reg4544[(2'h2):(2'h2)]) * (reg4511 + forvar4556[(1'h0):(1'h0)])))
                    begin
                      reg7111 <= (reg4385 ^~ $unsigned($signed((reg7038 & (8'h9d)))));
                      reg7112 <= $signed((~^($unsigned(forvar4520) ^~ $signed((8'hac)))));
                      reg7113 <= $signed((~((reg7025 ? reg7080 : reg4490) ?
                          (~^reg7034) : (reg7088 == reg4404))));
                    end
                  else
                    begin
                      reg7111 <= $signed((!($unsigned(reg4490) && {(8'ha4)})));
                    end
                end
              else
                begin
                  for (forvar7104 = (1'h0); (forvar7104 < (1'h0)); forvar7104 = (forvar7104 + (1'h1)))
                    begin
                      reg7105 <= reg4416[(3'h7):(2'h2)];
                    end
                  if (($unsigned(reg7099[(4'hf):(3'h6)]) ?
                      ((8'ha4) ?
                          {reg7041} : {$signed((8'hba))}) : $signed(((~&forvar7069) ?
                          {reg4422} : $unsigned(reg4506)))))
                    begin
                      reg7106 <= $unsigned($unsigned(((reg4444 ?
                              reg7057 : reg4564) ?
                          $unsigned(reg4362) : (reg4525 ?
                              forvar4486 : (8'h9c)))));
                      reg7107 <= {(~$signed((reg4430 || forvar4518)))};
                      reg7108 <= reg4425[(3'h4):(3'h4)];
                      reg7109 <= $signed($signed((8'hac)));
                    end
                  else
                    begin
                      reg7106 <= {((reg7045[(3'h6):(2'h3)] ?
                                  $unsigned(reg7045) : reg4373[(2'h2):(2'h2)]) ?
                              reg4508[(4'h8):(4'h8)] : (reg4435 ?
                                  reg4362[(4'ha):(3'h5)] : reg4396[(5'h10):(4'ha)]))};
                    end
                  reg7110 <= (reg4512[(4'ha):(2'h3)] ?
                      ({reg7050} >> (8'haf)) : $unsigned(forvar4561));
                  reg7111 <= $signed(forvar7037[(4'hd):(4'h9)]);
                end
              if ((~$signed(reg4350[(1'h1):(1'h0)])))
                begin
                  if (reg4499)
                    begin
                      reg7114 <= {reg7073[(4'he):(4'h9)]};
                      reg7115 <= (|{forvar7069[(3'h6):(2'h3)]});
                      reg7116 <= (&$unsigned($unsigned((~&forvar7023))));
                    end
                  else
                    begin
                      reg7114 <= ((^$unsigned(((8'hb9) ?
                          reg4511 : reg4477))) != {(forvar4412[(2'h2):(1'h1)] ?
                              (|reg7022) : reg4424[(3'h5):(1'h0)])});
                      reg7115 <= (8'ha1);
                      reg7116 <= (+({(forvar4459 ~^ (8'hb7))} > (|(|reg7105))));
                    end
                  if ($signed(reg7013))
                    begin
                      reg7117 <= {(+forvar7069[(4'hb):(4'ha)])};
                      reg7118 <= $unsigned($unsigned((forvar4344[(4'ha):(3'h7)] ?
                          (reg4412 <<< reg7101) : $unsigned(reg4458))));
                      reg7119 <= $unsigned(reg4353[(4'h8):(3'h5)]);
                    end
                  else
                    begin
                      reg7117 <= (reg7040[(4'h8):(3'h7)] ?
                          $unsigned(reg4395) : ($signed($signed(reg4540)) <<< ($signed(forvar4476) ?
                              (reg4438 >> reg4373) : $signed((8'hb4)))));
                    end
                  for (forvar7120 = (1'h0); (forvar7120 < (1'h1)); forvar7120 = (forvar7120 + (1'h1)))
                    begin
                      reg7121 <= (|(-reg7033[(3'h7):(2'h2)]));
                      reg7122 <= reg4410;
                      reg7123 <= ((~$unsigned((reg7057 ? (8'hae) : reg4418))) ?
                          reg4470[(2'h2):(2'h2)] : ($signed($unsigned(reg4538)) ?
                              reg7039[(1'h1):(1'h1)] : (((8'ha0) ?
                                  reg4376 : reg7083) >>> (forvar4403 ?
                                  reg4429 : reg4428))));
                    end
                end
              else
                begin
                  if ((({$signed(reg4362)} ?
                      (-(~|reg4453)) : forvar4500[(2'h3):(2'h3)]) && reg4442[(2'h2):(2'h2)]))
                    begin
                      reg7114 <= (~($signed((-(8'hb2))) >= ({reg4516} < reg7046)));
                      reg7115 <= (+({$unsigned(reg4435)} ?
                          ($unsigned((8'ha0)) >= reg4487[(3'h4):(3'h4)]) : (reg4548[(1'h0):(1'h0)] ?
                              reg7025[(2'h2):(2'h2)] : $signed(forvar4457))));
                      reg7116 <= reg4450;
                      reg7117 <= {$unsigned(reg4428[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg7114 <= ($signed((reg7031 ?
                              $signed(reg4441) : (-reg4514))) ?
                          ($signed($signed(reg4539)) && $signed($signed(forvar7104))) : (8'ha2));
                      reg7115 <= $unsigned(((forvar4475[(3'h4):(3'h4)] ?
                          reg4534[(1'h1):(1'h0)] : (forvar7071 ?
                              reg7065 : forvar7033)) >>> (!((8'had) || reg7097))));
                    end
                  if ($unsigned((~&(^((8'hab) ? reg4370 : reg7076)))))
                    begin
                      reg7118 <= ($signed({$signed(reg7070)}) ?
                          forvar7040[(4'hb):(4'h9)] : (forvar4506 & $signed((reg4555 ?
                              reg7052 : reg4493))));
                    end
                  else
                    begin
                      reg7118 <= {(reg4540[(1'h1):(1'h1)] >>> (^~{reg4388}))};
                    end
                end
              if ($unsigned($signed(reg7050[(2'h3):(2'h2)])))
                begin
                  reg7124 <= $unsigned(reg4455[(1'h0):(1'h0)]);
                  reg7125 <= $signed($signed(reg4543[(2'h3):(1'h1)]));
                end
              else
                begin
                  if (reg4526)
                    begin
                      reg7124 <= (($signed(forvar7087[(3'h4):(2'h2)]) ?
                          ($unsigned((8'hb5)) <<< $signed(reg7016)) : $unsigned(reg4407)) < $signed($signed(reg7060[(2'h3):(2'h2)])));
                    end
                  else
                    begin
                      reg7124 <= $signed((((forvar4391 ?
                          forvar7120 : wire4341) * reg7100) & wire4339));
                      reg7125 <= $unsigned((8'hba));
                    end
                  for (forvar7126 = (1'h0); (forvar7126 < (1'h0)); forvar7126 = (forvar7126 + (1'h1)))
                    begin
                      reg7127 <= ($unsigned((8'hab)) && (({reg4359} ?
                              $unsigned(reg4405) : reg4522[(3'h6):(1'h0)]) ?
                          $signed(((8'ha9) || forvar4427)) : reg4483[(1'h1):(1'h0)]));
                      reg7128 <= $signed($unsigned((|reg7030)));
                      reg7129 <= {reg4384};
                    end
                end
              for (forvar7130 = (1'h0); (forvar7130 < (1'h1)); forvar7130 = (forvar7130 + (1'h1)))
                begin
                  if (reg4471)
                    begin
                      reg7131 <= forvar4467[(4'hc):(1'h0)];
                    end
                  else
                    begin
                      reg7131 <= (8'hb8);
                      reg7132 <= reg4357[(1'h1):(1'h0)];
                      reg7133 <= ((reg7092[(3'h7):(3'h4)] ? reg4400 : reg4515) ?
                          reg4345 : $signed($signed((reg4439 ^~ reg4569))));
                      reg7134 <= $unsigned(({reg7025[(2'h2):(2'h2)]} > ($unsigned(reg7076) > (~|reg4539))));
                    end
                  for (forvar7135 = (1'h0); (forvar7135 < (2'h3)); forvar7135 = (forvar7135 + (1'h1)))
                    begin
                      reg7136 <= $signed(reg4516[(3'h4):(2'h3)]);
                      reg7137 <= $signed(forvar7044[(3'h4):(3'h4)]);
                      reg7138 <= $unsigned($signed($signed(((8'hb6) ?
                          reg7136 : (8'ha6)))));
                      reg7139 <= reg7067[(4'ha):(3'h4)];
                    end
                  for (forvar7140 = (1'h0); (forvar7140 < (2'h3)); forvar7140 = (forvar7140 + (1'h1)))
                    begin
                      reg7141 <= $signed({reg4361});
                      reg7142 <= reg7118[(4'hc):(1'h0)];
                      reg7143 <= reg7042[(2'h2):(1'h0)];
                      reg7144 <= (~&$signed($unsigned({(8'ha0)})));
                    end
                end
            end
          else
            begin
              for (forvar7104 = (1'h0); (forvar7104 < (2'h2)); forvar7104 = (forvar7104 + (1'h1)))
                begin
                  reg7105 <= (-reg7026);
                  for (forvar7106 = (1'h0); (forvar7106 < (1'h1)); forvar7106 = (forvar7106 + (1'h1)))
                    begin
                      reg7107 <= $unsigned($signed($signed((reg4388 ?
                          reg4461 : reg4383))));
                      reg7108 <= $signed((+$signed(forvar4567[(1'h1):(1'h1)])));
                      reg7109 <= {forvar4522};
                      reg7110 <= $unsigned($signed(forvar4506));
                    end
                end
              for (forvar7111 = (1'h0); (forvar7111 < (2'h3)); forvar7111 = (forvar7111 + (1'h1)))
                begin
                  for (forvar7112 = (1'h0); (forvar7112 < (2'h2)); forvar7112 = (forvar7112 + (1'h1)))
                    begin
                      reg7113 <= reg7072;
                      reg7114 <= reg7045;
                    end
                  reg7115 <= reg4544[(1'h1):(1'h1)];
                  reg7116 <= reg4458[(2'h2):(2'h2)];
                  if ((reg4417 >> reg7091[(3'h5):(3'h4)]))
                    begin
                      reg7117 <= forvar4535[(2'h2):(1'h0)];
                      reg7118 <= $signed({{(reg7119 ? reg4525 : reg7085)}});
                      reg7119 <= reg7088;
                    end
                  else
                    begin
                      reg7117 <= reg4465[(1'h1):(1'h0)];
                      reg7118 <= $unsigned($signed($unsigned(((8'hae) <<< reg4378))));
                      reg7119 <= $signed((forvar7089 >= $signed((~^forvar7069))));
                      reg7120 <= ((((~|reg4381) ?
                          reg4522[(2'h3):(2'h2)] : $unsigned(reg7070)) | $unsigned($signed(wire4338))) >>> $signed(reg7028));
                    end
                end
              for (forvar7121 = (1'h0); (forvar7121 < (2'h2)); forvar7121 = (forvar7121 + (1'h1)))
                begin
                  reg7122 <= ($signed(forvar4423[(4'h9):(1'h1)]) < (8'ha2));
                  for (forvar7123 = (1'h0); (forvar7123 < (2'h2)); forvar7123 = (forvar7123 + (1'h1)))
                    begin
                      reg7124 <= $signed($unsigned(($signed(forvar4401) > (8'hb0))));
                      reg7125 <= (8'hb9);
                      reg7126 <= (&reg7087);
                      reg7127 <= ((((reg4428 ?
                                  reg4441 : forvar4520) & forvar4568) ?
                              reg4447[(2'h3):(1'h0)] : forvar4509[(4'hd):(4'hb)]) ?
                          $unsigned(wire4338[(3'h4):(3'h4)]) : reg7035[(2'h3):(1'h1)]);
                    end
                  if ((reg7022 <= reg7131[(2'h2):(2'h2)]))
                    begin
                      reg7128 <= (8'ha0);
                      reg7129 <= (reg4395[(1'h0):(1'h0)] ~^ reg7036);
                    end
                  else
                    begin
                      reg7128 <= reg4445;
                    end
                  reg7130 <= {{$unsigned((&forvar4467))}};
                end
              if (forvar4538)
                begin
                  for (forvar7131 = (1'h0); (forvar7131 < (1'h1)); forvar7131 = (forvar7131 + (1'h1)))
                    begin
                      reg7132 <= (reg4412[(1'h1):(1'h1)] ?
                          reg4371 : reg7097[(3'h5):(2'h2)]);
                      reg7133 <= reg7128[(3'h7):(3'h6)];
                      reg7134 <= ((({reg7020} ^ (8'ha7)) ^ $signed(reg4434[(4'h8):(3'h6)])) ?
                          ((-(~^reg4424)) ?
                              forvar7068 : ((reg4463 ?
                                  reg4487 : (8'ha3)) - reg7022)) : reg4384);
                      reg7135 <= (!((^$signed(reg7075)) ?
                          forvar7094[(1'h1):(1'h1)] : {(reg4370 >= forvar4546)}));
                    end
                  for (forvar7136 = (1'h0); (forvar7136 < (1'h0)); forvar7136 = (forvar7136 + (1'h1)))
                    begin
                      reg7137 <= ({{{reg4482}}} ?
                          ({(reg4474 ? (8'h9d) : reg7076)} ?
                              reg7136[(1'h1):(1'h1)] : $signed((reg4352 ^ forvar4345))) : $signed(({forvar4522} > $unsigned(reg7059))));
                    end
                  for (forvar7138 = (1'h0); (forvar7138 < (2'h2)); forvar7138 = (forvar7138 + (1'h1)))
                    begin
                      reg7139 <= (!(&$signed(reg7024[(1'h0):(1'h0)])));
                      reg7140 <= (8'ha0);
                      reg7141 <= $signed($unsigned(reg7128));
                      reg7142 <= reg4483;
                    end
                  for (forvar7143 = (1'h0); (forvar7143 < (1'h0)); forvar7143 = (forvar7143 + (1'h1)))
                    begin
                      reg7144 <= ({$unsigned((8'ha2))} >= (8'ha7));
                      reg7145 <= (~^$unsigned((^~reg4470)));
                    end
                end
              else
                begin
                  for (forvar7131 = (1'h0); (forvar7131 < (1'h0)); forvar7131 = (forvar7131 + (1'h1)))
                    begin
                      reg7132 <= (~|((~^$signed(reg7053)) ?
                          (-wire4341[(3'h6):(2'h2)]) : reg4430));
                      reg7133 <= (reg4402[(2'h3):(2'h3)] >= (((-reg4492) && (reg4345 ?
                          reg4409 : reg7082)) ~^ $signed((-reg7078))));
                      reg7134 <= (reg7066[(3'h4):(2'h3)] || reg4396[(3'h4):(3'h4)]);
                      reg7135 <= reg4565;
                    end
                  for (forvar7136 = (1'h0); (forvar7136 < (1'h0)); forvar7136 = (forvar7136 + (1'h1)))
                    begin
                      reg7137 <= (((-(!reg4552)) > reg7082) ?
                          reg7095 : $unsigned(($unsigned(forvar4504) ?
                              (forvar4408 ?
                                  reg4429 : reg4391) : (|forvar7130))));
                    end
                  reg7138 <= ($signed(($signed(reg4371) > (forvar4344 ?
                          reg4455 : reg4370))) ?
                      $signed(wire4571) : ({(reg4423 || reg4431)} && reg7141[(3'h5):(1'h1)]));
                  for (forvar7139 = (1'h0); (forvar7139 < (1'h1)); forvar7139 = (forvar7139 + (1'h1)))
                    begin
                      reg7140 <= reg4359;
                    end
                end
            end
          reg7146 <= forvar7087;
        end
      else
        begin
          if (reg4507)
            begin
              for (forvar7086 = (1'h0); (forvar7086 < (1'h0)); forvar7086 = (forvar7086 + (1'h1)))
                begin
                  for (forvar7087 = (1'h0); (forvar7087 < (2'h3)); forvar7087 = (forvar7087 + (1'h1)))
                    begin
                      reg7088 <= $signed($unsigned(($unsigned(forvar4386) ?
                          $unsigned(reg7015) : forvar4374[(3'h4):(1'h1)])));
                      reg7089 <= reg7099;
                    end
                  for (forvar7090 = (1'h0); (forvar7090 < (2'h3)); forvar7090 = (forvar7090 + (1'h1)))
                    begin
                      reg7091 <= forvar4359[(3'h6):(2'h3)];
                    end
                  if ((~^(((forvar4459 ?
                      reg4480 : reg4413) - forvar7089) && $signed(forvar4485[(4'h8):(3'h6)]))))
                    begin
                      reg7092 <= {((+(reg4433 << reg4503)) == (8'ha6))};
                      reg7093 <= $signed((forvar7030[(3'h5):(1'h0)] ?
                          ((8'hab) ?
                              reg4510 : (!reg4409)) : reg7066[(1'h0):(1'h0)]));
                      reg7094 <= forvar4356[(4'h9):(4'h8)];
                      reg7095 <= reg4559[(3'h7):(2'h3)];
                    end
                  else
                    begin
                      reg7092 <= (($signed({reg4506}) ?
                              (-reg7061) : ((^reg7145) * $signed(reg4422))) ?
                          (((forvar4350 ? reg7099 : reg4438) ?
                              reg7080 : reg4537) <= reg4515[(1'h1):(1'h1)]) : {((8'h9d) ?
                                  (reg7014 || reg4550) : reg7064[(1'h1):(1'h0)])});
                    end
                  if ((!$unsigned(((~|reg4417) ~^ $signed(reg7085)))))
                    begin
                      reg7096 <= ($signed($unsigned({reg7051})) ~^ reg4525);
                    end
                  else
                    begin
                      reg7096 <= forvar7048;
                      reg7097 <= ({(~^(reg4498 > forvar7071))} + $signed(((reg7029 << reg7115) ?
                          reg4505[(4'ha):(4'h9)] : (reg4459 ?
                              reg4447 : reg7015))));
                      reg7098 <= (+($signed(((8'had) || reg4531)) ?
                          (((8'ha8) ? forvar7120 : reg4470) ?
                              (reg7062 || forvar4386) : reg4524[(1'h0):(1'h0)]) : {(reg4483 ^~ reg4540)}));
                      reg7099 <= (reg4484 | $signed($signed((8'hb5))));
                    end
                end
              reg7100 <= $signed({wire7008[(3'h4):(1'h1)]});
            end
          else
            begin
              for (forvar7086 = (1'h0); (forvar7086 < (1'h0)); forvar7086 = (forvar7086 + (1'h1)))
                begin
                  for (forvar7087 = (1'h0); (forvar7087 < (2'h3)); forvar7087 = (forvar7087 + (1'h1)))
                    begin
                      reg7088 <= reg4360[(3'h6):(1'h0)];
                      reg7089 <= $signed((reg4545 ? reg4355 : reg4458));
                      reg7090 <= (reg4433[(1'h0):(1'h0)] ?
                          (&$unsigned($signed(reg4409))) : {forvar4554});
                    end
                  if ($signed((8'ha0)))
                    begin
                      reg7091 <= $signed($signed({forvar4374}));
                    end
                  else
                    begin
                      reg7091 <= ($signed($unsigned(((8'hb4) == reg4496))) ?
                          (reg4526[(2'h3):(1'h0)] - ($unsigned(forvar7011) ?
                              (+forvar7090) : (+reg4517))) : (^reg7125));
                      reg7092 <= reg7087;
                    end
                  for (forvar7093 = (1'h0); (forvar7093 < (2'h3)); forvar7093 = (forvar7093 + (1'h1)))
                    begin
                      reg7094 <= (~&reg4380);
                      reg7095 <= {reg7133};
                      reg7096 <= reg7024[(2'h2):(2'h2)];
                      reg7097 <= (^~$unsigned(reg7067));
                    end
                end
              if ((|(~|((-reg4447) - ((8'ha9) > reg4394)))))
                begin
                  for (forvar7098 = (1'h0); (forvar7098 < (2'h3)); forvar7098 = (forvar7098 + (1'h1)))
                    begin
                      reg7099 <= (!(^~(8'ha4)));
                      reg7100 <= (^~(reg7084 ? {{reg4550}} : reg4499));
                      reg7101 <= $unsigned($signed($unsigned((reg7145 ?
                          reg4471 : reg4399))));
                    end
                  if ((reg4531[(3'h5):(1'h1)] ?
                      reg4508 : forvar7104[(3'h4):(1'h0)]))
                    begin
                      reg7102 <= {forvar4346[(3'h7):(3'h7)]};
                    end
                  else
                    begin
                      reg7102 <= (reg4565 <<< reg4347);
                    end
                end
              else
                begin
                  reg7098 <= $signed(reg4493[(3'h6):(2'h3)]);
                  for (forvar7099 = (1'h0); (forvar7099 < (1'h1)); forvar7099 = (forvar7099 + (1'h1)))
                    begin
                      reg7100 <= forvar7123;
                      reg7101 <= (^~(((reg7112 ~^ reg7111) ?
                          forvar7090 : (reg4493 ?
                              reg4512 : reg7112)) < $unsigned((reg7118 ?
                          reg4460 : (8'ha6)))));
                      reg7102 <= reg7013[(1'h0):(1'h0)];
                    end
                end
            end
          if ((~&reg4431))
            begin
              for (forvar7103 = (1'h0); (forvar7103 < (1'h1)); forvar7103 = (forvar7103 + (1'h1)))
                begin
                  for (forvar7104 = (1'h0); (forvar7104 < (2'h2)); forvar7104 = (forvar7104 + (1'h1)))
                    begin
                      reg7105 <= $unsigned(forvar7047[(3'h4):(3'h4)]);
                    end
                  if ((^(((~|reg4416) || $signed((8'hb5))) ?
                      reg4365[(4'ha):(3'h6)] : reg7036[(2'h2):(2'h2)])))
                    begin
                      reg7106 <= (^((^~$unsigned((8'had))) > ($signed(reg4469) ?
                          (reg4358 ? reg4395 : reg4422) : (reg7086 ?
                              (8'ha6) : forvar4568))));
                    end
                  else
                    begin
                      reg7106 <= reg7032;
                      reg7107 <= ($signed((~((8'hb5) >> reg4413))) ?
                          $signed(reg4470) : ($signed(reg4548) ?
                              $unsigned(reg4429) : forvar4440));
                      reg7108 <= (^~$unsigned(forvar7040));
                      reg7109 <= ({{forvar7048[(4'hc):(1'h1)]}} > reg4460);
                    end
                  if (forvar4413[(2'h2):(2'h2)])
                    begin
                      reg7110 <= forvar4436;
                      reg7111 <= reg7060[(2'h3):(1'h1)];
                      reg7112 <= $unsigned(reg4497);
                      reg7113 <= ((reg4428[(1'h1):(1'h0)] ?
                              reg4427[(2'h3):(1'h1)] : (((8'ha4) ?
                                  reg7133 : (8'h9f)) != forvar7121[(1'h0):(1'h0)])) ?
                          {($signed(reg4514) ?
                                  $unsigned(wire4571) : (~|reg4390))} : (8'ha4));
                    end
                  else
                    begin
                      reg7110 <= (-forvar4567);
                    end
                end
            end
          else
            begin
              reg7103 <= $signed(($signed(forvar7090[(3'h6):(1'h0)]) ?
                  (forvar4422[(3'h6):(2'h2)] ?
                      (8'ha9) : $signed(reg7141)) : forvar4423[(3'h7):(3'h7)]));
              for (forvar7104 = (1'h0); (forvar7104 < (2'h3)); forvar7104 = (forvar7104 + (1'h1)))
                begin
                  reg7105 <= reg7073;
                  for (forvar7106 = (1'h0); (forvar7106 < (1'h1)); forvar7106 = (forvar7106 + (1'h1)))
                    begin
                      reg7107 <= $unsigned($signed(((reg4469 ?
                              forvar4485 : reg4380) ?
                          (forvar7138 << forvar4487) : (reg4345 ?
                              forvar7037 : reg4367))));
                    end
                end
            end
          if (forvar7044)
            begin
              for (forvar7114 = (1'h0); (forvar7114 < (2'h3)); forvar7114 = (forvar7114 + (1'h1)))
                begin
                  for (forvar7115 = (1'h0); (forvar7115 < (1'h1)); forvar7115 = (forvar7115 + (1'h1)))
                    begin
                      reg7116 <= (&$unsigned($unsigned({reg7124})));
                    end
                end
              if (reg4452)
                begin
                  reg7117 <= ((~^(reg4448[(1'h0):(1'h0)] ?
                          reg4356[(4'hb):(4'h9)] : (forvar7111 ?
                              forvar4345 : (8'hba)))) ?
                      $signed(((-forvar4518) ?
                          $signed(reg4463) : (~|reg7095))) : (reg4371[(3'h4):(1'h1)] >= (^~$signed(reg4438))));
                  for (forvar7118 = (1'h0); (forvar7118 < (1'h1)); forvar7118 = (forvar7118 + (1'h1)))
                    begin
                      reg7119 <= ((($unsigned(forvar7126) + $signed(reg4421)) << (reg7090[(1'h0):(1'h0)] * $signed((8'h9d)))) + $signed((~|(forvar7140 ?
                          reg4491 : (8'h9f)))));
                      reg7120 <= reg4392[(1'h1):(1'h0)];
                    end
                  for (forvar7121 = (1'h0); (forvar7121 < (2'h2)); forvar7121 = (forvar7121 + (1'h1)))
                    begin
                      reg7122 <= reg4400;
                    end
                end
              else
                begin
                  if ((reg4505[(3'h6):(2'h3)] ?
                      ($signed({forvar4344}) ?
                          reg4505 : forvar4459) : $signed($unsigned($signed((8'hb6))))))
                    begin
                      reg7117 <= reg7027[(2'h2):(1'h1)];
                      reg7118 <= $signed(reg7083[(3'h6):(3'h4)]);
                      reg7119 <= forvar4530[(1'h0):(1'h0)];
                      reg7120 <= reg7031;
                    end
                  else
                    begin
                      reg7117 <= $unsigned($unsigned(((^~(8'ha6)) ?
                          $signed(reg7119) : $unsigned((8'ha8)))));
                      reg7118 <= ((8'ha4) ?
                          $signed(((&reg7039) <<< reg4424[(2'h3):(2'h2)])) : (({(8'h9e)} ?
                              {forvar4542} : (8'ha2)) <<< $unsigned(forvar4547)));
                      reg7119 <= {(($unsigned(reg4548) ?
                              (~reg4421) : (reg7110 ?
                                  reg7083 : reg4396)) > $unsigned((reg4363 || reg4367)))};
                    end
                end
              reg7123 <= wire4343;
            end
          else
            begin
              for (forvar7114 = (1'h0); (forvar7114 < (2'h3)); forvar7114 = (forvar7114 + (1'h1)))
                begin
                  reg7115 <= forvar4459[(1'h0):(1'h0)];
                  for (forvar7116 = (1'h0); (forvar7116 < (1'h0)); forvar7116 = (forvar7116 + (1'h1)))
                    begin
                      reg7117 <= reg4497[(3'h4):(2'h2)];
                      reg7118 <= {reg7118};
                      reg7119 <= $unsigned(({(+reg4524)} && ($unsigned((8'ha1)) ?
                          {reg7135} : (!reg7121))));
                      reg7120 <= reg7113[(4'h9):(3'h5)];
                    end
                  for (forvar7121 = (1'h0); (forvar7121 < (2'h3)); forvar7121 = (forvar7121 + (1'h1)))
                    begin
                      reg7122 <= (^~reg7076);
                      reg7123 <= forvar4353[(3'h4):(2'h2)];
                      reg7124 <= reg7083;
                    end
                end
            end
          for (forvar7125 = (1'h0); (forvar7125 < (1'h1)); forvar7125 = (forvar7125 + (1'h1)))
            begin
              if ({$unsigned((reg7050[(2'h3):(2'h3)] ?
                      (forvar4401 ?
                          reg4480 : reg4446) : $unsigned(forvar4345)))})
                begin
                  for (forvar7126 = (1'h0); (forvar7126 < (2'h3)); forvar7126 = (forvar7126 + (1'h1)))
                    begin
                      reg7127 <= forvar4556[(1'h1):(1'h1)];
                      reg7128 <= $signed(reg4371[(3'h5):(2'h2)]);
                      reg7129 <= (~(+$signed($signed(reg4522))));
                    end
                  if ((forvar4352 ?
                      $unsigned(reg4345[(4'ha):(4'ha)]) : reg4347))
                    begin
                      reg7130 <= reg7013[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg7130 <= reg4386;
                      reg7131 <= (reg4410 ?
                          reg4361 : ($unsigned(forvar4346[(4'h8):(2'h3)]) ?
                              reg4514 : forvar4501[(4'hd):(4'h9)]));
                    end
                  reg7132 <= ({reg4526[(1'h1):(1'h1)]} ?
                      (~&$unsigned((|(8'hb1)))) : $unsigned(reg4432[(3'h6):(1'h1)]));
                end
              else
                begin
                  for (forvar7126 = (1'h0); (forvar7126 < (1'h0)); forvar7126 = (forvar7126 + (1'h1)))
                    begin
                      reg7127 <= ($signed($signed((^forvar4554))) && reg7139);
                      reg7128 <= {(!$unsigned($unsigned(forvar7140)))};
                    end
                  for (forvar7129 = (1'h0); (forvar7129 < (1'h1)); forvar7129 = (forvar7129 + (1'h1)))
                    begin
                      reg7130 <= reg4348;
                      reg7131 <= (((^$signed(reg4490)) ?
                              reg4375 : $unsigned(reg7016[(2'h2):(1'h0)])) ?
                          (forvar7116 - ((reg4529 ?
                              reg7095 : reg4390) == $signed(reg4451))) : (~^$unsigned({reg4448})));
                    end
                  for (forvar7132 = (1'h0); (forvar7132 < (1'h0)); forvar7132 = (forvar7132 + (1'h1)))
                    begin
                      reg7133 <= $unsigned(($signed({forvar4554}) ?
                          $unsigned($signed(reg4359)) : {reg7145}));
                    end
                  for (forvar7134 = (1'h0); (forvar7134 < (2'h2)); forvar7134 = (forvar7134 + (1'h1)))
                    begin
                      reg7135 <= reg4410[(2'h3):(1'h1)];
                      reg7136 <= reg7024[(1'h0):(1'h0)];
                      reg7137 <= $signed((reg4419 < $unsigned(reg4442[(2'h2):(1'h1)])));
                      reg7138 <= $unsigned($signed({{reg7081}}));
                    end
                end
              for (forvar7139 = (1'h0); (forvar7139 < (2'h3)); forvar7139 = (forvar7139 + (1'h1)))
                begin
                  if (reg4542)
                    begin
                      reg7140 <= $unsigned(reg7095);
                    end
                  else
                    begin
                      reg7140 <= ({$signed(forvar4464[(1'h0):(1'h0)])} <= $signed($unsigned((reg4531 ?
                          reg4469 : reg7019))));
                    end
                end
              for (forvar7141 = (1'h0); (forvar7141 < (2'h3)); forvar7141 = (forvar7141 + (1'h1)))
                begin
                  for (forvar7142 = (1'h0); (forvar7142 < (1'h0)); forvar7142 = (forvar7142 + (1'h1)))
                    begin
                      reg7143 <= {forvar7125};
                      reg7144 <= forvar4509;
                      reg7145 <= reg7135[(2'h3):(2'h3)];
                      reg7146 <= forvar4538[(4'hb):(4'h9)];
                    end
                end
              reg7147 <= $unsigned(((~(forvar4414 ?
                  (8'hb9) : reg4503)) <<< reg4485));
            end
        end
      if (forvar4347)
        begin
          if (reg7086[(4'hd):(3'h4)])
            begin
              for (forvar7148 = (1'h0); (forvar7148 < (1'h1)); forvar7148 = (forvar7148 + (1'h1)))
                begin
                  for (forvar7149 = (1'h0); (forvar7149 < (1'h0)); forvar7149 = (forvar7149 + (1'h1)))
                    begin
                      reg7150 <= (^(-$unsigned(reg4399[(4'ha):(3'h5)])));
                      reg7151 <= ((|(forvar4427 + $signed((8'hb4)))) ?
                          ((+(reg7124 ?
                              reg4521 : forvar4344)) ^ $signed(reg4349[(2'h2):(2'h2)])) : ((~|(reg7028 == reg7122)) ?
                              $unsigned($unsigned(reg7123)) : (^(reg7018 ?
                                  forvar4391 : reg4472))));
                    end
                end
              for (forvar7152 = (1'h0); (forvar7152 < (1'h0)); forvar7152 = (forvar7152 + (1'h1)))
                begin
                  if ((&{(8'ha4)}))
                    begin
                      reg7153 <= $unsigned(reg4512[(2'h3):(1'h0)]);
                      reg7154 <= ($unsigned({$unsigned(reg7026)}) ?
                          $unsigned(((reg7057 + forvar7048) & {forvar4475})) : $signed(({reg7113} ?
                              (reg7051 * (8'hba)) : reg4433[(3'h5):(1'h0)])));
                      reg7155 <= ($unsigned(reg7099[(4'hc):(2'h2)]) ?
                          $unsigned(forvar7125) : $signed(($unsigned(reg4536) >>> $signed(reg7043))));
                    end
                  else
                    begin
                      reg7153 <= reg4452[(4'ha):(4'ha)];
                      reg7154 <= $signed(reg4361[(1'h0):(1'h0)]);
                      reg7155 <= $unsigned({reg4356});
                      reg7156 <= reg7131[(1'h0):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar7148 = (1'h0); (forvar7148 < (1'h0)); forvar7148 = (forvar7148 + (1'h1)))
                begin
                  reg7149 <= reg4570[(3'h4):(3'h4)];
                end
              if ((reg4511 & forvar4459[(2'h2):(1'h0)]))
                begin
                  for (forvar7150 = (1'h0); (forvar7150 < (2'h2)); forvar7150 = (forvar7150 + (1'h1)))
                    begin
                      reg7151 <= reg4538;
                      reg7152 <= (reg4484[(2'h3):(2'h2)] <<< reg7097);
                    end
                  for (forvar7153 = (1'h0); (forvar7153 < (1'h0)); forvar7153 = (forvar7153 + (1'h1)))
                    begin
                      reg7154 <= $signed((-(|((8'ha6) ? reg7097 : reg7080))));
                      reg7155 <= ($unsigned(($signed(forvar7068) && $unsigned(reg4351))) & $unsigned($unsigned($unsigned(reg4489))));
                    end
                end
              else
                begin
                  if (reg4487)
                    begin
                      reg7150 <= (reg4497[(4'h9):(1'h0)] > (~^reg4349));
                      reg7151 <= {{(~(reg4565 <<< forvar4567))}};
                      reg7152 <= (~&(($unsigned(forvar4518) == (&forvar7104)) ?
                          $unsigned({reg7034}) : ($signed(reg4369) && (reg4376 ?
                              reg4345 : wire7006))));
                    end
                  else
                    begin
                      reg7150 <= ((8'ha2) ~^ reg4494[(3'h6):(2'h3)]);
                      reg7151 <= reg4517;
                      reg7152 <= (&((|(reg7081 ? (8'ha7) : forvar4364)) ?
                          reg7083[(3'h4):(1'h1)] : $unsigned($unsigned((8'ha8)))));
                      reg7153 <= ({$signed($signed(reg4537))} + reg4373);
                    end
                  for (forvar7154 = (1'h0); (forvar7154 < (2'h3)); forvar7154 = (forvar7154 + (1'h1)))
                    begin
                      reg7155 <= reg4511;
                      reg7156 <= $signed((-{reg7028[(2'h2):(1'h1)]}));
                      reg7157 <= (~&$unsigned(((8'haa) ?
                          $unsigned(reg4510) : $signed(reg7113))));
                      reg7158 <= ({$signed($signed((8'h9f)))} >= $unsigned(forvar4567[(3'h7):(2'h3)]));
                    end
                end
              for (forvar7159 = (1'h0); (forvar7159 < (1'h0)); forvar7159 = (forvar7159 + (1'h1)))
                begin
                  for (forvar7160 = (1'h0); (forvar7160 < (2'h2)); forvar7160 = (forvar7160 + (1'h1)))
                    begin
                      reg7161 <= (|$signed(reg4477[(4'hb):(1'h1)]));
                      reg7162 <= ((-{{reg4569}}) ^ ($signed($signed(reg7084)) ?
                          forvar7138[(2'h2):(1'h0)] : $signed(reg4418[(2'h3):(2'h2)])));
                    end
                  if ($unsigned(reg4519))
                    begin
                      reg7163 <= $signed((reg4381 | $signed((^~forvar4496))));
                      reg7164 <= {reg4512[(3'h6):(1'h0)]};
                    end
                  else
                    begin
                      reg7163 <= {$unsigned((~|(forvar7106 ?
                              reg7050 : reg7111)))};
                      reg7164 <= (!{(~^$unsigned(forvar7131))});
                    end
                  reg7165 <= reg7138;
                  if (((~$unsigned($unsigned((8'hb6)))) ?
                      (reg4468 && reg4442[(1'h0):(1'h0)]) : ($signed((+reg4400)) - (forvar7089 ~^ reg4360[(4'h9):(1'h1)]))))
                    begin
                      reg7166 <= forvar7012[(3'h6):(1'h0)];
                      reg7167 <= {$signed(reg4356[(4'h8):(4'h8)])};
                      reg7168 <= {$unsigned($unsigned(reg4461))};
                    end
                  else
                    begin
                      reg7166 <= $signed({((^reg4504) && ((8'hab) ?
                              reg4372 : reg7055))});
                    end
                end
            end
          if (reg4564[(1'h0):(1'h0)])
            begin
              for (forvar7169 = (1'h0); (forvar7169 < (1'h0)); forvar7169 = (forvar7169 + (1'h1)))
                begin
                  for (forvar7170 = (1'h0); (forvar7170 < (2'h2)); forvar7170 = (forvar7170 + (1'h1)))
                    begin
                      reg7171 <= reg4473;
                      reg7172 <= (8'hb0);
                    end
                  if ({{(^~(reg7078 ? reg4515 : forvar4440))}})
                    begin
                      reg7173 <= forvar4554[(2'h2):(1'h0)];
                      reg7174 <= (~^(~|{(reg7097 ? reg4431 : reg7067)}));
                      reg7175 <= (8'h9e);
                      reg7176 <= ((reg4425[(2'h2):(1'h0)] < forvar7141[(1'h1):(1'h0)]) ~^ (($signed(reg7040) ?
                              $signed((8'hb1)) : $unsigned(reg7018)) ?
                          $signed((~&reg4402)) : forvar7130[(4'h9):(2'h2)]));
                    end
                  else
                    begin
                      reg7173 <= (8'haf);
                      reg7174 <= reg4394;
                    end
                  if (($signed((8'hb2)) ^~ (reg7115[(2'h2):(1'h1)] ?
                      ($signed((8'haa)) ?
                          (+forvar7148) : (^~reg4424)) : $signed((reg4415 ~^ reg7066)))))
                    begin
                      reg7177 <= $signed($unsigned((-(~reg7090))));
                      reg7178 <= $signed(reg4351[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg7177 <= (^($unsigned({forvar7154}) - {reg4380[(4'h8):(3'h7)]}));
                      reg7178 <= {forvar4542[(1'h0):(1'h0)]};
                      reg7179 <= ((reg4435 ?
                          ((reg4543 - (8'hb0)) <= $signed(reg4509)) : reg4348[(1'h0):(1'h0)]) & $signed($unsigned($signed(reg7026))));
                    end
                  reg7180 <= (((^~(reg4359 ?
                      (8'ha8) : reg7105)) && reg7097) ^~ (reg7162 ?
                      ({reg7117} ?
                          (8'ha6) : (wire4338 ?
                              reg4399 : forvar4509)) : $unsigned((~^(8'hac)))));
                end
              for (forvar7181 = (1'h0); (forvar7181 < (2'h3)); forvar7181 = (forvar7181 + (1'h1)))
                begin
                  reg7182 <= forvar7169;
                end
              for (forvar7183 = (1'h0); (forvar7183 < (2'h2)); forvar7183 = (forvar7183 + (1'h1)))
                begin
                  if ((reg4504 ?
                      (reg7018 ^ forvar7121[(4'hb):(3'h4)]) : ($signed((reg7109 ?
                          reg7051 : forvar7154)) ^~ {{(8'hb1)}})))
                    begin
                      reg7184 <= forvar7125[(4'hb):(4'h9)];
                      reg7185 <= ($unsigned($signed((reg4453 <= (8'h9d)))) || (+($signed(forvar4506) ?
                          (forvar7111 ^ (8'hb3)) : reg4500[(3'h5):(3'h4)])));
                      reg7186 <= $signed($signed($unsigned({reg7152})));
                      reg7187 <= $unsigned(($signed((forvar4467 ^~ forvar4510)) ?
                          reg7092[(3'h6):(3'h6)] : $signed((8'ha6))));
                    end
                  else
                    begin
                      reg7184 <= (+reg7041[(2'h2):(1'h1)]);
                      reg7185 <= {$unsigned($signed(forvar7130[(4'he):(2'h3)]))};
                      reg7186 <= ((forvar4553[(1'h1):(1'h0)] >= $signed($unsigned(reg4345))) ?
                          ($unsigned((reg7136 <= reg4410)) ?
                              {(!reg7093)} : {$unsigned(forvar4368)}) : reg7164);
                    end
                  if ((reg7035[(3'h7):(1'h0)] ?
                      $unsigned(((reg4515 ?
                          reg7019 : reg7155) <= (forvar7123 && forvar7123))) : (+reg7066[(4'h9):(3'h7)])))
                    begin
                      reg7188 <= forvar4437[(4'ha):(4'ha)];
                    end
                  else
                    begin
                      reg7188 <= reg7114;
                      reg7189 <= (-$unsigned($signed($signed(reg7188))));
                    end
                end
              reg7190 <= (8'hb6);
            end
          else
            begin
              for (forvar7169 = (1'h0); (forvar7169 < (2'h2)); forvar7169 = (forvar7169 + (1'h1)))
                begin
                  reg7170 <= forvar4487;
                  reg7171 <= reg7173[(3'h5):(3'h4)];
                end
            end
          for (forvar7191 = (1'h0); (forvar7191 < (1'h0)); forvar7191 = (forvar7191 + (1'h1)))
            begin
              if (({wire4339[(2'h2):(1'h1)]} ?
                  (reg4489 * ((reg4540 - reg4501) > $unsigned(reg7031))) : reg7032[(3'h4):(2'h2)]))
                begin
                  if (($unsigned($signed($unsigned(reg4548))) ?
                      ({{reg7134}} || $signed(reg7138[(1'h0):(1'h0)])) : ((|forvar4423[(1'h0):(1'h0)]) ?
                          $signed((forvar4346 ^~ reg4550)) : reg4511)))
                    begin
                      reg7192 <= forvar4501[(4'h8):(3'h7)];
                      reg7193 <= $unsigned({(&(-forvar7047))});
                      reg7194 <= (8'hba);
                    end
                  else
                    begin
                      reg7192 <= wire7008[(2'h3):(2'h3)];
                      reg7193 <= (reg4441 | (+(reg7040[(3'h4):(2'h2)] << (^forvar7044))));
                      reg7194 <= ((({reg4560} - reg7133) ?
                              reg7140[(2'h2):(2'h2)] : ((forvar7129 ?
                                  forvar4527 : forvar4436) & $signed(reg4421))) ?
                          reg7111[(1'h1):(1'h1)] : forvar4412[(1'h0):(1'h0)]);
                      reg7195 <= ($signed((~&$unsigned(reg7119))) ?
                          (((|reg7136) ?
                                  (~|reg4438) : forvar7181[(2'h3):(1'h1)]) ?
                              {(reg4524 || reg4478)} : ((forvar7123 | reg4348) << reg7021[(4'h9):(1'h0)])) : (!((8'hae) >= (!(8'ha4)))));
                    end
                  for (forvar7196 = (1'h0); (forvar7196 < (1'h1)); forvar7196 = (forvar7196 + (1'h1)))
                    begin
                      reg7197 <= $signed(reg7134);
                      reg7198 <= $unsigned(forvar4369);
                    end
                end
              else
                begin
                  reg7192 <= $signed($signed(($unsigned(reg7070) + forvar7030)));
                  for (forvar7193 = (1'h0); (forvar7193 < (2'h2)); forvar7193 = (forvar7193 + (1'h1)))
                    begin
                      reg7194 <= wire7008[(1'h1):(1'h0)];
                      reg7195 <= reg4444[(3'h6):(3'h6)];
                      reg7196 <= (~|{reg4354[(1'h1):(1'h1)]});
                    end
                  if (($unsigned($signed(reg7096[(4'h9):(3'h6)])) ?
                      (+{$unsigned(reg4427)}) : ({(reg7072 | reg4491)} ?
                          ((reg4569 >= (8'ha4)) ?
                              reg4493 : (+forvar7098)) : $unsigned($signed((8'hb3))))))
                    begin
                      reg7197 <= (~^{forvar4454});
                      reg7198 <= (!(((&forvar4346) && $unsigned(forvar7068)) > reg4356));
                      reg7199 <= (8'hab);
                      reg7200 <= forvar7054[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg7197 <= $signed((((8'hb1) ?
                          (reg4524 ?
                              reg7086 : forvar7044) : $signed(reg7096)) ^~ (~&(reg7142 ?
                          reg7044 : (8'ha9)))));
                      reg7198 <= {$signed(reg7144)};
                      reg7199 <= ($signed(((reg7060 ? wire7009 : reg4410) ?
                              (^reg4523) : ((8'ha9) ? reg4537 : wire4340))) ?
                          $signed(forvar4346[(3'h7):(1'h0)]) : reg4434);
                    end
                end
              if ($unsigned(forvar7023))
                begin
                  reg7201 <= (-$signed({(&reg4379)}));
                  if (((forvar4504 >= $signed((reg4409 ?
                          (8'hab) : forvar7148))) ?
                      forvar7079[(2'h2):(1'h0)] : (8'hb2)))
                    begin
                      reg7202 <= $unsigned($signed((~^{reg4511})));
                      reg7203 <= ((($unsigned((8'h9c)) != (reg4358 && (8'ha3))) ?
                          (&reg7058[(4'h8):(4'h8)]) : reg4488) && forvar4476[(4'h9):(4'h8)]);
                    end
                  else
                    begin
                      reg7202 <= ($unsigned((reg4414[(2'h3):(1'h0)] ?
                          (-reg7197) : $unsigned((8'h9d)))) == ($unsigned((forvar4412 * forvar7099)) == {(^~reg4345)}));
                      reg7203 <= ($unsigned(($unsigned(reg7020) ?
                              (reg7158 ? (8'hb1) : reg4469) : forvar7129)) ?
                          {(~$signed(forvar4403))} : (~|(8'ha8)));
                      reg7204 <= ((forvar4554[(1'h0):(1'h0)] ^~ ($unsigned(reg7116) <= $unsigned(reg7133))) ?
                          (8'hac) : (~|reg7093[(4'hb):(3'h4)]));
                      reg7205 <= forvar4389;
                    end
                end
              else
                begin
                  for (forvar7201 = (1'h0); (forvar7201 < (1'h1)); forvar7201 = (forvar7201 + (1'h1)))
                    begin
                      reg7202 <= $signed(reg7064[(1'h0):(1'h0)]);
                      reg7203 <= $unsigned((~&reg7170));
                      reg7204 <= reg4396;
                    end
                  for (forvar7205 = (1'h0); (forvar7205 < (1'h0)); forvar7205 = (forvar7205 + (1'h1)))
                    begin
                      reg7206 <= $unsigned(($signed((reg4369 & reg4432)) >>> reg7140[(3'h5):(1'h1)]));
                    end
                  for (forvar7207 = (1'h0); (forvar7207 < (2'h2)); forvar7207 = (forvar7207 + (1'h1)))
                    begin
                      reg7208 <= $unsigned((-forvar7099[(1'h0):(1'h0)]));
                      reg7209 <= $signed($unsigned((+(forvar4561 ?
                          reg4486 : forvar4427))));
                    end
                  if (((8'hb7) ?
                      (reg7161[(2'h3):(2'h2)] || $unsigned((reg4551 ?
                          reg4442 : reg7151))) : $unsigned((forvar7181 || (~|reg7019)))))
                    begin
                      reg7210 <= {(($unsigned(forvar4344) ?
                              reg7199[(2'h2):(1'h1)] : forvar7149[(1'h1):(1'h1)]) < (~|reg7017[(3'h6):(2'h2)]))};
                      reg7211 <= reg4388;
                      reg7212 <= (~|$signed((-(^reg4428))));
                    end
                  else
                    begin
                      reg7210 <= (~|(reg4422[(4'h8):(1'h1)] ?
                          reg7202 : reg4471));
                      reg7211 <= (+forvar7037);
                    end
                end
              for (forvar7213 = (1'h0); (forvar7213 < (2'h2)); forvar7213 = (forvar7213 + (1'h1)))
                begin
                  for (forvar7214 = (1'h0); (forvar7214 < (1'h0)); forvar7214 = (forvar7214 + (1'h1)))
                    begin
                      reg7215 <= ($unsigned($unsigned($signed((8'hb1)))) ?
                          wire4571 : (-reg7055));
                      reg7216 <= reg4548[(1'h1):(1'h0)];
                      reg7217 <= ($signed((^((8'ha3) ? (8'ha1) : (8'hb9)))) ?
                          forvar7136[(3'h7):(1'h0)] : (reg7098[(3'h4):(1'h1)] >>> ({reg4521} <= reg7056[(1'h0):(1'h0)])));
                      reg7218 <= (({reg7123[(2'h3):(1'h1)]} ?
                              $unsigned((~&reg7179)) : ({forvar4350} || $signed(forvar7040))) ?
                          ((^~(8'ha8)) ?
                              reg7176 : $unsigned((reg4465 ?
                                  reg7105 : reg7215))) : $signed((|reg4421)));
                    end
                  for (forvar7219 = (1'h0); (forvar7219 < (1'h0)); forvar7219 = (forvar7219 + (1'h1)))
                    begin
                      reg7220 <= forvar4422;
                      reg7221 <= $signed($signed(($unsigned(forvar4464) ?
                          $signed((8'h9c)) : (~^forvar7193))));
                      reg7222 <= ((((reg7046 ? reg7052 : forvar7023) ?
                              (reg4491 > reg7154) : $signed(reg4414)) * reg7154[(3'h5):(1'h0)]) ?
                          (8'hab) : $signed((reg4354 - $signed(forvar7193))));
                    end
                  if ($signed((^~(^(reg7143 ? reg4523 : reg4531)))))
                    begin
                      reg7223 <= $signed((+$unsigned((forvar7219 > reg7126))));
                      reg7224 <= $signed(reg4392);
                      reg7225 <= reg4513;
                    end
                  else
                    begin
                      reg7223 <= (~(~$unsigned({reg4514})));
                      reg7224 <= (|((~&$signed(reg7089)) ?
                          $signed(reg4393) : (8'ha7)));
                      reg7225 <= (forvar4353[(4'h9):(3'h5)] && $unsigned((^~{reg7216})));
                      reg7226 <= (~|{reg7056});
                    end
                end
              for (forvar7227 = (1'h0); (forvar7227 < (2'h2)); forvar7227 = (forvar7227 + (1'h1)))
                begin
                  for (forvar7228 = (1'h0); (forvar7228 < (2'h3)); forvar7228 = (forvar7228 + (1'h1)))
                    begin
                      reg7229 <= reg7016[(1'h0):(1'h0)];
                      reg7230 <= forvar7023;
                      reg7231 <= {(~|((8'h9d) ?
                              (&(8'ha6)) : (reg7218 ~^ forvar7227)))};
                      reg7232 <= $unsigned((|((reg4543 & forvar4527) ?
                          {reg7218} : reg4519)));
                    end
                  if (($signed(({reg7138} != (forvar7098 & (8'ha9)))) > $unsigned($signed($signed(reg7083)))))
                    begin
                      reg7233 <= $signed($signed(reg7173[(3'h4):(1'h0)]));
                      reg7234 <= (~|(({forvar7079} ?
                          reg7165[(1'h0):(1'h0)] : $signed(reg4453)) >= $signed((~^reg4422))));
                    end
                  else
                    begin
                      reg7233 <= reg7107[(4'h8):(3'h6)];
                      reg7234 <= $signed($signed($unsigned((forvar4490 | (8'ha5)))));
                      reg7235 <= $signed(reg4485[(1'h0):(1'h0)]);
                      reg7236 <= reg4417;
                    end
                end
            end
          for (forvar7237 = (1'h0); (forvar7237 < (1'h0)); forvar7237 = (forvar7237 + (1'h1)))
            begin
              for (forvar7238 = (1'h0); (forvar7238 < (2'h2)); forvar7238 = (forvar7238 + (1'h1)))
                begin
                  reg7239 <= (reg7072[(4'h8):(1'h0)] ?
                      reg7133 : $unsigned(wire7008));
                end
            end
        end
      else
        begin
          for (forvar7148 = (1'h0); (forvar7148 < (2'h2)); forvar7148 = (forvar7148 + (1'h1)))
            begin
              if ((({(^(8'hb8))} ?
                  ((reg7172 ? reg4482 : forvar7071) ?
                      reg4347 : {reg4503}) : $unsigned((wire4340 ?
                      reg4390 : reg7060))) && {((reg4516 ?
                      forvar7121 : reg4460) < (~reg7155))}))
                begin
                  for (forvar7149 = (1'h0); (forvar7149 < (1'h0)); forvar7149 = (forvar7149 + (1'h1)))
                    begin
                      reg7150 <= reg4569;
                      reg7151 <= reg4501[(3'h4):(1'h0)];
                      reg7152 <= $unsigned((-($unsigned(reg7100) ?
                          (reg4392 & reg4533) : $signed(forvar4372))));
                      reg7153 <= reg4515[(3'h5):(1'h1)];
                    end
                  for (forvar7154 = (1'h0); (forvar7154 < (1'h0)); forvar7154 = (forvar7154 + (1'h1)))
                    begin
                      reg7155 <= reg4433;
                      reg7156 <= reg4410;
                      reg7157 <= ((($signed(forvar7154) ?
                              (reg7129 ?
                                  forvar7149 : (8'h9d)) : {reg7096}) < (reg7170 ?
                              reg4453 : (-reg4360))) ?
                          (~|(8'hba)) : reg7129[(3'h4):(2'h3)]);
                      reg7158 <= (wire7006[(1'h1):(1'h0)] == reg7028[(1'h1):(1'h1)]);
                    end
                end
              else
                begin
                  reg7149 <= $unsigned((+$signed(reg7161[(3'h4):(3'h4)])));
                  reg7150 <= $unsigned(reg7202[(4'hb):(4'ha)]);
                end
            end
        end
      reg7240 <= ((~^(+$unsigned(reg7147))) ?
          forvar7160 : $unsigned((reg7055[(3'h6):(1'h1)] <= (reg4362 <= forvar4558))));
      for (forvar7241 = (1'h0); (forvar7241 < (2'h3)); forvar7241 = (forvar7241 + (1'h1)))
        begin
          if (reg7187)
            begin
              if ($signed(($signed(forvar7135) >>> ($signed((8'hb2)) * forvar4510))))
                begin
                  if (forvar7227[(4'hb):(4'h8)])
                    begin
                      reg7242 <= (!$unsigned({((8'hb0) <<< reg7061)}));
                      reg7243 <= (~&$unsigned($unsigned(reg7102)));
                      reg7244 <= reg4499[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg7242 <= $signed((((forvar7159 ?
                          forvar4427 : reg4438) - $signed(forvar4501)) < $signed((reg4367 > (8'h9e)))));
                      reg7243 <= ($unsigned({$signed(reg7046)}) ?
                          $unsigned(reg4529) : $signed((reg7046[(3'h7):(3'h5)] ?
                              $signed((8'hab)) : (reg7234 >>> reg7014))));
                    end
                  for (forvar7245 = (1'h0); (forvar7245 < (1'h0)); forvar7245 = (forvar7245 + (1'h1)))
                    begin
                      reg7246 <= $signed((+reg7131[(4'he):(4'h8)]));
                      reg7247 <= {reg4350[(1'h1):(1'h0)]};
                    end
                  if (reg7233[(3'h5):(2'h2)])
                    begin
                      reg7248 <= reg7179;
                    end
                  else
                    begin
                      reg7248 <= (reg7088[(2'h3):(2'h3)] ?
                          (reg7168 * reg4443[(2'h2):(2'h2)]) : (reg7115 ?
                              (reg7031[(2'h3):(1'h0)] > reg4399) : reg7222));
                    end
                  for (forvar7249 = (1'h0); (forvar7249 < (2'h2)); forvar7249 = (forvar7249 + (1'h1)))
                    begin
                      reg7250 <= (($unsigned((reg7157 && reg7177)) >>> $unsigned(forvar7047[(2'h3):(1'h0)])) <<< ((|$unsigned(reg7100)) ?
                          (reg4493 ?
                              reg7106[(3'h5):(1'h0)] : reg7199[(4'ha):(3'h5)]) : forvar4459));
                      reg7251 <= $unsigned(((~^(~reg7042)) >> $signed((~reg4422))));
                      reg7252 <= (|$unsigned($unsigned($unsigned(reg4373))));
                    end
                end
              else
                begin
                  for (forvar7242 = (1'h0); (forvar7242 < (2'h2)); forvar7242 = (forvar7242 + (1'h1)))
                    begin
                      reg7243 <= (&$signed((((8'hb6) ?
                          forvar4504 : reg7140) > reg4543[(1'h1):(1'h1)])));
                      reg7244 <= forvar7118[(1'h1):(1'h0)];
                      reg7245 <= forvar7132;
                      reg7246 <= $unsigned(reg4536[(3'h6):(2'h3)]);
                    end
                  if (forvar7149)
                    begin
                      reg7247 <= (-(-(reg7206 << $signed((8'hb8)))));
                      reg7248 <= (!{{(forvar4504 && reg7046)}});
                      reg7249 <= $unsigned((8'ha6));
                    end
                  else
                    begin
                      reg7247 <= (+((reg7147[(3'h7):(1'h1)] <<< (forvar7138 ?
                          reg7230 : reg7100)) < (~|$unsigned(forvar7130))));
                      reg7248 <= (8'hb0);
                    end
                end
              for (forvar7253 = (1'h0); (forvar7253 < (2'h2)); forvar7253 = (forvar7253 + (1'h1)))
                begin
                  for (forvar7254 = (1'h0); (forvar7254 < (1'h0)); forvar7254 = (forvar7254 + (1'h1)))
                    begin
                      reg7255 <= (8'hb1);
                      reg7256 <= forvar7139;
                      reg7257 <= ($unsigned(forvar7104) ?
                          ((~&$unsigned(reg4499)) ?
                              reg7202 : $signed((forvar7111 ?
                                  (8'had) : reg4409))) : reg7193);
                    end
                end
            end
          else
            begin
              for (forvar7242 = (1'h0); (forvar7242 < (2'h3)); forvar7242 = (forvar7242 + (1'h1)))
                begin
                  if ((8'ha2))
                    begin
                      reg7243 <= (^~($unsigned(forvar7153) ?
                          forvar7098 : $signed(reg7164)));
                      reg7244 <= (8'hb9);
                    end
                  else
                    begin
                      reg7243 <= reg7106[(2'h2):(2'h2)];
                    end
                  if (reg7091)
                    begin
                      reg7245 <= reg4489;
                    end
                  else
                    begin
                      reg7245 <= wire4338;
                      reg7246 <= $unsigned($signed($signed((reg7016 ?
                          reg7245 : reg4398))));
                      reg7247 <= forvar4374;
                      reg7248 <= reg7230[(3'h6):(3'h5)];
                    end
                end
              if (((reg7205[(4'ha):(1'h0)] >>> ($unsigned((8'ha5)) ^ (reg4536 << reg4359))) ?
                  (8'hb7) : {reg4537[(2'h2):(1'h1)]}))
                begin
                  for (forvar7249 = (1'h0); (forvar7249 < (1'h1)); forvar7249 = (forvar7249 + (1'h1)))
                    begin
                      reg7250 <= (((forvar7181[(2'h2):(2'h2)] ?
                              $unsigned(reg4481) : (reg7055 ?
                                  reg4489 : reg4483)) ?
                          ((reg7093 ? forvar4568 : reg4565) ?
                              (reg4533 ?
                                  forvar7150 : reg7044) : forvar7079) : $unsigned(reg7042[(2'h2):(2'h2)])) << $signed($signed((^forvar7116))));
                      reg7251 <= $signed($unsigned($unsigned((reg4559 ?
                          reg4525 : forvar7112))));
                      reg7252 <= (&$signed((reg4465 ? (8'hb7) : {(8'ha0)})));
                    end
                end
              else
                begin
                  for (forvar7249 = (1'h0); (forvar7249 < (2'h2)); forvar7249 = (forvar7249 + (1'h1)))
                    begin
                      reg7250 <= $signed($signed(({reg7162} ^~ reg7030)));
                      reg7251 <= reg4491[(1'h0):(1'h0)];
                    end
                end
              if (reg4421[(4'ha):(3'h7)])
                begin
                  if ((~(reg4517 ? reg4487 : forvar4414[(1'h1):(1'h1)])))
                    begin
                      reg7253 <= ($signed($unsigned((~reg7141))) ?
                          (reg7062 <= (8'ha1)) : {reg7032[(3'h4):(1'h1)]});
                      reg7254 <= reg4386[(4'h8):(3'h4)];
                      reg7255 <= (8'ha4);
                      reg7256 <= $unsigned(((^~$signed(reg4543)) || reg4412[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg7253 <= reg4466;
                    end
                  for (forvar7257 = (1'h0); (forvar7257 < (2'h2)); forvar7257 = (forvar7257 + (1'h1)))
                    begin
                      reg7258 <= {$signed(((~|reg7101) ?
                              {reg7217} : (reg7017 ^ forvar7153)))};
                    end
                end
              else
                begin
                  for (forvar7253 = (1'h0); (forvar7253 < (2'h3)); forvar7253 = (forvar7253 + (1'h1)))
                    begin
                      reg7254 <= reg7136;
                      reg7255 <= {{reg7248}};
                      reg7256 <= reg4492[(2'h2):(1'h1)];
                    end
                  reg7257 <= $unsigned(reg7103[(4'h8):(3'h5)]);
                  if (reg4386[(1'h0):(1'h0)])
                    begin
                      reg7258 <= (8'hac);
                    end
                  else
                    begin
                      reg7258 <= $unsigned(((8'hb4) ?
                          ($signed(forvar4422) >>> (reg4540 == reg4429)) : $signed(reg7102[(2'h3):(1'h1)])));
                      reg7259 <= reg4549;
                    end
                end
            end
          for (forvar7260 = (1'h0); (forvar7260 < (1'h1)); forvar7260 = (forvar7260 + (1'h1)))
            begin
              for (forvar7261 = (1'h0); (forvar7261 < (2'h2)); forvar7261 = (forvar7261 + (1'h1)))
                begin
                  if ((~^$signed(forvar7170)))
                    begin
                      reg7262 <= (!((|(!forvar7098)) >>> {(reg7070 + reg4505)}));
                    end
                  else
                    begin
                      reg7262 <= reg4524;
                      reg7263 <= (+reg4433[(2'h3):(1'h1)]);
                    end
                  reg7264 <= {forvar4518};
                  if ((reg4354[(4'hd):(1'h0)] || {reg7061}))
                    begin
                      reg7265 <= reg7200[(2'h2):(2'h2)];
                      reg7266 <= forvar7241[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg7265 <= ((~^reg7198[(1'h0):(1'h0)]) != $signed($unsigned(forvar4500[(4'h8):(2'h2)])));
                      reg7266 <= $unsigned((forvar4542[(1'h1):(1'h1)] == ($signed(forvar7087) || reg7138)));
                      reg7267 <= reg7100[(2'h2):(1'h0)];
                    end
                  if ((reg7200[(2'h2):(2'h2)] ? reg4365 : {(8'ha2)}))
                    begin
                      reg7268 <= ((~&$unsigned(forvar4368)) + ($signed((^reg7172)) ?
                          (reg7151[(4'hd):(3'h6)] ?
                              (^reg7120) : reg4450) : forvar4467[(3'h7):(3'h4)]));
                      reg7269 <= reg7234[(2'h2):(2'h2)];
                      reg7270 <= $signed(($unsigned((+reg4444)) ?
                          reg7121[(4'h8):(1'h0)] : {reg4406[(1'h0):(1'h0)]}));
                      reg7271 <= {(8'ha2)};
                    end
                  else
                    begin
                      reg7268 <= reg4510[(1'h0):(1'h0)];
                      reg7269 <= ({((|reg7127) ?
                              (~^(8'h9c)) : {reg7131})} ^ (reg4375 << {$signed(reg7111)}));
                      reg7270 <= (+$signed((reg4508[(4'he):(2'h2)] ?
                          $unsigned(reg4511) : forvar7136)));
                    end
                end
              reg7272 <= (reg7045 ?
                  $signed(reg7184[(3'h7):(1'h0)]) : $signed((^(^~reg4539))));
              for (forvar7273 = (1'h0); (forvar7273 < (2'h3)); forvar7273 = (forvar7273 + (1'h1)))
                begin
                  reg7274 <= {(!reg7119)};
                  if (reg7026[(1'h0):(1'h0)])
                    begin
                      reg7275 <= {$signed($signed(((8'haf) <= (8'hb1))))};
                      reg7276 <= (^~(!reg7193));
                    end
                  else
                    begin
                      reg7275 <= forvar4364[(4'hc):(4'hc)];
                      reg7276 <= reg7184[(4'h9):(3'h4)];
                    end
                  if ($unsigned(reg4510))
                    begin
                      reg7277 <= ((forvar7237[(3'h7):(3'h6)] ?
                              forvar7260 : (-$unsigned(reg7083))) ?
                          $signed((+reg4466)) : (((^~(8'hb8)) ?
                                  $signed(reg4371) : (reg7073 == reg4407)) ?
                              reg4566[(3'h4):(1'h1)] : (~|(-reg4447))));
                      reg7278 <= ($unsigned((&reg4505[(4'hb):(2'h2)])) ^~ $unsigned((((8'hb7) ?
                              forvar4345 : reg4500) ?
                          reg4466 : forvar7103)));
                    end
                  else
                    begin
                      reg7277 <= reg7015;
                      reg7278 <= (reg4460 ^ $signed(forvar7033[(1'h0):(1'h0)]));
                    end
                end
            end
          for (forvar7279 = (1'h0); (forvar7279 < (1'h0)); forvar7279 = (forvar7279 + (1'h1)))
            begin
              for (forvar7280 = (1'h0); (forvar7280 < (2'h2)); forvar7280 = (forvar7280 + (1'h1)))
                begin
                  for (forvar7281 = (1'h0); (forvar7281 < (1'h1)); forvar7281 = (forvar7281 + (1'h1)))
                    begin
                      reg7282 <= $unsigned($signed(((reg4366 ?
                              reg7070 : reg4423) ?
                          reg4526[(2'h3):(2'h3)] : (reg7212 ?
                              forvar7010 : reg7135))));
                    end
                  if ((($unsigned(reg7052) ?
                          $signed($unsigned(reg4470)) : ((8'hb0) * (reg7132 <= reg7211))) ?
                      (($unsigned(reg7099) << $signed(reg4484)) ?
                          (~$signed((8'h9d))) : (reg4350[(2'h2):(1'h1)] ?
                              (reg7065 ?
                                  reg7230 : reg4504) : (reg4532 || forvar7139))) : ($signed((reg7099 != reg4388)) || forvar7241)))
                    begin
                      reg7283 <= reg4431;
                      reg7284 <= (({(~forvar4456)} ?
                          $signed(reg4494) : ((~^forvar7193) ?
                              forvar7149 : ((8'ha7) ?
                                  reg4450 : (8'hb6)))) || ({((8'ha3) <= reg4348)} >= $signed(forvar4386)));
                    end
                  else
                    begin
                      reg7283 <= (!$signed((|(forvar4568 ?
                          reg7050 : forvar4553))));
                      reg7284 <= (+{reg7120});
                    end
                end
              if ($signed((reg7057[(3'h4):(2'h3)] ?
                  ((+reg7102) >= (&reg4521)) : (|reg4390))))
                begin
                  for (forvar7285 = (1'h0); (forvar7285 < (2'h2)); forvar7285 = (forvar7285 + (1'h1)))
                    begin
                      reg7286 <= ({(|(forvar4547 + reg7113))} > (reg7028[(1'h1):(1'h0)] ?
                          ((|forvar4464) <= (forvar4530 | forvar4391)) : {reg7113}));
                    end
                  for (forvar7287 = (1'h0); (forvar7287 < (1'h0)); forvar7287 = (forvar7287 + (1'h1)))
                    begin
                      reg7288 <= reg4516[(2'h3):(1'h0)];
                      reg7289 <= forvar4530[(2'h2):(1'h0)];
                    end
                  for (forvar7290 = (1'h0); (forvar7290 < (2'h2)); forvar7290 = (forvar7290 + (1'h1)))
                    begin
                      reg7291 <= $unsigned({((&reg4413) ?
                              forvar7193 : $unsigned(reg7149))});
                      reg7292 <= reg4490;
                      reg7293 <= $signed(reg4358);
                      reg7294 <= (|{reg4345[(4'ha):(2'h3)]});
                    end
                end
              else
                begin
                  for (forvar7285 = (1'h0); (forvar7285 < (1'h0)); forvar7285 = (forvar7285 + (1'h1)))
                    begin
                      reg7286 <= ({forvar7285} << $signed({(^~reg7094)}));
                      reg7287 <= (8'ha7);
                      reg7288 <= (&forvar7121[(4'he):(1'h1)]);
                      reg7289 <= (~^forvar4500[(2'h3):(2'h3)]);
                    end
                  for (forvar7290 = (1'h0); (forvar7290 < (1'h1)); forvar7290 = (forvar7290 + (1'h1)))
                    begin
                      reg7291 <= $signed((~((|reg7193) ^ reg4351)));
                    end
                  reg7292 <= $signed($unsigned(($unsigned(reg4354) ?
                      forvar7213[(2'h2):(1'h1)] : (reg4410 ?
                          reg7028 : (8'hac)))));
                  for (forvar7293 = (1'h0); (forvar7293 < (2'h2)); forvar7293 = (forvar7293 + (1'h1)))
                    begin
                      reg7294 <= reg4506[(4'h8):(2'h3)];
                    end
                end
            end
          for (forvar7295 = (1'h0); (forvar7295 < (2'h2)); forvar7295 = (forvar7295 + (1'h1)))
            begin
              reg7296 <= $unsigned((&forvar7207));
              if ($signed($signed($unsigned($signed(reg4417)))))
                begin
                  for (forvar7297 = (1'h0); (forvar7297 < (1'h1)); forvar7297 = (forvar7297 + (1'h1)))
                    begin
                      reg7298 <= $signed((&($signed(reg4474) | $unsigned(reg7053))));
                    end
                  reg7299 <= ((&$unsigned($unsigned(reg4363))) * $signed(forvar4456[(2'h3):(1'h0)]));
                  for (forvar7300 = (1'h0); (forvar7300 < (1'h1)); forvar7300 = (forvar7300 + (1'h1)))
                    begin
                      reg7301 <= $signed($signed((|$unsigned(reg4371))));
                    end
                  for (forvar7302 = (1'h0); (forvar7302 < (2'h2)); forvar7302 = (forvar7302 + (1'h1)))
                    begin
                      reg7303 <= (~&$signed($signed($signed(reg4418))));
                      reg7304 <= ((^forvar4418[(1'h1):(1'h1)]) ^~ (((~&forvar4414) > (forvar7207 ^~ forvar7093)) ?
                          ((reg4563 ?
                              reg7115 : forvar4408) & reg4362[(4'ha):(3'h5)]) : ((~&(8'hb8)) ?
                              reg4544[(3'h4):(2'h2)] : {reg7045})));
                      reg7305 <= forvar7207[(4'h8):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar7297 = (1'h0); (forvar7297 < (1'h0)); forvar7297 = (forvar7297 + (1'h1)))
                    begin
                      reg7298 <= (!(((+reg7088) + {(8'hb2)}) ?
                          $unsigned((reg4399 ?
                              forvar4518 : forvar7242)) : ((reg4544 == reg7215) ~^ reg4411[(2'h3):(2'h3)])));
                    end
                  for (forvar7299 = (1'h0); (forvar7299 < (1'h0)); forvar7299 = (forvar7299 + (1'h1)))
                    begin
                      reg7300 <= $signed($signed(reg7187));
                      reg7301 <= {$unsigned($signed((reg4491 == forvar7093)))};
                      reg7302 <= ((reg7050 != $unsigned(reg7217)) <<< ((reg4369 <= $signed(forvar7201)) ^~ (&reg7036)));
                      reg7303 <= reg4506;
                    end
                end
              for (forvar7306 = (1'h0); (forvar7306 < (1'h1)); forvar7306 = (forvar7306 + (1'h1)))
                begin
                  for (forvar7307 = (1'h0); (forvar7307 < (2'h3)); forvar7307 = (forvar7307 + (1'h1)))
                    begin
                      reg7308 <= reg7236;
                      reg7309 <= forvar7281[(3'h5):(1'h0)];
                      reg7310 <= (~(~^($unsigned(reg7078) ?
                          {forvar4437} : $unsigned(forvar7120))));
                    end
                  for (forvar7311 = (1'h0); (forvar7311 < (1'h0)); forvar7311 = (forvar7311 + (1'h1)))
                    begin
                      reg7312 <= (8'ha5);
                      reg7313 <= $unsigned(forvar7143);
                      reg7314 <= $unsigned(forvar7159[(1'h0):(1'h0)]);
                    end
                end
              for (forvar7315 = (1'h0); (forvar7315 < (1'h0)); forvar7315 = (forvar7315 + (1'h1)))
                begin
                  if (reg4411)
                    begin
                      reg7316 <= forvar4520[(1'h1):(1'h0)];
                      reg7317 <= reg7226[(1'h0):(1'h0)];
                      reg7318 <= reg4373;
                    end
                  else
                    begin
                      reg7316 <= $signed({(8'hb0)});
                      reg7317 <= $unsigned({((-reg7284) ?
                              reg4378 : (reg7185 ? reg7236 : forvar7260))});
                      reg7318 <= reg7016[(2'h2):(1'h0)];
                      reg7319 <= ($unsigned(forvar4414) ?
                          $unsigned((((8'hb2) ~^ forvar7116) ?
                              $unsigned(reg4560) : (reg4480 ^ reg7212))) : $signed((^~reg7119[(2'h2):(2'h2)])));
                    end
                  for (forvar7320 = (1'h0); (forvar7320 < (2'h2)); forvar7320 = (forvar7320 + (1'h1)))
                    begin
                      reg7321 <= reg7066[(2'h2):(1'h0)];
                      reg7322 <= {(+(^~(reg4452 < forvar7191)))};
                      reg7323 <= (8'h9f);
                      reg7324 <= (forvar7306[(3'h4):(2'h3)] ?
                          $signed(forvar7115) : forvar4401);
                    end
                  if ((reg7178[(1'h0):(1'h0)] >>> $unsigned($signed(reg4446))))
                    begin
                      reg7325 <= (forvar7134[(1'h0):(1'h0)] ?
                          $unsigned(($unsigned(reg7223) >> {reg4445})) : $signed(reg7072));
                      reg7326 <= reg7323[(4'h8):(1'h0)];
                      reg7327 <= (&($unsigned((reg4562 ?
                          reg4552 : (8'h9d))) < reg4514));
                      reg7328 <= $unsigned($unsigned(({reg7097} ?
                          $unsigned(reg7030) : ((8'haf) ? (8'hac) : (8'hb7)))));
                    end
                  else
                    begin
                      reg7325 <= (reg7328 >> $unsigned(reg4499));
                      reg7326 <= $unsigned(reg7038[(3'h5):(1'h0)]);
                      reg7327 <= {({$unsigned(reg4523)} < reg7246[(1'h0):(1'h0)])};
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg7329 <= ((((reg4432 ~^ reg7289) ?
              $signed(reg4430) : reg7050[(3'h5):(1'h1)]) != (reg7050[(1'h0):(1'h0)] | ((8'ha0) ?
              reg4534 : reg4550))) ?
          {forvar4546[(4'h9):(3'h7)]} : reg7053);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module888  (y, clk, wire889, wire890, wire891, wire892, wire893);
  output wire [(32'he34):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire889;
  input wire [(5'h10):(1'h0)] wire890;
  input wire signed [(3'h5):(1'h0)] wire891;
  input wire signed [(2'h3):(1'h0)] wire892;
  input wire signed [(4'ha):(1'h0)] wire893;
  wire [(4'he):(1'h0)] wire4168;
  wire [(4'hf):(1'h0)] wire4167;
  wire [(3'h5):(1'h0)] wire4165;
  wire [(2'h3):(1'h0)] wire1758;
  reg [(3'h5):(1'h0)] reg1757 = (1'h0);
  reg [(3'h5):(1'h0)] reg1756 = (1'h0);
  reg [(4'hb):(1'h0)] reg1755 = (1'h0);
  reg [(2'h2):(1'h0)] reg1754 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1753 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1752 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1751 = (1'h0);
  reg [(4'h9):(1'h0)] reg1750 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1749 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1748 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1747 = (1'h0);
  wire [(4'hb):(1'h0)] wire1746;
  wire signed [(4'h8):(1'h0)] wire894;
  wire [(4'h9):(1'h0)] wire895;
  wire [(4'hd):(1'h0)] wire896;
  reg signed [(4'he):(1'h0)] forvar897 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar898 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg899 = (1'h0);
  reg [(4'hf):(1'h0)] reg900 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg901 = (1'h0);
  reg [(4'he):(1'h0)] forvar902 = (1'h0);
  reg [(3'h7):(1'h0)] reg903 = (1'h0);
  reg [(4'hb):(1'h0)] reg904 = (1'h0);
  reg [(3'h6):(1'h0)] reg905 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg906 = (1'h0);
  reg [(3'h7):(1'h0)] reg907 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg908 = (1'h0);
  reg [(2'h2):(1'h0)] reg909 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar910 = (1'h0);
  reg [(2'h2):(1'h0)] reg911 = (1'h0);
  reg [(3'h6):(1'h0)] reg912 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg910 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg913 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg914 = (1'h0);
  reg [(4'he):(1'h0)] reg915 = (1'h0);
  reg [(4'hd):(1'h0)] reg916 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg897 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar900 = (1'h0);
  reg [(4'hd):(1'h0)] reg902 = (1'h0);
  reg [(4'h8):(1'h0)] forvar908 = (1'h0);
  reg [(4'hb):(1'h0)] forvar909 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg917 = (1'h0);
  reg [(3'h4):(1'h0)] forvar917 = (1'h0);
  reg [(4'he):(1'h0)] reg918 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar919 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar920 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg921 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg922 = (1'h0);
  reg [(4'hb):(1'h0)] reg923 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg924 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg919 = (1'h0);
  reg [(4'hb):(1'h0)] reg920 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar921 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg926 = (1'h0);
  reg [(3'h7):(1'h0)] reg927 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg928 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar929 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar930 = (1'h0);
  reg [(4'he):(1'h0)] reg931 = (1'h0);
  reg [(4'hb):(1'h0)] reg932 = (1'h0);
  reg [(4'hd):(1'h0)] reg933 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg934 = (1'h0);
  reg [(4'hb):(1'h0)] reg935 = (1'h0);
  reg [(3'h6):(1'h0)] reg936 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg937 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar938 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg939 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg940 = (1'h0);
  reg [(3'h4):(1'h0)] forvar941 = (1'h0);
  reg [(4'hc):(1'h0)] forvar942 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg943 = (1'h0);
  reg [(4'he):(1'h0)] reg944 = (1'h0);
  reg [(4'h8):(1'h0)] reg945 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg946 = (1'h0);
  reg [(4'he):(1'h0)] reg947 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar918 = (1'h0);
  reg [(3'h4):(1'h0)] forvar923 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar932 = (1'h0);
  reg signed [(4'he):(1'h0)] reg938 = (1'h0);
  reg [(4'h9):(1'h0)] reg941 = (1'h0);
  reg signed [(4'he):(1'h0)] reg942 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar946 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg948 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg949 = (1'h0);
  reg [(2'h3):(1'h0)] reg950 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar951 = (1'h0);
  reg [(4'hf):(1'h0)] reg952 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar953 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg954 = (1'h0);
  reg [(4'ha):(1'h0)] reg955 = (1'h0);
  reg [(4'hb):(1'h0)] reg956 = (1'h0);
  reg [(4'he):(1'h0)] reg957 = (1'h0);
  reg [(3'h6):(1'h0)] reg958 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg959 = (1'h0);
  reg [(4'hf):(1'h0)] forvar960 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg961 = (1'h0);
  reg [(3'h4):(1'h0)] reg951 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar952 = (1'h0);
  reg [(3'h7):(1'h0)] reg953 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar962 = (1'h0);
  reg [(4'hd):(1'h0)] forvar963 = (1'h0);
  reg [(3'h5):(1'h0)] reg964 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg965 = (1'h0);
  reg [(4'hf):(1'h0)] reg966 = (1'h0);
  reg [(3'h6):(1'h0)] forvar967 = (1'h0);
  reg [(4'hf):(1'h0)] reg968 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar955 = (1'h0);
  reg [(4'h8):(1'h0)] reg960 = (1'h0);
  reg [(4'hf):(1'h0)] forvar958 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg963 = (1'h0);
  reg [(4'hc):(1'h0)] forvar964 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg967 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg969 = (1'h0);
  reg signed [(4'he):(1'h0)] reg970 = (1'h0);
  reg [(3'h6):(1'h0)] reg971 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar971 = (1'h0);
  reg [(4'hb):(1'h0)] reg972 = (1'h0);
  reg [(4'hd):(1'h0)] reg973 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar974 = (1'h0);
  reg [(4'hd):(1'h0)] reg975 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg976 = (1'h0);
  reg [(2'h2):(1'h0)] reg977 = (1'h0);
  reg [(3'h6):(1'h0)] forvar978 = (1'h0);
  reg [(4'hf):(1'h0)] reg979 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg980 = (1'h0);
  reg [(4'hd):(1'h0)] reg978 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar981 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg982 = (1'h0);
  reg [(4'hc):(1'h0)] reg983 = (1'h0);
  reg [(4'hb):(1'h0)] reg984 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg985 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg981 = (1'h0);
  reg [(3'h6):(1'h0)] forvar986 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg987 = (1'h0);
  reg [(3'h5):(1'h0)] reg988 = (1'h0);
  reg [(4'ha):(1'h0)] reg989 = (1'h0);
  reg [(3'h6):(1'h0)] reg990 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg986 = (1'h0);
  reg [(4'hc):(1'h0)] forvar987 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg991 = (1'h0);
  reg [(3'h5):(1'h0)] forvar982 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar984 = (1'h0);
  reg [(4'hf):(1'h0)] forvar992 = (1'h0);
  reg [(3'h4):(1'h0)] forvar993 = (1'h0);
  reg [(4'hd):(1'h0)] reg994 = (1'h0);
  reg [(3'h7):(1'h0)] reg995 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg996 = (1'h0);
  reg [(5'h10):(1'h0)] reg997 = (1'h0);
  reg [(4'hd):(1'h0)] forvar998 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg999 = (1'h0);
  reg [(3'h5):(1'h0)] reg1000 = (1'h0);
  wire [(3'h6):(1'h0)] wire1018;
  reg signed [(4'h9):(1'h0)] forvar1020 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1021 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1022 = (1'h0);
  reg [(3'h7):(1'h0)] reg1023 = (1'h0);
  reg [(3'h6):(1'h0)] reg1024 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1025 = (1'h0);
  reg [(4'h9):(1'h0)] reg1026 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1027 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1028 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1029 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1030 = (1'h0);
  reg [(4'hd):(1'h0)] reg1031 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1032 = (1'h0);
  reg [(2'h3):(1'h0)] reg1033 = (1'h0);
  reg [(3'h4):(1'h0)] reg1034 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1035 = (1'h0);
  reg [(2'h2):(1'h0)] reg1036 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1037 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1038 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1039 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1040 = (1'h0);
  reg [(5'h10):(1'h0)] reg1041 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1042 = (1'h0);
  reg [(4'hb):(1'h0)] reg1043 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1044 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1045 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1046 = (1'h0);
  reg [(4'hd):(1'h0)] reg1022 = (1'h0);
  reg [(4'h8):(1'h0)] reg1028 = (1'h0);
  reg [(4'hf):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1030 = (1'h0);
  reg [(3'h6):(1'h0)] reg1032 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1033 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1036 = (1'h0);
  reg [(4'h8):(1'h0)] reg1037 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1040 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1044 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1047 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1048 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1049 = (1'h0);
  reg [(4'h9):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1051 = (1'h0);
  reg [(4'hc):(1'h0)] reg1052 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1053 = (1'h0);
  reg [(4'he):(1'h0)] forvar1054 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1055 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1056 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1057 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1058 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1059 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1060 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1061 = (1'h0);
  reg [(3'h6):(1'h0)] reg1062 = (1'h0);
  reg [(4'hc):(1'h0)] reg1063 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1064 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1065 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1066 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1067 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1068 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1069 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1070 = (1'h0);
  reg [(4'hd):(1'h0)] reg1071 = (1'h0);
  reg [(3'h7):(1'h0)] reg1072 = (1'h0);
  reg [(4'ha):(1'h0)] reg1060 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1065 = (1'h0);
  reg [(3'h5):(1'h0)] reg1073 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1074 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1075 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1076 = (1'h0);
  reg [(4'h8):(1'h0)] reg1077 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1078 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1079 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1080 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1081 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1082 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1083 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1084 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1085 = (1'h0);
  reg [(4'ha):(1'h0)] reg1086 = (1'h0);
  reg [(4'h8):(1'h0)] reg1087 = (1'h0);
  reg [(4'he):(1'h0)] reg1088 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1089 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1090 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1091 = (1'h0);
  reg [(4'h8):(1'h0)] reg1092 = (1'h0);
  reg [(4'he):(1'h0)] reg1093 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1094 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1095 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1096 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1097 = (1'h0);
  reg [(3'h7):(1'h0)] reg1098 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1099 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1100 = (1'h0);
  reg [(4'he):(1'h0)] reg1101 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1102 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1103 = (1'h0);
  reg [(2'h3):(1'h0)] reg1104 = (1'h0);
  reg [(3'h4):(1'h0)] reg1105 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1106 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1107 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1108 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1109 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1110 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1111 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1112 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1113 = (1'h0);
  reg [(4'hd):(1'h0)] reg1103 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1104 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1107 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1108 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1109 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1112 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1114 = (1'h0);
  reg [(4'hd):(1'h0)] reg1115 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1116 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1117 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1118 = (1'h0);
  reg [(4'h9):(1'h0)] reg1119 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1120 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1121 = (1'h0);
  reg [(5'h10):(1'h0)] reg1122 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1123 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1124 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1078 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1125 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1126 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1127 = (1'h0);
  reg [(5'h10):(1'h0)] reg1128 = (1'h0);
  reg [(4'hb):(1'h0)] reg1129 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1130 = (1'h0);
  reg [(5'h10):(1'h0)] reg1131 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1132 = (1'h0);
  reg [(2'h3):(1'h0)] reg1133 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1134 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1135 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1136 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1137 = (1'h0);
  reg [(5'h10):(1'h0)] reg1127 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1130 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1138 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1139 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1140 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1141 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1142 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1143 = (1'h0);
  reg [(4'ha):(1'h0)] reg1144 = (1'h0);
  reg [(4'he):(1'h0)] forvar1145 = (1'h0);
  reg [(2'h2):(1'h0)] reg1146 = (1'h0);
  reg [(5'h10):(1'h0)] reg1143 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1147 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1148 = (1'h0);
  reg [(4'he):(1'h0)] reg1149 = (1'h0);
  reg [(3'h4):(1'h0)] reg1150 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1151 = (1'h0);
  reg [(3'h7):(1'h0)] reg1152 = (1'h0);
  reg [(4'h9):(1'h0)] reg1153 = (1'h0);
  reg [(3'h7):(1'h0)] reg1154 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1155 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1156 = (1'h0);
  reg [(4'hc):(1'h0)] reg1157 = (1'h0);
  reg [(4'ha):(1'h0)] reg1158 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1159 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1160 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1161 = (1'h0);
  reg [(4'h9):(1'h0)] reg1162 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1125 = (1'h0);
  reg [(4'ha):(1'h0)] reg1126 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1132 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1138 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1139 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1133 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1141 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1146 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1147 = (1'h0);
  reg [(3'h7):(1'h0)] reg1148 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1155 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1156 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1163 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1164 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1165 = (1'h0);
  reg [(4'h9):(1'h0)] reg1166 = (1'h0);
  reg [(3'h7):(1'h0)] reg1167 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1168 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1169 = (1'h0);
  reg [(4'hb):(1'h0)] reg1170 = (1'h0);
  reg [(4'h8):(1'h0)] reg1171 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1165 = (1'h0);
  reg [(4'hf):(1'h0)] reg1172 = (1'h0);
  reg [(3'h6):(1'h0)] reg1173 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1174 = (1'h0);
  reg [(3'h4):(1'h0)] reg1175 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1176 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1164 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1169 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1177 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1178 = (1'h0);
  reg [(4'hb):(1'h0)] reg1179 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1180 = (1'h0);
  reg [(4'h9):(1'h0)] reg1181 = (1'h0);
  reg [(4'h8):(1'h0)] reg1182 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1183 = (1'h0);
  reg [(4'hd):(1'h0)] reg1184 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1185 = (1'h0);
  reg [(4'h9):(1'h0)] reg1186 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1187 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1188 = (1'h0);
  reg [(4'hc):(1'h0)] reg1189 = (1'h0);
  reg [(4'hd):(1'h0)] reg1190 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1191 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1192 = (1'h0);
  reg [(3'h7):(1'h0)] reg1193 = (1'h0);
  reg [(2'h3):(1'h0)] reg1194 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1195 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1196 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1197 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1198 = (1'h0);
  reg [(4'hd):(1'h0)] reg1199 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1200 = (1'h0);
  reg [(3'h6):(1'h0)] reg1201 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1202 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1203 = (1'h0);
  reg [(3'h7):(1'h0)] reg1204 = (1'h0);
  reg [(3'h6):(1'h0)] reg1205 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1206 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1207 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1208 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1209 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1211 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1212 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1213 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1214 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1215 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1216 = (1'h0);
  reg [(3'h4):(1'h0)] reg1217 = (1'h0);
  wire [(3'h7):(1'h0)] wire1218;
  wire signed [(4'hf):(1'h0)] wire1744;
  assign y = {wire4168,
                 wire4167,
                 wire4165,
                 wire1758,
                 reg1757,
                 reg1756,
                 reg1755,
                 reg1754,
                 reg1753,
                 reg1752,
                 forvar1751,
                 reg1750,
                 forvar1749,
                 forvar1748,
                 forvar1747,
                 wire1746,
                 wire894,
                 wire895,
                 wire896,
                 forvar897,
                 forvar898,
                 reg899,
                 reg900,
                 reg901,
                 forvar902,
                 reg903,
                 reg904,
                 reg905,
                 reg906,
                 reg907,
                 reg908,
                 reg909,
                 forvar910,
                 reg911,
                 reg912,
                 reg910,
                 reg913,
                 reg914,
                 reg915,
                 reg916,
                 reg897,
                 forvar900,
                 reg902,
                 forvar908,
                 forvar909,
                 reg917,
                 forvar917,
                 reg918,
                 forvar919,
                 forvar920,
                 reg921,
                 reg922,
                 reg923,
                 reg924,
                 reg919,
                 reg920,
                 forvar921,
                 reg925,
                 reg926,
                 reg927,
                 reg928,
                 forvar929,
                 forvar930,
                 reg931,
                 reg932,
                 reg933,
                 reg934,
                 reg935,
                 reg936,
                 reg937,
                 forvar938,
                 reg939,
                 reg940,
                 forvar941,
                 forvar942,
                 reg943,
                 reg944,
                 reg945,
                 reg946,
                 reg947,
                 forvar918,
                 forvar923,
                 forvar932,
                 reg938,
                 reg941,
                 reg942,
                 forvar946,
                 reg948,
                 reg949,
                 reg950,
                 forvar951,
                 reg952,
                 forvar953,
                 reg954,
                 reg955,
                 reg956,
                 reg957,
                 reg958,
                 reg959,
                 forvar960,
                 reg961,
                 reg951,
                 forvar952,
                 reg953,
                 forvar962,
                 forvar963,
                 reg964,
                 reg965,
                 reg966,
                 forvar967,
                 reg968,
                 forvar955,
                 reg960,
                 forvar958,
                 reg963,
                 forvar964,
                 reg967,
                 reg969,
                 reg970,
                 reg971,
                 forvar971,
                 reg972,
                 reg973,
                 forvar974,
                 reg975,
                 reg976,
                 reg977,
                 forvar978,
                 reg979,
                 reg980,
                 reg978,
                 forvar981,
                 reg982,
                 reg983,
                 reg984,
                 reg985,
                 reg981,
                 forvar986,
                 reg987,
                 reg988,
                 reg989,
                 reg990,
                 reg986,
                 forvar987,
                 reg991,
                 forvar982,
                 forvar984,
                 forvar992,
                 forvar993,
                 reg994,
                 reg995,
                 reg996,
                 reg997,
                 forvar998,
                 reg999,
                 reg1000,
                 wire1018,
                 forvar1020,
                 forvar1021,
                 forvar1022,
                 reg1023,
                 reg1024,
                 reg1025,
                 reg1026,
                 reg1027,
                 forvar1028,
                 forvar1029,
                 reg1030,
                 reg1031,
                 forvar1032,
                 reg1033,
                 reg1034,
                 reg1035,
                 reg1036,
                 forvar1037,
                 forvar1038,
                 reg1039,
                 forvar1040,
                 reg1041,
                 reg1042,
                 reg1043,
                 reg1044,
                 reg1045,
                 reg1046,
                 reg1022,
                 reg1028,
                 reg1029,
                 forvar1030,
                 reg1032,
                 forvar1033,
                 forvar1036,
                 reg1037,
                 reg1040,
                 forvar1044,
                 forvar1047,
                 forvar1048,
                 forvar1049,
                 reg1050,
                 reg1051,
                 reg1052,
                 reg1053,
                 forvar1054,
                 forvar1055,
                 reg1056,
                 reg1057,
                 reg1058,
                 forvar1059,
                 forvar1060,
                 reg1061,
                 reg1062,
                 reg1063,
                 reg1064,
                 forvar1065,
                 reg1066,
                 reg1067,
                 reg1068,
                 reg1069,
                 reg1070,
                 reg1071,
                 reg1072,
                 reg1060,
                 reg1065,
                 reg1073,
                 forvar1074,
                 forvar1075,
                 reg1076,
                 reg1077,
                 reg1078,
                 reg1079,
                 forvar1080,
                 reg1081,
                 reg1082,
                 reg1083,
                 forvar1084,
                 forvar1085,
                 reg1086,
                 reg1087,
                 reg1088,
                 forvar1089,
                 reg1090,
                 forvar1091,
                 reg1092,
                 reg1093,
                 reg1094,
                 reg1095,
                 reg1096,
                 forvar1097,
                 reg1098,
                 reg1099,
                 reg1100,
                 reg1101,
                 reg1102,
                 forvar1103,
                 reg1104,
                 reg1105,
                 reg1106,
                 reg1107,
                 forvar1108,
                 reg1109,
                 reg1110,
                 reg1111,
                 forvar1112,
                 reg1113,
                 reg1103,
                 forvar1104,
                 forvar1107,
                 reg1108,
                 forvar1109,
                 reg1112,
                 reg1114,
                 reg1115,
                 reg1116,
                 forvar1117,
                 reg1118,
                 reg1119,
                 forvar1120,
                 reg1121,
                 reg1122,
                 reg1123,
                 reg1124,
                 forvar1078,
                 reg1125,
                 forvar1126,
                 forvar1127,
                 reg1128,
                 reg1129,
                 forvar1130,
                 reg1131,
                 reg1132,
                 reg1133,
                 reg1134,
                 reg1135,
                 reg1136,
                 reg1137,
                 reg1127,
                 reg1130,
                 forvar1138,
                 forvar1139,
                 reg1140,
                 forvar1141,
                 reg1142,
                 forvar1143,
                 reg1144,
                 forvar1145,
                 reg1146,
                 reg1143,
                 forvar1147,
                 forvar1148,
                 reg1149,
                 reg1150,
                 reg1151,
                 reg1152,
                 reg1153,
                 reg1154,
                 reg1155,
                 forvar1156,
                 reg1157,
                 reg1158,
                 forvar1159,
                 reg1160,
                 reg1161,
                 reg1162,
                 forvar1125,
                 reg1126,
                 forvar1132,
                 reg1138,
                 reg1139,
                 forvar1133,
                 reg1141,
                 reg1145,
                 forvar1146,
                 reg1147,
                 reg1148,
                 forvar1155,
                 reg1156,
                 forvar1163,
                 reg1164,
                 reg1165,
                 reg1166,
                 reg1167,
                 reg1168,
                 reg1169,
                 reg1170,
                 reg1171,
                 forvar1165,
                 reg1172,
                 reg1173,
                 reg1174,
                 reg1175,
                 reg1176,
                 forvar1164,
                 forvar1169,
                 forvar1177,
                 forvar1178,
                 reg1179,
                 reg1180,
                 reg1181,
                 reg1182,
                 reg1183,
                 reg1184,
                 forvar1185,
                 reg1186,
                 reg1187,
                 reg1188,
                 reg1189,
                 reg1190,
                 reg1191,
                 forvar1192,
                 reg1193,
                 reg1194,
                 reg1195,
                 reg1196,
                 reg1197,
                 reg1198,
                 reg1199,
                 reg1200,
                 reg1201,
                 forvar1202,
                 forvar1203,
                 reg1204,
                 reg1205,
                 reg1206,
                 forvar1207,
                 reg1208,
                 forvar1209,
                 reg1210,
                 reg1211,
                 reg1212,
                 reg1213,
                 reg1214,
                 forvar1215,
                 reg1216,
                 reg1217,
                 wire1218,
                 wire1744,
                 (1'h0)};
  assign wire894 = {$unsigned((&wire890[(2'h3):(2'h2)]))};
  assign wire895 = $signed(((|wire893[(4'h8):(4'h8)]) != {wire891}));
  assign wire896 = wire894[(2'h2):(1'h0)];
  always
    @(posedge clk) begin
      if (wire891[(2'h3):(1'h0)])
        begin
          for (forvar897 = (1'h0); (forvar897 < (2'h3)); forvar897 = (forvar897 + (1'h1)))
            begin
              if (wire896)
                begin
                  for (forvar898 = (1'h0); (forvar898 < (2'h3)); forvar898 = (forvar898 + (1'h1)))
                    begin
                      reg899 <= $signed($signed(({wire895} || (wire890 || forvar898))));
                    end
                end
              else
                begin
                  for (forvar898 = (1'h0); (forvar898 < (1'h1)); forvar898 = (forvar898 + (1'h1)))
                    begin
                      reg899 <= $signed($signed({$unsigned(wire889)}));
                      reg900 <= $unsigned(wire893);
                      reg901 <= (~&$signed(($signed(wire896) ?
                          {wire891} : (wire892 ? wire896 : reg899))));
                    end
                end
              for (forvar902 = (1'h0); (forvar902 < (2'h3)); forvar902 = (forvar902 + (1'h1)))
                begin
                  if (({$unsigned({wire891})} ^~ reg901[(1'h0):(1'h0)]))
                    begin
                      reg903 <= wire896;
                      reg904 <= $signed(($unsigned($unsigned(wire896)) - (wire895 ?
                          (^~wire889) : (wire894 ^~ wire890))));
                    end
                  else
                    begin
                      reg903 <= ((~|$signed($unsigned(reg901))) ~^ $signed({(wire894 ?
                              wire891 : wire891)}));
                    end
                  reg905 <= $unsigned({(~&forvar902)});
                  if (({($signed(forvar897) & (forvar898 ?
                              wire896 : wire893))} ?
                      wire891[(3'h5):(3'h4)] : wire889))
                    begin
                      reg906 <= wire889;
                    end
                  else
                    begin
                      reg906 <= ((reg904[(3'h6):(1'h1)] && wire896[(4'hc):(3'h6)]) ?
                          ($signed(forvar897) ?
                              wire894 : ({wire894} >= $signed(wire889))) : (~(((8'hb3) ?
                                  wire896 : reg904) ?
                              forvar902 : wire893[(3'h4):(1'h1)])));
                      reg907 <= $unsigned(reg906);
                    end
                  reg908 <= ($signed(wire896[(3'h4):(2'h2)]) ?
                      (-wire891[(3'h4):(1'h0)]) : $unsigned(reg903));
                end
              reg909 <= (+(-reg905[(3'h6):(3'h4)]));
              if (($unsigned($signed({forvar902})) * $signed((+(wire894 <<< wire889)))))
                begin
                  for (forvar910 = (1'h0); (forvar910 < (2'h2)); forvar910 = (forvar910 + (1'h1)))
                    begin
                      reg911 <= (reg905 ?
                          (wire894 ?
                              $unsigned((wire889 << reg903)) : $unsigned($signed(wire894))) : {$signed(wire894[(3'h7):(3'h7)])});
                    end
                  if ($unsigned(wire892))
                    begin
                      reg912 <= ((reg900[(1'h0):(1'h0)] ?
                          reg906 : (reg907 != (~&wire890))) | wire890[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg912 <= ((~^wire894[(3'h6):(3'h4)]) ?
                          ((reg909[(1'h0):(1'h0)] >>> (reg912 ?
                              reg906 : forvar902)) + ($unsigned(forvar910) > $unsigned(reg912))) : $unsigned(((wire895 ?
                                  forvar898 : reg912) ?
                              (~|(8'hba)) : reg903)));
                    end
                end
              else
                begin
                  if (($signed(reg899[(4'h9):(1'h0)]) & (^~((reg906 ?
                          reg900 : (8'haa)) ?
                      $signed(wire895) : $signed(forvar898)))))
                    begin
                      reg910 <= (8'haa);
                      reg911 <= ((((8'had) ?
                          (^~wire896) : (forvar898 && wire891)) ^~ $signed(reg901[(2'h2):(1'h0)])) ^~ (forvar902[(1'h0):(1'h0)] != $signed((wire892 << wire891))));
                      reg912 <= forvar898;
                    end
                  else
                    begin
                      reg910 <= (|forvar897);
                    end
                  if ($signed((reg901 | reg912[(3'h4):(1'h0)])))
                    begin
                      reg913 <= wire889[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg913 <= reg912[(1'h0):(1'h0)];
                    end
                  reg914 <= (8'hac);
                end
            end
          reg915 <= $unsigned((wire895[(4'h9):(3'h4)] ^ {$signed(reg912)}));
          reg916 <= ({$unsigned(reg913)} & ($signed((wire890 - forvar898)) + $unsigned((wire893 ?
              reg912 : wire895))));
        end
      else
        begin
          reg897 <= (wire893 ?
              (+(reg903 ^~ (forvar898 < forvar910))) : (({wire895} && (8'hac)) ?
                  ((reg899 ? reg905 : wire889) | (^~reg899)) : wire894));
          for (forvar898 = (1'h0); (forvar898 < (2'h3)); forvar898 = (forvar898 + (1'h1)))
            begin
              reg899 <= $unsigned($signed(({reg912} ?
                  (-wire891) : (~^(8'hba)))));
              if ($signed((|($unsigned(reg913) <<< (wire890 < reg913)))))
                begin
                  for (forvar900 = (1'h0); (forvar900 < (2'h2)); forvar900 = (forvar900 + (1'h1)))
                    begin
                      reg901 <= wire890[(1'h0):(1'h0)];
                    end
                  if ((($signed(reg909[(2'h2):(2'h2)]) == (!(reg897 <= reg915))) ?
                      wire890[(2'h2):(1'h0)] : (+((8'had) ?
                          reg900 : {reg908}))))
                    begin
                      reg902 <= $signed($unsigned(wire890[(1'h0):(1'h0)]));
                      reg903 <= $unsigned(({(~&(8'had))} && (8'hae)));
                      reg904 <= (!(~^$unsigned((|reg907))));
                      reg905 <= {((reg915 >>> (~&wire892)) ?
                              (^~reg909[(1'h0):(1'h0)]) : wire891[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg902 <= {reg914};
                      reg903 <= reg899[(1'h0):(1'h0)];
                    end
                  reg906 <= reg915[(3'h4):(1'h0)];
                end
              else
                begin
                  for (forvar900 = (1'h0); (forvar900 < (1'h1)); forvar900 = (forvar900 + (1'h1)))
                    begin
                      reg901 <= $unsigned({{(-reg897)}});
                      reg902 <= $signed({((reg914 || forvar910) * $signed(reg915))});
                      reg903 <= {$signed((8'ha2))};
                      reg904 <= (reg908[(5'h10):(3'h6)] > {(^~(~&reg902))});
                    end
                  reg905 <= $signed((^~forvar902));
                  if (wire896[(1'h0):(1'h0)])
                    begin
                      reg906 <= $signed(reg901[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg906 <= $signed($signed(reg914));
                      reg907 <= forvar910;
                    end
                end
            end
          for (forvar908 = (1'h0); (forvar908 < (2'h2)); forvar908 = (forvar908 + (1'h1)))
            begin
              if ({($signed(forvar902[(3'h4):(3'h4)]) - reg914[(1'h1):(1'h0)])})
                begin
                  reg909 <= (~|reg899);
                  for (forvar910 = (1'h0); (forvar910 < (1'h1)); forvar910 = (forvar910 + (1'h1)))
                    begin
                      reg911 <= wire890[(3'h5):(2'h3)];
                      reg912 <= (forvar897[(4'he):(3'h6)] ^ $signed(reg899[(4'hb):(3'h5)]));
                      reg913 <= ($signed((~^$signed(forvar902))) ?
                          forvar900 : {$unsigned((wire889 ?
                                  wire892 : (8'hba)))});
                      reg914 <= wire895[(2'h3):(2'h3)];
                    end
                  reg915 <= reg905;
                end
              else
                begin
                  for (forvar909 = (1'h0); (forvar909 < (2'h3)); forvar909 = (forvar909 + (1'h1)))
                    begin
                      reg910 <= ((^$signed(forvar909)) ?
                          {((~^reg900) && (~&reg904))} : reg905[(3'h4):(1'h1)]);
                      reg911 <= $signed({(reg911 >> $signed(reg901))});
                      reg912 <= (|($unsigned($signed(reg913)) ^~ (reg897[(3'h4):(1'h1)] ?
                          $signed((8'ha7)) : $unsigned((8'h9c)))));
                      reg913 <= forvar900;
                    end
                  reg914 <= ($signed($signed((reg909 == forvar898))) * (!((reg908 && wire893) ?
                      $unsigned((8'ha9)) : $signed(forvar902))));
                end
            end
        end
      if ($unsigned((^($signed(reg910) ?
          wire895[(3'h5):(1'h0)] : $signed(reg912)))))
        begin
          if (((^(^(reg909 ? reg897 : reg911))) || $signed({(~&forvar908)})))
            begin
              if (($signed((&$signed(reg913))) <<< reg905))
                begin
                  reg917 <= (((((8'hab) ^~ (8'hb4)) * $signed(reg902)) >>> reg906[(4'hb):(2'h2)]) ?
                      ($signed((reg904 * reg916)) ?
                          (!(^~(8'hab))) : $signed((wire894 - (8'h9f)))) : reg908);
                end
              else
                begin
                  for (forvar917 = (1'h0); (forvar917 < (2'h2)); forvar917 = (forvar917 + (1'h1)))
                    begin
                      reg918 <= (~^reg913);
                    end
                end
              for (forvar919 = (1'h0); (forvar919 < (1'h1)); forvar919 = (forvar919 + (1'h1)))
                begin
                  for (forvar920 = (1'h0); (forvar920 < (1'h0)); forvar920 = (forvar920 + (1'h1)))
                    begin
                      reg921 <= $signed($signed(reg897));
                      reg922 <= reg915[(1'h0):(1'h0)];
                      reg923 <= reg922[(3'h4):(1'h0)];
                      reg924 <= $signed(wire891[(1'h1):(1'h1)]);
                    end
                end
            end
          else
            begin
              if ((8'ha7))
                begin
                  for (forvar917 = (1'h0); (forvar917 < (1'h1)); forvar917 = (forvar917 + (1'h1)))
                    begin
                      reg918 <= ((~reg905[(3'h4):(2'h2)]) ^~ (&(~^forvar908[(4'h8):(2'h2)])));
                      reg919 <= (^~$signed($signed($signed(reg917))));
                    end
                  if ($signed(reg918[(4'he):(4'hd)]))
                    begin
                      reg920 <= (8'hb8);
                      reg921 <= reg902;
                      reg922 <= ((~(+(|reg904))) - reg905[(1'h0):(1'h0)]);
                      reg923 <= ((reg900[(4'hb):(3'h4)] & ((reg916 ?
                              reg913 : reg911) - $signed(reg912))) ?
                          wire891[(3'h4):(2'h3)] : reg924[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg920 <= (&(forvar908 && ($signed(reg921) ?
                          (reg919 ? reg921 : reg921) : (reg920 ?
                              forvar920 : forvar917))));
                      reg921 <= (~^(reg912[(2'h2):(2'h2)] ?
                          {$unsigned(reg916)} : (reg914 ?
                              reg921[(3'h6):(1'h1)] : (8'hac))));
                      reg922 <= (8'hba);
                    end
                end
              else
                begin
                  if (reg908)
                    begin
                      reg917 <= $signed($unsigned(($signed(forvar900) ?
                          wire894 : $unsigned(reg917))));
                      reg918 <= forvar909;
                      reg919 <= $unsigned({forvar919[(2'h3):(1'h0)]});
                      reg920 <= (wire890[(4'hb):(3'h7)] > (reg923[(4'ha):(1'h0)] ?
                          ($signed(reg908) ?
                              (reg918 + reg920) : $signed(reg901)) : $signed($signed(wire896))));
                    end
                  else
                    begin
                      reg917 <= $signed($unsigned(reg906));
                    end
                  for (forvar921 = (1'h0); (forvar921 < (1'h0)); forvar921 = (forvar921 + (1'h1)))
                    begin
                      reg922 <= wire894[(1'h1):(1'h1)];
                      reg923 <= (reg903 ?
                          reg923 : (!$signed($unsigned(reg902))));
                      reg924 <= ((wire893[(2'h2):(1'h1)] + $signed($unsigned((8'ha6)))) ?
                          reg902 : $signed(forvar917));
                    end
                  if (forvar909)
                    begin
                      reg925 <= $signed((~&reg904[(3'h7):(1'h0)]));
                      reg926 <= (($signed(reg906[(4'h9):(4'h8)]) >= ((reg904 ?
                                  reg899 : forvar909) ?
                              (reg901 ?
                                  reg914 : (8'haf)) : $unsigned(reg909))) ?
                          $signed($signed(reg920)) : $signed((~^reg918[(3'h5):(3'h4)])));
                      reg927 <= $signed($signed(($unsigned(reg911) <= {reg915})));
                      reg928 <= (({$unsigned(reg920)} || $signed($unsigned((8'ha7)))) & (~^($unsigned(wire892) ?
                          $unsigned(reg904) : (reg925 ^~ wire889))));
                    end
                  else
                    begin
                      reg925 <= reg897;
                      reg926 <= ((^(-{(8'h9e)})) <= reg905[(3'h6):(3'h5)]);
                      reg927 <= forvar897;
                      reg928 <= forvar920[(2'h2):(1'h1)];
                    end
                end
              for (forvar929 = (1'h0); (forvar929 < (1'h0)); forvar929 = (forvar929 + (1'h1)))
                begin
                  for (forvar930 = (1'h0); (forvar930 < (1'h0)); forvar930 = (forvar930 + (1'h1)))
                    begin
                      reg931 <= $signed(wire892);
                      reg932 <= forvar902;
                      reg933 <= wire894;
                    end
                  if ({{(wire896 + wire895)}})
                    begin
                      reg934 <= $unsigned($signed(((reg924 >> reg933) ?
                          reg918 : (^~reg933))));
                      reg935 <= {(((~^reg901) ? $unsigned((8'had)) : reg920) ?
                              reg897[(3'h7):(3'h6)] : ($signed(reg925) ?
                                  (~^reg900) : {reg928}))};
                      reg936 <= (!(-({reg921} ?
                          forvar920 : wire892[(2'h3):(2'h2)])));
                      reg937 <= (reg924[(1'h1):(1'h0)] ?
                          $signed($unsigned($signed(reg924))) : reg928);
                    end
                  else
                    begin
                      reg934 <= ((|reg915) ?
                          $unsigned(reg915[(4'h8):(4'h8)]) : (reg937[(2'h3):(1'h0)] ^ reg908[(4'h9):(2'h3)]));
                      reg935 <= forvar900[(3'h6):(3'h5)];
                      reg936 <= reg927[(3'h7):(2'h2)];
                      reg937 <= reg923[(3'h5):(3'h4)];
                    end
                  for (forvar938 = (1'h0); (forvar938 < (1'h1)); forvar938 = (forvar938 + (1'h1)))
                    begin
                      reg939 <= (8'ha2);
                      reg940 <= ($signed($unsigned($unsigned((8'hae)))) ~^ reg928);
                    end
                end
              for (forvar941 = (1'h0); (forvar941 < (1'h1)); forvar941 = (forvar941 + (1'h1)))
                begin
                  for (forvar942 = (1'h0); (forvar942 < (2'h2)); forvar942 = (forvar942 + (1'h1)))
                    begin
                      reg943 <= forvar929;
                      reg944 <= (8'h9c);
                      reg945 <= forvar919[(4'hd):(3'h5)];
                      reg946 <= $signed(((^(~wire892)) != (8'ha1)));
                    end
                end
            end
          reg947 <= $signed(((8'ha2) ^ (reg928[(1'h0):(1'h0)] ?
              (forvar938 ? (8'hac) : forvar938) : ((8'hb0) ?
                  (8'hb7) : reg944))));
        end
      else
        begin
          for (forvar917 = (1'h0); (forvar917 < (1'h1)); forvar917 = (forvar917 + (1'h1)))
            begin
              if ($unsigned(forvar900))
                begin
                  for (forvar918 = (1'h0); (forvar918 < (2'h3)); forvar918 = (forvar918 + (1'h1)))
                    begin
                      reg919 <= $unsigned($signed($unsigned((reg900 ?
                          reg946 : reg918))));
                      reg920 <= ((^~reg928) - reg917[(4'hf):(3'h6)]);
                      reg921 <= ($unsigned({reg915}) ?
                          $unsigned({reg915}) : ((~{reg934}) ?
                              $signed($unsigned(reg906)) : ({wire892} ?
                                  (reg908 > reg922) : (reg927 && reg918))));
                      reg922 <= wire894[(2'h2):(1'h0)];
                    end
                  if (($unsigned((8'hb6)) ?
                      reg901[(2'h2):(2'h2)] : $unsigned((|reg901))))
                    begin
                      reg923 <= $unsigned($signed(($unsigned(reg909) || (reg908 ^ reg908))));
                      reg924 <= (~|$unsigned($signed(reg915)));
                      reg925 <= (8'ha5);
                      reg926 <= $unsigned($unsigned((-(|reg911))));
                    end
                  else
                    begin
                      reg923 <= reg916[(3'h6):(3'h6)];
                      reg924 <= wire895[(3'h7):(3'h4)];
                      reg925 <= ($signed($unsigned(forvar902)) || ($unsigned(reg936[(2'h3):(2'h2)]) << reg913));
                      reg926 <= ($unsigned($signed($signed(forvar919))) ?
                          {reg904} : $unsigned(forvar938));
                    end
                  if (reg934[(1'h1):(1'h0)])
                    begin
                      reg927 <= (8'h9d);
                      reg928 <= $unsigned($unsigned((forvar917[(2'h3):(1'h0)] == (reg926 ?
                          (8'hae) : forvar938))));
                    end
                  else
                    begin
                      reg927 <= (+reg906);
                    end
                end
              else
                begin
                  reg918 <= (|(reg911[(1'h1):(1'h1)] ?
                      $unsigned(reg907) : reg927));
                  for (forvar919 = (1'h0); (forvar919 < (1'h1)); forvar919 = (forvar919 + (1'h1)))
                    begin
                      reg920 <= (+reg931);
                      reg921 <= reg931;
                      reg922 <= $unsigned((+(forvar938 ^ wire895[(4'h9):(3'h6)])));
                    end
                  for (forvar923 = (1'h0); (forvar923 < (1'h1)); forvar923 = (forvar923 + (1'h1)))
                    begin
                      reg924 <= (8'ha5);
                      reg925 <= {($unsigned((-wire889)) ?
                              ($unsigned(forvar929) >= {(8'h9c)}) : $signed((8'h9c)))};
                      reg926 <= forvar909;
                      reg927 <= (reg945[(3'h7):(3'h6)] ?
                          $signed(($signed((8'hb6)) ^~ reg910[(3'h4):(1'h0)])) : ((^$unsigned(reg919)) ?
                              $signed(((8'had) ~^ wire889)) : $signed($signed(reg926))));
                    end
                end
              for (forvar929 = (1'h0); (forvar929 < (2'h3)); forvar929 = (forvar929 + (1'h1)))
                begin
                  for (forvar930 = (1'h0); (forvar930 < (2'h2)); forvar930 = (forvar930 + (1'h1)))
                    begin
                      reg931 <= reg927;
                    end
                  for (forvar932 = (1'h0); (forvar932 < (2'h2)); forvar932 = (forvar932 + (1'h1)))
                    begin
                      reg933 <= $signed($signed((&(8'hb5))));
                      reg934 <= $unsigned((wire896[(4'hb):(3'h4)] > reg926));
                      reg935 <= (+$signed(({reg915} <<< (forvar908 - reg909))));
                      reg936 <= $signed(((|reg945[(3'h6):(3'h6)]) & {reg928[(3'h7):(1'h1)]}));
                    end
                  if ($signed($signed($signed((~forvar898)))))
                    begin
                      reg937 <= ((!reg906) ?
                          {$signed((8'ha5))} : (&reg905[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg937 <= $signed($unsigned({reg937}));
                      reg938 <= wire893;
                      reg939 <= reg897[(4'hc):(4'hc)];
                    end
                end
              if (($unsigned((~|forvar932)) ?
                  (($signed(reg940) << reg911) ^~ (^reg924[(4'ha):(3'h6)])) : reg925))
                begin
                  reg940 <= (reg904[(2'h2):(1'h0)] | $unsigned($unsigned($signed(reg908))));
                end
              else
                begin
                  if (reg905)
                    begin
                      reg940 <= $signed($unsigned($signed({(8'h9c)})));
                      reg941 <= (($signed((reg913 + reg897)) ^ (forvar897[(3'h7):(3'h7)] >> $signed(reg939))) && wire889[(3'h5):(2'h2)]);
                      reg942 <= {reg902};
                    end
                  else
                    begin
                      reg940 <= $signed(forvar908);
                      reg941 <= ((reg932[(3'h6):(2'h2)] ?
                              ((reg912 ? reg936 : wire890) ?
                                  reg921[(4'h8):(4'h8)] : ((8'hb0) ~^ (8'hae))) : $signed((reg935 ?
                                  (8'hb3) : reg939))) ?
                          $signed(reg935) : $unsigned($signed((~|reg909))));
                      reg942 <= $signed(forvar932[(4'h8):(1'h0)]);
                    end
                  if ($signed((~&reg926)))
                    begin
                      reg943 <= ((($signed(forvar918) ?
                          (^forvar902) : {(8'h9d)}) <<< (forvar929[(3'h6):(1'h1)] && wire896[(3'h7):(3'h7)])) + reg912);
                      reg944 <= reg945[(3'h6):(2'h3)];
                      reg945 <= forvar917[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg943 <= reg906[(1'h1):(1'h1)];
                    end
                  for (forvar946 = (1'h0); (forvar946 < (2'h3)); forvar946 = (forvar946 + (1'h1)))
                    begin
                      reg947 <= $signed((|($signed(forvar898) & forvar930)));
                      reg948 <= $unsigned({$signed(reg912[(2'h3):(1'h0)])});
                      reg949 <= {{forvar908}};
                      reg950 <= reg899[(4'h9):(4'h8)];
                    end
                end
            end
          if ((!reg897[(3'h5):(1'h0)]))
            begin
              if ($unsigned({(^(|wire889))}))
                begin
                  for (forvar951 = (1'h0); (forvar951 < (1'h0)); forvar951 = (forvar951 + (1'h1)))
                    begin
                      reg952 <= forvar920[(3'h6):(1'h1)];
                    end
                  for (forvar953 = (1'h0); (forvar953 < (1'h1)); forvar953 = (forvar953 + (1'h1)))
                    begin
                      reg954 <= ($unsigned(reg907[(3'h7):(2'h3)]) * ($signed((reg947 ?
                          (8'ha4) : (8'hb2))) <= {(^reg916)}));
                      reg955 <= ({reg924[(1'h1):(1'h1)]} ?
                          ($unsigned($signed(reg932)) ?
                              (|wire894[(1'h0):(1'h0)]) : reg911[(1'h0):(1'h0)]) : {(~(~^reg936))});
                      reg956 <= (8'hb3);
                      reg957 <= $unsigned(reg934[(4'h8):(2'h3)]);
                    end
                  if (((~reg949) ? wire889[(1'h1):(1'h1)] : reg948))
                    begin
                      reg958 <= $unsigned((~^$signed((+forvar902))));
                      reg959 <= ({$unsigned($unsigned(reg923))} && ($signed({wire890}) - reg897));
                    end
                  else
                    begin
                      reg958 <= (reg936 >= (reg956[(4'h9):(4'h8)] <= $signed(wire894)));
                      reg959 <= $signed(($unsigned((reg940 | reg950)) < (((8'ha1) && wire895) ?
                          reg905 : reg942)));
                    end
                  for (forvar960 = (1'h0); (forvar960 < (2'h3)); forvar960 = (forvar960 + (1'h1)))
                    begin
                      reg961 <= ((((reg906 ~^ forvar908) ?
                              (reg950 || reg947) : reg919[(4'ha):(4'h8)]) != wire893) ?
                          {$unsigned(wire895[(4'h8):(3'h7)])} : {{(reg932 ^~ (8'haf))}});
                    end
                end
              else
                begin
                  reg951 <= (^(~forvar942));
                  for (forvar952 = (1'h0); (forvar952 < (1'h0)); forvar952 = (forvar952 + (1'h1)))
                    begin
                      reg953 <= (reg943 <<< (~&({forvar917} ?
                          $signed(forvar910) : $unsigned(forvar960))));
                    end
                end
              for (forvar962 = (1'h0); (forvar962 < (1'h1)); forvar962 = (forvar962 + (1'h1)))
                begin
                  for (forvar963 = (1'h0); (forvar963 < (1'h1)); forvar963 = (forvar963 + (1'h1)))
                    begin
                      reg964 <= ((8'ha8) ?
                          (reg910 ?
                              ((-reg903) + $unsigned(reg926)) : ((~&(8'hb2)) | $unsigned(reg911))) : forvar951[(1'h0):(1'h0)]);
                      reg965 <= (~(~^$signed((reg916 != reg909))));
                    end
                  reg966 <= (~$signed(reg919));
                  for (forvar967 = (1'h0); (forvar967 < (2'h2)); forvar967 = (forvar967 + (1'h1)))
                    begin
                      reg968 <= $unsigned(($unsigned((~|forvar942)) >>> ((-reg944) * reg907)));
                    end
                end
            end
          else
            begin
              for (forvar951 = (1'h0); (forvar951 < (1'h1)); forvar951 = (forvar951 + (1'h1)))
                begin
                  reg952 <= reg902[(4'h8):(3'h5)];
                  for (forvar953 = (1'h0); (forvar953 < (2'h2)); forvar953 = (forvar953 + (1'h1)))
                    begin
                      reg954 <= $signed({{(reg946 ? reg951 : (8'hab))}});
                    end
                end
              if (($unsigned(((^reg905) ~^ reg897[(2'h3):(1'h1)])) > {(~^(reg935 >> forvar963))}))
                begin
                  for (forvar955 = (1'h0); (forvar955 < (1'h1)); forvar955 = (forvar955 + (1'h1)))
                    begin
                      reg956 <= {reg956[(4'hb):(1'h1)]};
                      reg957 <= (reg913 ~^ {$unsigned((+(8'ha0)))});
                      reg958 <= reg951[(1'h0):(1'h0)];
                      reg959 <= forvar963[(4'h8):(2'h3)];
                    end
                  reg960 <= forvar952[(1'h1):(1'h0)];
                end
              else
                begin
                  if (((~^reg909) ? reg950 : $unsigned(reg942)))
                    begin
                      reg955 <= reg904[(4'h8):(1'h1)];
                      reg956 <= $signed((&reg921));
                      reg957 <= $unsigned($signed($signed($signed(reg919))));
                    end
                  else
                    begin
                      reg955 <= ((forvar953[(1'h0):(1'h0)] ?
                          $signed(((8'ha9) & forvar960)) : (reg953[(2'h2):(1'h1)] << (reg927 != wire894))) & $unsigned((!$unsigned(forvar898))));
                    end
                  for (forvar958 = (1'h0); (forvar958 < (2'h3)); forvar958 = (forvar958 + (1'h1)))
                    begin
                      reg959 <= reg904;
                      reg960 <= ($signed(reg897) ?
                          (|(reg932[(4'h9):(2'h3)] * $unsigned(forvar920))) : {($signed((8'hb9)) ?
                                  $unsigned(reg945) : reg919[(4'ha):(4'h8)])});
                      reg961 <= (^$unsigned($unsigned($signed(forvar952))));
                    end
                  for (forvar962 = (1'h0); (forvar962 < (1'h0)); forvar962 = (forvar962 + (1'h1)))
                    begin
                      reg963 <= $signed((reg934 >= reg959[(3'h4):(3'h4)]));
                    end
                end
              for (forvar964 = (1'h0); (forvar964 < (2'h2)); forvar964 = (forvar964 + (1'h1)))
                begin
                  reg965 <= ($unsigned({reg957}) ?
                      {(~(reg953 | (8'hb6)))} : $unsigned($signed((forvar910 ?
                          reg945 : reg903))));
                  if ({wire895[(3'h5):(2'h3)]})
                    begin
                      reg966 <= wire895[(4'h8):(3'h7)];
                      reg967 <= reg963[(2'h3):(2'h2)];
                      reg968 <= $signed($signed(reg961[(1'h1):(1'h1)]));
                      reg969 <= {reg921[(4'hb):(1'h0)]};
                    end
                  else
                    begin
                      reg966 <= {(^$unsigned($signed(reg951)))};
                      reg967 <= $unsigned({$signed(reg915)});
                    end
                end
              if (reg907[(2'h2):(1'h1)])
                begin
                  if (($signed((|(+reg900))) ^~ ($unsigned({forvar897}) ?
                      $unsigned((reg945 ?
                          (8'hb2) : forvar909)) : $signed((reg907 || reg907)))))
                    begin
                      reg970 <= $unsigned(((^(reg933 ?
                          reg943 : reg936)) <= reg942[(2'h2):(1'h1)]));
                      reg971 <= ($unsigned(((-(8'hb9)) <<< $unsigned(reg905))) ?
                          (reg969[(3'h7):(2'h3)] * $signed({reg939})) : reg927);
                    end
                  else
                    begin
                      reg970 <= forvar918[(1'h1):(1'h0)];
                      reg971 <= $signed((~|$signed((reg970 ?
                          (8'hae) : forvar962))));
                    end
                end
              else
                begin
                  reg970 <= ($unsigned(((|reg905) < (reg940 & reg971))) ?
                      (reg955[(1'h1):(1'h0)] + $signed($unsigned(reg919))) : {{reg901[(1'h0):(1'h0)]}});
                  for (forvar971 = (1'h0); (forvar971 < (1'h0)); forvar971 = (forvar971 + (1'h1)))
                    begin
                      reg972 <= wire891;
                      reg973 <= (($unsigned((^reg936)) ?
                              $signed((reg968 == reg924)) : $unsigned(wire894)) ?
                          (|reg940[(2'h2):(2'h2)]) : $unsigned(forvar900[(4'h8):(2'h2)]));
                    end
                  for (forvar974 = (1'h0); (forvar974 < (1'h1)); forvar974 = (forvar974 + (1'h1)))
                    begin
                      reg975 <= ($unsigned(forvar958[(3'h5):(3'h5)]) + (($signed(wire896) == (~&reg968)) - reg971[(3'h4):(2'h2)]));
                      reg976 <= forvar967;
                      reg977 <= reg920[(3'h5):(2'h2)];
                    end
                end
            end
          if (reg946)
            begin
              if (reg947)
                begin
                  for (forvar978 = (1'h0); (forvar978 < (2'h3)); forvar978 = (forvar978 + (1'h1)))
                    begin
                      reg979 <= ((reg970[(3'h4):(2'h3)] == forvar963) + (($signed(reg938) + $unsigned(forvar953)) && ({(8'hae)} <<< forvar930)));
                      reg980 <= reg928;
                    end
                end
              else
                begin
                  reg978 <= (|{((^~reg916) ^~ (forvar897 ? reg904 : reg899))});
                end
              if (reg936)
                begin
                  for (forvar981 = (1'h0); (forvar981 < (1'h1)); forvar981 = (forvar981 + (1'h1)))
                    begin
                      reg982 <= ((8'ha5) & (((|reg916) ?
                              (reg978 && reg972) : reg897[(4'hc):(2'h3)]) ?
                          reg937 : $signed(forvar962[(1'h0):(1'h0)])));
                      reg983 <= (~^reg916);
                      reg984 <= {($unsigned(reg965[(2'h3):(1'h1)]) >>> wire893[(3'h4):(3'h4)])};
                      reg985 <= $signed((&reg946[(4'ha):(1'h0)]));
                    end
                end
              else
                begin
                  reg981 <= forvar971[(2'h2):(2'h2)];
                end
              if ($signed(wire896[(3'h5):(2'h2)]))
                begin
                  for (forvar986 = (1'h0); (forvar986 < (2'h3)); forvar986 = (forvar986 + (1'h1)))
                    begin
                      reg987 <= reg968[(4'h8):(3'h6)];
                      reg988 <= (-wire895);
                      reg989 <= (~|forvar960[(4'hc):(4'h8)]);
                    end
                  reg990 <= reg955[(2'h3):(1'h1)];
                end
              else
                begin
                  reg986 <= $unsigned(reg902);
                  for (forvar987 = (1'h0); (forvar987 < (1'h0)); forvar987 = (forvar987 + (1'h1)))
                    begin
                      reg988 <= $unsigned((|{(~&reg921)}));
                      reg989 <= ((~&$unsigned((~reg923))) ~^ $signed($unsigned(((8'ha8) >= reg931))));
                      reg990 <= ((reg910 ?
                              ($signed(wire893) ?
                                  $unsigned(reg958) : (-reg971)) : (reg973[(1'h1):(1'h1)] | {(8'hba)})) ?
                          $signed(forvar897[(2'h2):(1'h0)]) : (~$signed($signed(reg917))));
                    end
                  reg991 <= $unsigned((+forvar923));
                end
            end
          else
            begin
              for (forvar978 = (1'h0); (forvar978 < (1'h0)); forvar978 = (forvar978 + (1'h1)))
                begin
                  if (reg986)
                    begin
                      reg979 <= reg927;
                      reg980 <= forvar919[(4'h9):(2'h3)];
                      reg981 <= {(($signed(wire890) ?
                                  $signed(forvar932) : (forvar963 ?
                                      reg905 : wire893)) ?
                              (8'hba) : reg985[(2'h3):(2'h3)])};
                    end
                  else
                    begin
                      reg979 <= $signed((wire892[(2'h2):(1'h0)] != ($unsigned(forvar987) ?
                          reg976 : (~&reg900))));
                      reg980 <= ($unsigned($signed($signed(reg963))) == (~|(((8'hac) ?
                          forvar932 : forvar986) <<< $unsigned((8'hb9)))));
                      reg981 <= reg981;
                    end
                  for (forvar982 = (1'h0); (forvar982 < (1'h0)); forvar982 = (forvar982 + (1'h1)))
                    begin
                      reg983 <= ($signed((&(&forvar967))) ?
                          $signed((~^(~&reg972))) : (forvar953[(2'h2):(1'h1)] != reg933));
                    end
                  for (forvar984 = (1'h0); (forvar984 < (2'h2)); forvar984 = (forvar984 + (1'h1)))
                    begin
                      reg985 <= (~&reg900);
                      reg986 <= forvar962;
                      reg987 <= {{$unsigned((|reg910))}};
                    end
                end
            end
          for (forvar992 = (1'h0); (forvar992 < (1'h0)); forvar992 = (forvar992 + (1'h1)))
            begin
              for (forvar993 = (1'h0); (forvar993 < (1'h1)); forvar993 = (forvar993 + (1'h1)))
                begin
                  if ((reg980[(1'h1):(1'h1)] ?
                      $signed(reg988) : ((8'hae) ? (!(-reg959)) : (8'ha4))))
                    begin
                      reg994 <= reg943;
                      reg995 <= ((forvar962[(3'h6):(3'h5)] ?
                          {reg970[(2'h3):(1'h0)]} : forvar909) | ($signed(((8'h9c) ?
                          reg902 : reg943)) <= $signed((reg950 ?
                          reg978 : reg983))));
                      reg996 <= ($unsigned((~|$unsigned(reg950))) & (~(reg932[(3'h6):(1'h1)] == (8'ha9))));
                      reg997 <= (~^reg990);
                    end
                  else
                    begin
                      reg994 <= ($unsigned((+{reg965})) ?
                          reg906 : $unsigned(reg997));
                      reg995 <= {((|reg903) ?
                              $unsigned(reg957[(2'h2):(2'h2)]) : reg897)};
                    end
                  for (forvar998 = (1'h0); (forvar998 < (2'h2)); forvar998 = (forvar998 + (1'h1)))
                    begin
                      reg999 <= (^{(+(reg963 <= forvar909))});
                      reg1000 <= (^~($signed({reg942}) ?
                          reg958 : $unsigned(reg932[(2'h2):(1'h1)])));
                    end
                end
            end
        end
    end
  module1001 modinst1019 (.wire1004(reg899), .wire1005(forvar930), .wire1003(reg983), .y(wire1018), .clk(clk), .wire1002(reg959));
  always
    @(posedge clk) begin
      if ($signed((reg943 >> reg911)))
        begin
          for (forvar1020 = (1'h0); (forvar1020 < (1'h1)); forvar1020 = (forvar1020 + (1'h1)))
            begin
              for (forvar1021 = (1'h0); (forvar1021 < (1'h1)); forvar1021 = (forvar1021 + (1'h1)))
                begin
                  for (forvar1022 = (1'h0); (forvar1022 < (2'h2)); forvar1022 = (forvar1022 + (1'h1)))
                    begin
                      reg1023 <= $unsigned({((reg926 ? forvar962 : wire892) ?
                              forvar919[(3'h5):(1'h1)] : reg934)});
                    end
                  if ({reg916})
                    begin
                      reg1024 <= $unsigned((~&reg927[(3'h5):(1'h1)]));
                      reg1025 <= (((~^(-reg957)) ?
                          reg997 : (forvar909[(3'h7):(3'h4)] || (reg978 + reg908))) == ($unsigned($signed((8'h9d))) > $signed($unsigned(reg1023))));
                      reg1026 <= $unsigned((~&forvar984));
                      reg1027 <= (~$unsigned(({reg916} ?
                          {forvar963} : $unsigned(forvar929))));
                    end
                  else
                    begin
                      reg1024 <= reg919[(4'he):(4'h9)];
                    end
                end
              for (forvar1028 = (1'h0); (forvar1028 < (1'h1)); forvar1028 = (forvar1028 + (1'h1)))
                begin
                  for (forvar1029 = (1'h0); (forvar1029 < (2'h3)); forvar1029 = (forvar1029 + (1'h1)))
                    begin
                      reg1030 <= (^~(($signed(reg942) | (reg924 < forvar987)) ?
                          {wire892[(2'h3):(2'h3)]} : forvar930));
                      reg1031 <= $signed($unsigned(forvar1028));
                    end
                  for (forvar1032 = (1'h0); (forvar1032 < (1'h1)); forvar1032 = (forvar1032 + (1'h1)))
                    begin
                      reg1033 <= {forvar993[(2'h2):(1'h1)]};
                      reg1034 <= ((~&(~^$unsigned(reg960))) ?
                          wire892 : $signed({$unsigned(reg985)}));
                      reg1035 <= reg937;
                      reg1036 <= {reg936[(1'h1):(1'h0)]};
                    end
                end
            end
          for (forvar1037 = (1'h0); (forvar1037 < (2'h3)); forvar1037 = (forvar1037 + (1'h1)))
            begin
              for (forvar1038 = (1'h0); (forvar1038 < (2'h3)); forvar1038 = (forvar1038 + (1'h1)))
                begin
                  reg1039 <= (~(~&$unsigned(reg924)));
                end
              for (forvar1040 = (1'h0); (forvar1040 < (1'h0)); forvar1040 = (forvar1040 + (1'h1)))
                begin
                  if ({(8'ha5)})
                    begin
                      reg1041 <= forvar960;
                      reg1042 <= $signed(($signed((~reg953)) > (~^$unsigned(reg983))));
                      reg1043 <= ($signed(((forvar955 ?
                          reg952 : forvar920) <= (reg990 ?
                          (8'hb0) : wire893))) ^ reg981);
                      reg1044 <= (8'h9c);
                    end
                  else
                    begin
                      reg1041 <= (~^($signed((~^reg1044)) && {(reg968 ^~ (8'hb1))}));
                      reg1042 <= (^((8'hba) && wire893[(3'h5):(2'h3)]));
                      reg1043 <= ((^~(+{reg945})) == reg1036[(2'h2):(2'h2)]);
                      reg1044 <= {((-$signed(forvar952)) ?
                              forvar1029 : ((^forvar955) ? reg931 : reg1027))};
                    end
                end
            end
          reg1045 <= reg906[(2'h2):(1'h0)];
          reg1046 <= {$signed((forvar964[(4'hb):(2'h3)] | reg939[(1'h1):(1'h1)]))};
        end
      else
        begin
          for (forvar1020 = (1'h0); (forvar1020 < (1'h0)); forvar1020 = (forvar1020 + (1'h1)))
            begin
              if ($signed(reg963[(2'h2):(1'h0)]))
                begin
                  for (forvar1021 = (1'h0); (forvar1021 < (2'h3)); forvar1021 = (forvar1021 + (1'h1)))
                    begin
                      reg1022 <= $unsigned($unsigned((&(~^reg1023))));
                      reg1023 <= ((((reg976 ? (8'ha1) : forvar898) ^ (reg897 ?
                              wire889 : (8'hb1))) >= $unsigned($unsigned(forvar951))) ?
                          ((-(8'hb1)) | wire894) : (~^$unsigned((8'hae))));
                      reg1024 <= (~^($signed(reg906[(1'h1):(1'h0)]) ?
                          $unsigned(reg965[(3'h5):(3'h4)]) : $signed((reg965 != reg914))));
                      reg1025 <= reg918;
                    end
                  if ((8'hb1))
                    begin
                      reg1026 <= reg915[(3'h5):(1'h1)];
                      reg1027 <= ({reg905[(1'h1):(1'h0)]} ^~ (|(|(reg1027 >> reg969))));
                      reg1028 <= $signed((+$unsigned(forvar998[(2'h3):(1'h0)])));
                      reg1029 <= $signed($signed(reg940));
                    end
                  else
                    begin
                      reg1026 <= reg982[(3'h5):(1'h0)];
                      reg1027 <= reg952[(4'he):(2'h3)];
                    end
                  for (forvar1030 = (1'h0); (forvar1030 < (2'h2)); forvar1030 = (forvar1030 + (1'h1)))
                    begin
                      reg1031 <= reg1023;
                      reg1032 <= wire894;
                    end
                end
              else
                begin
                  for (forvar1021 = (1'h0); (forvar1021 < (1'h1)); forvar1021 = (forvar1021 + (1'h1)))
                    begin
                      reg1022 <= ((~&($signed(forvar998) ?
                              (+forvar1038) : $signed(forvar941))) ?
                          ($signed(reg976[(2'h2):(2'h2)]) > forvar953[(2'h2):(2'h2)]) : {wire891[(3'h5):(3'h4)]});
                    end
                end
              for (forvar1033 = (1'h0); (forvar1033 < (1'h0)); forvar1033 = (forvar1033 + (1'h1)))
                begin
                  reg1034 <= (reg928 != ($unsigned($signed(forvar1029)) ?
                      (!$unsigned(reg946)) : $signed((forvar941 ?
                          reg938 : reg940))));
                  reg1035 <= (((~&$unsigned(forvar932)) + reg978[(1'h1):(1'h0)]) ?
                      $signed(reg903) : $unsigned($unsigned($signed(reg908))));
                end
              for (forvar1036 = (1'h0); (forvar1036 < (2'h3)); forvar1036 = (forvar1036 + (1'h1)))
                begin
                  reg1037 <= (reg1022 | (forvar1021 ~^ reg953[(3'h5):(1'h0)]));
                  for (forvar1038 = (1'h0); (forvar1038 < (1'h0)); forvar1038 = (forvar1038 + (1'h1)))
                    begin
                      reg1039 <= {$signed(forvar929[(3'h5):(2'h3)])};
                    end
                  if ((forvar1029 ?
                      (~(&(forvar986 << forvar921))) : {(^(forvar921 ?
                              wire1018 : forvar946))}))
                    begin
                      reg1040 <= $signed($unsigned(wire894));
                      reg1041 <= (|$signed(((^~forvar902) >> $unsigned(reg922))));
                    end
                  else
                    begin
                      reg1040 <= ({reg937} < (reg1035 || (reg1045[(3'h5):(3'h5)] ?
                          reg1044[(3'h4):(2'h2)] : forvar974)));
                      reg1041 <= forvar919[(1'h0):(1'h0)];
                      reg1042 <= $unsigned(reg969[(1'h0):(1'h0)]);
                      reg1043 <= $signed({(~&forvar902)});
                    end
                  for (forvar1044 = (1'h0); (forvar1044 < (1'h1)); forvar1044 = (forvar1044 + (1'h1)))
                    begin
                      reg1045 <= (^~reg1034);
                    end
                end
            end
        end
      for (forvar1047 = (1'h0); (forvar1047 < (2'h3)); forvar1047 = (forvar1047 + (1'h1)))
        begin
          for (forvar1048 = (1'h0); (forvar1048 < (2'h2)); forvar1048 = (forvar1048 + (1'h1)))
            begin
              for (forvar1049 = (1'h0); (forvar1049 < (2'h2)); forvar1049 = (forvar1049 + (1'h1)))
                begin
                  reg1050 <= $signed(reg920);
                  if ($unsigned((($unsigned(reg906) ?
                          (reg918 ? (8'h9e) : reg912) : (8'hac)) ?
                      ((-reg1024) >> $unsigned(reg907)) : ((8'h9d) ?
                          (8'ha1) : reg1041[(4'h8):(3'h6)]))))
                    begin
                      reg1051 <= (reg1039 != $signed($signed((forvar981 ?
                          reg935 : reg900))));
                    end
                  else
                    begin
                      reg1051 <= forvar917[(3'h4):(2'h3)];
                      reg1052 <= $unsigned((^{reg982}));
                    end
                end
              reg1053 <= (reg908 ? (8'haf) : reg948[(2'h2):(1'h1)]);
              for (forvar1054 = (1'h0); (forvar1054 < (2'h3)); forvar1054 = (forvar1054 + (1'h1)))
                begin
                  for (forvar1055 = (1'h0); (forvar1055 < (1'h1)); forvar1055 = (forvar1055 + (1'h1)))
                    begin
                      reg1056 <= (|reg897);
                      reg1057 <= ((($unsigned(reg982) ?
                              (forvar1022 << reg917) : (forvar920 << (8'hb6))) & (reg987[(1'h1):(1'h1)] * (8'ha5))) ?
                          $signed(forvar981) : reg945[(1'h0):(1'h0)]);
                    end
                  reg1058 <= (forvar993 ^ ($signed($unsigned(forvar984)) ~^ {{forvar942}}));
                end
            end
          if ($unsigned($signed($signed($unsigned(wire1018)))))
            begin
              for (forvar1059 = (1'h0); (forvar1059 < (2'h3)); forvar1059 = (forvar1059 + (1'h1)))
                begin
                  for (forvar1060 = (1'h0); (forvar1060 < (2'h3)); forvar1060 = (forvar1060 + (1'h1)))
                    begin
                      reg1061 <= wire892[(2'h3):(2'h2)];
                      reg1062 <= {reg911[(1'h1):(1'h1)]};
                      reg1063 <= (reg1053 ? (8'hb1) : reg995);
                      reg1064 <= ((reg926[(4'h9):(3'h4)] > reg940) >>> (~^(-$signed(reg999))));
                    end
                  for (forvar1065 = (1'h0); (forvar1065 < (1'h1)); forvar1065 = (forvar1065 + (1'h1)))
                    begin
                      reg1066 <= reg1062;
                      reg1067 <= reg949;
                      reg1068 <= (((forvar1022 > (&(8'hb0))) ?
                          $unsigned((reg936 ?
                              reg934 : reg921)) : (-forvar960)) >> (($signed(forvar978) || $signed(reg1026)) << (~((8'hab) ?
                          forvar953 : forvar998))));
                      reg1069 <= (&(~^($unsigned(reg901) ~^ $unsigned(forvar993))));
                    end
                  reg1070 <= ($signed(reg999[(2'h2):(2'h2)]) << ($signed((~&reg920)) ~^ ($unsigned(forvar971) ?
                      reg926[(5'h10):(2'h3)] : (&reg942))));
                end
              reg1071 <= reg943[(4'he):(4'hb)];
              reg1072 <= $unsigned(reg1025);
            end
          else
            begin
              for (forvar1059 = (1'h0); (forvar1059 < (1'h0)); forvar1059 = (forvar1059 + (1'h1)))
                begin
                  if (reg917[(3'h7):(3'h4)])
                    begin
                      reg1060 <= $unsigned(reg911);
                      reg1061 <= ({(^~(|(8'ha8)))} - (8'h9d));
                      reg1062 <= reg934[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1060 <= forvar1030;
                      reg1061 <= $signed(forvar1065[(3'h4):(3'h4)]);
                      reg1062 <= $unsigned($unsigned($signed((~&(8'haa)))));
                    end
                  if ($unsigned($unsigned($signed($unsigned((8'hb4))))))
                    begin
                      reg1063 <= ((forvar1030 ^~ ((reg1058 ?
                              reg970 : reg919) >>> $signed((8'ha5)))) ?
                          reg1029[(3'h6):(3'h4)] : (($signed(reg1028) > $unsigned(reg926)) ?
                              ($signed(reg1044) || (~&forvar993)) : $signed((~^forvar992))));
                    end
                  else
                    begin
                      reg1063 <= (forvar962[(3'h5):(1'h0)] ?
                          forvar1040 : reg942);
                      reg1064 <= reg924[(1'h0):(1'h0)];
                      reg1065 <= (forvar967[(1'h1):(1'h0)] || $unsigned($signed(reg934[(4'h8):(4'h8)])));
                      reg1066 <= reg900[(2'h3):(1'h1)];
                    end
                end
            end
          reg1073 <= {$unsigned(((reg925 ^ forvar987) ?
                  ((8'hac) >>> (8'hb1)) : (forvar1022 != (8'ha2))))};
        end
      if ($signed($unsigned($unsigned($signed(reg1072)))))
        begin
          for (forvar1074 = (1'h0); (forvar1074 < (2'h3)); forvar1074 = (forvar1074 + (1'h1)))
            begin
              for (forvar1075 = (1'h0); (forvar1075 < (2'h2)); forvar1075 = (forvar1075 + (1'h1)))
                begin
                  if ((!reg899))
                    begin
                      reg1076 <= reg901;
                    end
                  else
                    begin
                      reg1076 <= $signed(reg1051[(1'h0):(1'h0)]);
                      reg1077 <= $signed(reg963);
                    end
                  if ((reg983[(4'h8):(1'h1)] ?
                      reg914[(1'h0):(1'h0)] : ($unsigned($unsigned(reg955)) ^~ {{reg991}})))
                    begin
                      reg1078 <= forvar986[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg1078 <= (~^(((reg1062 ? reg1032 : wire893) ?
                              forvar902[(4'h8):(2'h2)] : (reg960 * forvar1054)) ?
                          ((-reg940) || (reg999 >= reg964)) : (~^wire896[(2'h2):(2'h2)])));
                    end
                  reg1079 <= $signed($signed($unsigned($signed((8'ha3)))));
                  for (forvar1080 = (1'h0); (forvar1080 < (2'h3)); forvar1080 = (forvar1080 + (1'h1)))
                    begin
                      reg1081 <= ((~^forvar987[(4'hb):(3'h5)]) < (reg1046[(1'h0):(1'h0)] ?
                          $signed(reg946[(2'h2):(1'h1)]) : ((8'hb5) ?
                              reg1056 : (forvar981 >>> forvar992))));
                      reg1082 <= ($unsigned(reg939[(2'h3):(2'h3)]) >>> {(~&((8'h9d) ?
                              (8'ha2) : (8'ha9)))});
                      reg1083 <= $signed(reg964);
                    end
                end
              for (forvar1084 = (1'h0); (forvar1084 < (1'h1)); forvar1084 = (forvar1084 + (1'h1)))
                begin
                  for (forvar1085 = (1'h0); (forvar1085 < (1'h0)); forvar1085 = (forvar1085 + (1'h1)))
                    begin
                      reg1086 <= $unsigned($signed($signed(forvar910)));
                      reg1087 <= $signed(reg1062);
                    end
                end
            end
          reg1088 <= reg903;
          for (forvar1089 = (1'h0); (forvar1089 < (1'h1)); forvar1089 = (forvar1089 + (1'h1)))
            begin
              reg1090 <= reg983[(3'h4):(1'h1)];
              for (forvar1091 = (1'h0); (forvar1091 < (1'h1)); forvar1091 = (forvar1091 + (1'h1)))
                begin
                  if ((reg976[(1'h0):(1'h0)] ?
                      (forvar921[(4'h8):(3'h7)] >>> forvar962[(3'h7):(3'h4)]) : $signed(forvar1020[(1'h1):(1'h1)])))
                    begin
                      reg1092 <= forvar992;
                      reg1093 <= ($unsigned((reg1022 ?
                          ((8'h9c) ?
                              reg926 : reg931) : forvar998)) + reg1072[(2'h2):(1'h0)]);
                      reg1094 <= $signed($unsigned($signed($unsigned(reg909))));
                    end
                  else
                    begin
                      reg1092 <= (($signed($signed(forvar992)) ?
                              $signed((reg966 ?
                                  reg970 : reg944)) : (~$unsigned(forvar918))) ?
                          $signed((^~(reg990 * (8'haa)))) : $signed(reg1072));
                      reg1093 <= $signed({$unsigned(reg952)});
                      reg1094 <= ($signed(((|forvar971) == $signed(reg925))) ~^ reg902);
                      reg1095 <= $unsigned($signed((((8'ha2) && (8'hb3)) ?
                          $unsigned(reg1092) : (reg975 - reg922))));
                    end
                  reg1096 <= $signed((forvar1084[(3'h4):(3'h4)] <<< $signed((8'ha1))));
                  for (forvar1097 = (1'h0); (forvar1097 < (1'h1)); forvar1097 = (forvar1097 + (1'h1)))
                    begin
                      reg1098 <= (~^({(~^reg967)} | wire895[(2'h3):(2'h3)]));
                      reg1099 <= (8'had);
                      reg1100 <= (($signed(reg989) >= $signed($signed(reg997))) ^~ (reg973 == $signed($unsigned(forvar987))));
                    end
                  if ({$unsigned($signed($signed(reg987)))})
                    begin
                      reg1101 <= $unsigned(((wire1018[(2'h2):(1'h0)] <<< (~^reg934)) >= $unsigned((forvar946 || forvar1084))));
                      reg1102 <= forvar998;
                    end
                  else
                    begin
                      reg1101 <= $unsigned($unsigned($signed($signed(reg1036))));
                    end
                end
            end
          if ($signed(reg955[(3'h7):(3'h4)]))
            begin
              if ($signed(($signed({reg914}) || forvar974[(3'h6):(2'h2)])))
                begin
                  for (forvar1103 = (1'h0); (forvar1103 < (1'h1)); forvar1103 = (forvar1103 + (1'h1)))
                    begin
                      reg1104 <= $unsigned(reg1062[(1'h1):(1'h0)]);
                      reg1105 <= reg917[(3'h5):(3'h5)];
                      reg1106 <= (~&reg954[(4'h8):(1'h1)]);
                      reg1107 <= {$signed((~^forvar1048[(4'hb):(4'hb)]))};
                    end
                  for (forvar1108 = (1'h0); (forvar1108 < (1'h0)); forvar1108 = (forvar1108 + (1'h1)))
                    begin
                      reg1109 <= ((reg914[(1'h1):(1'h1)] ?
                          $unsigned(reg1088) : (8'ha4)) | ((^(reg912 + reg905)) ?
                          $unsigned((~&reg964)) : ((forvar1047 ?
                              (8'hb5) : reg905) < (reg994 ?
                              reg1098 : forvar902))));
                      reg1110 <= $unsigned(((~(forvar1091 ^ reg910)) >> ($signed((8'ha4)) && reg1094[(2'h2):(2'h2)])));
                      reg1111 <= (|(~|$signed((reg1088 & reg927))));
                    end
                  for (forvar1112 = (1'h0); (forvar1112 < (2'h2)); forvar1112 = (forvar1112 + (1'h1)))
                    begin
                      reg1113 <= forvar953[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  reg1103 <= (~({(forvar930 * wire893)} <<< ((^~forvar918) ?
                      (reg952 >>> (8'hb1)) : {reg956})));
                  if ($signed(({$signed(forvar1048)} | (((8'ha2) <<< reg1057) ?
                      (~reg1056) : $unsigned(reg913)))))
                    begin
                      reg1104 <= forvar971;
                      reg1105 <= {((~$signed(reg1083)) > ({(8'ha4)} ?
                              $signed(reg1083) : $unsigned(reg1024)))};
                    end
                  else
                    begin
                      reg1104 <= (~&$unsigned($signed($unsigned((8'had)))));
                      reg1105 <= (8'ha3);
                      reg1106 <= (~&reg1042[(1'h1):(1'h1)]);
                      reg1107 <= {reg921};
                    end
                end
            end
          else
            begin
              for (forvar1103 = (1'h0); (forvar1103 < (2'h3)); forvar1103 = (forvar1103 + (1'h1)))
                begin
                  for (forvar1104 = (1'h0); (forvar1104 < (1'h1)); forvar1104 = (forvar1104 + (1'h1)))
                    begin
                      reg1105 <= forvar1089;
                      reg1106 <= (8'ha6);
                    end
                end
              for (forvar1107 = (1'h0); (forvar1107 < (1'h1)); forvar1107 = (forvar1107 + (1'h1)))
                begin
                  reg1108 <= wire890;
                  for (forvar1109 = (1'h0); (forvar1109 < (1'h1)); forvar1109 = (forvar1109 + (1'h1)))
                    begin
                      reg1110 <= $unsigned(reg972[(4'hb):(4'hb)]);
                      reg1111 <= reg939[(3'h4):(2'h2)];
                      reg1112 <= reg1058;
                      reg1113 <= (~^reg940);
                    end
                  if ({(-wire894[(3'h7):(1'h0)])})
                    begin
                      reg1114 <= (((~(forvar987 ? reg1110 : forvar1059)) ?
                          $signed((forvar1074 ?
                              forvar1089 : reg1083)) : forvar1075[(3'h7):(3'h5)]) >= $unsigned(forvar986[(1'h0):(1'h0)]));
                      reg1115 <= forvar938;
                      reg1116 <= (reg1050 ?
                          (reg1111[(4'hb):(2'h2)] ?
                              ((forvar1060 ^~ reg988) ?
                                  $signed((8'hab)) : (reg939 ?
                                      reg900 : reg945)) : $unsigned(reg968[(2'h3):(2'h3)])) : ((|$signed(reg1034)) ?
                              forvar923 : (((8'hb6) ? (8'hb3) : wire893) ?
                                  (reg1045 - reg921) : reg928)));
                    end
                  else
                    begin
                      reg1114 <= (8'h9e);
                      reg1115 <= (~^reg1057);
                    end
                end
              for (forvar1117 = (1'h0); (forvar1117 < (1'h1)); forvar1117 = (forvar1117 + (1'h1)))
                begin
                  reg1118 <= {{((reg910 ? forvar1029 : reg916) ?
                              (reg963 ~^ reg1071) : {reg975})}};
                  reg1119 <= (+$unsigned(((8'hb0) ?
                      (8'hb1) : (reg916 | forvar1117))));
                  for (forvar1120 = (1'h0); (forvar1120 < (2'h3)); forvar1120 = (forvar1120 + (1'h1)))
                    begin
                      reg1121 <= forvar1097[(3'h4):(1'h1)];
                      reg1122 <= ({(8'ha9)} ?
                          (8'hac) : $unsigned((~(forvar1047 != reg975))));
                      reg1123 <= (($unsigned((+(8'haf))) ?
                              (-$signed(reg906)) : (reg906[(1'h0):(1'h0)] ?
                                  reg1032[(2'h3):(1'h1)] : {forvar1084})) ?
                          reg924[(2'h2):(2'h2)] : $signed(($signed(reg912) ?
                              $unsigned(reg969) : $signed((8'h9e)))));
                    end
                  reg1124 <= $unsigned(forvar1022);
                end
            end
        end
      else
        begin
          for (forvar1074 = (1'h0); (forvar1074 < (1'h0)); forvar1074 = (forvar1074 + (1'h1)))
            begin
              for (forvar1075 = (1'h0); (forvar1075 < (2'h3)); forvar1075 = (forvar1075 + (1'h1)))
                begin
                  if ($unsigned((forvar1021[(4'ha):(2'h3)] ?
                      ({reg947} ?
                          forvar1080[(4'hf):(4'hb)] : $unsigned(reg902)) : forvar923)))
                    begin
                      reg1076 <= $unsigned($unsigned((~&(+reg986))));
                    end
                  else
                    begin
                      reg1076 <= reg1062;
                      reg1077 <= reg955[(4'h9):(1'h0)];
                    end
                  for (forvar1078 = (1'h0); (forvar1078 < (2'h3)); forvar1078 = (forvar1078 + (1'h1)))
                    begin
                      reg1079 <= forvar1054;
                    end
                end
            end
        end
      if ({($unsigned(forvar974) ?
              $unsigned(reg1060) : (reg1116[(1'h0):(1'h0)] ^~ reg995[(1'h0):(1'h0)]))})
        begin
          reg1125 <= ($signed($unsigned(forvar1047)) ^ reg918[(1'h0):(1'h0)]);
          if ($signed(reg951[(2'h3):(1'h1)]))
            begin
              for (forvar1126 = (1'h0); (forvar1126 < (1'h0)); forvar1126 = (forvar1126 + (1'h1)))
                begin
                  for (forvar1127 = (1'h0); (forvar1127 < (2'h2)); forvar1127 = (forvar1127 + (1'h1)))
                    begin
                      reg1128 <= (~|reg1116[(1'h0):(1'h0)]);
                      reg1129 <= $signed((8'ha3));
                    end
                  for (forvar1130 = (1'h0); (forvar1130 < (2'h3)); forvar1130 = (forvar1130 + (1'h1)))
                    begin
                      reg1131 <= {(^~$unsigned((forvar971 && forvar910)))};
                      reg1132 <= forvar1037;
                      reg1133 <= wire894;
                      reg1134 <= (forvar1044 != (!((forvar1130 ?
                              forvar1065 : forvar897) ?
                          (reg956 - (8'hb7)) : reg1113)));
                    end
                  if ((($signed(reg946[(1'h1):(1'h0)]) <= {forvar1037[(1'h0):(1'h0)]}) ?
                      reg1035 : $signed($unsigned((~(8'ha9))))))
                    begin
                      reg1135 <= reg1099[(3'h4):(2'h3)];
                      reg1136 <= $unsigned(($signed(reg1042) ?
                          reg1065 : ($unsigned((8'ha0)) ?
                              (reg1110 != reg1100) : (forvar953 ?
                                  (8'hae) : reg904))));
                      reg1137 <= $signed($unsigned((reg1050[(4'h9):(1'h1)] ?
                          $signed(reg1037) : $unsigned(reg1046))));
                    end
                  else
                    begin
                      reg1135 <= {reg980};
                    end
                end
            end
          else
            begin
              if ({{((8'hb4) ? $unsigned(reg934) : $unsigned((8'haa)))}})
                begin
                  for (forvar1126 = (1'h0); (forvar1126 < (2'h2)); forvar1126 = (forvar1126 + (1'h1)))
                    begin
                      reg1127 <= (reg940 + ((^{reg1051}) ?
                          $signed((8'hb4)) : (8'haa)));
                      reg1128 <= ((forvar917[(2'h2):(1'h1)] ?
                          $signed($signed(forvar1120)) : forvar946[(1'h1):(1'h0)]) << (8'hb2));
                      reg1129 <= (forvar942 ^~ $unsigned($unsigned($signed(forvar917))));
                    end
                  if (({($signed(forvar923) ?
                              reg942[(2'h2):(1'h0)] : (+reg913))} ?
                      (((^forvar1047) ? (wire896 || forvar1022) : reg961) ?
                          {(reg1000 <<< reg908)} : (^~$unsigned(reg1070))) : reg907))
                    begin
                      reg1130 <= ($unsigned($signed((|reg968))) ^~ ($signed((&reg1137)) ?
                          ({reg1100} | {reg1078}) : {(~&reg1132)}));
                      reg1131 <= forvar1022;
                      reg1132 <= (^(-{(reg1131 ? forvar1112 : reg1096)}));
                    end
                  else
                    begin
                      reg1130 <= reg1136;
                      reg1131 <= $unsigned(forvar908[(1'h1):(1'h1)]);
                      reg1132 <= (forvar919 ?
                          wire891[(1'h0):(1'h0)] : $unsigned((+(reg907 << (8'h9f)))));
                      reg1133 <= $signed(forvar998[(4'h8):(2'h3)]);
                    end
                  if (($signed($signed(reg963[(1'h1):(1'h0)])) ?
                      $unsigned((&(forvar1029 << reg1087))) : {{$unsigned((8'hb1))}}))
                    begin
                      reg1134 <= $signed((reg939[(3'h6):(1'h1)] ?
                          {(reg937 || reg1115)} : ($signed(forvar1022) ?
                              reg983 : reg960[(1'h1):(1'h1)])));
                      reg1135 <= $unsigned(((-$signed(reg1028)) < (~&forvar1047[(4'h9):(2'h3)])));
                    end
                  else
                    begin
                      reg1134 <= ((reg1026[(2'h2):(1'h1)] ~^ ((8'h9e) < (reg991 ?
                              forvar998 : reg1135))) ?
                          $unsigned($unsigned(forvar1048)) : ((^((8'ha8) ?
                              (8'hb1) : reg1061)) ^~ (8'h9d)));
                      reg1135 <= $signed(reg954);
                      reg1136 <= (+(reg1096 || $signed($unsigned(forvar978))));
                      reg1137 <= (&reg1046);
                    end
                end
              else
                begin
                  for (forvar1126 = (1'h0); (forvar1126 < (1'h0)); forvar1126 = (forvar1126 + (1'h1)))
                    begin
                      reg1127 <= $unsigned((~^(reg1121[(1'h0):(1'h0)] == (~&reg936))));
                    end
                end
              for (forvar1138 = (1'h0); (forvar1138 < (2'h3)); forvar1138 = (forvar1138 + (1'h1)))
                begin
                  for (forvar1139 = (1'h0); (forvar1139 < (2'h2)); forvar1139 = (forvar1139 + (1'h1)))
                    begin
                      reg1140 <= $unsigned($signed(reg967[(2'h2):(1'h1)]));
                    end
                end
            end
          for (forvar1141 = (1'h0); (forvar1141 < (1'h0)); forvar1141 = (forvar1141 + (1'h1)))
            begin
              reg1142 <= (~|(&forvar917[(3'h4):(2'h2)]));
              if (((reg1069[(4'hd):(3'h6)] ?
                      $signed($signed(reg912)) : reg955) ?
                  $signed((+$signed(reg915))) : reg1052))
                begin
                  for (forvar1143 = (1'h0); (forvar1143 < (2'h2)); forvar1143 = (forvar1143 + (1'h1)))
                    begin
                      reg1144 <= ((~^reg972) ?
                          reg1083[(3'h6):(3'h6)] : {{reg907[(3'h5):(2'h2)]}});
                    end
                  for (forvar1145 = (1'h0); (forvar1145 < (2'h2)); forvar1145 = (forvar1145 + (1'h1)))
                    begin
                      reg1146 <= $unsigned((((reg1071 ?
                          (8'hb8) : reg1144) != (reg1058 >> (8'hba))) >= $unsigned(forvar951[(3'h4):(1'h0)])));
                    end
                end
              else
                begin
                  reg1143 <= reg1137;
                end
              for (forvar1147 = (1'h0); (forvar1147 < (1'h0)); forvar1147 = (forvar1147 + (1'h1)))
                begin
                  for (forvar1148 = (1'h0); (forvar1148 < (2'h2)); forvar1148 = (forvar1148 + (1'h1)))
                    begin
                      reg1149 <= reg968;
                      reg1150 <= ($signed($signed((forvar998 ?
                              (8'h9e) : reg975))) ?
                          reg1045 : reg1061[(3'h7):(3'h7)]);
                    end
                  if ({$unsigned(((forvar1060 ? reg1113 : reg1051) ?
                          $signed(reg921) : (forvar908 <<< (8'hae))))})
                    begin
                      reg1151 <= reg1111[(4'hc):(3'h6)];
                      reg1152 <= (8'hb6);
                    end
                  else
                    begin
                      reg1151 <= (-forvar900);
                      reg1152 <= $unsigned((forvar918 ?
                          ($unsigned(forvar993) ?
                              {reg917} : {forvar1078}) : reg989));
                      reg1153 <= ({wire891[(2'h3):(2'h3)]} >> (($unsigned(reg928) ?
                          (-(8'h9e)) : $signed(forvar974)) & ($signed(reg957) < reg937[(2'h3):(2'h2)])));
                    end
                  if ($signed((-(forvar1141 ? (~&(8'h9e)) : (~^reg986)))))
                    begin
                      reg1154 <= reg1122[(4'hf):(4'hd)];
                      reg1155 <= (~&((forvar1074 ?
                              $unsigned(reg1103) : (~|reg1108)) ?
                          $signed((|reg1030)) : reg1129));
                    end
                  else
                    begin
                      reg1154 <= forvar1020[(1'h1):(1'h1)];
                    end
                end
              for (forvar1156 = (1'h0); (forvar1156 < (1'h0)); forvar1156 = (forvar1156 + (1'h1)))
                begin
                  if (reg953)
                    begin
                      reg1157 <= ((~&({reg949} ?
                              (reg1042 >> forvar1143) : ((8'ha3) && reg1090))) ?
                          (|(forvar900[(1'h1):(1'h0)] < forvar932[(4'h8):(3'h6)])) : $unsigned($signed((!reg999))));
                      reg1158 <= (((!(8'haf)) | (-(|(8'ha3)))) ?
                          (+((~|(8'hb8)) <<< {reg996})) : $signed((~|reg969)));
                    end
                  else
                    begin
                      reg1157 <= reg945[(3'h6):(2'h3)];
                    end
                  for (forvar1159 = (1'h0); (forvar1159 < (2'h3)); forvar1159 = (forvar1159 + (1'h1)))
                    begin
                      reg1160 <= $signed(reg1153[(3'h4):(2'h2)]);
                      reg1161 <= $signed(((reg959 >>> forvar1038) ?
                          {$unsigned(reg933)} : {$signed(reg1061)}));
                      reg1162 <= reg955[(4'ha):(2'h3)];
                    end
                end
            end
        end
      else
        begin
          for (forvar1125 = (1'h0); (forvar1125 < (2'h2)); forvar1125 = (forvar1125 + (1'h1)))
            begin
              reg1126 <= (forvar946[(3'h7):(2'h2)] > reg1106[(4'ha):(1'h1)]);
              for (forvar1127 = (1'h0); (forvar1127 < (2'h3)); forvar1127 = (forvar1127 + (1'h1)))
                begin
                  if (($signed(forvar1109[(3'h7):(1'h0)]) >> $signed({reg984})))
                    begin
                      reg1128 <= ($signed(reg995) ^~ $unsigned(wire896[(3'h4):(2'h2)]));
                      reg1129 <= $unsigned(({$signed((8'ha8))} >> forvar1033[(2'h3):(1'h0)]));
                      reg1130 <= $unsigned(reg1062[(3'h5):(3'h5)]);
                      reg1131 <= forvar946[(4'hc):(2'h3)];
                    end
                  else
                    begin
                      reg1128 <= ({(~^((8'h9d) ~^ forvar958))} >= ($signed((forvar993 << reg994)) ?
                          ((+(8'h9d)) ?
                              $unsigned(forvar1022) : $unsigned(reg1150)) : (^~(reg935 <<< (8'hae)))));
                      reg1129 <= ($unsigned(reg972) - ($signed(reg1086[(2'h3):(1'h1)]) || $signed((~^reg1098))));
                    end
                end
            end
          if ($signed(reg1124))
            begin
              for (forvar1132 = (1'h0); (forvar1132 < (1'h1)); forvar1132 = (forvar1132 + (1'h1)))
                begin
                  if (((({(8'hac)} == (~|(8'hb8))) ?
                      forvar908 : reg1107[(2'h2):(1'h1)]) != $unsigned({forvar1033[(1'h0):(1'h0)]})))
                    begin
                      reg1133 <= $signed(reg1078[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1133 <= $unsigned($unsigned(reg1111[(2'h2):(1'h0)]));
                      reg1134 <= forvar1126[(3'h4):(1'h1)];
                      reg1135 <= reg936;
                      reg1136 <= $unsigned(forvar958[(4'hc):(3'h4)]);
                    end
                  reg1137 <= (&reg938[(4'hc):(3'h5)]);
                  reg1138 <= (^~((~^(reg907 ? forvar1029 : reg973)) ?
                      {reg969} : {(~&reg1103)}));
                  reg1139 <= (($unsigned($unsigned(forvar1054)) ?
                      (&(^~reg1111)) : $unsigned(reg1130[(2'h2):(2'h2)])) - reg1040[(1'h0):(1'h0)]);
                end
              reg1140 <= forvar930;
            end
          else
            begin
              for (forvar1132 = (1'h0); (forvar1132 < (2'h3)); forvar1132 = (forvar1132 + (1'h1)))
                begin
                  for (forvar1133 = (1'h0); (forvar1133 < (1'h1)); forvar1133 = (forvar1133 + (1'h1)))
                    begin
                      reg1134 <= (forvar992[(4'hf):(2'h3)] << (!(reg1137 ~^ $unsigned(reg965))));
                      reg1135 <= (forvar1159[(2'h2):(2'h2)] + reg1137);
                      reg1136 <= forvar1103[(1'h1):(1'h0)];
                      reg1137 <= (reg1082[(3'h5):(1'h1)] ?
                          (!forvar920) : ($unsigned((reg1024 ?
                              forvar1097 : reg1122)) >= {(forvar932 ?
                                  reg1136 : reg1034)}));
                    end
                  reg1138 <= $unsigned($signed((~$unsigned(reg1127))));
                  for (forvar1139 = (1'h0); (forvar1139 < (2'h3)); forvar1139 = (forvar1139 + (1'h1)))
                    begin
                      reg1140 <= {$signed(forvar1120[(4'h9):(2'h2)])};
                      reg1141 <= ($signed(forvar898) ^~ $unsigned($signed({reg1023})));
                      reg1142 <= $unsigned($unsigned($signed({reg1072})));
                    end
                  if ({({(8'hb8)} ? forvar1029 : reg899[(3'h4):(1'h1)])})
                    begin
                      reg1143 <= $unsigned((reg1137[(3'h6):(2'h3)] == forvar1120[(4'ha):(2'h2)]));
                      reg1144 <= forvar1078;
                      reg1145 <= ($signed((wire890 << (!reg982))) ?
                          $unsigned(($signed(reg978) < (reg1083 ^~ reg1119))) : (~($signed((8'hb3)) != (reg1149 ?
                              reg899 : reg1161))));
                    end
                  else
                    begin
                      reg1143 <= reg999[(1'h1):(1'h0)];
                      reg1144 <= (~|(~&reg991[(4'ha):(2'h3)]));
                      reg1145 <= (((~&forvar1022[(2'h2):(1'h0)]) ?
                          reg978[(4'h8):(1'h1)] : reg1071[(3'h6):(1'h0)]) << (|($signed(reg912) ?
                          reg1076 : reg969[(1'h0):(1'h0)])));
                    end
                end
              for (forvar1146 = (1'h0); (forvar1146 < (2'h2)); forvar1146 = (forvar1146 + (1'h1)))
                begin
                  reg1147 <= $signed((forvar1048 ?
                      forvar1139[(4'ha):(4'h8)] : forvar1125[(2'h3):(2'h3)]));
                  if (wire895[(3'h6):(3'h4)])
                    begin
                      reg1148 <= $signed($signed(($signed(reg1023) ?
                          (forvar971 ?
                              reg1051 : reg1027) : forvar1085[(4'h8):(2'h2)])));
                    end
                  else
                    begin
                      reg1148 <= ((reg1045 || reg1135[(4'h8):(2'h2)]) <= (8'hb0));
                      reg1149 <= (8'haf);
                      reg1150 <= ((!$unsigned((^reg964))) ^ reg1086);
                    end
                  if ((&forvar902[(3'h5):(1'h0)]))
                    begin
                      reg1151 <= {$unsigned((reg1162 ?
                              (reg935 ? forvar1132 : reg1131) : reg1109))};
                      reg1152 <= (forvar1080[(1'h0):(1'h0)] ?
                          (reg897[(1'h0):(1'h0)] && {reg988[(2'h3):(1'h0)]}) : (reg960 ?
                              $unsigned((reg997 || reg931)) : $signed($signed(reg1090))));
                    end
                  else
                    begin
                      reg1151 <= $unsigned((~^(~^{forvar1139})));
                      reg1152 <= ((-(|(!forvar902))) ?
                          reg950 : {(forvar1028[(4'hd):(3'h4)] >> $unsigned(reg1024))});
                      reg1153 <= $unsigned((|($signed(reg1111) ?
                          {reg979} : ((8'ha9) || reg1057))));
                      reg1154 <= (~$unsigned((forvar900 ?
                          reg1150[(2'h2):(1'h0)] : $unsigned(reg1068))));
                    end
                  for (forvar1155 = (1'h0); (forvar1155 < (1'h1)); forvar1155 = (forvar1155 + (1'h1)))
                    begin
                      reg1156 <= $unsigned(forvar1133);
                      reg1157 <= $signed(forvar1120);
                      reg1158 <= forvar1059;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1163 = (1'h0); (forvar1163 < (2'h2)); forvar1163 = (forvar1163 + (1'h1)))
        begin
          if ({{reg1142[(2'h3):(1'h0)]}})
            begin
              if ($signed($unsigned($signed({forvar1078}))))
                begin
                  if ({(+(((8'hba) == (8'hb0)) < forvar1030[(4'hb):(4'ha)]))})
                    begin
                      reg1164 <= $unsigned($signed(reg970));
                      reg1165 <= $signed((((forvar982 < forvar1065) ?
                          (reg1079 ?
                              reg1083 : reg956) : $unsigned(reg1077)) < forvar921[(1'h1):(1'h1)]));
                      reg1166 <= (8'h9d);
                      reg1167 <= reg1060;
                    end
                  else
                    begin
                      reg1164 <= $unsigned($signed((~|$signed(forvar1065))));
                      reg1165 <= reg1061[(3'h4):(2'h3)];
                    end
                  if ((^forvar932))
                    begin
                      reg1168 <= ($unsigned(((!(8'hb0)) - forvar1125[(1'h1):(1'h1)])) ?
                          $signed($unsigned((forvar919 && wire895))) : $signed(reg938));
                      reg1169 <= (($unsigned($signed((8'ha2))) ?
                          (8'ha6) : forvar1155[(4'ha):(2'h2)]) <= forvar1022);
                      reg1170 <= ($signed(reg1138[(3'h5):(2'h2)]) >>> reg960[(4'h8):(4'h8)]);
                      reg1171 <= (($signed($unsigned(reg1057)) >= ($signed(reg928) & $signed((8'hb3)))) < $unsigned((&(reg1035 ?
                          reg1147 : reg1102))));
                    end
                  else
                    begin
                      reg1168 <= $signed({((8'ha5) ?
                              ((8'hae) ?
                                  forvar897 : forvar920) : $unsigned(reg1130))});
                      reg1169 <= (-(({reg1132} ?
                          (forvar1028 ?
                              forvar1108 : forvar1156) : (forvar897 <= forvar1033)) ^ reg1052[(3'h6):(1'h1)]));
                      reg1170 <= ((|wire892[(1'h1):(1'h0)]) == reg1154);
                    end
                end
              else
                begin
                  reg1164 <= reg1103[(2'h2):(1'h0)];
                  for (forvar1165 = (1'h0); (forvar1165 < (2'h3)); forvar1165 = (forvar1165 + (1'h1)))
                    begin
                      reg1166 <= (~^$unsigned({$unsigned(reg1157)}));
                      reg1167 <= (&reg975);
                      reg1168 <= (!reg1111);
                      reg1169 <= (!$signed((+(forvar910 && forvar955))));
                    end
                  if ((($unsigned($unsigned(reg1140)) >>> $signed((forvar992 == reg1067))) ?
                      $unsigned(((forvar958 ?
                          forvar918 : reg1140) >>> $unsigned((8'haa)))) : {(8'ha1)}))
                    begin
                      reg1170 <= (reg954 ?
                          reg921 : $unsigned((^((8'ha5) <= reg971))));
                      reg1171 <= forvar1085;
                    end
                  else
                    begin
                      reg1170 <= (($unsigned(forvar918[(1'h0):(1'h0)]) ^~ $signed(reg927[(2'h3):(1'h1)])) ^~ forvar910);
                      reg1171 <= $signed(((reg1168[(3'h7):(3'h7)] < forvar1091[(2'h3):(1'h1)]) && ((-reg1028) ?
                          reg925 : (^forvar919))));
                      reg1172 <= $signed($unsigned(($signed(reg999) << {forvar1155})));
                    end
                  if ($unsigned(reg919[(3'h5):(3'h5)]))
                    begin
                      reg1173 <= ($unsigned(({(8'hb8)} ?
                              $signed(forvar1107) : reg902)) ?
                          reg926 : ($unsigned((!reg1042)) ?
                              (-(&reg1028)) : (reg1154 ?
                                  $unsigned(reg1165) : (reg996 ?
                                      reg1044 : reg1171))));
                      reg1174 <= {{{(^reg1033)}}};
                      reg1175 <= (-(((+reg948) ?
                          forvar1130[(4'h8):(1'h0)] : (8'hb8)) >> $unsigned(((8'hb9) < reg1039))));
                    end
                  else
                    begin
                      reg1173 <= reg1051;
                      reg1174 <= $unsigned((-(8'hb0)));
                      reg1175 <= reg1136;
                      reg1176 <= (^forvar1107);
                    end
                end
            end
          else
            begin
              for (forvar1164 = (1'h0); (forvar1164 < (2'h3)); forvar1164 = (forvar1164 + (1'h1)))
                begin
                  if (forvar1036[(4'hb):(3'h4)])
                    begin
                      reg1165 <= reg1064[(2'h2):(1'h0)];
                      reg1166 <= forvar1139;
                      reg1167 <= {$signed($unsigned(((8'ha9) ?
                              (8'h9f) : reg931)))};
                      reg1168 <= $signed((8'h9d));
                    end
                  else
                    begin
                      reg1165 <= ({$unsigned(reg911[(1'h0):(1'h0)])} ?
                          (^{reg954}) : (^~reg914));
                      reg1166 <= (($unsigned(reg1033[(2'h2):(2'h2)]) << forvar919[(2'h2):(2'h2)]) <<< $unsigned((+{forvar992})));
                      reg1167 <= ((~^(~&$signed(forvar1109))) ?
                          ($signed((~^(8'hae))) >> $signed((reg1053 > forvar918))) : (((|forvar1130) ?
                              $unsigned(forvar938) : forvar942[(4'h8):(4'h8)]) ^~ reg1146));
                      reg1168 <= $signed(reg1104);
                    end
                end
              if ((&(!reg971[(1'h1):(1'h1)])))
                begin
                  for (forvar1169 = (1'h0); (forvar1169 < (2'h2)); forvar1169 = (forvar1169 + (1'h1)))
                    begin
                      reg1170 <= ((forvar953 ^ (&forvar1055[(4'h8):(2'h2)])) << $signed({$unsigned(reg934)}));
                      reg1171 <= $signed(($signed(reg1105) ^~ (reg1033[(1'h1):(1'h1)] ?
                          (!forvar1059) : (reg1051 >>> reg1025))));
                      reg1172 <= ($unsigned((&(reg907 ?
                          (8'hb5) : reg1022))) > (^~($unsigned(wire891) + (reg1123 >= reg1132))));
                    end
                  if ($unsigned((((~|reg1137) * $unsigned(reg1058)) ?
                      $unsigned((reg948 ?
                          reg964 : reg980)) : $signed((reg1065 > forvar946)))))
                    begin
                      reg1173 <= reg1030;
                      reg1174 <= (8'ha8);
                      reg1175 <= $unsigned($signed(forvar1020));
                    end
                  else
                    begin
                      reg1173 <= ({{(forvar1133 ?
                                  reg1093 : reg1165)}} ~^ (~|(~^wire894[(1'h1):(1'h1)])));
                      reg1174 <= $signed(reg1095);
                      reg1175 <= $signed(reg918);
                    end
                  reg1176 <= $unsigned(forvar941);
                end
              else
                begin
                  if ($signed(reg911))
                    begin
                      reg1169 <= ($unsigned(reg1107[(1'h0):(1'h0)]) ?
                          forvar984[(3'h5):(3'h4)] : reg1062);
                      reg1170 <= {{reg1152}};
                      reg1171 <= $signed(reg902);
                      reg1172 <= (($unsigned((reg953 > reg908)) ?
                              reg1098 : (~|(forvar952 ^~ (8'hab)))) ?
                          forvar998[(4'h8):(2'h3)] : $unsigned($signed(reg1139)));
                    end
                  else
                    begin
                      reg1169 <= (reg1105[(2'h3):(1'h1)] ?
                          (reg1099 ?
                              ((8'haa) ?
                                  (reg961 && reg1039) : (8'hb6)) : (forvar1048[(2'h3):(1'h0)] ?
                                  (8'hb6) : (~reg938))) : $signed(reg937[(1'h1):(1'h1)]));
                      reg1170 <= $unsigned((forvar902[(3'h4):(3'h4)] ~^ (8'hb7)));
                      reg1171 <= {(+forvar1089)};
                    end
                end
              for (forvar1177 = (1'h0); (forvar1177 < (1'h0)); forvar1177 = (forvar1177 + (1'h1)))
                begin
                  for (forvar1178 = (1'h0); (forvar1178 < (2'h2)); forvar1178 = (forvar1178 + (1'h1)))
                    begin
                      reg1179 <= $unsigned({forvar987});
                      reg1180 <= (reg1112 ?
                          $unsigned((reg904[(1'h0):(1'h0)] ?
                              (!reg1157) : {forvar1143})) : ((~^((8'hb3) >>> reg987)) ?
                              ($unsigned(reg1077) != $unsigned(reg1155)) : (-$unsigned((8'hb8)))));
                      reg1181 <= forvar1091;
                    end
                  if ($unsigned($signed(reg975)))
                    begin
                      reg1182 <= {$signed($signed($signed(reg910)))};
                      reg1183 <= ($signed((reg1138 <<< (forvar1126 ?
                              reg988 : reg905))) ?
                          (~|$unsigned((8'hb0))) : (^(!reg1165)));
                    end
                  else
                    begin
                      reg1182 <= {reg901[(1'h1):(1'h0)]};
                      reg1183 <= $unsigned((~&$signed($unsigned((8'h9c)))));
                      reg1184 <= ((~^((reg939 ? forvar902 : reg1103) ?
                              ((8'hb7) && forvar1089) : (!forvar1040))) ?
                          reg1136 : $signed(((^~forvar900) <<< (forvar1060 << reg1044))));
                    end
                  for (forvar1185 = (1'h0); (forvar1185 < (2'h2)); forvar1185 = (forvar1185 + (1'h1)))
                    begin
                      reg1186 <= ((8'ha6) || {((reg1156 ^~ forvar1049) ?
                              (~|forvar1074) : $signed(reg1106))});
                      reg1187 <= {(8'h9c)};
                    end
                  if ((~^reg1133[(1'h1):(1'h1)]))
                    begin
                      reg1188 <= ($unsigned($signed(reg1069)) != reg1035);
                      reg1189 <= reg1105;
                    end
                  else
                    begin
                      reg1188 <= $signed(reg1135);
                      reg1189 <= (-{forvar942});
                      reg1190 <= (forvar953[(1'h0):(1'h0)] ?
                          (($unsigned(reg1100) | ((8'hb9) <<< (8'hb7))) ?
                              ((&reg1034) | reg1100) : $signed($signed(reg1157))) : $signed($signed((forvar1044 != reg1158))));
                    end
                end
            end
          if (forvar1145)
            begin
              if (reg983)
                begin
                  reg1191 <= (-forvar897[(1'h0):(1'h0)]);
                  for (forvar1192 = (1'h0); (forvar1192 < (2'h3)); forvar1192 = (forvar1192 + (1'h1)))
                    begin
                      reg1193 <= ($signed({reg990[(3'h4):(3'h4)]}) ?
                          $unsigned((^(reg949 ?
                              reg1098 : reg1098))) : ((forvar1097 ?
                              reg1044[(4'h9):(2'h2)] : reg1046) != reg945[(1'h0):(1'h0)]));
                      reg1194 <= reg966;
                      reg1195 <= reg1109;
                      reg1196 <= forvar1049;
                    end
                  if (reg975)
                    begin
                      reg1197 <= $signed((((reg1044 | reg914) << (-reg918)) != (forvar958[(3'h7):(2'h2)] ?
                          (|forvar898) : (8'ha6))));
                      reg1198 <= (~&($signed($signed(forvar1109)) && $signed((reg980 ?
                          reg1079 : reg1134))));
                      reg1199 <= reg1043;
                      reg1200 <= $signed($signed({reg1147}));
                    end
                  else
                    begin
                      reg1197 <= reg915[(3'h4):(1'h1)];
                      reg1198 <= (~|({(forvar1075 != reg1154)} + reg966));
                    end
                  reg1201 <= forvar908;
                end
              else
                begin
                  if ($signed($signed((~$signed(reg955)))))
                    begin
                      reg1191 <= ($unsigned((8'ha8)) ?
                          reg1101 : reg1121[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg1191 <= reg1155;
                    end
                end
              for (forvar1202 = (1'h0); (forvar1202 < (2'h2)); forvar1202 = (forvar1202 + (1'h1)))
                begin
                  for (forvar1203 = (1'h0); (forvar1203 < (1'h0)); forvar1203 = (forvar1203 + (1'h1)))
                    begin
                      reg1204 <= forvar1202[(1'h1):(1'h0)];
                      reg1205 <= (^~$unsigned(reg1028));
                      reg1206 <= (reg1033[(2'h3):(2'h3)] ?
                          (((&reg1149) * (&reg1070)) > reg955[(1'h0):(1'h0)]) : {$signed((reg1051 + (8'ha9)))});
                    end
                  for (forvar1207 = (1'h0); (forvar1207 < (1'h0)); forvar1207 = (forvar1207 + (1'h1)))
                    begin
                      reg1208 <= $signed(reg1143);
                    end
                end
              for (forvar1209 = (1'h0); (forvar1209 < (2'h3)); forvar1209 = (forvar1209 + (1'h1)))
                begin
                  reg1210 <= (^reg1208);
                  if ({forvar1125[(3'h4):(2'h3)]})
                    begin
                      reg1211 <= $signed($unsigned(((~|forvar908) < reg1044)));
                      reg1212 <= reg1206;
                    end
                  else
                    begin
                      reg1211 <= $unsigned((8'h9c));
                      reg1212 <= (8'h9e);
                    end
                  if ((((~|$signed(reg950)) >>> (!$signed(reg936))) * (8'ha6)))
                    begin
                      reg1213 <= reg1142;
                    end
                  else
                    begin
                      reg1213 <= {reg1175};
                      reg1214 <= ($signed((&(reg935 <= reg1143))) ?
                          reg951 : {wire893});
                    end
                  for (forvar1215 = (1'h0); (forvar1215 < (2'h2)); forvar1215 = (forvar1215 + (1'h1)))
                    begin
                      reg1216 <= $unsigned((((+reg1193) == $signed(reg986)) == wire894[(3'h6):(3'h4)]));
                    end
                end
              reg1217 <= reg1027[(1'h1):(1'h1)];
            end
          else
            begin
              reg1191 <= (^~({$unsigned(reg939)} | $signed(forvar1177[(1'h1):(1'h0)])));
            end
        end
    end
  assign wire1218 = $signed(forvar1143[(4'hc):(3'h7)]);
  module1219 modinst1745 (.wire1224(reg1071), .wire1222(forvar897), .wire1220(reg1130), .clk(clk), .wire1223(reg954), .y(wire1744), .wire1221(reg1093));
  assign wire1746 = reg956;
  always
    @(posedge clk) begin
      for (forvar1747 = (1'h0); (forvar1747 < (2'h2)); forvar1747 = (forvar1747 + (1'h1)))
        begin
          for (forvar1748 = (1'h0); (forvar1748 < (2'h2)); forvar1748 = (forvar1748 + (1'h1)))
            begin
              for (forvar1749 = (1'h0); (forvar1749 < (1'h0)); forvar1749 = (forvar1749 + (1'h1)))
                begin
                  reg1750 <= $unsigned(reg924);
                  for (forvar1751 = (1'h0); (forvar1751 < (1'h0)); forvar1751 = (forvar1751 + (1'h1)))
                    begin
                      reg1752 <= (reg1077 ^ $signed(((forvar960 ?
                          wire1746 : forvar1060) == (reg958 || reg936))));
                      reg1753 <= (reg1057 >> ($unsigned((^~reg1057)) <= $signed((8'hb8))));
                      reg1754 <= reg923[(1'h0):(1'h0)];
                    end
                  reg1755 <= (+reg1134);
                end
              reg1756 <= {(({forvar1159} ?
                          forvar1078 : (forvar1054 ? reg1127 : reg1046)) ?
                      reg976 : (reg952[(4'hc):(4'h9)] && wire891))};
              reg1757 <= (forvar951 ? reg922 : $signed(reg903));
            end
        end
    end
  assign wire1758 = ({(((8'ha5) ^ reg988) ~^ reg1125)} ?
                        (!$signed({(8'ha6)})) : {forvar938});
  module1759 modinst4166 (.y(wire4165), .wire1763(reg973), .wire1762(reg902), .wire1761(reg1082), .wire1760(reg928), .clk(clk));
  assign wire4167 = $signed((reg924[(4'ha):(3'h4)] ?
                        ((reg967 ? reg1081 : reg1112) ?
                            $signed(reg1145) : ((8'ha5) ?
                                reg1138 : reg1083)) : $signed($unsigned(forvar1143))));
  assign wire4168 = reg988;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1759  (y, clk, wire1763, wire1762, wire1761, wire1760);
  output wire [(32'h23aa):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire1763;
  input wire [(4'h9):(1'h0)] wire1762;
  input wire signed [(4'hf):(1'h0)] wire1761;
  input wire [(5'h10):(1'h0)] wire1760;
  wire signed [(4'h9):(1'h0)] wire4164;
  reg [(3'h6):(1'h0)] reg4163 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4156 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4154 = (1'h0);
  reg [(4'hf):(1'h0)] reg4152 = (1'h0);
  reg [(3'h5):(1'h0)] reg4162 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4161 = (1'h0);
  reg [(3'h7):(1'h0)] reg4160 = (1'h0);
  reg [(3'h7):(1'h0)] reg4159 = (1'h0);
  reg [(4'hc):(1'h0)] reg4158 = (1'h0);
  reg [(5'h10):(1'h0)] reg4157 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4156 = (1'h0);
  reg [(4'he):(1'h0)] reg4155 = (1'h0);
  reg [(4'h8):(1'h0)] reg4154 = (1'h0);
  reg [(3'h4):(1'h0)] reg4153 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4152 = (1'h0);
  reg [(4'hb):(1'h0)] reg4151 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4150 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4149 = (1'h0);
  reg [(4'h8):(1'h0)] reg4148 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4147 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4146 = (1'h0);
  reg [(4'he):(1'h0)] reg4145 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4144 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4143 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4142 = (1'h0);
  reg [(2'h3):(1'h0)] reg4141 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4140 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4139 = (1'h0);
  reg [(4'hb):(1'h0)] reg4138 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4137 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4136 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4135 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4134 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4133 = (1'h0);
  reg [(2'h2):(1'h0)] reg4122 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4132 = (1'h0);
  reg [(3'h4):(1'h0)] reg4131 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4128 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4130 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4129 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4128 = (1'h0);
  reg [(2'h2):(1'h0)] reg4127 = (1'h0);
  reg [(4'hf):(1'h0)] reg4126 = (1'h0);
  reg [(2'h3):(1'h0)] reg4125 = (1'h0);
  reg [(4'he):(1'h0)] reg4124 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4123 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4122 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4121 = (1'h0);
  reg [(5'h10):(1'h0)] reg4120 = (1'h0);
  reg [(3'h6):(1'h0)] reg4119 = (1'h0);
  reg [(3'h5):(1'h0)] reg4118 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4117 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4116 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4116 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4115 = (1'h0);
  reg [(4'hb):(1'h0)] reg4114 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4113 = (1'h0);
  reg [(4'h8):(1'h0)] reg4112 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4111 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4110 = (1'h0);
  reg [(4'h8):(1'h0)] reg4098 = (1'h0);
  reg [(5'h10):(1'h0)] reg4093 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4090 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4103 = (1'h0);
  reg [(3'h7):(1'h0)] reg4109 = (1'h0);
  reg [(4'he):(1'h0)] reg4108 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4107 = (1'h0);
  reg [(4'hb):(1'h0)] reg4106 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4105 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4104 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4103 = (1'h0);
  reg [(3'h4):(1'h0)] reg4102 = (1'h0);
  reg [(5'h10):(1'h0)] reg4101 = (1'h0);
  reg [(2'h2):(1'h0)] reg4100 = (1'h0);
  reg [(4'hb):(1'h0)] reg4099 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4098 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4097 = (1'h0);
  reg [(3'h6):(1'h0)] reg4096 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4095 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4094 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4093 = (1'h0);
  reg [(3'h6):(1'h0)] reg4092 = (1'h0);
  reg [(2'h2):(1'h0)] reg4091 = (1'h0);
  reg [(3'h7):(1'h0)] reg4090 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4086 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4084 = (1'h0);
  reg [(4'ha):(1'h0)] reg4082 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4078 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4089 = (1'h0);
  reg [(5'h10):(1'h0)] reg4088 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4087 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4086 = (1'h0);
  reg [(4'h9):(1'h0)] reg4085 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4084 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4083 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4082 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4081 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4080 = (1'h0);
  reg [(5'h10):(1'h0)] reg4079 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4078 = (1'h0);
  reg [(3'h7):(1'h0)] reg4077 = (1'h0);
  reg [(2'h3):(1'h0)] reg4076 = (1'h0);
  reg [(3'h4):(1'h0)] reg4075 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4074 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4073 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4072 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4071 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4070 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4069 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4068 = (1'h0);
  reg [(4'h9):(1'h0)] reg4067 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4066 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4065 = (1'h0);
  reg [(4'hc):(1'h0)] reg4064 = (1'h0);
  reg [(4'h9):(1'h0)] reg4063 = (1'h0);
  reg [(4'hd):(1'h0)] reg4062 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4061 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4060 = (1'h0);
  reg [(4'hb):(1'h0)] reg4059 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4058 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4057 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4056 = (1'h0);
  reg [(4'hd):(1'h0)] reg4055 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4054 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4053 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4052 = (1'h0);
  reg [(4'hc):(1'h0)] reg4051 = (1'h0);
  reg [(4'ha):(1'h0)] reg4050 = (1'h0);
  reg [(3'h7):(1'h0)] reg4049 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4048 = (1'h0);
  reg [(4'hc):(1'h0)] reg4047 = (1'h0);
  reg [(4'hd):(1'h0)] reg4046 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4045 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4044 = (1'h0);
  reg [(3'h7):(1'h0)] reg4043 = (1'h0);
  reg [(4'hd):(1'h0)] reg4042 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4041 = (1'h0);
  reg [(4'h8):(1'h0)] reg4040 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4027 = (1'h0);
  reg [(3'h4):(1'h0)] reg4039 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4038 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4037 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4036 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4035 = (1'h0);
  reg [(2'h3):(1'h0)] reg4034 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4033 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4032 = (1'h0);
  reg [(2'h3):(1'h0)] reg4031 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4030 = (1'h0);
  reg [(4'hc):(1'h0)] reg4029 = (1'h0);
  reg [(2'h3):(1'h0)] reg4028 = (1'h0);
  reg [(4'hc):(1'h0)] reg4026 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4027 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4026 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4025 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4024 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4023 = (1'h0);
  reg [(4'hd):(1'h0)] reg4022 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4021 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4020 = (1'h0);
  wire [(3'h7):(1'h0)] wire4019;
  wire signed [(4'hb):(1'h0)] wire3601;
  reg signed [(4'hf):(1'h0)] reg3493 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3491 = (1'h0);
  reg [(3'h7):(1'h0)] reg3489 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3486 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3483 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3477 = (1'h0);
  reg [(4'he):(1'h0)] forvar3476 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3501 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3500 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3499 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3498 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3497 = (1'h0);
  reg [(4'he):(1'h0)] reg3496 = (1'h0);
  reg [(2'h3):(1'h0)] reg3495 = (1'h0);
  reg [(4'hf):(1'h0)] reg3494 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3493 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3492 = (1'h0);
  reg [(3'h4):(1'h0)] reg3491 = (1'h0);
  reg [(2'h3):(1'h0)] reg3490 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3489 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3488 = (1'h0);
  reg [(4'hb):(1'h0)] reg3487 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3486 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3485 = (1'h0);
  reg [(4'h9):(1'h0)] reg3484 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3483 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3482 = (1'h0);
  reg [(4'he):(1'h0)] reg3473 = (1'h0);
  reg [(2'h2):(1'h0)] reg3481 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3480 = (1'h0);
  reg [(2'h3):(1'h0)] reg3479 = (1'h0);
  reg [(2'h2):(1'h0)] reg3478 = (1'h0);
  reg [(4'hf):(1'h0)] reg3477 = (1'h0);
  reg [(4'hc):(1'h0)] reg3476 = (1'h0);
  reg [(4'hd):(1'h0)] reg3475 = (1'h0);
  reg [(4'hc):(1'h0)] reg3474 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3473 = (1'h0);
  reg [(2'h2):(1'h0)] reg3472 = (1'h0);
  reg [(2'h3):(1'h0)] reg3471 = (1'h0);
  reg [(5'h10):(1'h0)] reg3470 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3469 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3466 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3464 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3461 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3468 = (1'h0);
  reg [(4'h9):(1'h0)] reg3467 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3466 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3465 = (1'h0);
  reg [(4'ha):(1'h0)] reg3464 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3463 = (1'h0);
  reg [(5'h10):(1'h0)] reg3462 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3461 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3460 = (1'h0);
  reg [(2'h2):(1'h0)] reg3459 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3458 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3457 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3456 = (1'h0);
  reg [(4'he):(1'h0)] reg3455 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3454 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3453 = (1'h0);
  reg [(3'h5):(1'h0)] reg3452 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3451 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3450 = (1'h0);
  reg [(4'ha):(1'h0)] reg3449 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3448 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3447 = (1'h0);
  reg [(2'h3):(1'h0)] reg3446 = (1'h0);
  reg [(4'ha):(1'h0)] reg3445 = (1'h0);
  reg [(4'h9):(1'h0)] reg3444 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3443 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3442 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3441 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3428 = (1'h0);
  reg [(2'h3):(1'h0)] reg3440 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3439 = (1'h0);
  reg [(4'he):(1'h0)] reg3438 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3437 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3436 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3435 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3434 = (1'h0);
  reg [(3'h6):(1'h0)] reg3433 = (1'h0);
  reg [(4'h9):(1'h0)] reg3432 = (1'h0);
  reg [(4'h9):(1'h0)] reg3431 = (1'h0);
  reg [(4'hf):(1'h0)] reg3430 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3429 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3428 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3427 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3426 = (1'h0);
  reg [(4'hc):(1'h0)] reg3425 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3424 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3423 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3422 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3421 = (1'h0);
  reg [(2'h2):(1'h0)] reg3420 = (1'h0);
  reg [(4'hb):(1'h0)] reg3419 = (1'h0);
  reg [(3'h5):(1'h0)] reg3418 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3417 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3416 = (1'h0);
  reg [(4'hd):(1'h0)] reg3415 = (1'h0);
  reg [(3'h4):(1'h0)] reg3414 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3413 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3408 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3412 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3411 = (1'h0);
  reg [(3'h4):(1'h0)] reg3410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3409 = (1'h0);
  reg [(4'he):(1'h0)] reg3408 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3407 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3404 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3402 = (1'h0);
  reg [(3'h5):(1'h0)] reg3401 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3395 = (1'h0);
  reg [(4'h8):(1'h0)] reg3406 = (1'h0);
  reg [(4'ha):(1'h0)] reg3405 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3404 = (1'h0);
  reg [(4'hc):(1'h0)] reg3403 = (1'h0);
  reg [(5'h10):(1'h0)] reg3402 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3401 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3400 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3399 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3398 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3397 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3396 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3395 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3394 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3393 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3382 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3392 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3391 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3390 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3389 = (1'h0);
  reg [(4'ha):(1'h0)] reg3388 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3387 = (1'h0);
  reg [(2'h2):(1'h0)] reg3386 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3385 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3384 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3383 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3382 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3381 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3367 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3365 = (1'h0);
  reg [(4'hd):(1'h0)] reg3363 = (1'h0);
  reg [(3'h4):(1'h0)] reg3362 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3361 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3380 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3379 = (1'h0);
  reg [(5'h10):(1'h0)] reg3378 = (1'h0);
  reg [(3'h5):(1'h0)] reg3377 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3376 = (1'h0);
  reg [(4'hb):(1'h0)] reg3375 = (1'h0);
  reg [(4'hf):(1'h0)] reg3374 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3372 = (1'h0);
  reg [(2'h3):(1'h0)] reg3373 = (1'h0);
  reg [(3'h7):(1'h0)] reg3372 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3371 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3370 = (1'h0);
  reg [(4'hb):(1'h0)] reg3369 = (1'h0);
  reg [(4'hf):(1'h0)] reg3368 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3367 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3366 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3365 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3364 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3363 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3362 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3361 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3360 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3359 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3358 = (1'h0);
  reg [(2'h2):(1'h0)] reg3357 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3356 = (1'h0);
  reg [(2'h2):(1'h0)] reg3355 = (1'h0);
  reg [(4'h9):(1'h0)] reg3354 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3353 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3352 = (1'h0);
  reg [(3'h6):(1'h0)] reg3351 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3350 = (1'h0);
  reg [(3'h6):(1'h0)] reg3349 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3348 = (1'h0);
  reg [(4'he):(1'h0)] reg3347 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3346 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3345 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3344 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3343 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3342 = (1'h0);
  reg [(3'h4):(1'h0)] reg3341 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3340 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3339 = (1'h0);
  reg [(4'h8):(1'h0)] reg3338 = (1'h0);
  reg [(4'hf):(1'h0)] reg3337 = (1'h0);
  reg [(4'h8):(1'h0)] reg3336 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3335 = (1'h0);
  reg [(4'h8):(1'h0)] reg3334 = (1'h0);
  reg [(2'h2):(1'h0)] reg3333 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3332 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3331 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3330 = (1'h0);
  reg [(3'h4):(1'h0)] reg3329 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3328 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3327 = (1'h0);
  reg [(3'h5):(1'h0)] reg3326 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3325 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3324 = (1'h0);
  reg [(3'h6):(1'h0)] reg3323 = (1'h0);
  reg [(4'hd):(1'h0)] reg3322 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3321 = (1'h0);
  reg [(4'hc):(1'h0)] reg3320 = (1'h0);
  reg [(2'h2):(1'h0)] reg3319 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3318 = (1'h0);
  reg [(4'hf):(1'h0)] reg3317 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3316 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3315 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3314 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3313 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3312 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3311 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3310 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3309 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3308 = (1'h0);
  reg [(3'h5):(1'h0)] reg3307 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3306 = (1'h0);
  reg [(2'h3):(1'h0)] reg3305 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3304 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3303 = (1'h0);
  reg [(3'h7):(1'h0)] reg3302 = (1'h0);
  reg [(4'h8):(1'h0)] reg3301 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3300 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3299 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3298 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3297 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3296 = (1'h0);
  reg [(4'h8):(1'h0)] reg3295 = (1'h0);
  reg [(3'h4):(1'h0)] reg3294 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3293 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3292 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3291 = (1'h0);
  reg [(4'hd):(1'h0)] reg3290 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3289 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3288 = (1'h0);
  reg [(4'ha):(1'h0)] reg3287 = (1'h0);
  reg [(4'he):(1'h0)] forvar3285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3284 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3283 = (1'h0);
  reg [(4'hb):(1'h0)] reg3280 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3274 = (1'h0);
  reg [(4'h8):(1'h0)] reg3286 = (1'h0);
  reg [(3'h4):(1'h0)] reg3285 = (1'h0);
  reg [(4'he):(1'h0)] forvar3284 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3283 = (1'h0);
  reg [(5'h10):(1'h0)] reg3282 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3281 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3280 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3279 = (1'h0);
  reg [(3'h6):(1'h0)] reg3278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3277 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3276 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3275 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3274 = (1'h0);
  reg [(4'he):(1'h0)] reg3273 = (1'h0);
  reg [(4'ha):(1'h0)] reg3272 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3271 = (1'h0);
  reg [(4'ha):(1'h0)] reg3270 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3269 = (1'h0);
  reg [(4'ha):(1'h0)] reg3268 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3267 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3266 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3265 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3264 = (1'h0);
  reg [(4'hc):(1'h0)] reg3263 = (1'h0);
  reg [(4'hf):(1'h0)] reg3262 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3261 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3260 = (1'h0);
  reg [(3'h7):(1'h0)] reg3259 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3258 = (1'h0);
  reg [(3'h6):(1'h0)] reg3257 = (1'h0);
  reg [(2'h3):(1'h0)] reg3256 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3255 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3254 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3253 = (1'h0);
  reg [(4'h9):(1'h0)] reg3237 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3232 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3231 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3228 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3224 = (1'h0);
  reg [(4'ha):(1'h0)] reg3252 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3251 = (1'h0);
  reg [(4'h9):(1'h0)] reg3250 = (1'h0);
  reg [(2'h2):(1'h0)] reg3249 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3248 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3247 = (1'h0);
  reg [(4'he):(1'h0)] reg3246 = (1'h0);
  reg [(2'h3):(1'h0)] reg3245 = (1'h0);
  reg [(4'h8):(1'h0)] reg3244 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3243 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3242 = (1'h0);
  reg [(3'h5):(1'h0)] reg3241 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3240 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3239 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3238 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3237 = (1'h0);
  reg [(4'he):(1'h0)] reg3236 = (1'h0);
  reg [(4'hf):(1'h0)] reg3235 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3234 = (1'h0);
  reg [(4'h8):(1'h0)] reg3233 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3232 = (1'h0);
  reg [(2'h3):(1'h0)] reg3231 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3230 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3229 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3228 = (1'h0);
  reg [(4'he):(1'h0)] reg3227 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3226 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3225 = (1'h0);
  reg [(4'he):(1'h0)] forvar3224 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3223 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3205 = (1'h0);
  reg [(3'h6):(1'h0)] reg3200 = (1'h0);
  reg [(4'hd):(1'h0)] reg3222 = (1'h0);
  reg [(4'h8):(1'h0)] reg3221 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3220 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3219 = (1'h0);
  reg [(4'hb):(1'h0)] reg3217 = (1'h0);
  reg [(2'h3):(1'h0)] reg3215 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3218 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3217 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3216 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3215 = (1'h0);
  reg [(3'h5):(1'h0)] reg3214 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3213 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3212 = (1'h0);
  reg [(4'hb):(1'h0)] reg3211 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3210 = (1'h0);
  reg [(4'ha):(1'h0)] reg3209 = (1'h0);
  reg [(3'h6):(1'h0)] reg3208 = (1'h0);
  reg [(4'hc):(1'h0)] reg3203 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3207 = (1'h0);
  reg [(3'h6):(1'h0)] reg3206 = (1'h0);
  reg [(4'h8):(1'h0)] reg3205 = (1'h0);
  reg [(4'hf):(1'h0)] reg3204 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3203 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3202 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3201 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3200 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3199 = (1'h0);
  reg [(2'h3):(1'h0)] reg3198 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3197 = (1'h0);
  reg [(4'h9):(1'h0)] reg3196 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3195 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3194 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3193 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3192 = (1'h0);
  reg [(3'h5):(1'h0)] reg3191 = (1'h0);
  reg [(4'hb):(1'h0)] reg3190 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3189 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3188 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3187 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3186 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3185 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3184 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3183 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire3182;
  reg [(4'ha):(1'h0)] reg3181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3177 = (1'h0);
  reg [(3'h7):(1'h0)] reg3180 = (1'h0);
  reg [(4'hb):(1'h0)] reg3179 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3178 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3177 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3176 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3175 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3174 = (1'h0);
  reg [(2'h2):(1'h0)] reg3173 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3172 = (1'h0);
  reg [(4'h9):(1'h0)] reg3171 = (1'h0);
  reg [(4'h9):(1'h0)] reg3170 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3169 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3168 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3167 = (1'h0);
  reg [(3'h7):(1'h0)] reg3166 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3165 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3164 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3163 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3120 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3112 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3110 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3109 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3108 = (1'h0);
  reg [(4'he):(1'h0)] reg3103 = (1'h0);
  reg [(3'h5):(1'h0)] reg3101 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3095 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3091 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3162 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3161 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3160 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3159 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3158 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3157 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3156 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3155 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3154 = (1'h0);
  reg [(2'h2):(1'h0)] reg3153 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3152 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3151 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3150 = (1'h0);
  reg [(4'hc):(1'h0)] reg3149 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3148 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3147 = (1'h0);
  reg [(3'h4):(1'h0)] reg3143 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3142 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3141 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3139 = (1'h0);
  reg [(5'h10):(1'h0)] reg3146 = (1'h0);
  reg [(4'hf):(1'h0)] reg3145 = (1'h0);
  reg [(4'hf):(1'h0)] reg3144 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3143 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3142 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3141 = (1'h0);
  reg [(4'ha):(1'h0)] reg3140 = (1'h0);
  reg [(4'ha):(1'h0)] reg3139 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3138 = (1'h0);
  reg [(4'hb):(1'h0)] reg3130 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3137 = (1'h0);
  reg [(4'ha):(1'h0)] reg3136 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3135 = (1'h0);
  reg [(4'hc):(1'h0)] reg3134 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3133 = (1'h0);
  reg [(4'h9):(1'h0)] reg3132 = (1'h0);
  reg [(3'h4):(1'h0)] reg3131 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3130 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3129 = (1'h0);
  reg [(3'h6):(1'h0)] reg3128 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3127 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3126 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3125 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3124 = (1'h0);
  reg [(4'hd):(1'h0)] reg3123 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3122 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3121 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3120 = (1'h0);
  reg [(4'hf):(1'h0)] reg3119 = (1'h0);
  reg [(4'h8):(1'h0)] reg3118 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3117 = (1'h0);
  reg [(2'h2):(1'h0)] reg3116 = (1'h0);
  reg [(4'h8):(1'h0)] reg3115 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3114 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3113 = (1'h0);
  reg [(3'h6):(1'h0)] reg3112 = (1'h0);
  reg [(4'hd):(1'h0)] reg3111 = (1'h0);
  reg [(4'h8):(1'h0)] reg3110 = (1'h0);
  reg [(3'h6):(1'h0)] reg3109 = (1'h0);
  reg [(4'hb):(1'h0)] reg3108 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3107 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3106 = (1'h0);
  reg [(4'he):(1'h0)] reg3105 = (1'h0);
  reg [(3'h5):(1'h0)] reg3104 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3103 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3102 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3101 = (1'h0);
  reg [(4'h9):(1'h0)] reg3100 = (1'h0);
  reg [(3'h6):(1'h0)] reg3099 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3098 = (1'h0);
  reg [(4'hb):(1'h0)] reg3097 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3096 = (1'h0);
  reg [(3'h5):(1'h0)] reg3095 = (1'h0);
  reg [(3'h7):(1'h0)] reg3094 = (1'h0);
  reg [(3'h6):(1'h0)] reg3093 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3092 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3091 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3090 = (1'h0);
  reg [(4'h8):(1'h0)] reg3089 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3088 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3087 = (1'h0);
  reg [(4'hb):(1'h0)] reg3086 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3084 = (1'h0);
  reg [(4'h8):(1'h0)] reg3081 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3085 = (1'h0);
  reg [(2'h3):(1'h0)] reg3084 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3083 = (1'h0);
  reg [(2'h2):(1'h0)] reg3082 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3081 = (1'h0);
  reg [(4'h9):(1'h0)] reg3080 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3079 = (1'h0);
  reg [(4'h8):(1'h0)] reg3078 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3077 = (1'h0);
  reg [(4'hd):(1'h0)] reg3076 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3075 = (1'h0);
  reg [(4'hd):(1'h0)] reg3074 = (1'h0);
  reg [(2'h2):(1'h0)] reg3073 = (1'h0);
  reg [(3'h7):(1'h0)] reg3072 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3071 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3070 = (1'h0);
  reg [(3'h5):(1'h0)] reg3069 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3068 = (1'h0);
  reg [(4'he):(1'h0)] reg3067 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3066 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3065 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3064 = (1'h0);
  reg [(2'h3):(1'h0)] reg3063 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3062 = (1'h0);
  reg [(4'he):(1'h0)] forvar3061 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3060 = (1'h0);
  reg [(4'h8):(1'h0)] reg3052 = (1'h0);
  reg [(4'hc):(1'h0)] reg3047 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3059 = (1'h0);
  reg [(3'h4):(1'h0)] reg3058 = (1'h0);
  reg [(3'h7):(1'h0)] reg3057 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3056 = (1'h0);
  reg [(4'h8):(1'h0)] reg3055 = (1'h0);
  reg [(4'h8):(1'h0)] reg3054 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3053 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3052 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3051 = (1'h0);
  reg [(4'he):(1'h0)] reg3050 = (1'h0);
  reg [(3'h4):(1'h0)] reg3049 = (1'h0);
  reg [(4'ha):(1'h0)] reg3048 = (1'h0);
  reg [(4'he):(1'h0)] forvar3047 = (1'h0);
  reg [(4'hc):(1'h0)] reg3046 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3045 = (1'h0);
  reg [(4'ha):(1'h0)] reg3044 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3043 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3033 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3027 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3011 = (1'h0);
  reg [(4'he):(1'h0)] forvar3006 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3029 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3042 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3041 = (1'h0);
  reg [(4'h8):(1'h0)] reg3040 = (1'h0);
  reg [(4'ha):(1'h0)] reg3039 = (1'h0);
  reg [(4'hb):(1'h0)] reg3038 = (1'h0);
  reg [(4'h9):(1'h0)] reg3037 = (1'h0);
  reg [(5'h10):(1'h0)] reg3036 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3035 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3034 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3033 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3032 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3031 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3030 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3029 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3028 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3022 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3021 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3017 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3010 = (1'h0);
  reg [(3'h4):(1'h0)] reg3016 = (1'h0);
  reg [(4'hd):(1'h0)] reg3012 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3009 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3007 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3004 = (1'h0);
  reg [(4'hf):(1'h0)] reg3027 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3026 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3025 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3024 = (1'h0);
  reg [(2'h2):(1'h0)] reg3023 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3022 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3021 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3020 = (1'h0);
  reg [(4'hb):(1'h0)] reg3019 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3018 = (1'h0);
  reg [(5'h10):(1'h0)] reg3017 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3016 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3015 = (1'h0);
  reg [(4'hd):(1'h0)] reg3014 = (1'h0);
  reg [(4'h9):(1'h0)] reg3013 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3012 = (1'h0);
  reg [(3'h7):(1'h0)] reg3011 = (1'h0);
  reg [(3'h7):(1'h0)] reg3010 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3009 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3008 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3007 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3005 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3006 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3005 = (1'h0);
  reg [(3'h4):(1'h0)] reg3004 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire3003;
  wire [(4'h9):(1'h0)] wire3002;
  reg [(4'ha):(1'h0)] forvar2966 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2964 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2963 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2959 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2958 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2950 = (1'h0);
  reg [(4'he):(1'h0)] forvar2945 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2944 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2978 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2974 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2970 = (1'h0);
  reg [(3'h7):(1'h0)] reg2969 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2968 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3001 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3000 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2999 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2998 = (1'h0);
  reg [(3'h7):(1'h0)] reg2997 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2996 = (1'h0);
  reg [(4'hd):(1'h0)] reg2995 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2994 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2993 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2992 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2991 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2990 = (1'h0);
  reg [(2'h3):(1'h0)] reg2989 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2988 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2987 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2986 = (1'h0);
  reg [(4'hc):(1'h0)] reg2983 = (1'h0);
  reg [(4'hd):(1'h0)] reg2985 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2984 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2983 = (1'h0);
  reg [(4'hc):(1'h0)] reg2982 = (1'h0);
  reg [(4'ha):(1'h0)] reg2981 = (1'h0);
  reg [(5'h10):(1'h0)] reg2980 = (1'h0);
  reg [(4'hb):(1'h0)] reg2979 = (1'h0);
  reg [(4'he):(1'h0)] reg2978 = (1'h0);
  reg [(4'ha):(1'h0)] reg2977 = (1'h0);
  reg [(4'ha):(1'h0)] reg2976 = (1'h0);
  reg [(2'h2):(1'h0)] reg2975 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2974 = (1'h0);
  reg [(4'h9):(1'h0)] reg2973 = (1'h0);
  reg [(2'h3):(1'h0)] reg2972 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2971 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2970 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2969 = (1'h0);
  reg [(4'he):(1'h0)] forvar2968 = (1'h0);
  reg [(2'h2):(1'h0)] reg2967 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2966 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2965 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2964 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2963 = (1'h0);
  reg [(4'hc):(1'h0)] reg2962 = (1'h0);
  reg [(3'h6):(1'h0)] reg2961 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2960 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2959 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2958 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2957 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2956 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2955 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2953 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2948 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2947 = (1'h0);
  reg [(2'h3):(1'h0)] reg2943 = (1'h0);
  reg [(4'hb):(1'h0)] reg2955 = (1'h0);
  reg [(4'ha):(1'h0)] reg2954 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2953 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2952 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2951 = (1'h0);
  reg [(3'h6):(1'h0)] reg2950 = (1'h0);
  reg [(5'h10):(1'h0)] reg2949 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2948 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2947 = (1'h0);
  reg [(4'hc):(1'h0)] reg2946 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2945 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2944 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2943 = (1'h0);
  reg [(4'h9):(1'h0)] reg2942 = (1'h0);
  reg [(3'h5):(1'h0)] reg2941 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2940 = (1'h0);
  reg [(3'h4):(1'h0)] reg2939 = (1'h0);
  reg [(3'h5):(1'h0)] reg2938 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2937 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2931 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2936 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2935 = (1'h0);
  reg [(3'h7):(1'h0)] reg2934 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2933 = (1'h0);
  reg [(3'h4):(1'h0)] reg2932 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2931 = (1'h0);
  reg [(4'hd):(1'h0)] reg2930 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2919 = (1'h0);
  reg [(4'hb):(1'h0)] reg2927 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2925 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2922 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2920 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2929 = (1'h0);
  reg [(4'hc):(1'h0)] reg2928 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2927 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2926 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2925 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2917 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2924 = (1'h0);
  reg [(3'h6):(1'h0)] reg2923 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2922 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2921 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2920 = (1'h0);
  reg [(4'he):(1'h0)] reg2919 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2918 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2917 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2916 = (1'h0);
  reg [(4'h9):(1'h0)] reg2915 = (1'h0);
  reg [(4'hf):(1'h0)] reg2914 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2913 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2912 = (1'h0);
  reg [(4'hd):(1'h0)] reg2911 = (1'h0);
  reg [(4'hf):(1'h0)] reg2910 = (1'h0);
  reg [(3'h6):(1'h0)] reg2909 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2908 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2907 = (1'h0);
  reg [(4'h8):(1'h0)] reg2906 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2905 = (1'h0);
  reg [(4'hd):(1'h0)] reg2904 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2902 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2897 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2903 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2902 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2901 = (1'h0);
  reg [(3'h5):(1'h0)] reg2900 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2899 = (1'h0);
  reg [(4'hf):(1'h0)] reg2898 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2897 = (1'h0);
  reg [(3'h4):(1'h0)] reg2896 = (1'h0);
  reg [(4'ha):(1'h0)] reg2895 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2894 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2893 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2892 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2891 = (1'h0);
  reg [(4'hb):(1'h0)] reg2890 = (1'h0);
  reg [(4'hd):(1'h0)] reg2889 = (1'h0);
  reg [(4'hc):(1'h0)] reg2888 = (1'h0);
  reg [(3'h5):(1'h0)] reg2887 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2886 = (1'h0);
  reg [(3'h5):(1'h0)] reg2885 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2884 = (1'h0);
  reg [(3'h4):(1'h0)] reg2883 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2882 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2881 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2879 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2878 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2876 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2873 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2868 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2862 = (1'h0);
  reg [(4'hb):(1'h0)] reg2880 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2879 = (1'h0);
  reg [(4'hc):(1'h0)] reg2878 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2877 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2876 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2872 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2871 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2866 = (1'h0);
  reg [(4'hd):(1'h0)] reg2865 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2861 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2860 = (1'h0);
  reg [(3'h7):(1'h0)] reg2875 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2874 = (1'h0);
  reg [(5'h10):(1'h0)] reg2873 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2872 = (1'h0);
  reg [(3'h4):(1'h0)] reg2871 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2870 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2869 = (1'h0);
  reg [(4'h9):(1'h0)] reg2868 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2867 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2866 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2865 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2864 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2863 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2862 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2861 = (1'h0);
  reg [(4'he):(1'h0)] forvar2860 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2793 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2790 = (1'h0);
  reg [(3'h4):(1'h0)] reg2781 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2778 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2777 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2776 = (1'h0);
  reg [(4'hf):(1'h0)] reg2775 = (1'h0);
  reg [(2'h3):(1'h0)] reg2858 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2850 = (1'h0);
  reg [(3'h4):(1'h0)] reg2859 = (1'h0);
  reg [(4'he):(1'h0)] forvar2858 = (1'h0);
  reg [(3'h4):(1'h0)] reg2857 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2856 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2855 = (1'h0);
  reg [(4'hb):(1'h0)] reg2854 = (1'h0);
  reg [(2'h3):(1'h0)] reg2853 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2852 = (1'h0);
  reg [(2'h2):(1'h0)] reg2851 = (1'h0);
  reg [(3'h4):(1'h0)] reg2850 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2849 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2842 = (1'h0);
  reg [(4'h8):(1'h0)] reg2838 = (1'h0);
  reg [(4'hb):(1'h0)] reg2848 = (1'h0);
  reg [(4'h8):(1'h0)] reg2847 = (1'h0);
  reg [(4'h8):(1'h0)] reg2846 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2845 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2844 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2843 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2842 = (1'h0);
  reg [(2'h2):(1'h0)] reg2841 = (1'h0);
  reg [(4'hd):(1'h0)] reg2840 = (1'h0);
  reg [(3'h4):(1'h0)] reg2839 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2838 = (1'h0);
  reg [(4'hc):(1'h0)] reg2837 = (1'h0);
  reg [(3'h4):(1'h0)] reg2836 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2835 = (1'h0);
  reg [(3'h6):(1'h0)] reg2834 = (1'h0);
  reg [(2'h2):(1'h0)] reg2833 = (1'h0);
  reg [(4'h9):(1'h0)] reg2832 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2831 = (1'h0);
  reg [(2'h2):(1'h0)] reg2830 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2829 = (1'h0);
  reg [(4'hd):(1'h0)] reg2828 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2827 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2826 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2825 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2824 = (1'h0);
  reg [(3'h4):(1'h0)] reg2823 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2822 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2821 = (1'h0);
  reg [(4'hb):(1'h0)] reg2820 = (1'h0);
  reg [(4'ha):(1'h0)] reg2819 = (1'h0);
  reg [(4'h9):(1'h0)] reg2818 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2817 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2816 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2815 = (1'h0);
  reg [(4'hc):(1'h0)] reg2814 = (1'h0);
  reg [(3'h5):(1'h0)] reg2813 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2812 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2811 = (1'h0);
  reg [(4'hc):(1'h0)] reg2810 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2809 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2808 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2807 = (1'h0);
  reg [(4'hd):(1'h0)] reg2803 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2801 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2799 = (1'h0);
  reg [(4'h8):(1'h0)] reg2798 = (1'h0);
  reg [(4'he):(1'h0)] reg2806 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2805 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2804 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2803 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2802 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2801 = (1'h0);
  reg [(4'h8):(1'h0)] reg2800 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2799 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2798 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2797 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2796 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2795 = (1'h0);
  reg [(4'h9):(1'h0)] reg2794 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2793 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2792 = (1'h0);
  reg [(5'h10):(1'h0)] reg2791 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2790 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2783 = (1'h0);
  reg [(4'hd):(1'h0)] reg2789 = (1'h0);
  reg [(3'h7):(1'h0)] reg2788 = (1'h0);
  reg [(2'h3):(1'h0)] reg2787 = (1'h0);
  reg [(4'hf):(1'h0)] reg2786 = (1'h0);
  reg [(4'h8):(1'h0)] reg2785 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2784 = (1'h0);
  reg [(3'h4):(1'h0)] reg2783 = (1'h0);
  reg [(5'h10):(1'h0)] reg2782 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2781 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2780 = (1'h0);
  reg [(3'h5):(1'h0)] reg2779 = (1'h0);
  reg [(4'ha):(1'h0)] reg2778 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2777 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2776 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2775 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2774 = (1'h0);
  reg [(4'hb):(1'h0)] reg2773 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2772 = (1'h0);
  reg [(2'h3):(1'h0)] reg2771 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2770 = (1'h0);
  reg [(4'hb):(1'h0)] reg2769 = (1'h0);
  reg [(4'hb):(1'h0)] reg2768 = (1'h0);
  reg [(4'hb):(1'h0)] reg2767 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2766 = (1'h0);
  reg [(2'h2):(1'h0)] reg2765 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2764 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2755 = (1'h0);
  reg [(3'h7):(1'h0)] reg2763 = (1'h0);
  reg [(2'h3):(1'h0)] reg2762 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2761 = (1'h0);
  reg [(4'hf):(1'h0)] reg2760 = (1'h0);
  reg [(4'h9):(1'h0)] reg2759 = (1'h0);
  reg [(4'h9):(1'h0)] reg2758 = (1'h0);
  reg [(2'h2):(1'h0)] reg2757 = (1'h0);
  reg [(3'h4):(1'h0)] reg2756 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2755 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2754 = (1'h0);
  wire [(4'ha):(1'h0)] wire2753;
  wire [(4'hc):(1'h0)] wire2752;
  wire [(4'hb):(1'h0)] wire2751;
  wire signed [(3'h6):(1'h0)] wire2749;
  wire [(4'ha):(1'h0)] wire4017;
  assign y = {wire4164,
                 reg4163,
                 reg4156,
                 forvar4154,
                 reg4152,
                 reg4162,
                 reg4161,
                 reg4160,
                 reg4159,
                 reg4158,
                 reg4157,
                 forvar4156,
                 reg4155,
                 reg4154,
                 reg4153,
                 forvar4152,
                 reg4151,
                 reg4150,
                 forvar4149,
                 reg4148,
                 reg4147,
                 reg4146,
                 reg4145,
                 forvar4144,
                 reg4143,
                 reg4142,
                 reg4141,
                 reg4140,
                 reg4139,
                 reg4138,
                 reg4137,
                 reg4136,
                 reg4135,
                 forvar4134,
                 forvar4133,
                 reg4122,
                 reg4132,
                 reg4131,
                 reg4128,
                 reg4130,
                 reg4129,
                 forvar4128,
                 reg4127,
                 reg4126,
                 reg4125,
                 reg4124,
                 forvar4123,
                 forvar4122,
                 reg4121,
                 reg4120,
                 reg4119,
                 reg4118,
                 reg4117,
                 forvar4116,
                 reg4116,
                 reg4115,
                 reg4114,
                 forvar4113,
                 reg4112,
                 forvar4111,
                 forvar4110,
                 reg4098,
                 reg4093,
                 forvar4090,
                 reg4103,
                 reg4109,
                 reg4108,
                 forvar4107,
                 reg4106,
                 reg4105,
                 reg4104,
                 forvar4103,
                 reg4102,
                 reg4101,
                 reg4100,
                 reg4099,
                 forvar4098,
                 reg4097,
                 reg4096,
                 reg4095,
                 reg4094,
                 forvar4093,
                 reg4092,
                 reg4091,
                 reg4090,
                 reg4086,
                 forvar4084,
                 reg4082,
                 reg4078,
                 reg4089,
                 reg4088,
                 reg4087,
                 forvar4086,
                 reg4085,
                 reg4084,
                 reg4083,
                 forvar4082,
                 reg4081,
                 reg4080,
                 reg4079,
                 forvar4078,
                 reg4077,
                 reg4076,
                 reg4075,
                 forvar4074,
                 reg4073,
                 reg4072,
                 reg4071,
                 reg4070,
                 reg4069,
                 reg4068,
                 reg4067,
                 reg4066,
                 reg4065,
                 reg4064,
                 reg4063,
                 reg4062,
                 reg4061,
                 reg4060,
                 reg4059,
                 forvar4058,
                 reg4057,
                 reg4056,
                 reg4055,
                 reg4054,
                 forvar4053,
                 forvar4052,
                 reg4051,
                 reg4050,
                 reg4049,
                 reg4048,
                 reg4047,
                 reg4046,
                 forvar4045,
                 forvar4044,
                 reg4043,
                 reg4042,
                 forvar4041,
                 reg4040,
                 forvar4027,
                 reg4039,
                 reg4038,
                 forvar4037,
                 reg4036,
                 reg4035,
                 reg4034,
                 reg4033,
                 forvar4032,
                 reg4031,
                 reg4030,
                 reg4029,
                 reg4028,
                 reg4026,
                 reg4027,
                 forvar4026,
                 reg4025,
                 reg4024,
                 reg4023,
                 reg4022,
                 forvar4021,
                 forvar4020,
                 wire4019,
                 wire3601,
                 reg3493,
                 forvar3491,
                 reg3489,
                 forvar3486,
                 forvar3483,
                 forvar3477,
                 forvar3476,
                 reg3501,
                 forvar3500,
                 reg3499,
                 reg3498,
                 reg3497,
                 reg3496,
                 reg3495,
                 reg3494,
                 forvar3493,
                 forvar3492,
                 reg3491,
                 reg3490,
                 forvar3489,
                 reg3488,
                 reg3487,
                 reg3486,
                 reg3485,
                 reg3484,
                 reg3483,
                 forvar3482,
                 reg3473,
                 reg3481,
                 reg3480,
                 reg3479,
                 reg3478,
                 reg3477,
                 reg3476,
                 reg3475,
                 reg3474,
                 forvar3473,
                 reg3472,
                 reg3471,
                 reg3470,
                 reg3469,
                 forvar3466,
                 forvar3464,
                 reg3461,
                 reg3468,
                 reg3467,
                 reg3466,
                 reg3465,
                 reg3464,
                 reg3463,
                 reg3462,
                 forvar3461,
                 forvar3460,
                 reg3459,
                 reg3458,
                 forvar3457,
                 reg3456,
                 reg3455,
                 reg3454,
                 forvar3453,
                 reg3452,
                 forvar3451,
                 forvar3450,
                 reg3449,
                 reg3448,
                 reg3447,
                 reg3446,
                 reg3445,
                 reg3444,
                 reg3443,
                 reg3442,
                 forvar3441,
                 reg3428,
                 reg3440,
                 reg3439,
                 reg3438,
                 forvar3437,
                 reg3436,
                 reg3435,
                 reg3434,
                 reg3433,
                 reg3432,
                 reg3431,
                 reg3430,
                 reg3429,
                 forvar3428,
                 forvar3427,
                 forvar3426,
                 reg3425,
                 forvar3424,
                 reg3423,
                 forvar3422,
                 reg3421,
                 reg3420,
                 reg3419,
                 reg3418,
                 reg3417,
                 forvar3416,
                 reg3415,
                 reg3414,
                 forvar3413,
                 forvar3408,
                 reg3412,
                 reg3411,
                 reg3410,
                 reg3409,
                 reg3408,
                 reg3407,
                 reg3404,
                 forvar3402,
                 reg3401,
                 forvar3395,
                 reg3406,
                 reg3405,
                 forvar3404,
                 reg3403,
                 reg3402,
                 forvar3401,
                 reg3400,
                 reg3399,
                 reg3398,
                 forvar3397,
                 reg3396,
                 reg3395,
                 forvar3394,
                 reg3393,
                 forvar3382,
                 reg3392,
                 reg3391,
                 forvar3390,
                 reg3389,
                 reg3388,
                 reg3387,
                 reg3386,
                 reg3385,
                 reg3384,
                 reg3383,
                 reg3382,
                 forvar3381,
                 forvar3367,
                 reg3365,
                 reg3363,
                 reg3362,
                 forvar3361,
                 reg3380,
                 forvar3379,
                 reg3378,
                 reg3377,
                 reg3376,
                 reg3375,
                 reg3374,
                 forvar3372,
                 reg3373,
                 reg3372,
                 reg3371,
                 reg3370,
                 reg3369,
                 reg3368,
                 reg3367,
                 reg3366,
                 forvar3365,
                 reg3364,
                 forvar3363,
                 forvar3362,
                 reg3361,
                 reg3360,
                 forvar3359,
                 reg3358,
                 reg3357,
                 forvar3356,
                 reg3355,
                 reg3354,
                 reg3353,
                 reg3352,
                 reg3351,
                 forvar3350,
                 reg3349,
                 forvar3348,
                 reg3347,
                 forvar3346,
                 reg3345,
                 forvar3344,
                 forvar3343,
                 reg3342,
                 reg3341,
                 reg3340,
                 reg3339,
                 reg3338,
                 reg3337,
                 reg3336,
                 reg3335,
                 reg3334,
                 reg3333,
                 forvar3332,
                 reg3331,
                 reg3330,
                 reg3329,
                 reg3328,
                 forvar3327,
                 reg3326,
                 forvar3325,
                 forvar3324,
                 reg3323,
                 reg3322,
                 forvar3321,
                 reg3320,
                 reg3319,
                 reg3318,
                 reg3317,
                 reg3316,
                 reg3315,
                 reg3314,
                 reg3313,
                 forvar3312,
                 forvar3311,
                 reg3310,
                 reg3309,
                 forvar3308,
                 reg3307,
                 reg3306,
                 reg3305,
                 reg3304,
                 forvar3303,
                 reg3302,
                 reg3301,
                 reg3300,
                 reg3299,
                 reg3298,
                 forvar3297,
                 forvar3296,
                 reg3295,
                 reg3294,
                 forvar3293,
                 forvar3292,
                 reg3291,
                 reg3290,
                 reg3289,
                 forvar3288,
                 reg3287,
                 forvar3285,
                 reg3284,
                 forvar3283,
                 reg3280,
                 reg3274,
                 reg3286,
                 reg3285,
                 forvar3284,
                 reg3283,
                 reg3282,
                 reg3281,
                 forvar3280,
                 reg3279,
                 reg3278,
                 reg3277,
                 reg3276,
                 forvar3275,
                 forvar3274,
                 reg3273,
                 reg3272,
                 forvar3271,
                 reg3270,
                 reg3269,
                 reg3268,
                 reg3267,
                 forvar3266,
                 forvar3265,
                 reg3264,
                 reg3263,
                 reg3262,
                 reg3261,
                 forvar3260,
                 reg3259,
                 reg3258,
                 reg3257,
                 reg3256,
                 forvar3255,
                 forvar3254,
                 forvar3253,
                 reg3237,
                 reg3232,
                 forvar3231,
                 reg3228,
                 reg3224,
                 reg3252,
                 reg3251,
                 reg3250,
                 reg3249,
                 reg3248,
                 forvar3247,
                 reg3246,
                 reg3245,
                 reg3244,
                 reg3243,
                 forvar3242,
                 reg3241,
                 forvar3240,
                 reg3239,
                 reg3238,
                 forvar3237,
                 reg3236,
                 reg3235,
                 reg3234,
                 reg3233,
                 forvar3232,
                 reg3231,
                 reg3230,
                 reg3229,
                 forvar3228,
                 reg3227,
                 reg3226,
                 reg3225,
                 forvar3224,
                 forvar3223,
                 forvar3205,
                 reg3200,
                 reg3222,
                 reg3221,
                 forvar3220,
                 reg3219,
                 reg3217,
                 reg3215,
                 reg3218,
                 forvar3217,
                 reg3216,
                 forvar3215,
                 reg3214,
                 forvar3213,
                 reg3212,
                 reg3211,
                 forvar3210,
                 reg3209,
                 reg3208,
                 reg3203,
                 reg3207,
                 reg3206,
                 reg3205,
                 reg3204,
                 forvar3203,
                 reg3202,
                 reg3201,
                 forvar3200,
                 reg3199,
                 reg3198,
                 reg3197,
                 reg3196,
                 reg3195,
                 forvar3194,
                 reg3193,
                 reg3192,
                 reg3191,
                 reg3190,
                 reg3189,
                 reg3188,
                 forvar3187,
                 forvar3186,
                 reg3185,
                 forvar3184,
                 forvar3183,
                 wire3182,
                 reg3181,
                 reg3177,
                 reg3180,
                 reg3179,
                 reg3178,
                 forvar3177,
                 reg3176,
                 reg3175,
                 reg3174,
                 reg3173,
                 reg3172,
                 reg3171,
                 reg3170,
                 reg3169,
                 forvar3168,
                 reg3167,
                 reg3166,
                 forvar3165,
                 forvar3164,
                 forvar3163,
                 reg3120,
                 forvar3112,
                 forvar3110,
                 forvar3109,
                 forvar3108,
                 reg3103,
                 reg3101,
                 forvar3095,
                 reg3091,
                 reg3162,
                 reg3161,
                 reg3160,
                 reg3159,
                 reg3158,
                 forvar3157,
                 reg3156,
                 reg3155,
                 reg3154,
                 reg3153,
                 forvar3152,
                 forvar3151,
                 reg3150,
                 reg3149,
                 reg3148,
                 reg3147,
                 reg3143,
                 forvar3142,
                 reg3141,
                 forvar3139,
                 reg3146,
                 reg3145,
                 reg3144,
                 forvar3143,
                 reg3142,
                 forvar3141,
                 reg3140,
                 reg3139,
                 reg3138,
                 reg3130,
                 reg3137,
                 reg3136,
                 forvar3135,
                 reg3134,
                 reg3133,
                 reg3132,
                 reg3131,
                 forvar3130,
                 reg3129,
                 reg3128,
                 reg3127,
                 reg3126,
                 forvar3125,
                 reg3124,
                 reg3123,
                 forvar3122,
                 reg3121,
                 forvar3120,
                 reg3119,
                 reg3118,
                 reg3117,
                 reg3116,
                 reg3115,
                 forvar3114,
                 reg3113,
                 reg3112,
                 reg3111,
                 reg3110,
                 reg3109,
                 reg3108,
                 reg3107,
                 reg3106,
                 reg3105,
                 reg3104,
                 forvar3103,
                 forvar3102,
                 forvar3101,
                 reg3100,
                 reg3099,
                 reg3098,
                 reg3097,
                 reg3096,
                 reg3095,
                 reg3094,
                 reg3093,
                 reg3092,
                 forvar3091,
                 forvar3090,
                 reg3089,
                 reg3088,
                 forvar3087,
                 reg3086,
                 forvar3084,
                 reg3081,
                 reg3085,
                 reg3084,
                 reg3083,
                 reg3082,
                 forvar3081,
                 reg3080,
                 reg3079,
                 reg3078,
                 reg3077,
                 reg3076,
                 forvar3075,
                 reg3074,
                 reg3073,
                 reg3072,
                 reg3071,
                 forvar3070,
                 reg3069,
                 reg3068,
                 reg3067,
                 forvar3066,
                 reg3065,
                 reg3064,
                 reg3063,
                 reg3062,
                 forvar3061,
                 forvar3060,
                 reg3052,
                 reg3047,
                 reg3059,
                 reg3058,
                 reg3057,
                 forvar3056,
                 reg3055,
                 reg3054,
                 reg3053,
                 forvar3052,
                 reg3051,
                 reg3050,
                 reg3049,
                 reg3048,
                 forvar3047,
                 reg3046,
                 forvar3045,
                 reg3044,
                 forvar3043,
                 forvar3033,
                 forvar3027,
                 forvar3011,
                 forvar3006,
                 reg3029,
                 reg3042,
                 forvar3041,
                 reg3040,
                 reg3039,
                 reg3038,
                 reg3037,
                 reg3036,
                 reg3035,
                 reg3034,
                 reg3033,
                 reg3032,
                 reg3031,
                 reg3030,
                 forvar3029,
                 forvar3028,
                 forvar3022,
                 reg3021,
                 forvar3017,
                 forvar3010,
                 reg3016,
                 reg3012,
                 reg3009,
                 forvar3007,
                 forvar3004,
                 reg3027,
                 reg3026,
                 reg3025,
                 reg3024,
                 reg3023,
                 reg3022,
                 forvar3021,
                 reg3020,
                 reg3019,
                 reg3018,
                 reg3017,
                 forvar3016,
                 reg3015,
                 reg3014,
                 reg3013,
                 forvar3012,
                 reg3011,
                 reg3010,
                 forvar3009,
                 reg3008,
                 reg3007,
                 forvar3005,
                 reg3006,
                 reg3005,
                 reg3004,
                 wire3003,
                 wire3002,
                 forvar2966,
                 forvar2964,
                 reg2963,
                 forvar2959,
                 forvar2958,
                 forvar2950,
                 forvar2945,
                 reg2944,
                 forvar2978,
                 forvar2974,
                 forvar2970,
                 reg2969,
                 reg2968,
                 reg3001,
                 reg3000,
                 reg2999,
                 reg2998,
                 reg2997,
                 reg2996,
                 reg2995,
                 reg2994,
                 forvar2993,
                 reg2992,
                 reg2991,
                 forvar2990,
                 reg2989,
                 reg2988,
                 reg2987,
                 reg2986,
                 reg2983,
                 reg2985,
                 reg2984,
                 forvar2983,
                 reg2982,
                 reg2981,
                 reg2980,
                 reg2979,
                 reg2978,
                 reg2977,
                 reg2976,
                 reg2975,
                 reg2974,
                 reg2973,
                 reg2972,
                 reg2971,
                 reg2970,
                 forvar2969,
                 forvar2968,
                 reg2967,
                 reg2966,
                 reg2965,
                 reg2964,
                 forvar2963,
                 reg2962,
                 reg2961,
                 reg2960,
                 reg2959,
                 reg2958,
                 reg2957,
                 reg2956,
                 forvar2955,
                 reg2953,
                 reg2948,
                 reg2947,
                 reg2943,
                 reg2955,
                 reg2954,
                 forvar2953,
                 reg2952,
                 reg2951,
                 reg2950,
                 reg2949,
                 forvar2948,
                 forvar2947,
                 reg2946,
                 reg2945,
                 forvar2944,
                 forvar2943,
                 reg2942,
                 reg2941,
                 reg2940,
                 reg2939,
                 reg2938,
                 reg2937,
                 forvar2931,
                 reg2936,
                 reg2935,
                 reg2934,
                 reg2933,
                 reg2932,
                 reg2931,
                 reg2930,
                 forvar2919,
                 reg2927,
                 reg2925,
                 forvar2922,
                 reg2920,
                 reg2929,
                 reg2928,
                 forvar2927,
                 reg2926,
                 forvar2925,
                 reg2917,
                 reg2924,
                 reg2923,
                 reg2922,
                 reg2921,
                 forvar2920,
                 reg2919,
                 reg2918,
                 forvar2917,
                 reg2916,
                 reg2915,
                 reg2914,
                 reg2913,
                 forvar2912,
                 reg2911,
                 reg2910,
                 reg2909,
                 forvar2908,
                 reg2907,
                 reg2906,
                 reg2905,
                 reg2904,
                 forvar2902,
                 reg2897,
                 reg2903,
                 reg2902,
                 reg2901,
                 reg2900,
                 forvar2899,
                 reg2898,
                 forvar2897,
                 reg2896,
                 reg2895,
                 reg2894,
                 reg2893,
                 forvar2892,
                 forvar2891,
                 reg2890,
                 reg2889,
                 reg2888,
                 reg2887,
                 forvar2886,
                 reg2885,
                 reg2884,
                 reg2883,
                 reg2882,
                 reg2881,
                 reg2879,
                 forvar2878,
                 reg2876,
                 forvar2873,
                 forvar2868,
                 forvar2862,
                 reg2880,
                 forvar2879,
                 reg2878,
                 reg2877,
                 forvar2876,
                 reg2872,
                 forvar2871,
                 forvar2866,
                 reg2865,
                 forvar2861,
                 reg2860,
                 reg2875,
                 reg2874,
                 reg2873,
                 forvar2872,
                 reg2871,
                 reg2870,
                 reg2869,
                 reg2868,
                 reg2867,
                 reg2866,
                 forvar2865,
                 reg2864,
                 reg2863,
                 reg2862,
                 reg2861,
                 forvar2860,
                 reg2793,
                 reg2790,
                 reg2781,
                 forvar2778,
                 forvar2777,
                 reg2776,
                 reg2775,
                 reg2858,
                 forvar2850,
                 reg2859,
                 forvar2858,
                 reg2857,
                 reg2856,
                 forvar2855,
                 reg2854,
                 reg2853,
                 reg2852,
                 reg2851,
                 reg2850,
                 forvar2849,
                 reg2842,
                 reg2838,
                 reg2848,
                 reg2847,
                 reg2846,
                 reg2845,
                 forvar2844,
                 reg2843,
                 forvar2842,
                 reg2841,
                 reg2840,
                 reg2839,
                 forvar2838,
                 reg2837,
                 reg2836,
                 reg2835,
                 reg2834,
                 reg2833,
                 reg2832,
                 reg2831,
                 reg2830,
                 forvar2829,
                 reg2828,
                 reg2827,
                 forvar2826,
                 reg2825,
                 reg2824,
                 reg2823,
                 forvar2822,
                 forvar2821,
                 reg2820,
                 reg2819,
                 reg2818,
                 reg2817,
                 reg2816,
                 reg2815,
                 reg2814,
                 reg2813,
                 reg2812,
                 reg2811,
                 reg2810,
                 forvar2809,
                 forvar2808,
                 reg2807,
                 reg2803,
                 forvar2801,
                 forvar2799,
                 reg2798,
                 reg2806,
                 reg2805,
                 reg2804,
                 forvar2803,
                 reg2802,
                 reg2801,
                 reg2800,
                 reg2799,
                 forvar2798,
                 forvar2797,
                 reg2796,
                 reg2795,
                 reg2794,
                 forvar2793,
                 reg2792,
                 reg2791,
                 forvar2790,
                 forvar2783,
                 reg2789,
                 reg2788,
                 reg2787,
                 reg2786,
                 reg2785,
                 reg2784,
                 reg2783,
                 reg2782,
                 forvar2781,
                 reg2780,
                 reg2779,
                 reg2778,
                 reg2777,
                 forvar2776,
                 forvar2775,
                 forvar2774,
                 reg2773,
                 reg2772,
                 reg2771,
                 forvar2770,
                 reg2769,
                 reg2768,
                 reg2767,
                 reg2766,
                 reg2765,
                 forvar2764,
                 reg2755,
                 reg2763,
                 reg2762,
                 reg2761,
                 reg2760,
                 reg2759,
                 reg2758,
                 reg2757,
                 reg2756,
                 forvar2755,
                 forvar2754,
                 wire2753,
                 wire2752,
                 wire2751,
                 wire2749,
                 wire4017,
                 (1'h0)};
  module1764 modinst2750 (wire2749, clk, wire1763, wire1762, wire1760, wire1761);
  assign wire2751 = ((wire1762 ?
                            (^wire1762) : ($signed(wire1762) || $unsigned((8'h9c)))) ?
                        (~&(~{wire1763})) : $unsigned($unsigned($unsigned(wire1760))));
  assign wire2752 = wire1760;
  assign wire2753 = {($signed((8'ha3)) ?
                            (wire1762 - {wire1760}) : ((&wire1760) ~^ ((8'hb1) ?
                                (8'h9e) : (8'ha8))))};
  always
    @(posedge clk) begin
      for (forvar2754 = (1'h0); (forvar2754 < (1'h1)); forvar2754 = (forvar2754 + (1'h1)))
        begin
          if (wire1762[(3'h7):(3'h4)])
            begin
              if ((($unsigned($signed(forvar2754)) ^ ({wire2749} ?
                      $signed(wire2751) : $signed((8'ha1)))) ?
                  ((|(wire1763 > wire1760)) ^~ (-((8'hb0) != wire2749))) : (($unsigned(wire1760) != ((8'hb3) ?
                      wire2749 : wire2751)) | wire2749[(3'h4):(2'h3)])))
                begin
                  for (forvar2755 = (1'h0); (forvar2755 < (2'h3)); forvar2755 = (forvar2755 + (1'h1)))
                    begin
                      reg2756 <= {wire2751};
                      reg2757 <= (~({$unsigned(wire1763)} >= {$signed(wire1761)}));
                      reg2758 <= wire1760[(3'h7):(2'h3)];
                    end
                  if ((8'ha2))
                    begin
                      reg2759 <= forvar2754;
                      reg2760 <= (&((~|((8'h9e) ? wire1760 : reg2757)) ?
                          wire1762 : reg2756[(3'h4):(3'h4)]));
                    end
                  else
                    begin
                      reg2759 <= (wire2749 ? $signed(wire1762) : (8'hae));
                      reg2760 <= (~^((wire2752[(2'h2):(2'h2)] ?
                          {forvar2754} : $signed(reg2756)) <= ({reg2757} == (!wire2749))));
                      reg2761 <= (^$unsigned(reg2759[(1'h0):(1'h0)]));
                      reg2762 <= {$signed(wire1760[(4'h8):(2'h3)])};
                    end
                  reg2763 <= $signed((($signed(reg2761) << (forvar2755 < wire2749)) ?
                      (~&(^~wire2751)) : forvar2754[(1'h1):(1'h1)]));
                end
              else
                begin
                  reg2755 <= (wire2752 - $signed((~|$unsigned((8'had)))));
                end
              for (forvar2764 = (1'h0); (forvar2764 < (1'h1)); forvar2764 = (forvar2764 + (1'h1)))
                begin
                  if ({($signed(((8'haa) && (8'hb3))) ?
                          reg2756[(1'h1):(1'h0)] : (!$unsigned(wire1763)))})
                    begin
                      reg2765 <= $unsigned(((reg2762[(1'h1):(1'h1)] >> reg2755[(3'h4):(1'h1)]) ?
                          forvar2755 : $signed(reg2760[(4'hf):(3'h7)])));
                      reg2766 <= $unsigned($unsigned(($unsigned(wire2751) & (wire2751 || forvar2764))));
                      reg2767 <= (reg2758 & (8'ha6));
                    end
                  else
                    begin
                      reg2765 <= ((($unsigned((8'had)) ?
                                  {reg2757} : wire2753[(4'ha):(4'h8)]) ?
                              {((8'ha9) ?
                                      reg2759 : (8'hba))} : wire2753[(4'h9):(3'h5)]) ?
                          ($signed((~&reg2767)) ?
                              ($signed((8'hba)) ?
                                  (&reg2760) : (wire2753 == (8'ha8))) : $unsigned($unsigned(wire1760))) : (((|reg2765) >> forvar2754) ?
                              wire2749 : reg2765));
                      reg2766 <= {(((reg2760 ?
                              reg2762 : forvar2764) ^~ wire2752) > ($unsigned(wire2753) ^~ (~^reg2758)))};
                    end
                  reg2768 <= (~reg2755[(3'h4):(1'h1)]);
                end
              reg2769 <= wire1763;
              if ((^~wire1760[(3'h7):(3'h5)]))
                begin
                  for (forvar2770 = (1'h0); (forvar2770 < (2'h3)); forvar2770 = (forvar2770 + (1'h1)))
                    begin
                      reg2771 <= {$signed((~|wire2753[(2'h3):(2'h3)]))};
                      reg2772 <= reg2771[(2'h2):(1'h1)];
                      reg2773 <= wire2751;
                    end
                end
              else
                begin
                  for (forvar2770 = (1'h0); (forvar2770 < (2'h2)); forvar2770 = (forvar2770 + (1'h1)))
                    begin
                      reg2771 <= $unsigned((reg2759 && reg2755));
                      reg2772 <= reg2762[(2'h2):(2'h2)];
                      reg2773 <= reg2758;
                    end
                end
            end
          else
            begin
              for (forvar2755 = (1'h0); (forvar2755 < (1'h1)); forvar2755 = (forvar2755 + (1'h1)))
                begin
                  if (($signed(wire1762) >> reg2765))
                    begin
                      reg2756 <= ($unsigned($unsigned($unsigned(reg2758))) & wire2751[(3'h7):(3'h6)]);
                      reg2757 <= reg2769[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg2756 <= (8'hb3);
                      reg2757 <= wire1761[(4'he):(2'h3)];
                      reg2758 <= $unsigned($signed((wire2752 ?
                          $signed((8'h9c)) : $signed(reg2762))));
                    end
                end
              reg2759 <= ($signed((((8'ha6) >>> (8'ha6)) ?
                      (reg2757 * wire2753) : (^~wire2749))) ?
                  $signed($signed(reg2771[(1'h1):(1'h0)])) : (8'had));
            end
        end
      if ($unsigned((~$unsigned($unsigned(wire2753)))))
        begin
          for (forvar2774 = (1'h0); (forvar2774 < (1'h0)); forvar2774 = (forvar2774 + (1'h1)))
            begin
              for (forvar2775 = (1'h0); (forvar2775 < (1'h0)); forvar2775 = (forvar2775 + (1'h1)))
                begin
                  for (forvar2776 = (1'h0); (forvar2776 < (2'h3)); forvar2776 = (forvar2776 + (1'h1)))
                    begin
                      reg2777 <= (($signed((forvar2754 * wire1762)) >= (8'h9c)) ^ ($unsigned((|forvar2764)) > $unsigned(forvar2776[(3'h7):(3'h4)])));
                      reg2778 <= ($signed($unsigned((-forvar2774))) ?
                          $signed(forvar2754[(1'h0):(1'h0)]) : $signed(wire2753[(1'h0):(1'h0)]));
                    end
                  if (wire2751[(1'h0):(1'h0)])
                    begin
                      reg2779 <= (reg2769 ^~ (reg2756 << (reg2758[(3'h4):(2'h2)] != $unsigned(forvar2775))));
                    end
                  else
                    begin
                      reg2779 <= forvar2775;
                      reg2780 <= $unsigned(reg2773[(3'h4):(1'h1)]);
                    end
                  for (forvar2781 = (1'h0); (forvar2781 < (2'h3)); forvar2781 = (forvar2781 + (1'h1)))
                    begin
                      reg2782 <= (((~&(wire2751 ? reg2767 : wire1761)) ?
                              ((forvar2764 ? (8'hb5) : reg2766) ?
                                  (wire1763 && reg2765) : reg2778) : reg2769[(1'h0):(1'h0)]) ?
                          $unsigned((forvar2781[(4'hb):(2'h2)] || (reg2766 > wire1760))) : ((reg2769 ?
                              (forvar2764 <= reg2759) : (reg2768 && forvar2764)) != ({reg2771} | $unsigned(reg2768))));
                    end
                end
              if (forvar2781[(3'h4):(1'h0)])
                begin
                  if ((8'ha1))
                    begin
                      reg2783 <= $unsigned(wire1760[(4'he):(1'h1)]);
                      reg2784 <= $unsigned(((~&reg2771[(1'h1):(1'h0)]) || $unsigned({wire2751})));
                      reg2785 <= ($signed($unsigned($signed(reg2773))) ?
                          $unsigned(((reg2765 || forvar2774) | $unsigned((8'ha4)))) : reg2779[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg2783 <= {$unsigned($signed((~^reg2773)))};
                      reg2784 <= $unsigned($unsigned((^~(reg2761 ?
                          reg2763 : reg2755))));
                      reg2785 <= $signed((|$unsigned($signed((8'h9f)))));
                    end
                  if ((-wire2752[(4'hc):(4'hb)]))
                    begin
                      reg2786 <= $unsigned($signed(($unsigned(reg2777) ~^ $signed(reg2763))));
                      reg2787 <= reg2766[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg2786 <= ($unsigned($signed($unsigned(reg2757))) ?
                          ($unsigned($signed(wire2753)) >= (~^$unsigned(reg2757))) : (((reg2780 * reg2766) >>> $unsigned((8'hac))) <<< reg2785[(2'h2):(1'h0)]));
                      reg2787 <= reg2784;
                    end
                  reg2788 <= $unsigned((8'ha8));
                  reg2789 <= {$signed(forvar2755)};
                end
              else
                begin
                  for (forvar2783 = (1'h0); (forvar2783 < (1'h0)); forvar2783 = (forvar2783 + (1'h1)))
                    begin
                      reg2784 <= reg2755[(2'h2):(2'h2)];
                      reg2785 <= (&($unsigned((reg2763 ?
                          forvar2770 : forvar2776)) - (~^reg2758[(3'h7):(3'h4)])));
                      reg2786 <= (reg2785 && reg2765);
                      reg2787 <= (~|reg2763[(3'h7):(1'h0)]);
                    end
                end
              for (forvar2790 = (1'h0); (forvar2790 < (1'h1)); forvar2790 = (forvar2790 + (1'h1)))
                begin
                  if ($signed(reg2767))
                    begin
                      reg2791 <= reg2769;
                      reg2792 <= (forvar2770 ?
                          ($unsigned((reg2763 ?
                              reg2786 : wire1762)) & $signed((wire1763 << reg2761))) : $unsigned($signed(reg2783)));
                    end
                  else
                    begin
                      reg2791 <= reg2768[(4'ha):(3'h7)];
                      reg2792 <= (^{$signed($unsigned((8'hb6)))});
                    end
                end
            end
          for (forvar2793 = (1'h0); (forvar2793 < (1'h1)); forvar2793 = (forvar2793 + (1'h1)))
            begin
              reg2794 <= ((($signed((8'hba)) << (reg2762 | reg2783)) || $unsigned((reg2768 ?
                      reg2755 : forvar2755))) ?
                  forvar2790[(3'h4):(3'h4)] : (((reg2783 ~^ forvar2790) ?
                      $signed(reg2756) : (reg2789 ?
                          forvar2776 : forvar2793)) ~^ ($unsigned(wire2753) < $signed(reg2760))));
              reg2795 <= reg2762;
              reg2796 <= $signed($unsigned(reg2765[(1'h1):(1'h1)]));
            end
          for (forvar2797 = (1'h0); (forvar2797 < (2'h2)); forvar2797 = (forvar2797 + (1'h1)))
            begin
              if (reg2769[(1'h1):(1'h0)])
                begin
                  for (forvar2798 = (1'h0); (forvar2798 < (2'h2)); forvar2798 = (forvar2798 + (1'h1)))
                    begin
                      reg2799 <= ($unsigned($unsigned(((8'h9c) ~^ forvar2798))) ?
                          forvar2770[(2'h3):(2'h2)] : $signed((~&reg2792[(1'h1):(1'h0)])));
                      reg2800 <= $signed($signed((~(&(8'ha4)))));
                      reg2801 <= $signed((($unsigned(reg2783) - (~|reg2757)) ?
                          $signed((forvar2770 >> reg2765)) : {{forvar2790}}));
                      reg2802 <= ((((8'h9c) ?
                                  $signed((8'h9d)) : (reg2777 ?
                                      (8'hae) : wire1760)) ?
                              $signed((~reg2778)) : $unsigned($signed(wire1763))) ?
                          $unsigned(($unsigned(reg2788) << $unsigned(forvar2783))) : ($signed($signed(reg2796)) ?
                              forvar2798 : (^~$unsigned(forvar2774))));
                    end
                  for (forvar2803 = (1'h0); (forvar2803 < (1'h0)); forvar2803 = (forvar2803 + (1'h1)))
                    begin
                      reg2804 <= $unsigned($signed({(&reg2758)}));
                      reg2805 <= reg2758[(3'h7):(3'h5)];
                      reg2806 <= ((+$unsigned($signed(reg2794))) || reg2792[(3'h7):(3'h7)]);
                    end
                end
              else
                begin
                  reg2798 <= $unsigned(({reg2768} ?
                      (~&{wire1761}) : (~&(wire1763 ? reg2806 : (8'h9e)))));
                  for (forvar2799 = (1'h0); (forvar2799 < (1'h0)); forvar2799 = (forvar2799 + (1'h1)))
                    begin
                      reg2800 <= reg2772;
                    end
                  for (forvar2801 = (1'h0); (forvar2801 < (2'h3)); forvar2801 = (forvar2801 + (1'h1)))
                    begin
                      reg2802 <= reg2761;
                      reg2803 <= reg2806;
                    end
                  if ($signed($signed($signed($unsigned(forvar2797)))))
                    begin
                      reg2804 <= $signed((($signed(reg2761) ?
                              $unsigned(reg2804) : (|reg2763)) ?
                          $signed($unsigned(reg2791)) : {$signed(reg2804)}));
                      reg2805 <= wire2749[(3'h4):(2'h2)];
                      reg2806 <= {wire2753};
                      reg2807 <= $signed(($unsigned(reg2758) ?
                          reg2765[(2'h2):(2'h2)] : $signed($signed(reg2762))));
                    end
                  else
                    begin
                      reg2804 <= (^~(^~((reg2806 ? reg2757 : reg2800) ?
                          {(8'ha5)} : (8'haa))));
                      reg2805 <= (($unsigned((forvar2801 ?
                          (8'hac) : forvar2801)) | $signed(reg2802[(4'hc):(4'hb)])) || (reg2773[(1'h0):(1'h0)] < ((~&wire2753) > (reg2756 ?
                          reg2785 : reg2763))));
                      reg2806 <= reg2778[(1'h0):(1'h0)];
                    end
                end
              for (forvar2808 = (1'h0); (forvar2808 < (2'h3)); forvar2808 = (forvar2808 + (1'h1)))
                begin
                  for (forvar2809 = (1'h0); (forvar2809 < (2'h2)); forvar2809 = (forvar2809 + (1'h1)))
                    begin
                      reg2810 <= ((forvar2793 ?
                          $unsigned((|forvar2790)) : $signed({wire2751})) <<< (($unsigned(forvar2755) ?
                              $unsigned(reg2765) : (reg2772 ^~ reg2763)) ?
                          $unsigned($unsigned(reg2765)) : (~&(|reg2805))));
                      reg2811 <= (~^$signed($signed((reg2799 ^~ forvar2783))));
                      reg2812 <= (((!wire1760[(3'h6):(3'h6)]) <= reg2806[(2'h2):(2'h2)]) ?
                          (((forvar2798 ? reg2759 : reg2798) ?
                                  wire2753 : $signed(reg2811)) ?
                              ($signed(forvar2790) ?
                                  reg2757[(1'h0):(1'h0)] : reg2783) : ($unsigned(forvar2774) >>> reg2777[(2'h3):(1'h0)])) : wire2749);
                      reg2813 <= {reg2799};
                    end
                  if ((~|reg2786))
                    begin
                      reg2814 <= $unsigned((!{forvar2783}));
                      reg2815 <= $unsigned(((&(+forvar2776)) == forvar2790));
                    end
                  else
                    begin
                      reg2814 <= ((~|((~|reg2762) ?
                              (~&reg2791) : $unsigned(reg2801))) ?
                          ($signed($unsigned(reg2814)) ?
                              ((reg2811 ?
                                  reg2771 : forvar2783) >> (forvar2775 <<< (8'hb5))) : (forvar2776 + $signed(forvar2793))) : (~|$unsigned(forvar2793)));
                    end
                  if ((~|$unsigned(reg2794[(3'h7):(3'h7)])))
                    begin
                      reg2816 <= $unsigned(reg2799);
                      reg2817 <= (^reg2780[(2'h3):(1'h1)]);
                      reg2818 <= ((~(((8'hab) ?
                          reg2759 : reg2756) + $signed(reg2811))) << (~(forvar2764[(3'h7):(2'h2)] ?
                          $unsigned(reg2758) : (~|reg2779))));
                    end
                  else
                    begin
                      reg2816 <= reg2760[(4'hb):(4'h8)];
                      reg2817 <= reg2799;
                    end
                  if ($unsigned(((!(^~reg2772)) ?
                      reg2807 : reg2796[(2'h3):(1'h0)])))
                    begin
                      reg2819 <= reg2784;
                      reg2820 <= reg2762[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2819 <= $unsigned((((forvar2809 ?
                              reg2778 : wire2749) > (^forvar2801)) ?
                          reg2784 : $unsigned($unsigned(reg2802))));
                    end
                end
              for (forvar2821 = (1'h0); (forvar2821 < (2'h2)); forvar2821 = (forvar2821 + (1'h1)))
                begin
                  for (forvar2822 = (1'h0); (forvar2822 < (2'h3)); forvar2822 = (forvar2822 + (1'h1)))
                    begin
                      reg2823 <= (forvar2790[(2'h3):(1'h0)] ?
                          reg2818 : reg2791[(2'h2):(1'h0)]);
                      reg2824 <= $signed((+reg2787));
                      reg2825 <= ((8'ha0) >= (^((~wire2753) ?
                          $unsigned((8'hb2)) : (reg2789 && reg2779))));
                    end
                  for (forvar2826 = (1'h0); (forvar2826 < (1'h0)); forvar2826 = (forvar2826 + (1'h1)))
                    begin
                      reg2827 <= (((~|(forvar2793 == forvar2801)) ?
                          (wire2751[(1'h0):(1'h0)] ?
                              (~reg2825) : (~&(8'hae))) : $unsigned((reg2816 ?
                              forvar2781 : reg2805))) != forvar2776[(3'h7):(1'h1)]);
                      reg2828 <= forvar2821;
                    end
                  for (forvar2829 = (1'h0); (forvar2829 < (2'h2)); forvar2829 = (forvar2829 + (1'h1)))
                    begin
                      reg2830 <= ((8'hb2) ?
                          {$unsigned((reg2816 ?
                                  forvar2797 : reg2792))} : {(~$unsigned(reg2773))});
                      reg2831 <= ($signed(reg2795) >= ((reg2806 && reg2789) ~^ reg2777[(3'h6):(3'h5)]));
                      reg2832 <= {$signed($signed({wire1760}))};
                      reg2833 <= wire2751;
                    end
                  if (($unsigned($signed($signed(reg2788))) && $signed(((reg2755 ?
                          reg2759 : forvar2821) ?
                      forvar2826[(3'h5):(2'h2)] : $unsigned(forvar2793)))))
                    begin
                      reg2834 <= $signed((reg2817[(1'h1):(1'h1)] != $unsigned(reg2768)));
                      reg2835 <= {$signed({(~forvar2808)})};
                      reg2836 <= reg2786[(3'h7):(3'h5)];
                      reg2837 <= ($signed(((wire2753 <= (8'ha6)) ?
                          reg2778 : (-reg2828))) <= forvar2774[(4'h8):(3'h5)]);
                    end
                  else
                    begin
                      reg2834 <= {$signed({forvar2809})};
                      reg2835 <= forvar2755;
                    end
                end
              if (((~|(^$signed(reg2788))) + reg2802[(1'h1):(1'h1)]))
                begin
                  for (forvar2838 = (1'h0); (forvar2838 < (1'h1)); forvar2838 = (forvar2838 + (1'h1)))
                    begin
                      reg2839 <= forvar2799;
                      reg2840 <= $signed(reg2779[(2'h3):(1'h1)]);
                      reg2841 <= (((^(^forvar2808)) ?
                              $signed($unsigned((8'hb2))) : reg2810[(4'h8):(4'h8)]) ?
                          (reg2817[(2'h2):(1'h1)] ?
                              $signed($unsigned(reg2762)) : wire2753[(4'h8):(2'h3)]) : {reg2794[(3'h4):(2'h2)]});
                    end
                  for (forvar2842 = (1'h0); (forvar2842 < (1'h0)); forvar2842 = (forvar2842 + (1'h1)))
                    begin
                      reg2843 <= $unsigned(forvar2770[(1'h1):(1'h0)]);
                    end
                  for (forvar2844 = (1'h0); (forvar2844 < (2'h3)); forvar2844 = (forvar2844 + (1'h1)))
                    begin
                      reg2845 <= (reg2817[(1'h1):(1'h0)] ?
                          (&(8'ha4)) : ((~^(reg2789 >= reg2819)) >>> {$unsigned(forvar2829)}));
                      reg2846 <= forvar2798[(2'h2):(1'h1)];
                      reg2847 <= $unsigned((+(!(^forvar2755))));
                      reg2848 <= ($unsigned(((forvar2842 ? reg2769 : reg2836) ?
                          $unsigned(reg2835) : $unsigned(reg2803))) * (forvar2774[(2'h3):(2'h2)] ~^ $unsigned(reg2810)));
                    end
                end
              else
                begin
                  if ($unsigned($unsigned(reg2765[(2'h2):(1'h0)])))
                    begin
                      reg2838 <= ($signed(reg2771[(1'h1):(1'h0)]) ?
                          $signed({(&(8'hb4))}) : ((+(8'ha7)) == ((reg2840 ?
                                  forvar2797 : reg2830) ?
                              (reg2836 ?
                                  reg2789 : reg2759) : $unsigned(reg2815))));
                      reg2839 <= wire1761;
                      reg2840 <= (&(~^(~|(reg2810 != reg2783))));
                    end
                  else
                    begin
                      reg2838 <= ((+(wire1762[(3'h5):(3'h4)] < reg2805[(3'h4):(1'h1)])) ?
                          reg2836 : reg2813[(3'h5):(3'h4)]);
                    end
                  if ($signed((~&$unsigned((^reg2782)))))
                    begin
                      reg2841 <= (8'ha4);
                    end
                  else
                    begin
                      reg2841 <= (($signed($signed(reg2840)) ?
                              $unsigned((forvar2793 ?
                                  (8'hae) : reg2819)) : reg2833) ?
                          (|(~&(reg2796 - forvar2798))) : $signed({{reg2836}}));
                      reg2842 <= reg2820[(3'h4):(2'h2)];
                    end
                end
            end
          for (forvar2849 = (1'h0); (forvar2849 < (1'h0)); forvar2849 = (forvar2849 + (1'h1)))
            begin
              if ($signed((-forvar2803)))
                begin
                  if ((((-reg2779[(1'h0):(1'h0)]) ?
                          (~|(forvar2754 ? reg2800 : reg2824)) : (|reg2815)) ?
                      ((reg2756[(2'h2):(1'h0)] ~^ (reg2777 ?
                              (8'hb3) : forvar2801)) ?
                          {(&(8'ha7))} : ((forvar2754 ? reg2777 : (8'ha6)) ?
                              $unsigned(reg2836) : $signed(reg2773))) : reg2800))
                    begin
                      reg2850 <= (~({(reg2825 ? reg2803 : forvar2755)} ?
                          ((reg2798 ?
                              reg2837 : forvar2774) > $signed(reg2795)) : $unsigned(reg2798)));
                    end
                  else
                    begin
                      reg2850 <= (reg2832 ? (reg2836 >> reg2780) : wire1762);
                      reg2851 <= {(reg2791 - forvar2783[(2'h3):(1'h1)])};
                    end
                  if ($signed(reg2773))
                    begin
                      reg2852 <= {reg2805};
                      reg2853 <= ($unsigned({{(8'hb6)}}) ?
                          ((+{reg2840}) ^~ ($signed(reg2836) * forvar2776[(4'h8):(3'h5)])) : $signed((8'hb9)));
                      reg2854 <= ({(~&(^reg2779))} - ($unsigned($unsigned(reg2817)) ?
                          (~|(reg2840 ?
                              reg2771 : (8'hb2))) : $unsigned((reg2815 ?
                              (8'hb4) : wire1760))));
                    end
                  else
                    begin
                      reg2852 <= $unsigned((~$unsigned(reg2823[(1'h0):(1'h0)])));
                      reg2853 <= reg2839[(2'h2):(2'h2)];
                      reg2854 <= reg2811;
                    end
                  for (forvar2855 = (1'h0); (forvar2855 < (1'h0)); forvar2855 = (forvar2855 + (1'h1)))
                    begin
                      reg2856 <= ($unsigned(forvar2801[(2'h3):(1'h1)]) ?
                          (~^($unsigned(reg2782) ?
                              {(8'had)} : $signed(reg2778))) : reg2825);
                      reg2857 <= (($unsigned((-reg2782)) ?
                          $unsigned(reg2761) : reg2785[(3'h6):(3'h4)]) ^~ ((^~((8'hb6) | (8'hb7))) << ((~|reg2810) < ((8'ha2) ?
                          reg2766 : reg2820))));
                    end
                  for (forvar2858 = (1'h0); (forvar2858 < (1'h0)); forvar2858 = (forvar2858 + (1'h1)))
                    begin
                      reg2859 <= reg2762[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar2850 = (1'h0); (forvar2850 < (2'h3)); forvar2850 = (forvar2850 + (1'h1)))
                    begin
                      reg2851 <= reg2807;
                      reg2852 <= (reg2837 ?
                          (reg2843[(1'h0):(1'h0)] ?
                              (!$signed(reg2814)) : ((^~reg2765) - reg2857[(1'h0):(1'h0)])) : (reg2801 == $signed(((8'had) ?
                              reg2813 : reg2802))));
                      reg2853 <= ({forvar2821} ?
                          {($unsigned(forvar2797) - $unsigned(forvar2821))} : $unsigned(((reg2810 ?
                              reg2815 : reg2772) ~^ $unsigned(reg2792))));
                      reg2854 <= (({(forvar2781 ?
                                  reg2859 : reg2852)} && ((!forvar2850) ?
                              reg2831 : (8'h9e))) ?
                          forvar2858[(2'h2):(1'h0)] : (reg2801[(4'h8):(4'h8)] ?
                              (8'h9c) : ($signed(forvar2790) & reg2847)));
                    end
                  for (forvar2855 = (1'h0); (forvar2855 < (1'h1)); forvar2855 = (forvar2855 + (1'h1)))
                    begin
                      reg2856 <= $signed($signed((forvar2829[(4'h9):(4'h9)] == reg2789[(3'h4):(3'h4)])));
                      reg2857 <= (8'hab);
                      reg2858 <= ((reg2834 ?
                              forvar2776[(4'h9):(4'h9)] : ((&reg2771) | (reg2803 ?
                                  forvar2844 : reg2815))) ?
                          ((8'ha9) << {reg2780[(3'h7):(1'h0)]}) : (reg2755 ?
                              reg2817 : reg2769));
                    end
                end
            end
        end
      else
        begin
          for (forvar2774 = (1'h0); (forvar2774 < (2'h3)); forvar2774 = (forvar2774 + (1'h1)))
            begin
              reg2775 <= $signed($unsigned(reg2800));
            end
          reg2776 <= $unsigned($unsigned($signed(reg2850[(3'h4):(2'h2)])));
          for (forvar2777 = (1'h0); (forvar2777 < (2'h3)); forvar2777 = (forvar2777 + (1'h1)))
            begin
              if ($signed((~$signed((forvar2849 == reg2816)))))
                begin
                  reg2778 <= ((^~$signed($signed(reg2828))) ?
                      ((!$unsigned(reg2837)) >= ($unsigned(reg2768) ?
                          forvar2844 : $signed(forvar2858))) : $unsigned(reg2806[(4'hb):(3'h5)]));
                end
              else
                begin
                  for (forvar2778 = (1'h0); (forvar2778 < (1'h0)); forvar2778 = (forvar2778 + (1'h1)))
                    begin
                      reg2779 <= $unsigned({$signed({wire2753})});
                      reg2780 <= ($signed($signed($signed(wire2752))) || ($unsigned($unsigned(reg2834)) ?
                          reg2773[(3'h7):(3'h4)] : reg2794));
                      reg2781 <= forvar2838;
                      reg2782 <= reg2800;
                    end
                  if ($unsigned($unsigned((forvar2822[(1'h0):(1'h0)] * ((8'hb9) <= forvar2801)))))
                    begin
                      reg2783 <= {(~^{reg2786[(4'hc):(4'h9)]})};
                      reg2784 <= reg2776;
                      reg2785 <= ($unsigned({(reg2838 + reg2759)}) >>> ((~$signed((8'haa))) ~^ ($unsigned(reg2786) << $unsigned(forvar2764))));
                    end
                  else
                    begin
                      reg2783 <= $signed({reg2810});
                      reg2784 <= (({$signed((8'hb0))} > ($signed(reg2858) * reg2784[(4'h8):(3'h4)])) >>> (((+(8'hb9)) ?
                          (8'ha6) : ((8'hb7) ?
                              reg2763 : reg2837)) & (|$unsigned(reg2798))));
                      reg2785 <= {$signed((-$unsigned(forvar2803)))};
                      reg2786 <= reg2761;
                    end
                  if ((reg2763[(2'h2):(2'h2)] != (reg2812 ?
                      $unsigned((!reg2841)) : (8'ha9))))
                    begin
                      reg2787 <= (reg2851[(2'h2):(1'h0)] ?
                          $signed(reg2850) : (forvar2790 ^~ forvar2829[(2'h2):(1'h1)]));
                      reg2788 <= $signed((8'h9d));
                    end
                  else
                    begin
                      reg2787 <= forvar2850;
                    end
                  if (reg2775)
                    begin
                      reg2789 <= ($unsigned(((forvar2790 >= reg2815) >= $unsigned(reg2845))) ^ {reg2803});
                    end
                  else
                    begin
                      reg2789 <= reg2830[(1'h0):(1'h0)];
                      reg2790 <= forvar2797[(3'h7):(2'h3)];
                      reg2791 <= $signed(forvar2849);
                      reg2792 <= ((((|reg2816) || (^forvar2770)) ?
                              reg2767[(1'h1):(1'h0)] : (reg2853[(1'h0):(1'h0)] ?
                                  (^reg2815) : (8'hab))) ?
                          (((forvar2764 ?
                                  reg2801 : reg2789) <<< (reg2767 >= (8'ha9))) ?
                              reg2842[(1'h1):(1'h0)] : ((+reg2803) >> {reg2806})) : (-$unsigned((!reg2794))));
                    end
                end
              reg2793 <= ((-reg2847[(3'h4):(2'h2)]) ?
                  (&$signed((~reg2815))) : reg2859);
            end
        end
      if (forvar2799[(1'h0):(1'h0)])
        begin
          if (((~|($unsigned(reg2833) ?
              reg2758[(3'h7):(1'h1)] : (reg2820 ?
                  reg2778 : wire2753))) >> $unsigned({(reg2831 ~^ reg2825)})))
            begin
              for (forvar2860 = (1'h0); (forvar2860 < (2'h3)); forvar2860 = (forvar2860 + (1'h1)))
                begin
                  if (($unsigned((~reg2833[(1'h1):(1'h0)])) > (+reg2813[(3'h4):(2'h2)])))
                    begin
                      reg2861 <= $unsigned((reg2854 > reg2800[(3'h5):(3'h4)]));
                      reg2862 <= $unsigned($unsigned((forvar2770[(2'h3):(2'h2)] + $signed(forvar2808))));
                      reg2863 <= reg2789[(4'hd):(2'h2)];
                      reg2864 <= (!($signed(reg2814[(4'h9):(3'h7)]) ?
                          ($signed(forvar2844) && (wire1762 ?
                              reg2782 : wire2749)) : $unsigned($signed(reg2841))));
                    end
                  else
                    begin
                      reg2861 <= {$unsigned($unsigned((-forvar2850)))};
                      reg2862 <= ((((8'ha2) >> $signed(reg2830)) ?
                          reg2836 : (+$signed(reg2831))) || forvar2793);
                      reg2863 <= (~&(($unsigned(reg2801) >>> forvar2821) ?
                          (&(&(8'h9c))) : (-(~|(8'had)))));
                    end
                  for (forvar2865 = (1'h0); (forvar2865 < (1'h0)); forvar2865 = (forvar2865 + (1'h1)))
                    begin
                      reg2866 <= $unsigned(reg2838);
                      reg2867 <= (reg2837[(1'h0):(1'h0)] ?
                          (~^reg2864[(2'h3):(1'h0)]) : (~&forvar2801[(4'hd):(4'h8)]));
                    end
                  if (({(!$signed((8'hba)))} | $signed($unsigned({reg2866}))))
                    begin
                      reg2868 <= {reg2856};
                      reg2869 <= reg2818[(1'h1):(1'h0)];
                      reg2870 <= $signed((reg2820[(4'hb):(1'h0)] & (reg2760[(4'hf):(4'h9)] == (reg2837 || (8'hb3)))));
                      reg2871 <= reg2842[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2868 <= ((8'haf) << (|$unsigned(reg2804)));
                      reg2869 <= $unsigned((forvar2799 ?
                          $unsigned(reg2831[(2'h2):(1'h1)]) : reg2771[(1'h0):(1'h0)]));
                      reg2870 <= $signed(forvar2822[(2'h2):(2'h2)]);
                      reg2871 <= ((8'h9d) ^ $unsigned(($unsigned(reg2793) ^~ reg2796[(1'h1):(1'h0)])));
                    end
                  for (forvar2872 = (1'h0); (forvar2872 < (2'h3)); forvar2872 = (forvar2872 + (1'h1)))
                    begin
                      reg2873 <= reg2771[(1'h1):(1'h0)];
                      reg2874 <= {(reg2851 ? (8'ha8) : {(reg2856 >= (8'hab))})};
                      reg2875 <= reg2778;
                    end
                end
            end
          else
            begin
              reg2860 <= (($signed((^reg2850)) - ((reg2788 ^~ (8'ha3)) > (!reg2818))) || forvar2865[(3'h5):(1'h0)]);
              for (forvar2861 = (1'h0); (forvar2861 < (2'h2)); forvar2861 = (forvar2861 + (1'h1)))
                begin
                  if ($unsigned($unsigned(reg2824[(1'h1):(1'h0)])))
                    begin
                      reg2862 <= ($signed(wire2749) * reg2837);
                      reg2863 <= $unsigned(reg2776);
                      reg2864 <= ((((forvar2776 ? reg2847 : reg2843) ?
                          reg2846[(4'h8):(3'h6)] : $signed((8'h9f))) <<< forvar2829[(2'h2):(2'h2)]) == reg2859[(2'h3):(2'h2)]);
                      reg2865 <= $unsigned((reg2757[(2'h2):(1'h1)] ?
                          (8'ha7) : ($signed(reg2798) ? reg2819 : (|reg2838))));
                    end
                  else
                    begin
                      reg2862 <= {{$signed((forvar2781 ? reg2769 : reg2839))}};
                      reg2863 <= forvar2838[(2'h3):(1'h1)];
                      reg2864 <= (reg2846[(4'h8):(1'h0)] ?
                          $unsigned($unsigned((reg2784 ?
                              reg2870 : forvar2801))) : (~&$signed(reg2761)));
                    end
                  for (forvar2866 = (1'h0); (forvar2866 < (2'h2)); forvar2866 = (forvar2866 + (1'h1)))
                    begin
                      reg2867 <= $unsigned(((((8'h9d) ? reg2840 : forvar2781) ?
                          forvar2774[(4'ha):(2'h3)] : {forvar2775}) > ((reg2791 + (8'hab)) ?
                          (reg2813 == forvar2774) : ((8'hb7) ?
                              reg2835 : reg2824))));
                      reg2868 <= ($signed($signed(reg2848[(4'h9):(1'h0)])) ?
                          $signed({$signed(reg2861)}) : ($unsigned($unsigned(forvar2842)) ?
                              $unsigned({reg2800}) : reg2815[(3'h4):(1'h0)]));
                      reg2869 <= forvar2764[(4'h8):(1'h1)];
                      reg2870 <= ($unsigned(forvar2808) ?
                          $unsigned((forvar2770[(2'h3):(1'h0)] >> $signed(reg2783))) : {(8'ha7)});
                    end
                  for (forvar2871 = (1'h0); (forvar2871 < (1'h1)); forvar2871 = (forvar2871 + (1'h1)))
                    begin
                      reg2872 <= (forvar2844[(4'hb):(3'h5)] ?
                          ((reg2787 ?
                              (reg2772 >= reg2810) : forvar2860[(1'h1):(1'h1)]) + ($signed(forvar2809) ~^ reg2842)) : reg2792[(4'h9):(3'h5)]);
                      reg2873 <= (^(^((&reg2862) ?
                          $signed(reg2865) : $unsigned(wire2749))));
                      reg2874 <= ((^$unsigned(forvar2764[(3'h5):(3'h5)])) ?
                          (reg2776 & ((reg2869 && wire2752) << $signed(reg2801))) : reg2850[(2'h2):(1'h1)]);
                      reg2875 <= forvar2822;
                    end
                  for (forvar2876 = (1'h0); (forvar2876 < (2'h3)); forvar2876 = (forvar2876 + (1'h1)))
                    begin
                      reg2877 <= ((|(-reg2781)) ?
                          $unsigned($unsigned(reg2843)) : (reg2781[(1'h0):(1'h0)] ?
                              reg2834 : ($signed(reg2839) ?
                                  (reg2871 ?
                                      reg2796 : (8'ha8)) : reg2854[(4'hb):(4'hb)])));
                    end
                end
              reg2878 <= ((^~reg2773) & $unsigned((^{reg2811})));
            end
          for (forvar2879 = (1'h0); (forvar2879 < (1'h1)); forvar2879 = (forvar2879 + (1'h1)))
            begin
              reg2880 <= ((~reg2816[(1'h1):(1'h0)]) ^ $unsigned($unsigned(reg2877)));
            end
        end
      else
        begin
          for (forvar2860 = (1'h0); (forvar2860 < (1'h0)); forvar2860 = (forvar2860 + (1'h1)))
            begin
              for (forvar2861 = (1'h0); (forvar2861 < (1'h0)); forvar2861 = (forvar2861 + (1'h1)))
                begin
                  for (forvar2862 = (1'h0); (forvar2862 < (1'h1)); forvar2862 = (forvar2862 + (1'h1)))
                    begin
                      reg2863 <= (-reg2838[(3'h5):(1'h0)]);
                      reg2864 <= reg2865;
                    end
                  for (forvar2865 = (1'h0); (forvar2865 < (1'h1)); forvar2865 = (forvar2865 + (1'h1)))
                    begin
                      reg2866 <= (~reg2838[(2'h3):(2'h2)]);
                    end
                  reg2867 <= (reg2877[(2'h3):(1'h1)] ?
                      $unsigned(((~&reg2791) | $signed(reg2810))) : $unsigned(((reg2858 ?
                          reg2785 : reg2819) ~^ (!reg2865))));
                  for (forvar2868 = (1'h0); (forvar2868 < (2'h3)); forvar2868 = (forvar2868 + (1'h1)))
                    begin
                      reg2869 <= (^~{(reg2864[(3'h4):(3'h4)] ^~ $unsigned(reg2768))});
                      reg2870 <= {(^(-(reg2848 <= reg2847)))};
                      reg2871 <= ($unsigned(reg2852) ~^ {reg2877[(3'h6):(2'h3)]});
                    end
                end
              for (forvar2872 = (1'h0); (forvar2872 < (1'h0)); forvar2872 = (forvar2872 + (1'h1)))
                begin
                  for (forvar2873 = (1'h0); (forvar2873 < (2'h3)); forvar2873 = (forvar2873 + (1'h1)))
                    begin
                      reg2874 <= (($signed($unsigned(forvar2862)) ?
                              reg2864 : reg2798[(2'h2):(2'h2)]) ?
                          reg2853 : $unsigned(((forvar2860 || reg2803) ?
                              $signed((8'hb5)) : $unsigned(reg2861))));
                      reg2875 <= $unsigned(((-(forvar2844 != (8'had))) > ($unsigned(forvar2801) ?
                          reg2811[(3'h4):(2'h3)] : {reg2786})));
                      reg2876 <= (~{reg2838[(3'h4):(1'h1)]});
                      reg2877 <= reg2792;
                    end
                  for (forvar2878 = (1'h0); (forvar2878 < (2'h3)); forvar2878 = (forvar2878 + (1'h1)))
                    begin
                      reg2879 <= $signed($signed({(!reg2781)}));
                      reg2880 <= ((^(!$signed(reg2842))) ?
                          (reg2860 ?
                              forvar2783[(4'hb):(4'h9)] : reg2759[(3'h7):(2'h3)]) : $signed($signed(forvar2862)));
                      reg2881 <= {$unsigned($signed(reg2836[(2'h2):(1'h0)]))};
                      reg2882 <= {$signed($unsigned(reg2843))};
                    end
                  if (((($signed(reg2856) ?
                          reg2858[(2'h2):(1'h0)] : ((8'h9c) ?
                              reg2853 : reg2818)) || (8'ha1)) ?
                      wire1761 : reg2758))
                    begin
                      reg2883 <= $unsigned($signed(({reg2766} ?
                          {forvar2879} : (reg2833 ? (8'hac) : forvar2866))));
                      reg2884 <= $unsigned($unsigned(($unsigned(reg2840) ?
                          (reg2863 & forvar2838) : (-reg2756))));
                      reg2885 <= (^~(!reg2803));
                    end
                  else
                    begin
                      reg2883 <= (^(8'hb8));
                      reg2884 <= (~(^reg2767[(1'h0):(1'h0)]));
                    end
                  for (forvar2886 = (1'h0); (forvar2886 < (2'h2)); forvar2886 = (forvar2886 + (1'h1)))
                    begin
                      reg2887 <= (((reg2869[(3'h6):(2'h2)] <= $unsigned(reg2852)) ?
                          $signed((!(8'ha2))) : (|forvar2822[(4'hb):(4'ha)])) == {(|reg2869)});
                      reg2888 <= (8'hb9);
                      reg2889 <= reg2781;
                      reg2890 <= reg2854;
                    end
                end
            end
          if ($signed(wire2753[(1'h0):(1'h0)]))
            begin
              for (forvar2891 = (1'h0); (forvar2891 < (2'h2)); forvar2891 = (forvar2891 + (1'h1)))
                begin
                  for (forvar2892 = (1'h0); (forvar2892 < (1'h1)); forvar2892 = (forvar2892 + (1'h1)))
                    begin
                      reg2893 <= ($unsigned(reg2888[(3'h6):(3'h6)]) != (~^$signed((~reg2843))));
                      reg2894 <= $unsigned(($signed(wire1761) ?
                          (~^(reg2873 + reg2876)) : $unsigned({reg2836})));
                      reg2895 <= ($signed(($unsigned(reg2818) ?
                          (+forvar2858) : (8'hb9))) <<< $signed((+$signed(forvar2777))));
                      reg2896 <= reg2816[(2'h2):(1'h1)];
                    end
                  for (forvar2897 = (1'h0); (forvar2897 < (1'h0)); forvar2897 = (forvar2897 + (1'h1)))
                    begin
                      reg2898 <= reg2766[(4'hc):(1'h1)];
                    end
                end
              for (forvar2899 = (1'h0); (forvar2899 < (1'h0)); forvar2899 = (forvar2899 + (1'h1)))
                begin
                  if (({$unsigned($signed(reg2813))} ?
                      ((&$signed(forvar2778)) ?
                          wire2749[(1'h0):(1'h0)] : $signed($signed(reg2787))) : (reg2831[(1'h0):(1'h0)] == forvar2850)))
                    begin
                      reg2900 <= reg2839;
                      reg2901 <= reg2841;
                    end
                  else
                    begin
                      reg2900 <= $signed(({(~reg2843)} ?
                          ((reg2816 <= reg2834) ?
                              (-reg2768) : ((8'ha7) * reg2858)) : ((reg2791 ^ forvar2858) ?
                              reg2867[(4'hc):(1'h1)] : $unsigned(forvar2844))));
                      reg2901 <= ((8'hb7) ?
                          (~(~^(^reg2867))) : (|(forvar2764 << (|reg2831))));
                      reg2902 <= {$unsigned((^$unsigned((8'haf))))};
                      reg2903 <= ($signed(reg2756) ?
                          forvar2891[(3'h4):(1'h1)] : $signed(reg2790));
                    end
                end
            end
          else
            begin
              for (forvar2891 = (1'h0); (forvar2891 < (2'h2)); forvar2891 = (forvar2891 + (1'h1)))
                begin
                  for (forvar2892 = (1'h0); (forvar2892 < (2'h2)); forvar2892 = (forvar2892 + (1'h1)))
                    begin
                      reg2893 <= reg2772;
                      reg2894 <= (forvar2886 >= $signed(reg2769[(3'h6):(2'h3)]));
                      reg2895 <= ($signed($signed(forvar2799)) ?
                          $unsigned($unsigned((forvar2798 ?
                              (8'hac) : reg2859))) : (^(reg2845[(1'h0):(1'h0)] ?
                              $unsigned(forvar2799) : reg2893)));
                      reg2896 <= (~reg2859);
                    end
                  if (((forvar2809 ?
                      (~^forvar2790[(2'h2):(1'h0)]) : (reg2802[(3'h7):(2'h3)] ^ {reg2839})) >> reg2861[(1'h1):(1'h0)]))
                    begin
                      reg2897 <= ((wire2753 ?
                              {(forvar2892 ?
                                      reg2796 : forvar2850)} : $unsigned(reg2902)) ?
                          ({$unsigned(forvar2799)} ?
                              forvar2861 : reg2881[(4'hc):(4'h8)]) : $signed((forvar2808 ?
                              $signed((8'hab)) : (&reg2804))));
                      reg2898 <= (-$unsigned(((~|reg2792) | $signed(reg2888))));
                    end
                  else
                    begin
                      reg2897 <= $signed(($unsigned($unsigned(reg2837)) ?
                          ({(8'ha9)} ?
                              reg2798[(3'h6):(2'h2)] : $signed(forvar2797)) : ((forvar2862 | forvar2855) ?
                              reg2878 : (~|reg2860))));
                      reg2898 <= $signed((8'had));
                    end
                  for (forvar2899 = (1'h0); (forvar2899 < (2'h3)); forvar2899 = (forvar2899 + (1'h1)))
                    begin
                      reg2900 <= $signed((!$signed({(8'h9e)})));
                      reg2901 <= (~|($signed(reg2767) ^~ $unsigned(wire1762)));
                    end
                end
              for (forvar2902 = (1'h0); (forvar2902 < (1'h0)); forvar2902 = (forvar2902 + (1'h1)))
                begin
                  if ($signed((~|($signed(reg2866) > forvar2770[(1'h0):(1'h0)]))))
                    begin
                      reg2903 <= (~|$signed($signed((forvar2860 ?
                          reg2861 : forvar2879))));
                      reg2904 <= $unsigned(((reg2873 << (reg2895 ?
                          reg2845 : reg2758)) | reg2858));
                      reg2905 <= ((&$signed((reg2847 ? reg2865 : forvar2829))) ?
                          $signed({{reg2792}}) : $unsigned(reg2769));
                      reg2906 <= (((+reg2846[(1'h1):(1'h1)]) && $unsigned((forvar2897 ?
                              reg2837 : reg2852))) ?
                          $signed((8'ha3)) : reg2785);
                    end
                  else
                    begin
                      reg2903 <= (-((~|reg2878[(4'hb):(2'h2)]) ?
                          forvar2860[(4'ha):(3'h6)] : $unsigned(((8'ha0) ?
                              forvar2821 : forvar2858))));
                      reg2904 <= $signed($signed($unsigned((forvar2860 ?
                          reg2814 : forvar2892))));
                      reg2905 <= reg2867;
                    end
                  reg2907 <= reg2825[(3'h6):(3'h5)];
                  for (forvar2908 = (1'h0); (forvar2908 < (1'h0)); forvar2908 = (forvar2908 + (1'h1)))
                    begin
                      reg2909 <= ($signed(reg2814[(4'h9):(4'h9)]) ?
                          ((~&(reg2772 >>> reg2783)) != ({wire1761} ?
                              (^reg2806) : reg2856)) : $unsigned($signed($unsigned(forvar2873))));
                    end
                  reg2910 <= reg2818;
                end
              reg2911 <= $unsigned((8'ha3));
              for (forvar2912 = (1'h0); (forvar2912 < (1'h0)); forvar2912 = (forvar2912 + (1'h1)))
                begin
                  if ($signed(((reg2862[(1'h1):(1'h0)] & (8'hb6)) <<< $unsigned((forvar2861 ?
                      forvar2868 : reg2894)))))
                    begin
                      reg2913 <= $signed(reg2865[(4'hc):(2'h3)]);
                      reg2914 <= forvar2871;
                      reg2915 <= {((~&reg2807) + reg2859[(2'h2):(1'h0)])};
                    end
                  else
                    begin
                      reg2913 <= reg2832;
                      reg2914 <= $signed({((8'hb9) > (reg2868 != reg2803))});
                    end
                end
            end
          reg2916 <= reg2825[(1'h0):(1'h0)];
          if ($signed((((reg2862 || (8'hb5)) ? {reg2843} : $signed(reg2758)) ?
              (reg2761 ? {reg2812} : (reg2902 != forvar2822)) : (reg2780 ?
                  reg2831 : forvar2822[(4'hb):(4'hb)]))))
            begin
              if (reg2910)
                begin
                  for (forvar2917 = (1'h0); (forvar2917 < (2'h3)); forvar2917 = (forvar2917 + (1'h1)))
                    begin
                      reg2918 <= $unsigned(reg2881[(5'h10):(3'h5)]);
                      reg2919 <= $unsigned(reg2765[(1'h1):(1'h0)]);
                    end
                  for (forvar2920 = (1'h0); (forvar2920 < (2'h3)); forvar2920 = (forvar2920 + (1'h1)))
                    begin
                      reg2921 <= ($unsigned($unsigned((reg2841 && reg2767))) ^~ forvar2778[(3'h7):(3'h6)]);
                      reg2922 <= (^~($unsigned($signed(forvar2912)) >>> (-(reg2785 ?
                          reg2831 : reg2900))));
                    end
                  if (((~|(-(reg2835 ? reg2866 : reg2840))) ?
                      reg2831[(3'h7):(2'h2)] : forvar2776))
                    begin
                      reg2923 <= (+(($signed(forvar2866) ?
                              (-reg2802) : (8'ha1)) ?
                          reg2835 : $signed((reg2921 != reg2889))));
                    end
                  else
                    begin
                      reg2923 <= reg2914[(3'h5):(3'h5)];
                      reg2924 <= forvar2899[(3'h5):(2'h2)];
                    end
                end
              else
                begin
                  if (reg2907)
                    begin
                      reg2917 <= (reg2791 + (+((forvar2764 ?
                              forvar2826 : forvar2902) ?
                          $signed(forvar2770) : (reg2887 ?
                              reg2859 : reg2815))));
                      reg2918 <= (~$signed($signed($unsigned(forvar2868))));
                      reg2919 <= (~|(forvar2842 ?
                          $unsigned($unsigned(reg2802)) : (reg2803[(3'h4):(3'h4)] ?
                              forvar2793[(3'h5):(2'h3)] : (!reg2815))));
                    end
                  else
                    begin
                      reg2917 <= $unsigned(((8'ha1) ?
                          $signed((reg2799 <= reg2884)) : $unsigned((forvar2858 ?
                              forvar2764 : forvar2764))));
                      reg2918 <= $signed(($signed($signed(reg2807)) <= $signed((reg2786 < reg2800))));
                    end
                end
              for (forvar2925 = (1'h0); (forvar2925 < (2'h2)); forvar2925 = (forvar2925 + (1'h1)))
                begin
                  reg2926 <= (forvar2842 * ($signed(reg2803) ?
                      reg2903[(1'h1):(1'h1)] : $unsigned((~^reg2919))));
                  for (forvar2927 = (1'h0); (forvar2927 < (1'h1)); forvar2927 = (forvar2927 + (1'h1)))
                    begin
                      reg2928 <= ((-$signed((reg2902 ?
                          reg2787 : forvar2775))) >= $unsigned($signed($unsigned(reg2910))));
                      reg2929 <= ((-reg2882) ?
                          {((reg2820 ?
                                  (8'hb8) : reg2790) < $signed(wire1762))} : reg2772[(1'h0):(1'h0)]);
                    end
                end
            end
          else
            begin
              if ($signed((~^reg2803)))
                begin
                  for (forvar2917 = (1'h0); (forvar2917 < (2'h2)); forvar2917 = (forvar2917 + (1'h1)))
                    begin
                      reg2918 <= ((((forvar2801 >> reg2805) ?
                              {(8'ha6)} : $unsigned(forvar2891)) ?
                          (~(reg2802 ?
                              reg2762 : reg2793)) : $unsigned(reg2828)) <<< (^~$unsigned((^~reg2768))));
                      reg2919 <= (forvar2774 ^~ ((|(reg2796 < forvar2873)) ?
                          {forvar2844[(3'h7):(3'h6)]} : forvar2860));
                      reg2920 <= ($signed($unsigned($unsigned((8'hac)))) ^~ (~&{(reg2868 || reg2863)}));
                      reg2921 <= {{($signed((8'hb4)) ?
                                  (~|reg2787) : forvar2822)}};
                    end
                  for (forvar2922 = (1'h0); (forvar2922 < (2'h3)); forvar2922 = (forvar2922 + (1'h1)))
                    begin
                      reg2923 <= (&reg2824);
                    end
                  if ({$signed($signed(reg2884))})
                    begin
                      reg2924 <= $signed((forvar2850 >>> reg2838[(3'h4):(2'h2)]));
                      reg2925 <= (($unsigned(reg2765) ?
                          $signed((-forvar2873)) : ($signed(reg2900) && (reg2917 <<< reg2870))) ~^ reg2776[(4'ha):(3'h5)]);
                      reg2926 <= {$signed($unsigned({reg2807}))};
                      reg2927 <= ((((reg2783 < (8'hae)) ~^ (+reg2916)) << (~|$unsigned(forvar2801))) < ($signed(reg2874) ^~ {forvar2770[(1'h0):(1'h0)]}));
                    end
                  else
                    begin
                      reg2924 <= ({{reg2882}} ?
                          ($unsigned($signed(forvar2793)) ?
                              reg2814 : (~|forvar2764[(3'h5):(1'h1)])) : {reg2813[(2'h2):(1'h1)]});
                      reg2925 <= forvar2776;
                    end
                end
              else
                begin
                  reg2917 <= reg2762;
                  reg2918 <= ($signed($unsigned((~|reg2890))) ?
                      ($unsigned($signed(reg2916)) + ((forvar2922 ?
                          reg2786 : reg2902) >= $unsigned(wire1762))) : reg2870);
                  for (forvar2919 = (1'h0); (forvar2919 < (2'h3)); forvar2919 = (forvar2919 + (1'h1)))
                    begin
                      reg2920 <= ($signed(reg2835[(4'ha):(3'h5)]) ?
                          $unsigned($unsigned((~^forvar2808))) : (-(~&reg2846)));
                      reg2921 <= forvar2850;
                      reg2922 <= ($signed((((8'h9f) * forvar2849) && (reg2803 ?
                              forvar2873 : (8'hb3)))) ?
                          reg2910[(4'hc):(2'h2)] : $unsigned(($unsigned(forvar2808) ?
                              reg2807[(1'h0):(1'h0)] : (reg2788 ?
                                  (8'hac) : forvar2860))));
                    end
                end
              if ($signed(reg2833[(2'h2):(1'h1)]))
                begin
                  reg2928 <= {reg2865[(3'h4):(2'h3)]};
                  if ($signed((+(!reg2878[(3'h4):(1'h0)]))))
                    begin
                      reg2929 <= reg2802;
                      reg2930 <= (&((reg2919[(4'hb):(1'h1)] < (^reg2877)) ?
                          (reg2875[(3'h4):(2'h3)] ?
                              (!reg2915) : reg2834) : (reg2906 ?
                              (~|reg2903) : {reg2864})));
                      reg2931 <= forvar2886;
                      reg2932 <= $signed($unsigned(reg2790[(3'h7):(3'h7)]));
                    end
                  else
                    begin
                      reg2929 <= {$signed((reg2868[(4'h8):(4'h8)] ?
                              reg2914 : $signed(forvar2891)))};
                      reg2930 <= reg2784[(2'h2):(2'h2)];
                    end
                  if ({($signed($unsigned(reg2866)) < {reg2928})})
                    begin
                      reg2933 <= (($signed((reg2860 >= reg2827)) == $signed($signed(forvar2822))) & (&$unsigned((forvar2801 != reg2864))));
                      reg2934 <= (-forvar2876);
                    end
                  else
                    begin
                      reg2933 <= $signed($signed(((^reg2934) ?
                          reg2839[(1'h0):(1'h0)] : $unsigned((8'ha3)))));
                      reg2934 <= ({((~|forvar2822) ?
                              reg2872 : (reg2836 >= wire1760))} > $unsigned($unsigned((reg2852 ?
                          reg2811 : reg2923))));
                      reg2935 <= reg2866[(1'h0):(1'h0)];
                      reg2936 <= reg2935;
                    end
                end
              else
                begin
                  if (reg2876)
                    begin
                      reg2928 <= ((~&(reg2781 ?
                          reg2828 : (reg2769 ^ reg2925))) < (^$signed(((8'hae) > reg2904))));
                      reg2929 <= $signed(wire2752[(2'h3):(2'h2)]);
                      reg2930 <= forvar2868[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg2928 <= $unsigned($signed((reg2931[(2'h2):(1'h0)] ^ reg2787[(1'h1):(1'h1)])));
                      reg2929 <= reg2775;
                      reg2930 <= (|$signed(((reg2889 ?
                          reg2823 : reg2805) - ((8'hb5) ? reg2922 : (8'ha5)))));
                    end
                  for (forvar2931 = (1'h0); (forvar2931 < (1'h0)); forvar2931 = (forvar2931 + (1'h1)))
                    begin
                      reg2932 <= reg2807[(3'h6):(3'h4)];
                      reg2933 <= reg2796[(2'h2):(1'h1)];
                      reg2934 <= reg2901[(4'h9):(1'h0)];
                    end
                  if ($unsigned(reg2857[(1'h1):(1'h1)]))
                    begin
                      reg2935 <= ($unsigned((~|forvar2861[(2'h3):(2'h3)])) << (reg2926[(3'h7):(3'h5)] ?
                          ((reg2805 ? reg2933 : reg2842) ?
                              reg2757[(2'h2):(2'h2)] : $unsigned(forvar2829)) : $signed(reg2925[(2'h2):(1'h1)])));
                      reg2936 <= (reg2907[(1'h1):(1'h1)] ?
                          (reg2911[(3'h5):(1'h1)] ?
                              ((~^reg2795) == {reg2910}) : {reg2793[(2'h2):(2'h2)]}) : $signed((reg2921 ?
                              reg2840[(4'h8):(1'h0)] : {reg2875})));
                      reg2937 <= (+wire1763);
                      reg2938 <= wire2753;
                    end
                  else
                    begin
                      reg2935 <= $signed(reg2792);
                      reg2936 <= reg2814;
                      reg2937 <= forvar2755[(4'hc):(2'h3)];
                      reg2938 <= $signed(((reg2884[(2'h2):(1'h1)] << (&(8'hb8))) ~^ (8'had)));
                    end
                  if (($unsigned((|$signed(reg2905))) ?
                      {$signed((^~reg2870))} : forvar2776[(3'h5):(3'h5)]))
                    begin
                      reg2939 <= forvar2764;
                    end
                  else
                    begin
                      reg2939 <= reg2790[(2'h3):(1'h0)];
                      reg2940 <= $unsigned($signed({(reg2778 ?
                              reg2833 : (8'hb2))}));
                      reg2941 <= reg2788;
                    end
                end
              reg2942 <= (reg2823 ^~ (reg2889[(3'h7):(3'h4)] ?
                  (reg2937[(2'h3):(2'h3)] ~^ (+reg2810)) : (&reg2828)));
            end
        end
      if (reg2773)
        begin
          if (reg2926[(4'hc):(4'h8)])
            begin
              for (forvar2943 = (1'h0); (forvar2943 < (2'h3)); forvar2943 = (forvar2943 + (1'h1)))
                begin
                  for (forvar2944 = (1'h0); (forvar2944 < (1'h1)); forvar2944 = (forvar2944 + (1'h1)))
                    begin
                      reg2945 <= ((forvar2920 ?
                              (reg2902[(1'h1):(1'h0)] ?
                                  $signed(forvar2944) : reg2919) : $unsigned(reg2915)) ?
                          $unsigned($signed($signed(reg2807))) : ((((8'haf) - reg2923) ?
                                  $unsigned(reg2863) : (~^wire2751)) ?
                              ($unsigned(reg2882) <<< (reg2805 && (8'ha8))) : forvar2902[(3'h5):(1'h0)]));
                      reg2946 <= (!$unsigned($unsigned($unsigned(reg2814))));
                    end
                end
              for (forvar2947 = (1'h0); (forvar2947 < (1'h1)); forvar2947 = (forvar2947 + (1'h1)))
                begin
                  for (forvar2948 = (1'h0); (forvar2948 < (2'h2)); forvar2948 = (forvar2948 + (1'h1)))
                    begin
                      reg2949 <= $unsigned(reg2917);
                      reg2950 <= (((&$signed(reg2900)) ?
                          $signed($signed(reg2859)) : ((^~(8'ha9)) ?
                              (reg2890 ?
                                  forvar2809 : forvar2821) : reg2881[(1'h0):(1'h0)])) + $unsigned(($unsigned(forvar2858) ?
                          (reg2919 + reg2766) : (~reg2884))));
                      reg2951 <= ((^(~|(^~(8'hb8)))) ?
                          reg2864 : ($signed((!reg2814)) | ((reg2888 ~^ forvar2897) ?
                              (reg2813 ?
                                  reg2841 : reg2827) : reg2921[(1'h1):(1'h0)])));
                      reg2952 <= (8'ha9);
                    end
                end
              for (forvar2953 = (1'h0); (forvar2953 < (1'h1)); forvar2953 = (forvar2953 + (1'h1)))
                begin
                  if (((((~|reg2862) ? $signed(reg2883) : $signed(reg2932)) ?
                          ((forvar2886 ?
                              reg2888 : reg2870) & reg2832[(3'h5):(1'h1)]) : $unsigned((reg2773 ?
                              reg2863 : wire2751))) ?
                      ((~(&forvar2855)) ?
                          reg2850[(3'h4):(2'h2)] : (-$signed(forvar2902))) : {$unsigned(forvar2774[(3'h5):(3'h5)])}))
                    begin
                      reg2954 <= $unsigned({$unsigned(reg2767)});
                      reg2955 <= $unsigned(((^~$signed(forvar2948)) ^~ $unsigned((wire1761 * reg2882))));
                    end
                  else
                    begin
                      reg2954 <= {$signed((reg2813[(3'h4):(3'h4)] >>> reg2942[(4'h9):(2'h3)]))};
                      reg2955 <= ({((&(8'hb3)) <= $signed(reg2858))} ?
                          $signed((|reg2939)) : $unsigned({(forvar2821 ?
                                  reg2942 : reg2884)}));
                    end
                end
            end
          else
            begin
              reg2943 <= $signed($signed(((^~reg2930) ? (8'hb2) : {reg2913})));
              for (forvar2944 = (1'h0); (forvar2944 < (2'h3)); forvar2944 = (forvar2944 + (1'h1)))
                begin
                  if (reg2775[(4'he):(4'he)])
                    begin
                      reg2945 <= (~^$unsigned(reg2842));
                      reg2946 <= (((forvar2871 ?
                          {(8'ha1)} : $signed((8'ha7))) ^ {$signed((8'hb0))}) - $signed($signed(reg2871[(3'h4):(2'h2)])));
                      reg2947 <= forvar2944;
                    end
                  else
                    begin
                      reg2945 <= (^$signed(($unsigned(reg2865) != $signed((8'h9e)))));
                      reg2946 <= forvar2842;
                      reg2947 <= ($unsigned(forvar2899) ?
                          ($unsigned((8'hac)) ?
                              reg2837[(3'h6):(3'h4)] : forvar2776) : {(~&(reg2762 ?
                                  reg2868 : reg2819))});
                      reg2948 <= (~^(8'hab));
                    end
                  if ((-reg2895))
                    begin
                      reg2949 <= {(((!reg2955) >>> forvar2822) ^~ $signed((reg2932 != reg2875)))};
                      reg2950 <= {$unsigned($signed($signed((8'ha0))))};
                      reg2951 <= ($signed({(-(8'h9c))}) >>> (($signed(reg2773) ?
                              reg2794 : (8'ha1)) ?
                          {$unsigned(reg2760)} : (!wire2749)));
                    end
                  else
                    begin
                      reg2949 <= $unsigned(reg2943[(2'h2):(1'h1)]);
                      reg2950 <= ((!{(^forvar2868)}) ?
                          $signed($unsigned(reg2888[(2'h2):(2'h2)])) : reg2916);
                      reg2951 <= ({forvar2774} <<< reg2857[(2'h3):(1'h1)]);
                    end
                  if (reg2884[(1'h0):(1'h0)])
                    begin
                      reg2952 <= reg2837[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg2952 <= {(~&$signed($signed(reg2793)))};
                      reg2953 <= reg2904;
                      reg2954 <= {(forvar2755 ?
                              (reg2794[(4'h9):(3'h5)] >= $unsigned(reg2785)) : (reg2928[(3'h6):(1'h1)] == (^forvar2809)))};
                    end
                end
              if ((forvar2808[(4'ha):(4'ha)] ?
                  $signed(($unsigned(reg2924) ?
                      forvar2943[(2'h2):(1'h1)] : reg2901[(2'h3):(1'h1)])) : (({reg2788} ?
                      (!reg2910) : reg2833[(1'h0):(1'h0)]) - $signed($unsigned(reg2778)))))
                begin
                  for (forvar2955 = (1'h0); (forvar2955 < (1'h1)); forvar2955 = (forvar2955 + (1'h1)))
                    begin
                      reg2956 <= ((!reg2911[(2'h3):(2'h2)]) ?
                          ((reg2939[(2'h3):(2'h3)] ?
                                  reg2772[(3'h6):(1'h0)] : (-reg2771)) ?
                              $unsigned(reg2907[(1'h0):(1'h0)]) : forvar2892[(4'ha):(4'ha)]) : (reg2795 + (reg2775 ^~ forvar2908)));
                      reg2957 <= (!(^~(+(reg2758 != reg2874))));
                      reg2958 <= forvar2793[(2'h2):(1'h0)];
                    end
                  if (reg2812)
                    begin
                      reg2959 <= (~&{forvar2793});
                      reg2960 <= ((forvar2919 ?
                              $unsigned(reg2911) : reg2931[(2'h2):(2'h2)]) ?
                          $unsigned(reg2890[(3'h5):(2'h2)]) : {($unsigned((8'ha1)) ?
                                  $signed(reg2758) : (8'hb6))});
                    end
                  else
                    begin
                      reg2959 <= (|((~|(reg2890 ?
                          reg2812 : reg2914)) ^~ $unsigned((reg2772 ?
                          reg2931 : reg2883))));
                      reg2960 <= $signed((^~{(|reg2803)}));
                      reg2961 <= (8'hb5);
                      reg2962 <= reg2918[(3'h4):(3'h4)];
                    end
                  for (forvar2963 = (1'h0); (forvar2963 < (1'h1)); forvar2963 = (forvar2963 + (1'h1)))
                    begin
                      reg2964 <= reg2887[(3'h4):(2'h3)];
                      reg2965 <= (~|(($unsigned(reg2879) ?
                              (reg2911 >= forvar2778) : {(8'ha4)}) ?
                          reg2877 : $unsigned(((8'ha9) < reg2805))));
                      reg2966 <= {(!forvar2899[(1'h0):(1'h0)])};
                      reg2967 <= ($unsigned((forvar2826[(3'h5):(3'h5)] ?
                          $signed(forvar2947) : (!forvar2878))) && (($unsigned(reg2765) ?
                          (|reg2823) : (8'ha2)) >= (reg2838 >>> (^reg2818))));
                    end
                end
              else
                begin
                  for (forvar2955 = (1'h0); (forvar2955 < (2'h2)); forvar2955 = (forvar2955 + (1'h1)))
                    begin
                      reg2956 <= (+$unsigned(reg2951));
                    end
                  reg2957 <= $signed($unsigned(($unsigned(reg2806) + reg2890[(4'h9):(2'h3)])));
                end
            end
          if ($signed(forvar2876[(2'h3):(1'h1)]))
            begin
              for (forvar2968 = (1'h0); (forvar2968 < (2'h3)); forvar2968 = (forvar2968 + (1'h1)))
                begin
                  for (forvar2969 = (1'h0); (forvar2969 < (1'h1)); forvar2969 = (forvar2969 + (1'h1)))
                    begin
                      reg2970 <= (+(~&$signed((reg2967 != reg2949))));
                      reg2971 <= reg2781[(2'h3):(2'h3)];
                      reg2972 <= reg2971;
                      reg2973 <= ($unsigned((reg2848[(4'h8):(3'h4)] ^ forvar2920)) ?
                          (reg2927[(3'h7):(2'h3)] ^~ reg2937) : $unsigned($unsigned((forvar2797 + reg2934))));
                    end
                  if (reg2941)
                    begin
                      reg2974 <= (((-$signed(reg2796)) < ($unsigned(reg2961) ^ (reg2814 ?
                          reg2903 : (8'ha9)))) ^~ $unsigned(forvar2912));
                      reg2975 <= forvar2872;
                      reg2976 <= (-(reg2820[(4'ha):(1'h1)] ?
                          reg2910[(4'hb):(2'h2)] : (~$signed(reg2946))));
                    end
                  else
                    begin
                      reg2974 <= forvar2799[(1'h0):(1'h0)];
                      reg2975 <= (reg2940[(4'hc):(3'h4)] <= $signed((^(~|reg2953))));
                      reg2976 <= (^~{(reg2879[(1'h0):(1'h0)] ?
                              (forvar2919 ?
                                  reg2798 : reg2771) : (reg2880 >= reg2870))});
                      reg2977 <= ({(8'hab)} ?
                          $unsigned({{reg2860}}) : reg2825[(2'h3):(2'h2)]);
                    end
                  reg2978 <= (reg2903 & (!(&forvar2799[(1'h1):(1'h1)])));
                  if ($unsigned((&{((8'hb5) << reg2918)})))
                    begin
                      reg2979 <= (~^$unsigned((reg2792 & reg2946)));
                      reg2980 <= $unsigned($signed($unsigned(reg2783)));
                      reg2981 <= reg2756[(1'h1):(1'h0)];
                      reg2982 <= (reg2952[(4'ha):(4'h8)] ?
                          forvar2891[(3'h6):(3'h6)] : (~^(~&(forvar2799 ?
                              (8'hb9) : forvar2897))));
                    end
                  else
                    begin
                      reg2979 <= $signed($signed((|$signed(forvar2858))));
                      reg2980 <= $signed($signed(((forvar2793 ?
                          reg2904 : forvar2850) >= $signed((8'h9d)))));
                    end
                end
              if ($unsigned((^reg2924[(4'hc):(4'hc)])))
                begin
                  for (forvar2983 = (1'h0); (forvar2983 < (1'h1)); forvar2983 = (forvar2983 + (1'h1)))
                    begin
                      reg2984 <= reg2867;
                    end
                  reg2985 <= $signed($signed($signed(reg2914[(4'hd):(1'h0)])));
                end
              else
                begin
                  reg2983 <= $unsigned((~|$unsigned({forvar2868})));
                  if ((8'ha6))
                    begin
                      reg2984 <= $signed($signed($unsigned((~^(8'h9f)))));
                      reg2985 <= $unsigned({(8'had)});
                      reg2986 <= ({$unsigned(reg2806)} ~^ reg2933[(4'h8):(3'h5)]);
                      reg2987 <= (forvar2876 ?
                          $signed($unsigned($unsigned(reg2793))) : reg2840[(3'h5):(3'h4)]);
                    end
                  else
                    begin
                      reg2984 <= $signed((~((~^wire1761) ?
                          $unsigned(reg2845) : $unsigned((8'hae)))));
                    end
                  reg2988 <= (~^reg2798[(1'h1):(1'h1)]);
                  reg2989 <= (-(forvar2969 ?
                      ((~&reg2802) >> (reg2933 && reg2812)) : $unsigned((reg2795 ?
                          reg2972 : reg2960))));
                end
              for (forvar2990 = (1'h0); (forvar2990 < (1'h0)); forvar2990 = (forvar2990 + (1'h1)))
                begin
                  if ($signed($unsigned(reg2906)))
                    begin
                      reg2991 <= ($signed($unsigned(((8'ha8) ?
                              reg2777 : reg2784))) ?
                          (^~reg2763) : $unsigned(reg2917[(3'h7):(3'h5)]));
                    end
                  else
                    begin
                      reg2991 <= forvar2919;
                      reg2992 <= reg2765[(1'h0):(1'h0)];
                    end
                  for (forvar2993 = (1'h0); (forvar2993 < (1'h1)); forvar2993 = (forvar2993 + (1'h1)))
                    begin
                      reg2994 <= ((8'hb5) ?
                          reg2794[(4'h8):(3'h6)] : $signed((+{(8'ha4)})));
                      reg2995 <= reg2785;
                      reg2996 <= (!((~{(8'hb7)}) ?
                          (wire2752 ?
                              $unsigned(reg2903) : (~^reg2919)) : $unsigned($signed(forvar2868))));
                    end
                  if ((^~$signed((+$unsigned((8'haa))))))
                    begin
                      reg2997 <= {(&reg2793[(1'h0):(1'h0)])};
                      reg2998 <= reg2869[(3'h4):(3'h4)];
                      reg2999 <= $signed(forvar2917[(3'h6):(2'h3)]);
                      reg3000 <= $signed(($signed($unsigned(forvar2844)) ?
                          ((reg2769 ? (8'h9c) : reg2765) ?
                              {reg2830} : (reg2772 << reg2769)) : ($unsigned(reg2830) >> $unsigned(reg2958))));
                    end
                  else
                    begin
                      reg2997 <= (|(reg2974[(3'h7):(1'h0)] ?
                          $unsigned(reg2763) : (reg2795 ?
                              ((8'hb1) + reg2904) : (reg2828 && (8'hb0)))));
                      reg2998 <= $signed(reg2777);
                      reg2999 <= $unsigned(($signed(reg2950) > ($unsigned(reg2939) & (reg2843 <<< reg2962))));
                      reg3000 <= $unsigned($signed(forvar2797[(3'h4):(1'h0)]));
                    end
                end
              reg3001 <= (forvar2944[(4'hd):(3'h6)] >> {($unsigned(wire1760) && (reg2889 ?
                      reg2979 : forvar2844))});
            end
          else
            begin
              reg2968 <= $unsigned(reg2985);
              if ({($unsigned((reg2786 ~^ reg2975)) ?
                      ((reg2798 != reg2777) ?
                          (reg2771 && (8'hb2)) : forvar2963) : reg2998[(3'h5):(1'h1)])})
                begin
                  reg2969 <= ($signed((~{(8'hb9)})) ?
                      {{(8'ha9)}} : (~&forvar2944[(1'h0):(1'h0)]));
                  for (forvar2970 = (1'h0); (forvar2970 < (2'h3)); forvar2970 = (forvar2970 + (1'h1)))
                    begin
                      reg2971 <= $unsigned(reg2847[(3'h7):(3'h7)]);
                      reg2972 <= reg2887[(1'h0):(1'h0)];
                      reg2973 <= (~&$unsigned((~|reg2933)));
                    end
                  for (forvar2974 = (1'h0); (forvar2974 < (2'h2)); forvar2974 = (forvar2974 + (1'h1)))
                    begin
                      reg2975 <= {(~|$unsigned((-forvar2797)))};
                      reg2976 <= (~^forvar2822);
                      reg2977 <= $unsigned((forvar2963[(3'h5):(3'h5)] ?
                          reg2794[(4'h8):(3'h5)] : ($unsigned(forvar2912) | (reg2975 << reg2983))));
                    end
                end
              else
                begin
                  for (forvar2969 = (1'h0); (forvar2969 < (2'h3)); forvar2969 = (forvar2969 + (1'h1)))
                    begin
                      reg2970 <= reg2919;
                      reg2971 <= {{forvar2908}};
                      reg2972 <= (!$signed(reg2825));
                    end
                end
              for (forvar2978 = (1'h0); (forvar2978 < (1'h1)); forvar2978 = (forvar2978 + (1'h1)))
                begin
                  if ($unsigned((8'hb0)))
                    begin
                      reg2979 <= (-(((forvar2925 <<< reg2958) ?
                          reg2835[(4'hb):(3'h5)] : (forvar2793 ?
                              reg2813 : reg2880)) && $signed(forvar2879[(3'h5):(2'h3)])));
                      reg2980 <= reg2807;
                      reg2981 <= reg2775;
                    end
                  else
                    begin
                      reg2979 <= (!(reg2863[(2'h3):(1'h1)] << reg2997[(1'h1):(1'h1)]));
                      reg2980 <= {reg2974[(4'ha):(4'ha)]};
                      reg2981 <= (((reg2777 ?
                              forvar2790 : {(8'haf)}) << ((wire2751 && reg2806) * (~&(8'hb0)))) ?
                          reg2847[(1'h0):(1'h0)] : $signed((reg2830[(1'h1):(1'h1)] ?
                              reg2782[(3'h4):(1'h1)] : {reg2896})));
                      reg2982 <= $unsigned($unsigned($signed($unsigned(forvar2897))));
                    end
                end
            end
        end
      else
        begin
          for (forvar2943 = (1'h0); (forvar2943 < (1'h1)); forvar2943 = (forvar2943 + (1'h1)))
            begin
              if ({(~^(wire1760[(4'ha):(3'h6)] > (reg2948 ?
                      forvar2797 : reg2882)))})
                begin
                  if ({{($unsigned(wire2749) >= {reg2767})}})
                    begin
                      reg2944 <= $unsigned($unsigned(reg2799[(3'h6):(2'h3)]));
                      reg2945 <= $unsigned($signed($unsigned((!reg2924))));
                      reg2946 <= {($signed($unsigned(reg2916)) ?
                              (forvar2953[(1'h0):(1'h0)] > (reg2841 ?
                                  (8'ha9) : reg2999)) : reg2791[(5'h10):(2'h3)])};
                    end
                  else
                    begin
                      reg2944 <= forvar2983;
                      reg2945 <= (-wire2752[(3'h5):(3'h4)]);
                      reg2946 <= forvar2876[(2'h3):(1'h1)];
                      reg2947 <= reg2939;
                    end
                  if (reg2976)
                    begin
                      reg2948 <= {($signed(reg2924[(3'h7):(2'h2)]) ?
                              $unsigned({(8'hb1)}) : {(forvar2797 <= reg2879)})};
                      reg2949 <= ($unsigned(($unsigned(forvar2897) ?
                          (&forvar2919) : $unsigned(reg2994))) << (((reg2979 ?
                                  reg2777 : reg2817) ?
                              reg2926[(3'h6):(2'h3)] : reg2885[(3'h5):(1'h1)]) ?
                          $unsigned($unsigned((8'hb4))) : {reg2951[(3'h5):(2'h3)]}));
                      reg2950 <= reg2762[(1'h0):(1'h0)];
                      reg2951 <= reg2863[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg2948 <= {reg2967};
                    end
                  reg2952 <= reg2798[(2'h2):(2'h2)];
                end
              else
                begin
                  reg2944 <= $unsigned((^reg2858[(1'h0):(1'h0)]));
                  for (forvar2945 = (1'h0); (forvar2945 < (2'h3)); forvar2945 = (forvar2945 + (1'h1)))
                    begin
                      reg2946 <= reg2968;
                      reg2947 <= {$signed((~|$unsigned(reg2960)))};
                      reg2948 <= reg2756;
                      reg2949 <= forvar2871[(4'hb):(4'ha)];
                    end
                  for (forvar2950 = (1'h0); (forvar2950 < (1'h1)); forvar2950 = (forvar2950 + (1'h1)))
                    begin
                      reg2951 <= (~$signed($unsigned($signed(reg2832))));
                      reg2952 <= $signed((|$signed(reg2865[(4'hc):(4'hc)])));
                      reg2953 <= (reg2812[(2'h2):(1'h0)] ?
                          ($signed(wire2753) <= (^~$unsigned(forvar2993))) : (reg2950[(2'h2):(2'h2)] << $unsigned({forvar2797})));
                      reg2954 <= $unsigned(reg2981);
                    end
                  for (forvar2955 = (1'h0); (forvar2955 < (2'h3)); forvar2955 = (forvar2955 + (1'h1)))
                    begin
                      reg2956 <= reg2901[(3'h5):(2'h3)];
                      reg2957 <= $unsigned(({$signed(reg2860)} ?
                          (reg2907 ?
                              $signed(reg2921) : {reg2843}) : ($unsigned((8'ha5)) ?
                              (~|reg2799) : $unsigned(reg2780))));
                    end
                end
              for (forvar2958 = (1'h0); (forvar2958 < (1'h1)); forvar2958 = (forvar2958 + (1'h1)))
                begin
                  for (forvar2959 = (1'h0); (forvar2959 < (1'h1)); forvar2959 = (forvar2959 + (1'h1)))
                    begin
                      reg2960 <= forvar2993[(1'h1):(1'h1)];
                      reg2961 <= $signed(reg2937);
                      reg2962 <= $signed(($signed($signed(reg2997)) * reg2801));
                      reg2963 <= {(~{(reg2884 ? reg2952 : reg2807)})};
                    end
                end
              for (forvar2964 = (1'h0); (forvar2964 < (1'h1)); forvar2964 = (forvar2964 + (1'h1)))
                begin
                  reg2965 <= ((|(8'hb1)) ^ (~$unsigned($signed((8'hb1)))));
                  for (forvar2966 = (1'h0); (forvar2966 < (2'h3)); forvar2966 = (forvar2966 + (1'h1)))
                    begin
                      reg2967 <= reg2762[(1'h1):(1'h0)];
                      reg2968 <= $unsigned({({reg2977} ?
                              $signed(forvar2948) : forvar2945[(3'h4):(1'h0)])});
                      reg2969 <= (~&reg2958[(1'h0):(1'h0)]);
                      reg2970 <= forvar2953[(4'h8):(4'h8)];
                    end
                end
            end
          reg2971 <= forvar2969[(1'h0):(1'h0)];
        end
    end
  assign wire3002 = reg2868[(3'h6):(3'h4)];
  assign wire3003 = reg2790[(3'h5):(3'h4)];
  always
    @(posedge clk) begin
      if ($signed(reg2843))
        begin
          if (((&reg2804) ~^ (-reg2936[(2'h2):(2'h2)])))
            begin
              reg3004 <= (forvar2858 ?
                  $signed(reg2909[(1'h1):(1'h0)]) : ($signed({reg2870}) ?
                      (+$unsigned((8'hb3))) : (reg2922[(1'h0):(1'h0)] < $unsigned(forvar2920))));
              if ({$unsigned((-forvar2849[(2'h2):(2'h2)]))})
                begin
                  if ((^~$signed(reg2985[(4'hd):(3'h6)])))
                    begin
                      reg3005 <= reg2929;
                      reg3006 <= (wire3002 << $signed((&$unsigned(forvar2798))));
                    end
                  else
                    begin
                      reg3005 <= reg2905;
                      reg3006 <= $signed(($signed($signed(reg2799)) ?
                          forvar2943[(1'h0):(1'h0)] : reg2811[(4'h8):(3'h5)]));
                    end
                end
              else
                begin
                  for (forvar3005 = (1'h0); (forvar3005 < (2'h2)); forvar3005 = (forvar3005 + (1'h1)))
                    begin
                      reg3006 <= forvar2822[(2'h3):(2'h3)];
                      reg3007 <= $unsigned($unsigned((~$signed(reg2937))));
                      reg3008 <= $unsigned({reg2810[(4'h8):(3'h5)]});
                    end
                  for (forvar3009 = (1'h0); (forvar3009 < (2'h3)); forvar3009 = (forvar3009 + (1'h1)))
                    begin
                      reg3010 <= ((^~reg2867[(3'h4):(2'h3)]) ?
                          ((|(-reg2806)) != reg2997[(1'h0):(1'h0)]) : (forvar2950[(1'h0):(1'h0)] & (-(~^reg2955))));
                      reg3011 <= reg2827;
                    end
                  for (forvar3012 = (1'h0); (forvar3012 < (1'h0)); forvar3012 = (forvar3012 + (1'h1)))
                    begin
                      reg3013 <= (&((reg2787[(1'h0):(1'h0)] ?
                              ((8'haf) ? reg2982 : (8'hac)) : (reg2866 ?
                                  forvar2793 : forvar2764)) ?
                          (reg2869 ?
                              (reg2989 ?
                                  reg2961 : reg2944) : forvar2861) : $signed((8'hae))));
                      reg3014 <= ((reg2846[(2'h3):(2'h2)] != reg2823) ?
                          $signed(reg2814[(4'h8):(3'h4)]) : ((reg2945 ?
                                  (wire3002 >>> reg2923) : reg2864[(1'h0):(1'h0)]) ?
                              ((-reg2848) >>> $unsigned(reg2924)) : ((8'ha3) ?
                                  ((8'ha6) - (8'h9e)) : (reg2878 ?
                                      forvar2927 : (8'hb6)))));
                      reg3015 <= (~^$unsigned({(|reg2865)}));
                    end
                  for (forvar3016 = (1'h0); (forvar3016 < (2'h3)); forvar3016 = (forvar3016 + (1'h1)))
                    begin
                      reg3017 <= (!($unsigned(forvar2953) - reg2897));
                      reg3018 <= (^~$unsigned($signed((forvar2917 ?
                          reg2951 : forvar2799))));
                      reg3019 <= $unsigned((~|(forvar3012 && $signed(reg2955))));
                      reg3020 <= (reg2971[(1'h1):(1'h1)] != wire2753[(2'h2):(1'h0)]);
                    end
                end
              for (forvar3021 = (1'h0); (forvar3021 < (1'h1)); forvar3021 = (forvar3021 + (1'h1)))
                begin
                  reg3022 <= ((~(8'ha0)) ^ (-(reg2977 ?
                      $signed(wire2752) : {reg2965})));
                  reg3023 <= ($unsigned($signed(reg2967)) <<< (~|$signed(reg3013[(2'h3):(2'h3)])));
                  if ($unsigned(reg3007[(3'h5):(1'h0)]))
                    begin
                      reg3024 <= forvar2891;
                    end
                  else
                    begin
                      reg3024 <= (!reg2848[(3'h7):(2'h2)]);
                      reg3025 <= wire1762;
                      reg3026 <= forvar2862;
                      reg3027 <= reg3026;
                    end
                end
            end
          else
            begin
              for (forvar3004 = (1'h0); (forvar3004 < (2'h2)); forvar3004 = (forvar3004 + (1'h1)))
                begin
                  if ((+forvar2917[(2'h3):(1'h1)]))
                    begin
                      reg3005 <= (($unsigned((reg3018 ? reg2980 : wire1762)) ?
                              (reg2766[(4'h9):(3'h5)] ?
                                  $signed(reg2962) : $signed((8'hb0))) : (^(^~reg3007))) ?
                          $signed(reg2869) : ((+{wire2752}) | (~&(|reg3011))));
                      reg3006 <= ({(^~$signed(reg2983))} ?
                          $signed($signed((reg2756 && (8'hb7)))) : $unsigned($unsigned($unsigned(reg2870))));
                    end
                  else
                    begin
                      reg3005 <= {(reg2876[(2'h2):(2'h2)] ^ ((^~reg3024) ?
                              $signed(forvar2755) : $unsigned(reg2919)))};
                      reg3006 <= $unsigned(reg2913);
                    end
                  for (forvar3007 = (1'h0); (forvar3007 < (2'h3)); forvar3007 = (forvar3007 + (1'h1)))
                    begin
                      reg3008 <= $signed(forvar2950);
                    end
                  reg3009 <= ((~&(^(reg2914 ?
                      reg2812 : forvar2897))) == (reg3008 >>> forvar3012[(3'h7):(2'h3)]));
                end
              if ((reg2901[(4'hb):(3'h4)] > {reg3013}))
                begin
                  if (reg2960)
                    begin
                      reg3010 <= ($unsigned(($signed(forvar2948) <= (~&(8'h9d)))) ?
                          $unsigned((+(forvar3021 ?
                              reg2929 : (8'ha2)))) : (reg2804 == $signed(forvar2770)));
                      reg3011 <= reg2781;
                    end
                  else
                    begin
                      reg3010 <= {($signed($unsigned((8'hb6))) ^~ $signed((-reg2989)))};
                    end
                  reg3012 <= reg2962;
                  if (wire2753)
                    begin
                      reg3013 <= $unsigned(($signed($signed(forvar2774)) >>> forvar2899[(1'h0):(1'h0)]));
                      reg3014 <= $unsigned((reg3007 && reg2970[(3'h6):(3'h5)]));
                      reg3015 <= (|$unsigned($signed((+forvar2969))));
                      reg3016 <= $unsigned(forvar2866[(3'h4):(1'h1)]);
                    end
                  else
                    begin
                      reg3013 <= $unsigned(forvar2963);
                      reg3014 <= reg2862;
                      reg3015 <= $signed($signed(reg2902[(1'h1):(1'h1)]));
                      reg3016 <= $signed($unsigned(((wire1762 >> forvar2821) * (~^reg2947))));
                    end
                end
              else
                begin
                  for (forvar3010 = (1'h0); (forvar3010 < (2'h3)); forvar3010 = (forvar3010 + (1'h1)))
                    begin
                      reg3011 <= $signed(reg2998);
                      reg3012 <= $signed((&reg2977[(3'h4):(1'h0)]));
                      reg3013 <= forvar2844[(3'h5):(3'h5)];
                    end
                end
              for (forvar3017 = (1'h0); (forvar3017 < (2'h3)); forvar3017 = (forvar3017 + (1'h1)))
                begin
                  if ($signed(reg2795))
                    begin
                      reg3018 <= (-reg2915[(3'h5):(2'h2)]);
                      reg3019 <= (+((+forvar2878) + forvar2879[(2'h3):(2'h2)]));
                      reg3020 <= {forvar3005};
                    end
                  else
                    begin
                      reg3018 <= forvar2801;
                      reg3019 <= ((-(^(forvar3021 ?
                          reg2824 : reg2998))) >> $unsigned((~|$unsigned(forvar2963))));
                      reg3020 <= reg2841;
                      reg3021 <= $unsigned((~^(!(reg2762 == reg2773))));
                    end
                end
              for (forvar3022 = (1'h0); (forvar3022 < (2'h2)); forvar3022 = (forvar3022 + (1'h1)))
                begin
                  if ((8'ha4))
                    begin
                      reg3023 <= reg2835;
                      reg3024 <= $signed((8'h9f));
                      reg3025 <= $signed(((8'hb8) * reg2979));
                    end
                  else
                    begin
                      reg3023 <= $unsigned(($signed(reg2890[(4'h9):(2'h3)]) == (~{reg2928})));
                    end
                end
            end
          if ({(~&((forvar2866 ?
                  forvar2774 : reg2927) <= (reg2951 ~^ forvar2783)))})
            begin
              for (forvar3028 = (1'h0); (forvar3028 < (2'h3)); forvar3028 = (forvar3028 + (1'h1)))
                begin
                  for (forvar3029 = (1'h0); (forvar3029 < (1'h0)); forvar3029 = (forvar3029 + (1'h1)))
                    begin
                      reg3030 <= $signed(((8'haf) >= ((~^(8'h9f)) >= reg2779[(3'h5):(2'h3)])));
                      reg3031 <= (reg2786[(1'h0):(1'h0)] ?
                          (^reg2793[(3'h4):(2'h2)]) : (forvar2922 ?
                              wire2753 : ({reg2798} ?
                                  $signed(forvar2865) : (~reg2866))));
                    end
                  reg3032 <= $signed(reg2957);
                  if (((!({reg2973} ?
                      reg2936[(4'ha):(2'h2)] : reg2980[(4'hf):(4'hf)])) >>> reg2851[(2'h2):(2'h2)]))
                    begin
                      reg3033 <= $unsigned($unsigned({reg3031}));
                    end
                  else
                    begin
                      reg3033 <= (8'ha1);
                      reg3034 <= {forvar2872};
                      reg3035 <= (|((reg2898[(2'h3):(1'h1)] ?
                          $unsigned(reg2983) : reg2795) << reg2979[(4'ha):(4'h9)]));
                      reg3036 <= forvar2969;
                    end
                  if (forvar2865)
                    begin
                      reg3037 <= (8'ha8);
                      reg3038 <= $signed(reg3004[(1'h1):(1'h1)]);
                      reg3039 <= forvar2919[(4'ha):(4'ha)];
                    end
                  else
                    begin
                      reg3037 <= ((+reg2961) ?
                          reg2787 : reg2871[(1'h1):(1'h1)]);
                      reg3038 <= $signed({$unsigned((+forvar2860))});
                      reg3039 <= $unsigned((reg2799 ^~ reg2884));
                      reg3040 <= (~^forvar2944[(4'he):(4'hc)]);
                    end
                end
              for (forvar3041 = (1'h0); (forvar3041 < (2'h3)); forvar3041 = (forvar3041 + (1'h1)))
                begin
                  if ((&$signed(($unsigned(reg2932) ^ reg3015[(1'h0):(1'h0)]))))
                    begin
                      reg3042 <= forvar2969[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg3042 <= ((~|$signed((reg2805 || (8'hb7)))) * $signed((reg2780[(1'h1):(1'h1)] > (~^reg2994))));
                    end
                end
            end
          else
            begin
              for (forvar3028 = (1'h0); (forvar3028 < (1'h0)); forvar3028 = (forvar3028 + (1'h1)))
                begin
                  if (reg2799)
                    begin
                      reg3029 <= $unsigned(($signed((+wire1763)) ?
                          (-(-forvar2781)) : $unsigned((8'hb8))));
                      reg3030 <= reg2782[(4'hf):(3'h4)];
                      reg3031 <= $signed(((8'hb3) ?
                          {(reg2850 ? reg2896 : forvar3009)} : reg2888));
                    end
                  else
                    begin
                      reg3029 <= (((~(+reg2945)) ?
                          reg2900 : $signed({reg3035})) >>> (|($unsigned((8'hb1)) ?
                          $unsigned(wire1763) : $unsigned(reg2803))));
                      reg3030 <= $unsigned($signed(reg2861[(1'h0):(1'h0)]));
                    end
                end
              reg3032 <= (&(^(~|((8'ha4) ? forvar2860 : reg2836))));
            end
        end
      else
        begin
          for (forvar3004 = (1'h0); (forvar3004 < (2'h2)); forvar3004 = (forvar3004 + (1'h1)))
            begin
              for (forvar3005 = (1'h0); (forvar3005 < (1'h0)); forvar3005 = (forvar3005 + (1'h1)))
                begin
                  for (forvar3006 = (1'h0); (forvar3006 < (2'h2)); forvar3006 = (forvar3006 + (1'h1)))
                    begin
                      reg3007 <= reg2976[(2'h2):(1'h1)];
                      reg3008 <= {$signed(reg2858)};
                      reg3009 <= reg3031[(2'h3):(1'h0)];
                      reg3010 <= ($signed($signed((reg2857 >>> forvar2955))) ?
                          (!(~|(reg2980 >= reg3018))) : reg2963);
                    end
                  for (forvar3011 = (1'h0); (forvar3011 < (1'h1)); forvar3011 = (forvar3011 + (1'h1)))
                    begin
                      reg3012 <= (reg3034 > ((reg2956[(4'hd):(4'ha)] - {forvar3004}) ?
                          (&(reg2938 ? wire2749 : reg2854)) : {{forvar2829}}));
                      reg3013 <= ((&reg3032) ?
                          reg2903[(1'h0):(1'h0)] : $unsigned(reg2798));
                    end
                  if ($signed((|$signed((^reg2916)))))
                    begin
                      reg3014 <= $signed((reg2893[(2'h2):(1'h0)] || $signed(reg2850[(1'h0):(1'h0)])));
                      reg3015 <= (reg2983 ?
                          reg2979[(3'h6):(1'h0)] : $signed(reg2935[(2'h3):(1'h1)]));
                      reg3016 <= (|reg2885);
                    end
                  else
                    begin
                      reg3014 <= (reg2949[(4'ha):(2'h3)] & {$unsigned((forvar2922 >>> reg2838))});
                      reg3015 <= reg2875;
                      reg3016 <= {$unsigned(({forvar3011} ?
                              (|reg2781) : $signed((8'hb9))))};
                    end
                  if ({wire1761})
                    begin
                      reg3017 <= (^~$signed({(reg2945 ? reg2950 : reg2868)}));
                      reg3018 <= $signed((^reg3033));
                      reg3019 <= {(reg2758 ?
                              reg2951[(1'h1):(1'h0)] : (~|reg3015[(2'h2):(2'h2)]))};
                      reg3020 <= ({reg2885[(1'h1):(1'h0)]} < (~wire1760));
                    end
                  else
                    begin
                      reg3017 <= (~|(+reg3027));
                      reg3018 <= ({reg2810} * reg2933[(2'h3):(2'h2)]);
                      reg3019 <= ({{(forvar2948 * reg2915)}} ?
                          reg2791[(4'h8):(3'h4)] : (-($signed(reg2998) ?
                              $unsigned(forvar3029) : forvar3028)));
                    end
                end
              for (forvar3021 = (1'h0); (forvar3021 < (1'h0)); forvar3021 = (forvar3021 + (1'h1)))
                begin
                  for (forvar3022 = (1'h0); (forvar3022 < (1'h0)); forvar3022 = (forvar3022 + (1'h1)))
                    begin
                      reg3023 <= (-((^~{forvar2822}) ? reg3024 : forvar2778));
                      reg3024 <= (8'hb8);
                      reg3025 <= ((($unsigned(reg3000) & reg2945) ?
                              $signed(forvar2947[(3'h6):(3'h4)]) : (reg2778 ?
                                  ((8'haa) ? (8'ha0) : (8'ha0)) : (+reg2923))) ?
                          (!($signed((8'ha0)) + (reg2876 ?
                              reg2823 : reg2878))) : {(~&{(8'hab)})});
                    end
                  reg3026 <= (($signed($signed((8'h9f))) ?
                      ((~&reg2973) && $signed(reg3040)) : ((~&(8'ha6)) || $signed(reg2807))) << $signed((((8'hb4) | reg2757) ?
                      $unsigned(reg2884) : (-forvar2879))));
                end
              for (forvar3027 = (1'h0); (forvar3027 < (1'h1)); forvar3027 = (forvar3027 + (1'h1)))
                begin
                  for (forvar3028 = (1'h0); (forvar3028 < (2'h2)); forvar3028 = (forvar3028 + (1'h1)))
                    begin
                      reg3029 <= $signed((((~|reg2934) ^ $signed(reg2971)) && ((^reg2852) ?
                          (~^reg2970) : {reg2811})));
                      reg3030 <= reg2989[(1'h0):(1'h0)];
                      reg3031 <= $unsigned((~|{(reg2840 ?
                              reg2910 : forvar3012)}));
                      reg3032 <= ($signed(reg2878) ?
                          forvar2764 : $unsigned($signed((&(8'ha7)))));
                    end
                  for (forvar3033 = (1'h0); (forvar3033 < (2'h2)); forvar3033 = (forvar3033 + (1'h1)))
                    begin
                      reg3034 <= (~$signed($unsigned($unsigned(reg2864))));
                      reg3035 <= $signed($signed((&reg2872[(2'h2):(2'h2)])));
                      reg3036 <= forvar2919[(4'hb):(4'h8)];
                    end
                end
            end
        end
      for (forvar3043 = (1'h0); (forvar3043 < (2'h3)); forvar3043 = (forvar3043 + (1'h1)))
        begin
          reg3044 <= (^reg2941[(1'h0):(1'h0)]);
          for (forvar3045 = (1'h0); (forvar3045 < (2'h2)); forvar3045 = (forvar3045 + (1'h1)))
            begin
              reg3046 <= $unsigned($unsigned(((reg2768 ? reg2794 : reg2865) ?
                  (8'hb0) : reg2793[(3'h4):(2'h2)])));
              if (forvar3028[(1'h0):(1'h0)])
                begin
                  for (forvar3047 = (1'h0); (forvar3047 < (2'h3)); forvar3047 = (forvar3047 + (1'h1)))
                    begin
                      reg3048 <= $unsigned((((~&(8'haa)) ?
                          $signed(reg2813) : reg2967) >= ((forvar2978 ?
                          reg2934 : reg2854) <<< $unsigned(reg2922))));
                      reg3049 <= $signed(forvar2873[(2'h3):(2'h3)]);
                      reg3050 <= forvar3005[(2'h2):(1'h1)];
                      reg3051 <= (~reg2901);
                    end
                  for (forvar3052 = (1'h0); (forvar3052 < (2'h2)); forvar3052 = (forvar3052 + (1'h1)))
                    begin
                      reg3053 <= {(($unsigned(reg3050) - (-reg3012)) ?
                              ($unsigned(reg2869) ?
                                  forvar2866[(3'h5):(3'h4)] : forvar2927) : (^(wire3003 << (8'ha7))))};
                      reg3054 <= $signed((reg2953[(3'h7):(3'h4)] ?
                          $unsigned((~&reg2879)) : $signed(reg3030[(3'h7):(3'h4)])));
                      reg3055 <= {reg2852};
                    end
                  for (forvar3056 = (1'h0); (forvar3056 < (1'h0)); forvar3056 = (forvar3056 + (1'h1)))
                    begin
                      reg3057 <= $signed(({reg2893} ?
                          $signed((reg3020 & reg3021)) : reg2918[(2'h2):(1'h0)]));
                      reg3058 <= $signed(((forvar3041 ~^ reg2983) != {reg2914}));
                      reg3059 <= (~^(~&$signed($unsigned(forvar2878))));
                    end
                end
              else
                begin
                  reg3047 <= reg2916;
                  if (forvar3017[(3'h5):(2'h2)])
                    begin
                      reg3048 <= ((~$unsigned(wire2753[(4'h8):(2'h3)])) * {$unsigned($signed(forvar3005))});
                      reg3049 <= reg2893[(2'h3):(2'h2)];
                      reg3050 <= (($unsigned($unsigned((8'hb8))) ?
                          $signed($unsigned(reg2992)) : reg3012) & $unsigned((reg2761 ?
                          (reg2856 != (8'hb9)) : ((8'hb4) ?
                              forvar2950 : reg3048))));
                    end
                  else
                    begin
                      reg3048 <= $unsigned((($unsigned(forvar3012) || $signed(forvar2902)) & reg2997[(3'h5):(1'h0)]));
                    end
                  reg3051 <= $signed($unsigned((reg2801 && (reg2998 ?
                      (8'hb0) : reg2885))));
                  if (($signed(reg2949[(4'hb):(2'h3)]) <= $signed(reg2923)))
                    begin
                      reg3052 <= (^~(reg2972[(1'h1):(1'h0)] != {(-reg2801)}));
                    end
                  else
                    begin
                      reg3052 <= (~^$signed({reg2939}));
                      reg3053 <= ($unsigned((|$signed(reg2932))) ?
                          reg2825 : $unsigned($signed(forvar2849[(4'h8):(2'h3)])));
                    end
                end
              for (forvar3060 = (1'h0); (forvar3060 < (2'h3)); forvar3060 = (forvar3060 + (1'h1)))
                begin
                  for (forvar3061 = (1'h0); (forvar3061 < (1'h1)); forvar3061 = (forvar3061 + (1'h1)))
                    begin
                      reg3062 <= reg3000;
                      reg3063 <= (reg2896 ?
                          (8'hab) : (|(forvar2958[(2'h2):(1'h0)] > $unsigned((8'hb4)))));
                      reg3064 <= (&$signed({$unsigned((8'ha4))}));
                      reg3065 <= {$unsigned(($signed(reg2794) ?
                              reg2889 : (8'haa)))};
                    end
                  for (forvar3066 = (1'h0); (forvar3066 < (1'h1)); forvar3066 = (forvar3066 + (1'h1)))
                    begin
                      reg3067 <= ((~&$signed((reg2984 ? reg2995 : (8'ha6)))) ?
                          forvar2963 : reg2945);
                      reg3068 <= forvar3027;
                      reg3069 <= ($unsigned(($unsigned(reg2941) ?
                          (!reg3012) : {forvar3009})) - $signed(forvar3007[(1'h0):(1'h0)]));
                    end
                  for (forvar3070 = (1'h0); (forvar3070 < (2'h2)); forvar3070 = (forvar3070 + (1'h1)))
                    begin
                      reg3071 <= $signed((~reg3042[(1'h0):(1'h0)]));
                      reg3072 <= ($unsigned({forvar2862[(4'h8):(3'h5)]}) ?
                          {(~^(reg2782 ?
                                  forvar3045 : forvar2861))} : $unsigned(reg2762));
                      reg3073 <= (+($unsigned(wire2753) ?
                          reg3000[(2'h2):(2'h2)] : ($signed(reg2858) + reg2907[(1'h0):(1'h0)])));
                      reg3074 <= {({forvar2925} ?
                              ($signed(forvar2777) || forvar2891) : (&reg2924))};
                    end
                  for (forvar3075 = (1'h0); (forvar3075 < (1'h0)); forvar3075 = (forvar3075 + (1'h1)))
                    begin
                      reg3076 <= (^~reg2958[(2'h3):(2'h2)]);
                      reg3077 <= reg2907[(1'h1):(1'h0)];
                      reg3078 <= (forvar3005 ^~ $signed($unsigned((reg2879 + reg3073))));
                      reg3079 <= (forvar2897 >> reg2795[(3'h6):(1'h0)]);
                    end
                end
              if ((8'hb8))
                begin
                  reg3080 <= forvar2917;
                  for (forvar3081 = (1'h0); (forvar3081 < (1'h0)); forvar3081 = (forvar3081 + (1'h1)))
                    begin
                      reg3082 <= (+(+$unsigned(forvar2978)));
                      reg3083 <= ($signed(reg2760[(4'h9):(4'h8)]) > (forvar2755 != ($unsigned(reg2814) ?
                          (forvar2826 && reg2941) : $signed(forvar2891))));
                      reg3084 <= $unsigned($signed(forvar2808));
                      reg3085 <= (!forvar2899[(3'h6):(1'h0)]);
                    end
                end
              else
                begin
                  if ($unsigned($signed((~^(reg3009 != reg2873)))))
                    begin
                      reg3080 <= $signed(forvar2964);
                    end
                  else
                    begin
                      reg3080 <= (~|{reg2759[(3'h4):(1'h1)]});
                      reg3081 <= $signed(reg2783);
                      reg3082 <= ($unsigned({((8'hae) ? reg2758 : reg3013)}) ?
                          (^~(~(8'hb6))) : $unsigned(reg2806));
                      reg3083 <= (((forvar3066 || (&reg2789)) & $signed((~^(8'hac)))) ?
                          reg3047[(4'hb):(1'h0)] : (((reg3085 ?
                              reg3053 : reg3054) != $signed((8'h9f))) != {(reg3044 ?
                                  reg2995 : (8'haf))}));
                    end
                  for (forvar3084 = (1'h0); (forvar3084 < (2'h3)); forvar3084 = (forvar3084 + (1'h1)))
                    begin
                      reg3085 <= reg2773[(2'h3):(1'h0)];
                      reg3086 <= (~$unsigned((((8'had) <<< forvar2855) << (^~forvar3021))));
                    end
                end
            end
          for (forvar3087 = (1'h0); (forvar3087 < (1'h0)); forvar3087 = (forvar3087 + (1'h1)))
            begin
              reg3088 <= reg2857[(2'h3):(1'h0)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg3089 <= {reg2943[(2'h3):(1'h1)]};
      if ((($signed(forvar3060) != (8'hb2)) & (-((~&reg2927) ?
          (!(8'hac)) : ((8'hb9) ^~ reg3009)))))
        begin
          for (forvar3090 = (1'h0); (forvar3090 < (2'h3)); forvar3090 = (forvar3090 + (1'h1)))
            begin
              for (forvar3091 = (1'h0); (forvar3091 < (2'h2)); forvar3091 = (forvar3091 + (1'h1)))
                begin
                  if ($unsigned($unsigned(forvar2892)))
                    begin
                      reg3092 <= reg2915;
                      reg3093 <= (+(~^(forvar2850 ~^ (reg2782 & reg2776))));
                      reg3094 <= {(($signed((8'hb2)) < $unsigned(forvar3029)) - $unsigned($unsigned(reg2983)))};
                      reg3095 <= $unsigned($signed($unsigned((wire1762 ^ reg2763))));
                    end
                  else
                    begin
                      reg3092 <= $unsigned(reg3073[(2'h2):(1'h0)]);
                      reg3093 <= (|forvar2955);
                      reg3094 <= {$unsigned((&(8'h9c)))};
                      reg3095 <= $signed(reg2755);
                    end
                  reg3096 <= $unsigned((^reg3077[(3'h5):(2'h2)]));
                  if ((8'ha4))
                    begin
                      reg3097 <= forvar3010;
                      reg3098 <= $signed($signed(reg2980));
                      reg3099 <= $signed(($unsigned(forvar2922) ?
                          {{forvar3005}} : ((+reg2832) | (reg3012 ?
                              reg2876 : reg3088))));
                      reg3100 <= (8'hb8);
                    end
                  else
                    begin
                      reg3097 <= $unsigned($signed((reg2992[(4'ha):(3'h4)] ?
                          reg3071[(4'ha):(3'h5)] : reg2957)));
                      reg3098 <= reg2864;
                      reg3099 <= reg3089[(3'h4):(3'h4)];
                    end
                end
            end
          for (forvar3101 = (1'h0); (forvar3101 < (2'h3)); forvar3101 = (forvar3101 + (1'h1)))
            begin
              for (forvar3102 = (1'h0); (forvar3102 < (1'h1)); forvar3102 = (forvar3102 + (1'h1)))
                begin
                  for (forvar3103 = (1'h0); (forvar3103 < (2'h3)); forvar3103 = (forvar3103 + (1'h1)))
                    begin
                      reg3104 <= reg2887;
                      reg3105 <= {(+((forvar2842 && forvar2990) > (~reg3046)))};
                      reg3106 <= wire2752[(3'h7):(3'h6)];
                    end
                  if (((8'ha6) >> $signed(reg3100[(3'h7):(1'h1)])))
                    begin
                      reg3107 <= {$unsigned(((reg2786 < reg3098) ?
                              $signed((8'ha4)) : $signed(reg3055)))};
                      reg3108 <= $unsigned((forvar2774[(3'h7):(3'h7)] ^ wire1760));
                      reg3109 <= {{((reg3083 ? reg3044 : forvar2809) ?
                                  forvar2777[(3'h4):(2'h2)] : (+forvar2920))}};
                      reg3110 <= forvar2945[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3107 <= ((reg2943[(1'h1):(1'h1)] ?
                              $signed((&reg3085)) : reg3036[(3'h5):(3'h4)]) ?
                          $signed($signed($unsigned(reg2854))) : (~{$signed(reg2888)}));
                      reg3108 <= (((+(reg2878 ~^ reg2956)) ?
                              (reg2812[(2'h2):(2'h2)] ?
                                  reg3073 : (~&reg2945)) : ((forvar2829 < forvar2948) ?
                                  $unsigned((8'ha2)) : forvar3090)) ?
                          reg3099 : {$unsigned($signed(reg2943))});
                      reg3109 <= (forvar2770[(2'h3):(2'h2)] ?
                          reg3085[(3'h7):(3'h6)] : $signed(forvar2912[(3'h7):(2'h2)]));
                      reg3110 <= reg3014[(1'h1):(1'h1)];
                    end
                  if (((~|(~|(reg2980 <<< reg3050))) << $unsigned((~|$signed(reg2834)))))
                    begin
                      reg3111 <= (($unsigned(forvar3027) << (~|(&reg2927))) >> forvar2959);
                    end
                  else
                    begin
                      reg3111 <= (^reg2919);
                    end
                  if ($signed($unsigned($signed((+forvar3066)))))
                    begin
                      reg3112 <= reg2786[(3'h7):(3'h5)];
                      reg3113 <= $signed(forvar2876);
                    end
                  else
                    begin
                      reg3112 <= reg2882;
                    end
                end
              for (forvar3114 = (1'h0); (forvar3114 < (2'h2)); forvar3114 = (forvar3114 + (1'h1)))
                begin
                  reg3115 <= forvar3114[(4'ha):(4'h8)];
                  if (forvar2775[(3'h4):(3'h4)])
                    begin
                      reg3116 <= reg2811;
                    end
                  else
                    begin
                      reg3116 <= (((-(&reg2979)) ~^ $unsigned(forvar3009)) ~^ (|reg2813));
                      reg3117 <= reg3107[(2'h3):(2'h2)];
                      reg3118 <= (~|(forvar3017[(1'h0):(1'h0)] ?
                          {reg2977[(4'h8):(3'h7)]} : reg3109));
                      reg3119 <= ((($unsigned((8'hac)) >= forvar3075[(1'h0):(1'h0)]) ?
                              $signed({reg2772}) : reg2975[(1'h1):(1'h0)]) ?
                          (-$signed($unsigned(reg2782))) : (^~reg2988));
                    end
                  for (forvar3120 = (1'h0); (forvar3120 < (1'h0)); forvar3120 = (forvar3120 + (1'h1)))
                    begin
                      reg3121 <= forvar2958[(2'h2):(2'h2)];
                    end
                  for (forvar3122 = (1'h0); (forvar3122 < (2'h3)); forvar3122 = (forvar3122 + (1'h1)))
                    begin
                      reg3123 <= {(^(^(&forvar2826)))};
                      reg3124 <= $signed({$signed(reg3083)});
                    end
                end
            end
          for (forvar3125 = (1'h0); (forvar3125 < (2'h3)); forvar3125 = (forvar3125 + (1'h1)))
            begin
              if ($unsigned((8'hb7)))
                begin
                  if ($signed((8'ha7)))
                    begin
                      reg3126 <= reg2931[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg3126 <= ($signed(reg2825[(3'h4):(2'h2)]) ?
                          $unsigned(($unsigned(forvar2953) ?
                              $unsigned(reg2890) : forvar2919[(2'h3):(2'h2)])) : reg3076);
                      reg3127 <= {($unsigned({reg3095}) >= ((forvar2797 & reg2966) * reg3044[(4'ha):(3'h4)]))};
                      reg3128 <= {(($signed(forvar2908) ^~ forvar3056[(2'h2):(1'h0)]) != (forvar3103 + wire2749))};
                      reg3129 <= reg3073;
                    end
                  for (forvar3130 = (1'h0); (forvar3130 < (1'h0)); forvar3130 = (forvar3130 + (1'h1)))
                    begin
                      reg3131 <= $signed($signed(((reg2835 != reg2964) ?
                          (reg2967 ?
                              reg2969 : forvar2775) : forvar3070[(1'h0):(1'h0)])));
                      reg3132 <= ((+((reg3082 ? reg3123 : (8'haa)) >> (reg3115 ?
                          reg2777 : reg2991))) && reg2880);
                      reg3133 <= ($signed(reg2986) ?
                          $signed(($signed(reg2937) >> (reg2977 ?
                              wire3002 : forvar2917))) : $signed(((reg3015 - reg2978) < {reg2830})));
                      reg3134 <= reg2812[(3'h4):(1'h0)];
                    end
                  for (forvar3135 = (1'h0); (forvar3135 < (1'h1)); forvar3135 = (forvar3135 + (1'h1)))
                    begin
                      reg3136 <= ($signed($unsigned($unsigned(reg3059))) < $unsigned(forvar2959));
                      reg3137 <= $unsigned(reg3007[(3'h4):(2'h2)]);
                    end
                end
              else
                begin
                  if ($unsigned($signed(reg2989[(2'h2):(2'h2)])))
                    begin
                      reg3126 <= reg2894;
                      reg3127 <= {({$unsigned(forvar3061)} ?
                              (~|reg3039[(4'h9):(3'h6)]) : forvar3135[(3'h6):(3'h4)])};
                    end
                  else
                    begin
                      reg3126 <= $unsigned(($unsigned((reg2915 <<< reg2968)) ?
                          (~^$signed(reg2773)) : $signed((!reg3058))));
                      reg3127 <= {$signed($signed($unsigned((8'hae))))};
                      reg3128 <= $unsigned($unsigned((~^reg3113[(1'h1):(1'h1)])));
                      reg3129 <= (|reg2923[(2'h2):(1'h1)]);
                    end
                  if ((~^forvar2958))
                    begin
                      reg3130 <= ((((+reg2832) != {reg2983}) >> {{(8'h9f)}}) ?
                          reg2783 : $signed({{(8'ha5)}}));
                    end
                  else
                    begin
                      reg3130 <= ((forvar3006 ?
                              ((^forvar2978) ?
                                  (reg3121 ?
                                      reg3016 : reg2896) : (reg3064 ^~ wire2753)) : ({reg2947} ?
                                  (reg2786 ~^ reg2762) : {reg2799})) ?
                          {($unsigned((8'haa)) >= reg2994)} : $signed(forvar3103));
                    end
                  reg3131 <= forvar2777[(2'h3):(1'h0)];
                end
              if (forvar2799[(3'h4):(3'h4)])
                begin
                  if ((-reg2772))
                    begin
                      reg3138 <= $signed(forvar2855);
                    end
                  else
                    begin
                      reg3138 <= {(&{$signed(reg3032)})};
                      reg3139 <= (&forvar2868[(3'h4):(1'h1)]);
                      reg3140 <= forvar2947;
                    end
                  for (forvar3141 = (1'h0); (forvar3141 < (1'h0)); forvar3141 = (forvar3141 + (1'h1)))
                    begin
                      reg3142 <= ($unsigned($signed(reg2883)) ^~ (reg2794[(2'h3):(2'h2)] << reg2842[(2'h2):(2'h2)]));
                    end
                  for (forvar3143 = (1'h0); (forvar3143 < (2'h3)); forvar3143 = (forvar3143 + (1'h1)))
                    begin
                      reg3144 <= $signed($unsigned(($unsigned(reg2992) ?
                          reg3011 : reg3068[(1'h0):(1'h0)])));
                      reg3145 <= ($signed(reg2988[(3'h7):(1'h0)]) ^~ (&((~^(8'hb6)) ^ (forvar2917 >= forvar2755))));
                      reg3146 <= (reg3012 == $unsigned(reg2921[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  reg3138 <= ($unsigned({$signed(reg3138)}) ?
                      $unsigned($unsigned($unsigned(reg2898))) : reg2833);
                  for (forvar3139 = (1'h0); (forvar3139 < (2'h2)); forvar3139 = (forvar3139 + (1'h1)))
                    begin
                      reg3140 <= reg3117[(4'h8):(3'h7)];
                      reg3141 <= (forvar2947[(1'h0):(1'h0)] ?
                          (-(!forvar2925[(3'h7):(2'h3)])) : forvar2803[(4'hb):(4'h9)]);
                    end
                  for (forvar3142 = (1'h0); (forvar3142 < (2'h2)); forvar3142 = (forvar3142 + (1'h1)))
                    begin
                      reg3143 <= reg3082;
                      reg3144 <= $unsigned({{$unsigned(reg2837)}});
                      reg3145 <= reg2788;
                      reg3146 <= reg2994;
                    end
                  if (reg3025[(1'h0):(1'h0)])
                    begin
                      reg3147 <= {($unsigned((|reg2840)) ?
                              ($signed(reg2783) <= reg2874) : $unsigned($unsigned((8'hb8))))};
                      reg3148 <= (!(-$unsigned((reg2840 ?
                          forvar2821 : forvar2902))));
                      reg3149 <= {forvar2925};
                      reg3150 <= {reg3094};
                    end
                  else
                    begin
                      reg3147 <= $unsigned(((~&reg3136[(3'h6):(1'h0)]) + $signed(reg3040[(2'h2):(1'h1)])));
                      reg3148 <= reg3095[(3'h5):(1'h0)];
                      reg3149 <= reg2806;
                    end
                end
              for (forvar3151 = (1'h0); (forvar3151 < (2'h2)); forvar3151 = (forvar3151 + (1'h1)))
                begin
                  for (forvar3152 = (1'h0); (forvar3152 < (2'h3)); forvar3152 = (forvar3152 + (1'h1)))
                    begin
                      reg3153 <= ($signed({(^reg3031)}) & $signed(((reg3068 <= reg2981) ?
                          reg2831 : $unsigned((8'hae)))));
                      reg3154 <= reg3093;
                      reg3155 <= $signed(reg2918);
                      reg3156 <= (reg3077[(4'hd):(2'h2)] ^ ($unsigned(forvar3091) ~^ $signed((reg3081 ?
                          wire2753 : reg3037))));
                    end
                  for (forvar3157 = (1'h0); (forvar3157 < (2'h3)); forvar3157 = (forvar3157 + (1'h1)))
                    begin
                      reg3158 <= reg2953;
                      reg3159 <= ($unsigned($signed(reg2905[(1'h1):(1'h0)])) && (~$unsigned($signed(reg3097))));
                      reg3160 <= (forvar2872[(4'hb):(3'h6)] - (forvar2891 >> (reg2913[(1'h0):(1'h0)] ?
                          (^~reg2893) : (reg2827 ? reg2964 : reg2835))));
                    end
                  reg3161 <= $signed(((|(~|forvar2822)) || ($signed(reg2815) == (^reg3034))));
                end
              reg3162 <= (8'haa);
            end
        end
      else
        begin
          for (forvar3090 = (1'h0); (forvar3090 < (2'h2)); forvar3090 = (forvar3090 + (1'h1)))
            begin
              if ($signed(reg2835))
                begin
                  if (reg2790)
                    begin
                      reg3091 <= $signed({$unsigned((~|reg2773))});
                    end
                  else
                    begin
                      reg3091 <= ({{forvar2849}} * (8'hb8));
                      reg3092 <= (((reg3109 <= ((8'ha3) << reg3018)) && $signed($signed(reg2940))) ?
                          (reg3062 ?
                              $signed({forvar2947}) : ($signed((8'ha9)) ?
                                  $signed((8'hb2)) : ((8'hb5) + forvar2990))) : (~^($signed((8'ha9)) ?
                              {reg2945} : $unsigned(reg2881))));
                      reg3093 <= $unsigned(forvar3142);
                      reg3094 <= reg2972;
                    end
                  for (forvar3095 = (1'h0); (forvar3095 < (2'h2)); forvar3095 = (forvar3095 + (1'h1)))
                    begin
                      reg3096 <= (-((~&forvar2964) < (8'hb7)));
                      reg3097 <= $signed((~&($signed(reg2888) ?
                          (~reg3069) : $unsigned(reg2957))));
                    end
                  if (((((forvar2912 ? reg3155 : reg2868) ?
                          $signed(reg3093) : (+(8'ha0))) ?
                      ((reg2762 << reg2884) & reg2980) : (~$unsigned((8'haa)))) > ($unsigned(reg2801) & ({(8'hb2)} | {reg2998}))))
                    begin
                      reg3098 <= {(^~(reg2796 ?
                              $signed(reg3130) : $signed(reg3076)))};
                      reg3099 <= (forvar2871[(4'hc):(3'h7)] ?
                          $unsigned(reg2914) : reg2942);
                      reg3100 <= reg3162[(2'h3):(1'h1)];
                      reg3101 <= (($signed(reg3116[(1'h1):(1'h1)]) << reg3115[(3'h5):(2'h2)]) <<< (~|reg3032));
                    end
                  else
                    begin
                      reg3098 <= {$unsigned((forvar3005[(1'h0):(1'h0)] ?
                              (reg2783 >= forvar3033) : (reg3001 ^~ reg2834)))};
                      reg3099 <= (~|$signed({reg2831[(3'h7):(3'h5)]}));
                      reg3100 <= ($signed(forvar3056[(1'h0):(1'h0)]) ~^ ((8'hb9) ^ forvar2793[(3'h6):(2'h3)]));
                      reg3101 <= (reg3067[(1'h1):(1'h0)] >>> (^~((&wire3003) ^~ reg2943)));
                    end
                end
              else
                begin
                  for (forvar3091 = (1'h0); (forvar3091 < (1'h0)); forvar3091 = (forvar3091 + (1'h1)))
                    begin
                      reg3092 <= ($signed(reg2867) + (({reg2836} << (~^forvar3029)) <= reg2858[(1'h0):(1'h0)]));
                    end
                end
              for (forvar3102 = (1'h0); (forvar3102 < (2'h3)); forvar3102 = (forvar3102 + (1'h1)))
                begin
                  if (($unsigned(reg2967) ?
                      $signed(($signed(forvar2953) ?
                          (forvar2955 ? reg2782 : reg3097) : (reg2777 ?
                              reg3131 : wire1761))) : ((reg2904[(4'hb):(3'h7)] * (8'h9e)) ?
                          (reg2944[(3'h4):(2'h2)] <= reg3150) : reg2902)))
                    begin
                      reg3103 <= (+forvar2781[(3'h7):(3'h7)]);
                      reg3104 <= {((wire2753 ?
                              $signed((8'ha6)) : $signed(forvar2919)) - $unsigned($unsigned(reg2877)))};
                    end
                  else
                    begin
                      reg3103 <= (((~|reg3054) ?
                              ({reg2980} | reg2839) : forvar3012) ?
                          {$unsigned(forvar3070)} : (reg2863 >= reg2784));
                      reg3104 <= ($signed($signed((reg3020 ?
                              forvar3009 : reg2868))) ?
                          (((^reg3031) >> $signed(forvar2963)) ?
                              (~^$signed(reg3080)) : $unsigned((reg3078 - (8'ha7)))) : ($unsigned(((8'hb4) || reg3129)) ?
                              reg2800[(3'h4):(1'h0)] : {(~reg2876)}));
                      reg3105 <= (|reg3104);
                      reg3106 <= (8'ha6);
                    end
                end
            end
          reg3107 <= (+(((-forvar2922) ? reg2995[(1'h0):(1'h0)] : (|reg3006)) ?
              ((reg3155 ^ reg2955) > $signed(reg3008)) : ($signed(reg2775) ?
                  $unsigned(reg2890) : $unsigned(forvar2978))));
          for (forvar3108 = (1'h0); (forvar3108 < (2'h3)); forvar3108 = (forvar3108 + (1'h1)))
            begin
              for (forvar3109 = (1'h0); (forvar3109 < (1'h1)); forvar3109 = (forvar3109 + (1'h1)))
                begin
                  for (forvar3110 = (1'h0); (forvar3110 < (2'h2)); forvar3110 = (forvar3110 + (1'h1)))
                    begin
                      reg3111 <= reg3073[(1'h1):(1'h1)];
                    end
                end
              for (forvar3112 = (1'h0); (forvar3112 < (2'h3)); forvar3112 = (forvar3112 + (1'h1)))
                begin
                  reg3113 <= reg2804[(2'h2):(2'h2)];
                  for (forvar3114 = (1'h0); (forvar3114 < (2'h3)); forvar3114 = (forvar3114 + (1'h1)))
                    begin
                      reg3115 <= (forvar3075[(1'h0):(1'h0)] ?
                          $unsigned((~&reg3149[(3'h7):(1'h1)])) : $unsigned((forvar3011 ?
                              (reg2995 ?
                                  forvar2838 : reg3159) : $signed((8'ha7)))));
                      reg3116 <= reg3156[(4'h9):(3'h6)];
                      reg3117 <= reg2810;
                      reg3118 <= (forvar2793[(4'h8):(3'h6)] ?
                          $unsigned($signed($unsigned(reg3148))) : (^~reg2857));
                    end
                end
              reg3119 <= reg3026;
              reg3120 <= ({($unsigned(reg2819) ?
                          (~^forvar3101) : (reg2896 << (8'h9d)))} ?
                  {($signed(forvar2872) >> ((8'ha2) ?
                          reg2812 : reg3158))} : ((8'hb0) >>> ({reg2937} >= reg3096)));
            end
          reg3121 <= $unsigned(reg2769);
        end
      for (forvar3163 = (1'h0); (forvar3163 < (2'h2)); forvar3163 = (forvar3163 + (1'h1)))
        begin
          for (forvar3164 = (1'h0); (forvar3164 < (1'h1)); forvar3164 = (forvar3164 + (1'h1)))
            begin
              for (forvar3165 = (1'h0); (forvar3165 < (2'h2)); forvar3165 = (forvar3165 + (1'h1)))
                begin
                  if (reg3013)
                    begin
                      reg3166 <= $signed((reg2868[(2'h2):(1'h0)] > (forvar2978[(2'h3):(1'h1)] - wire1760)));
                    end
                  else
                    begin
                      reg3166 <= (reg3098 + $unsigned(reg2938));
                    end
                end
              reg3167 <= (|(((reg2850 != forvar2868) <= (|reg2916)) <<< (~(reg3022 ?
                  reg2965 : reg3132))));
              for (forvar3168 = (1'h0); (forvar3168 < (1'h1)); forvar3168 = (forvar3168 + (1'h1)))
                begin
                  if ($signed(wire2751[(3'h7):(2'h2)]))
                    begin
                      reg3169 <= $signed($signed($unsigned(reg3084)));
                      reg3170 <= ($unsigned($unsigned($unsigned(forvar3043))) ^ ($unsigned(reg3091) ?
                          reg3017[(4'hd):(4'hd)] : forvar3016));
                      reg3171 <= (reg3004 ?
                          reg3023[(2'h2):(2'h2)] : $unsigned((^~(^reg2914))));
                      reg3172 <= $signed(($unsigned((~forvar2844)) ?
                          reg3099 : reg2953));
                    end
                  else
                    begin
                      reg3169 <= ((reg3172[(1'h1):(1'h1)] >> (reg3121[(4'hb):(4'ha)] | reg3059[(2'h2):(1'h0)])) ?
                          $unsigned($unsigned(reg2812[(2'h3):(2'h2)])) : {(+(~reg2956))});
                    end
                  if ($signed(((|(forvar2902 * forvar2908)) << (^{reg3073}))))
                    begin
                      reg3173 <= {(^(reg2839[(1'h0):(1'h0)] == (~&forvar3006)))};
                      reg3174 <= $signed((($unsigned(reg2964) ?
                              forvar2838 : $unsigned(forvar2968)) ?
                          ({reg2780} ?
                              wire1762 : (reg3024 ^ reg2784)) : $unsigned($unsigned(reg2757))));
                    end
                  else
                    begin
                      reg3173 <= ({(^~(|(8'hb1)))} > {reg2807});
                      reg3174 <= reg3111[(4'hd):(4'h8)];
                      reg3175 <= reg3172;
                      reg3176 <= reg2782;
                    end
                end
              if (((forvar2886[(2'h2):(1'h0)] * reg3072[(2'h2):(1'h0)]) & ($signed($signed(reg3158)) ?
                  (reg2869[(3'h7):(3'h7)] != (reg2938 ^ forvar3090)) : (forvar3109[(3'h5):(2'h3)] ?
                      (8'ha3) : (reg2798 ? (8'ha2) : (8'had))))))
                begin
                  for (forvar3177 = (1'h0); (forvar3177 < (1'h1)); forvar3177 = (forvar3177 + (1'h1)))
                    begin
                      reg3178 <= $unsigned($unsigned((reg3042[(1'h1):(1'h1)] || (-forvar2797))));
                      reg3179 <= forvar3029[(3'h5):(1'h1)];
                      reg3180 <= $unsigned($signed((~&(^reg2820))));
                    end
                end
              else
                begin
                  if ({$unsigned(reg3005)})
                    begin
                      reg3177 <= $signed($unsigned(reg2960[(2'h3):(2'h3)]));
                      reg3178 <= (($unsigned((forvar3016 == reg2982)) << (-$unsigned((8'hb0)))) <= (&forvar3163));
                    end
                  else
                    begin
                      reg3177 <= ((8'ha6) ?
                          ($signed((reg2804 ? reg2885 : (8'ha7))) ?
                              ($unsigned(forvar2925) ~^ (-reg2761)) : (-(forvar2803 && reg2992))) : (^~{$unsigned(forvar2876)}));
                      reg3178 <= $unsigned(reg3054[(1'h1):(1'h1)]);
                    end
                end
            end
        end
      reg3181 <= $signed((8'hb7));
    end
  assign wire3182 = $signed((((+forvar2783) ?
                        $signed((8'hb1)) : $unsigned(reg2762)) | reg3129[(4'h9):(4'h9)]));
  always
    @(posedge clk) begin
      for (forvar3183 = (1'h0); (forvar3183 < (1'h1)); forvar3183 = (forvar3183 + (1'h1)))
        begin
          for (forvar3184 = (1'h0); (forvar3184 < (2'h2)); forvar3184 = (forvar3184 + (1'h1)))
            begin
              reg3185 <= {(((8'ha1) <<< (~&(8'h9f))) || reg3176)};
            end
          for (forvar3186 = (1'h0); (forvar3186 < (2'h3)); forvar3186 = (forvar3186 + (1'h1)))
            begin
              for (forvar3187 = (1'h0); (forvar3187 < (1'h1)); forvar3187 = (forvar3187 + (1'h1)))
                begin
                  if (reg2784[(3'h4):(1'h1)])
                    begin
                      reg3188 <= (|reg2801);
                    end
                  else
                    begin
                      reg3188 <= ((!reg3073) >>> forvar2908[(4'hc):(3'h6)]);
                      reg3189 <= ({$unsigned(((8'hb1) ?
                              (8'hba) : reg2758))} + {reg3080});
                    end
                end
              if (reg3088[(4'h8):(4'h8)])
                begin
                  if ((forvar2912[(1'h1):(1'h0)] ^~ $signed($unsigned(reg2919))))
                    begin
                      reg3190 <= $unsigned((($unsigned(reg2873) ?
                          reg2958 : (reg2796 ?
                              wire1762 : reg2866)) >= reg3141));
                    end
                  else
                    begin
                      reg3190 <= (~&(^(8'hb0)));
                      reg3191 <= forvar2781[(4'hf):(1'h1)];
                      reg3192 <= reg3140;
                      reg3193 <= {{$unsigned(forvar3168[(1'h0):(1'h0)])}};
                    end
                  for (forvar3194 = (1'h0); (forvar3194 < (1'h1)); forvar3194 = (forvar3194 + (1'h1)))
                    begin
                      reg3195 <= reg2940;
                      reg3196 <= ($signed(($unsigned(reg2811) ?
                              reg2883[(1'h1):(1'h0)] : {reg2973})) ?
                          (!{$unsigned((8'ha8))}) : ({(reg2771 ?
                                  reg3032 : reg3108)} && (reg3008[(2'h3):(1'h0)] ?
                              $signed(reg3147) : (forvar2917 ?
                                  (8'had) : (8'ha1)))));
                      reg3197 <= $unsigned(($signed(((8'hb8) ?
                              (8'hb1) : (8'hb0))) ?
                          (reg2959[(2'h3):(2'h3)] ?
                              (forvar3165 >> reg3190) : (forvar3143 < forvar3102)) : ({forvar2803} ?
                              ((8'had) | (8'hab)) : forvar2790[(1'h1):(1'h1)])));
                      reg3198 <= (^~forvar3005);
                    end
                  reg3199 <= ($unsigned((forvar2970 ? (-reg3096) : reg3148)) ?
                      (($signed(reg2905) ? (!reg2885) : wire1762) ?
                          (8'ha6) : (!$unsigned(reg2948))) : $signed(reg2814[(3'h6):(3'h6)]));
                end
              else
                begin
                  reg3190 <= reg2920[(3'h7):(2'h3)];
                end
            end
          if (forvar3165[(3'h5):(3'h5)])
            begin
              if (reg2895[(1'h0):(1'h0)])
                begin
                  for (forvar3200 = (1'h0); (forvar3200 < (2'h2)); forvar3200 = (forvar3200 + (1'h1)))
                    begin
                      reg3201 <= $unsigned($unsigned((reg3195 ^~ (forvar2808 > reg3105))));
                      reg3202 <= ((~|($signed((8'hb8)) ?
                          (reg2996 ?
                              reg3166 : forvar3081) : $unsigned(forvar2886))) && $unsigned($unsigned($unsigned(reg2956))));
                    end
                  for (forvar3203 = (1'h0); (forvar3203 < (1'h1)); forvar3203 = (forvar3203 + (1'h1)))
                    begin
                      reg3204 <= reg2876[(2'h2):(1'h0)];
                    end
                  if ({($signed((reg2789 ? (8'hba) : forvar3045)) ?
                          (reg3195[(2'h2):(1'h1)] ?
                              {forvar2963} : (forvar2866 ?
                                  reg3039 : wire1762)) : forvar3186[(3'h4):(2'h3)])})
                    begin
                      reg3205 <= {(!($unsigned(reg2911) ?
                              reg2941[(3'h4):(1'h0)] : reg2788[(2'h2):(1'h1)]))};
                    end
                  else
                    begin
                      reg3205 <= forvar2902[(1'h1):(1'h0)];
                      reg3206 <= $unsigned((~((^forvar2764) ?
                          forvar2844 : forvar3090)));
                      reg3207 <= $unsigned($unsigned($unsigned((reg3116 ?
                          forvar2969 : reg2874))));
                    end
                end
              else
                begin
                  for (forvar3200 = (1'h0); (forvar3200 < (1'h1)); forvar3200 = (forvar3200 + (1'h1)))
                    begin
                      reg3201 <= (~(8'hb1));
                      reg3202 <= (^forvar3070[(1'h0):(1'h0)]);
                      reg3203 <= {(($unsigned(reg3174) + reg2851) ~^ reg3172[(1'h1):(1'h1)])};
                      reg3204 <= (reg2907[(1'h1):(1'h0)] ?
                          $unsigned(((forvar2764 >> reg2801) >= ((8'ha4) ?
                              reg3189 : reg2864))) : $unsigned((^(reg3189 ?
                              forvar2862 : reg3039))));
                    end
                  if (reg2980)
                    begin
                      reg3205 <= forvar2897;
                      reg3206 <= (reg2813 ?
                          ($signed(forvar2927) ?
                              $unsigned((+forvar2990)) : $signed(reg3118[(1'h0):(1'h0)])) : reg3190[(3'h6):(3'h4)]);
                      reg3207 <= ($signed(((reg2915 ? reg3202 : forvar3165) ?
                          reg2773[(1'h0):(1'h0)] : forvar3087)) > reg3204);
                      reg3208 <= $signed(($signed((8'hb4)) ?
                          ((reg3018 ?
                              forvar2899 : (8'hb2)) >> (reg2930 == reg3000)) : (8'ha6)));
                    end
                  else
                    begin
                      reg3205 <= (reg3144[(1'h0):(1'h0)] ?
                          (reg2824[(3'h4):(2'h3)] ?
                              ($unsigned(reg2966) >> (~reg2948)) : $unsigned($signed(reg2872))) : $unsigned((8'hb8)));
                    end
                  reg3209 <= $signed({$unsigned($unsigned(reg2810))});
                end
              for (forvar3210 = (1'h0); (forvar3210 < (1'h1)); forvar3210 = (forvar3210 + (1'h1)))
                begin
                  if (forvar2912[(2'h3):(1'h0)])
                    begin
                      reg3211 <= $unsigned($unsigned((reg3197 ?
                          wire1762 : $signed(reg3191))));
                      reg3212 <= $unsigned(($signed($unsigned(reg2934)) ?
                          reg2956[(4'h8):(1'h1)] : (8'hb8)));
                    end
                  else
                    begin
                      reg3211 <= $signed($unsigned(reg2914));
                    end
                  for (forvar3213 = (1'h0); (forvar3213 < (1'h0)); forvar3213 = (forvar3213 + (1'h1)))
                    begin
                      reg3214 <= ($signed((!$signed(reg3019))) | ((~&(reg2991 ?
                          reg2937 : forvar2970)) <= {reg3162[(4'h8):(3'h7)]}));
                    end
                end
              if ($unsigned($unsigned($unsigned((reg3017 ?
                  reg2997 : (8'hb9))))))
                begin
                  for (forvar3215 = (1'h0); (forvar3215 < (2'h3)); forvar3215 = (forvar3215 + (1'h1)))
                    begin
                      reg3216 <= (8'ha2);
                    end
                  for (forvar3217 = (1'h0); (forvar3217 < (2'h2)); forvar3217 = (forvar3217 + (1'h1)))
                    begin
                      reg3218 <= $signed(reg2901[(4'hb):(4'hb)]);
                    end
                end
              else
                begin
                  reg3215 <= (((reg2976[(1'h1):(1'h1)] ^~ reg2976[(3'h7):(1'h1)]) ?
                          $signed(((8'ha8) >>> reg2828)) : (~reg2877)) ?
                      reg2843[(3'h5):(1'h1)] : ($signed(reg2762[(2'h3):(2'h3)]) <= (reg3019[(4'ha):(3'h5)] ?
                          reg2801 : (reg2848 ? forvar3109 : reg2883))));
                  if ($signed(reg3156))
                    begin
                      reg3216 <= reg2854;
                      reg3217 <= $signed((($unsigned((8'ha6)) | $signed(forvar3033)) | (|(reg3112 != reg2932))));
                      reg3218 <= (~|$signed({{reg3180}}));
                    end
                  else
                    begin
                      reg3216 <= (~(&(reg3018[(2'h2):(2'h2)] < (forvar2966 ?
                          forvar3047 : reg2933))));
                      reg3217 <= (reg3042[(2'h3):(2'h3)] != (~^{(reg2884 > reg2784)}));
                    end
                  reg3219 <= {(forvar2860[(3'h4):(2'h3)] - (!reg2854))};
                  for (forvar3220 = (1'h0); (forvar3220 < (1'h1)); forvar3220 = (forvar3220 + (1'h1)))
                    begin
                      reg3221 <= (&((reg2893 ?
                              (^reg2853) : (reg2801 ? (8'hb1) : reg2982)) ?
                          (reg3131 ^ (-(8'hb7))) : (~^reg2864)));
                      reg3222 <= ((({forvar3184} ?
                                  $unsigned((8'ha1)) : (reg2919 ?
                                      reg2931 : reg3018)) ?
                              reg3119 : $unsigned($unsigned(reg3012))) ?
                          $unsigned(reg2852) : (8'h9f));
                    end
                end
            end
          else
            begin
              if ((reg3079[(3'h6):(1'h0)] || reg2937[(3'h7):(2'h2)]))
                begin
                  if ($signed($unsigned((~(reg3209 ? reg3053 : forvar2891)))))
                    begin
                      reg3200 <= ($signed(reg3099[(3'h5):(3'h5)]) <= forvar2774[(3'h5):(3'h4)]);
                    end
                  else
                    begin
                      reg3200 <= $unsigned(forvar2764[(3'h5):(1'h1)]);
                      reg3201 <= (~reg3016[(1'h0):(1'h0)]);
                      reg3202 <= $unsigned(reg3169);
                    end
                  reg3203 <= $unsigned(($signed({reg3216}) ?
                      reg3014 : (reg2832[(1'h1):(1'h1)] ~^ (reg3193 >> forvar3157))));
                end
              else
                begin
                  for (forvar3200 = (1'h0); (forvar3200 < (1'h0)); forvar3200 = (forvar3200 + (1'h1)))
                    begin
                      reg3201 <= {($unsigned(forvar2950) ?
                              ($signed(forvar3016) | reg2935[(3'h7):(1'h1)]) : forvar3139[(3'h5):(2'h2)])};
                      reg3202 <= $unsigned($unsigned({((8'hb6) ^~ (8'hb9))}));
                      reg3203 <= $unsigned(reg2902[(2'h2):(2'h2)]);
                      reg3204 <= $signed((reg3024 ?
                          (&$signed(reg3064)) : reg2763));
                    end
                  for (forvar3205 = (1'h0); (forvar3205 < (2'h3)); forvar3205 = (forvar3205 + (1'h1)))
                    begin
                      reg3206 <= (!reg2848);
                    end
                  if ((forvar2871[(2'h2):(1'h0)] <<< $signed(forvar2764)))
                    begin
                      reg3207 <= $unsigned(reg2771);
                      reg3208 <= {((forvar2970 & (&reg2800)) ?
                              {(reg3104 ?
                                      (8'hba) : reg2807)} : reg3113[(2'h2):(1'h1)])};
                      reg3209 <= reg2915[(4'h8):(3'h6)];
                    end
                  else
                    begin
                      reg3207 <= forvar2783;
                      reg3208 <= $signed(((~(forvar2860 ? reg3022 : reg2895)) ?
                          ((reg2799 ?
                              reg2978 : reg3156) - $unsigned((8'hac))) : reg3180));
                      reg3209 <= (((~|(reg2988 ? reg3059 : reg3192)) ?
                              ($signed((8'ha5)) ?
                                  (reg3039 ?
                                      (8'h9c) : reg2981) : {forvar3213}) : ($signed((8'hb3)) && reg3197[(1'h0):(1'h0)])) ?
                          (reg2806 ?
                              {(reg2932 - reg3065)} : $signed({reg2782})) : $signed(forvar2963[(3'h4):(2'h3)]));
                    end
                end
              for (forvar3210 = (1'h0); (forvar3210 < (1'h1)); forvar3210 = (forvar3210 + (1'h1)))
                begin
                  reg3211 <= ($signed($signed((reg2804 ?
                      reg2936 : reg2977))) && reg2942);
                  reg3212 <= forvar3183[(3'h4):(3'h4)];
                  for (forvar3213 = (1'h0); (forvar3213 < (2'h2)); forvar3213 = (forvar3213 + (1'h1)))
                    begin
                      reg3214 <= $unsigned(forvar2774);
                      reg3215 <= reg3046;
                    end
                end
              reg3216 <= ((!$unsigned($signed(forvar2886))) ^ (reg3109[(2'h2):(1'h0)] >>> $unsigned((reg2790 >>> forvar3045))));
            end
          if ((($signed((8'hb0)) != $unsigned($unsigned(forvar2983))) ?
              forvar2873[(2'h2):(2'h2)] : ((~^(reg3094 ?
                  reg3024 : forvar2860)) ^~ (-forvar3164[(3'h7):(1'h0)]))))
            begin
              for (forvar3223 = (1'h0); (forvar3223 < (1'h1)); forvar3223 = (forvar3223 + (1'h1)))
                begin
                  for (forvar3224 = (1'h0); (forvar3224 < (2'h3)); forvar3224 = (forvar3224 + (1'h1)))
                    begin
                      reg3225 <= reg2801[(4'ha):(4'h9)];
                      reg3226 <= reg3081[(3'h7):(3'h6)];
                      reg3227 <= $signed((8'hb6));
                    end
                  for (forvar3228 = (1'h0); (forvar3228 < (1'h1)); forvar3228 = (forvar3228 + (1'h1)))
                    begin
                      reg3229 <= reg2995[(3'h4):(2'h2)];
                      reg3230 <= (reg2866[(1'h0):(1'h0)] <= (8'hb8));
                      reg3231 <= (($signed((+(8'ha4))) ^ $unsigned((forvar2826 ?
                          reg2785 : (8'ha9)))) >= (8'hb5));
                    end
                  for (forvar3232 = (1'h0); (forvar3232 < (2'h3)); forvar3232 = (forvar3232 + (1'h1)))
                    begin
                      reg3233 <= ((reg3058 ?
                              ((reg3093 ?
                                  reg3048 : forvar3183) << wire2753[(1'h0):(1'h0)]) : $signed(((8'haa) ?
                                  forvar3130 : reg2757))) ?
                          reg3205 : $unsigned($unsigned($unsigned(reg2901))));
                      reg3234 <= ((~((forvar2866 ?
                          forvar2945 : reg2972) + reg2769[(4'hb):(1'h0)])) <<< $unsigned(reg3049[(2'h2):(1'h0)]));
                      reg3235 <= ($unsigned((8'ha8)) ?
                          (reg3189 ?
                              ($signed(reg2812) ?
                                  (forvar3164 ?
                                      reg2804 : (8'ha4)) : reg2778) : (^~reg2920[(2'h2):(2'h2)])) : forvar3056);
                      reg3236 <= ((-reg2980) <= reg3136[(1'h1):(1'h1)]);
                    end
                  for (forvar3237 = (1'h0); (forvar3237 < (1'h0)); forvar3237 = (forvar3237 + (1'h1)))
                    begin
                      reg3238 <= (~&reg2868);
                      reg3239 <= (^forvar3022[(2'h3):(1'h0)]);
                    end
                end
              for (forvar3240 = (1'h0); (forvar3240 < (2'h2)); forvar3240 = (forvar3240 + (1'h1)))
                begin
                  reg3241 <= {(^(reg3216[(1'h1):(1'h0)] + reg3174))};
                end
              if (reg2966)
                begin
                  for (forvar3242 = (1'h0); (forvar3242 < (2'h2)); forvar3242 = (forvar3242 + (1'h1)))
                    begin
                      reg3243 <= forvar3091;
                      reg3244 <= (~(&$unsigned($signed((8'ha9)))));
                      reg3245 <= {$unsigned(({reg3226} ?
                              {reg3005} : (forvar2959 ^~ forvar2855)))};
                      reg3246 <= forvar2974;
                    end
                  for (forvar3247 = (1'h0); (forvar3247 < (2'h3)); forvar3247 = (forvar3247 + (1'h1)))
                    begin
                      reg3248 <= reg2971[(1'h0):(1'h0)];
                    end
                  if (reg2916[(3'h6):(3'h4)])
                    begin
                      reg3249 <= $unsigned($unsigned(((reg3233 ?
                          (8'h9e) : reg3091) && $signed(reg3202))));
                      reg3250 <= {reg3158};
                      reg3251 <= reg2820[(3'h4):(2'h3)];
                      reg3252 <= reg3144;
                    end
                  else
                    begin
                      reg3249 <= $unsigned((($unsigned(forvar2876) >> $signed(reg2944)) ?
                          (-$signed(reg2768)) : reg3016[(2'h2):(1'h1)]));
                    end
                end
              else
                begin
                  for (forvar3242 = (1'h0); (forvar3242 < (2'h3)); forvar3242 = (forvar3242 + (1'h1)))
                    begin
                      reg3243 <= $signed($unsigned({{forvar2803}}));
                      reg3244 <= $unsigned($signed(reg3037[(3'h4):(1'h0)]));
                      reg3245 <= {(reg2931 + $signed(((8'h9e) ?
                              forvar3043 : forvar2950)))};
                    end
                end
            end
          else
            begin
              for (forvar3223 = (1'h0); (forvar3223 < (2'h2)); forvar3223 = (forvar3223 + (1'h1)))
                begin
                  if (((!{$unsigned(reg2802)}) * ((8'hb1) > $unsigned(reg2997))))
                    begin
                      reg3224 <= ((($signed(reg2851) - forvar2908) ?
                              ((reg2970 ^ reg2847) >= reg3016) : reg2854) ?
                          (^~(reg3058 + (forvar3052 >>> reg2918))) : (~(8'haa)));
                    end
                  else
                    begin
                      reg3224 <= reg3103;
                      reg3225 <= reg2818[(3'h5):(1'h0)];
                      reg3226 <= ((({forvar2855} ? forvar2801 : {(8'hb8)}) ?
                              ((reg3108 ?
                                  reg2904 : (8'hb5)) < (-(8'hb8))) : (((8'ha1) <<< forvar3184) || (-reg3044))) ?
                          ((8'ha9) + ({(8'h9f)} ?
                              (8'hb8) : (!reg2878))) : (~^((reg2793 << forvar3004) ?
                              $unsigned(reg2869) : (!(8'hb5)))));
                      reg3227 <= (($unsigned((reg3154 >> reg3000)) ?
                          (reg2889 ?
                              $unsigned(reg2816) : (forvar2892 * reg3058)) : reg2817) ^ reg3035[(3'h7):(3'h5)]);
                    end
                  if ((reg3010 ?
                      $signed($signed((reg2940 ^ reg2945))) : ({(reg3136 ?
                                  forvar3011 : (8'hba))} ?
                          (-reg2785[(1'h0):(1'h0)]) : {(8'hb8)})))
                    begin
                      reg3228 <= reg2986[(4'hd):(4'hb)];
                    end
                  else
                    begin
                      reg3228 <= $unsigned($signed({(-reg2884)}));
                      reg3229 <= reg3067[(4'hb):(4'hb)];
                      reg3230 <= (({reg3173} ?
                          ($signed(forvar2878) >> forvar2969) : forvar2927) << ($unsigned((~|forvar2899)) || (^~(~&forvar2865))));
                    end
                  for (forvar3231 = (1'h0); (forvar3231 < (2'h2)); forvar3231 = (forvar3231 + (1'h1)))
                    begin
                      reg3232 <= (reg2906[(3'h4):(1'h0)] ^ (reg3017[(3'h7):(2'h3)] & $signed((^(8'hb0)))));
                      reg3233 <= {forvar2945[(2'h2):(2'h2)]};
                      reg3234 <= $signed(reg2959[(1'h1):(1'h1)]);
                      reg3235 <= $signed((|$unsigned({(8'hb0)})));
                    end
                  if (reg3069)
                    begin
                      reg3236 <= forvar2781;
                    end
                  else
                    begin
                      reg3236 <= forvar3027;
                      reg3237 <= ((forvar2927[(3'h4):(1'h1)] ?
                          $signed(reg2903[(1'h0):(1'h0)]) : $signed((8'ha1))) > $signed($signed((&reg3040))));
                      reg3238 <= (((~|$signed(reg3232)) >>> (~|reg3113)) ?
                          (reg3080 ?
                              {(forvar2878 != reg3049)} : reg3216[(2'h3):(2'h3)]) : $unsigned((reg2788 ?
                              (reg3211 ?
                                  reg2917 : reg3169) : forvar2983[(4'h9):(1'h0)])));
                      reg3239 <= (reg3188 >> {($signed(reg3196) ^ $unsigned(reg3176))});
                    end
                end
            end
        end
      for (forvar3253 = (1'h0); (forvar3253 < (2'h3)); forvar3253 = (forvar3253 + (1'h1)))
        begin
          for (forvar3254 = (1'h0); (forvar3254 < (2'h2)); forvar3254 = (forvar3254 + (1'h1)))
            begin
              for (forvar3255 = (1'h0); (forvar3255 < (1'h0)); forvar3255 = (forvar3255 + (1'h1)))
                begin
                  reg3256 <= {reg2812};
                  if (($signed((reg3219 ?
                          (forvar2860 ?
                              forvar2897 : (8'had)) : (reg2935 < reg3031))) ?
                      $unsigned((reg3089[(2'h2):(2'h2)] ?
                          $unsigned(reg2923) : (reg2779 ~^ reg2801))) : $signed(reg3202[(3'h6):(2'h3)])))
                    begin
                      reg3257 <= {$unsigned(reg3174[(3'h6):(2'h2)])};
                      reg3258 <= $unsigned($unsigned(reg2949[(3'h6):(1'h1)]));
                      reg3259 <= $signed(($signed((reg2924 <= reg3229)) & reg3166));
                    end
                  else
                    begin
                      reg3257 <= {reg2868[(3'h6):(2'h2)]};
                      reg3258 <= $signed((+($unsigned(reg3077) ?
                          $unsigned(forvar2945) : ((8'had) | reg3173))));
                      reg3259 <= ((!reg3010) == reg2874);
                    end
                  for (forvar3260 = (1'h0); (forvar3260 < (2'h2)); forvar3260 = (forvar3260 + (1'h1)))
                    begin
                      reg3261 <= ($signed(((reg3154 >>> (8'ha1)) || reg3038)) | {((forvar2943 << forvar2803) ~^ (reg2798 ^~ forvar3135))});
                      reg3262 <= $signed((reg3238 > ((reg2786 + reg3128) ?
                          (forvar2754 ?
                              reg2950 : reg2765) : (forvar2862 >> reg2957))));
                      reg3263 <= {forvar3060[(4'h8):(4'h8)]};
                      reg3264 <= {(($unsigned(forvar2947) & {reg3256}) ?
                              $signed($signed(reg2971)) : {(reg3162 ?
                                      reg3104 : reg3058)})};
                    end
                end
              for (forvar3265 = (1'h0); (forvar3265 < (2'h3)); forvar3265 = (forvar3265 + (1'h1)))
                begin
                  for (forvar3266 = (1'h0); (forvar3266 < (2'h2)); forvar3266 = (forvar3266 + (1'h1)))
                    begin
                      reg3267 <= (reg3133[(3'h7):(1'h1)] ^ ($unsigned($unsigned(reg2957)) << reg3177[(3'h5):(2'h2)]));
                      reg3268 <= reg2816[(1'h0):(1'h0)];
                      reg3269 <= (~|reg2959);
                      reg3270 <= forvar3157;
                    end
                  for (forvar3271 = (1'h0); (forvar3271 < (1'h1)); forvar3271 = (forvar3271 + (1'h1)))
                    begin
                      reg3272 <= $unsigned(reg3166);
                      reg3273 <= $unsigned($unsigned($signed(((8'had) ~^ reg2830))));
                    end
                end
            end
          if (reg2790[(2'h2):(1'h0)])
            begin
              for (forvar3274 = (1'h0); (forvar3274 < (1'h0)); forvar3274 = (forvar3274 + (1'h1)))
                begin
                  for (forvar3275 = (1'h0); (forvar3275 < (1'h0)); forvar3275 = (forvar3275 + (1'h1)))
                    begin
                      reg3276 <= $signed((((~&reg3078) ?
                              (^~reg2924) : reg2781) ?
                          $unsigned((reg2864 ?
                              forvar2925 : (8'ha2))) : (reg2962[(4'hc):(3'h5)] ?
                              (forvar3114 ?
                                  reg3154 : reg2900) : $unsigned(reg3259))));
                      reg3277 <= reg2949;
                      reg3278 <= reg3149[(4'h8):(1'h1)];
                      reg3279 <= $unsigned($signed(($unsigned(reg3267) >>> reg2789)));
                    end
                  for (forvar3280 = (1'h0); (forvar3280 < (1'h0)); forvar3280 = (forvar3280 + (1'h1)))
                    begin
                      reg3281 <= (((&$unsigned((8'hba))) ?
                              reg2898[(4'h8):(3'h5)] : $unsigned((reg3098 + reg2991))) ?
                          $unsigned($unsigned({(8'haf)})) : $unsigned(((^(8'hb5)) + (reg3105 ?
                              reg3086 : (8'ha2)))));
                      reg3282 <= (~|{$signed((|reg3085))});
                      reg3283 <= ($signed($unsigned(reg3011[(1'h0):(1'h0)])) >= wire3002);
                    end
                end
              for (forvar3284 = (1'h0); (forvar3284 < (2'h2)); forvar3284 = (forvar3284 + (1'h1)))
                begin
                  reg3285 <= ((|(^~(~|(8'ha6)))) && (~&$unsigned(forvar2793)));
                  reg3286 <= $unsigned($signed($unsigned($signed(reg2885))));
                end
            end
          else
            begin
              reg3274 <= $unsigned($unsigned({((8'hac) - reg2794)}));
              for (forvar3275 = (1'h0); (forvar3275 < (2'h3)); forvar3275 = (forvar3275 + (1'h1)))
                begin
                  if ($signed($signed(forvar2944)))
                    begin
                      reg3276 <= {(-$signed($signed(reg2991)))};
                    end
                  else
                    begin
                      reg3276 <= (($unsigned($unsigned(reg2866)) < forvar2826) >= $unsigned($signed($signed(reg3154))));
                      reg3277 <= {(8'hb6)};
                      reg3278 <= forvar2990[(1'h1):(1'h1)];
                    end
                  if (reg3062)
                    begin
                      reg3279 <= ($signed(reg3126) ?
                          {($unsigned(forvar3011) ?
                                  (reg3243 << forvar3274) : $unsigned(reg2819))} : ((((8'hb2) != reg3160) < $signed(reg2782)) << $unsigned((reg3170 ~^ reg3097))));
                      reg3280 <= ($unsigned(($unsigned(reg2888) ^~ reg3055)) ?
                          $signed(forvar2829) : $unsigned(reg3077[(1'h1):(1'h0)]));
                      reg3281 <= (reg2789[(4'hc):(4'hc)] ?
                          (~$signed(forvar3152[(3'h7):(1'h0)])) : (~$signed($signed(reg2784))));
                      reg3282 <= reg2765;
                    end
                  else
                    begin
                      reg3279 <= $signed((-($unsigned(reg3067) ?
                          (~&reg2897) : (|forvar3017))));
                      reg3280 <= $signed({reg2915[(1'h0):(1'h0)]});
                      reg3281 <= (8'hae);
                    end
                  for (forvar3283 = (1'h0); (forvar3283 < (1'h0)); forvar3283 = (forvar3283 + (1'h1)))
                    begin
                      reg3284 <= (~^$unsigned($unsigned(reg3283)));
                    end
                end
              for (forvar3285 = (1'h0); (forvar3285 < (2'h2)); forvar3285 = (forvar3285 + (1'h1)))
                begin
                  if (reg3204[(4'h9):(3'h7)])
                    begin
                      reg3286 <= ((|$signed((wire3003 ?
                          reg2933 : reg3124))) && reg3068);
                      reg3287 <= (reg3100[(3'h4):(2'h3)] ^~ $unsigned(reg2851[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg3286 <= (forvar3255[(2'h3):(1'h1)] && (8'ha0));
                    end
                  for (forvar3288 = (1'h0); (forvar3288 < (2'h3)); forvar3288 = (forvar3288 + (1'h1)))
                    begin
                      reg3289 <= (~&((forvar2953 ?
                              $signed(forvar3151) : {forvar3187}) ?
                          (8'ha0) : (+$signed(reg3238))));
                      reg3290 <= $unsigned($signed((&$unsigned(reg2939))));
                    end
                end
              reg3291 <= (|reg2958[(1'h1):(1'h0)]);
            end
          for (forvar3292 = (1'h0); (forvar3292 < (2'h2)); forvar3292 = (forvar3292 + (1'h1)))
            begin
              for (forvar3293 = (1'h0); (forvar3293 < (2'h3)); forvar3293 = (forvar3293 + (1'h1)))
                begin
                  if ($unsigned($unsigned(forvar2783[(3'h6):(3'h4)])))
                    begin
                      reg3294 <= (8'ha8);
                    end
                  else
                    begin
                      reg3294 <= ((-$signed($unsigned(wire3003))) ?
                          (8'hac) : reg3113[(1'h1):(1'h1)]);
                      reg3295 <= $signed(reg3082);
                    end
                end
              for (forvar3296 = (1'h0); (forvar3296 < (1'h0)); forvar3296 = (forvar3296 + (1'h1)))
                begin
                  for (forvar3297 = (1'h0); (forvar3297 < (1'h0)); forvar3297 = (forvar3297 + (1'h1)))
                    begin
                      reg3298 <= forvar3027[(4'ha):(4'ha)];
                      reg3299 <= (($signed((^reg3034)) ?
                              reg3243[(1'h1):(1'h1)] : forvar3220) ?
                          (8'hb9) : reg2868);
                      reg3300 <= $signed(reg3193);
                    end
                  if ($signed({$signed($unsigned((8'hb7)))}))
                    begin
                      reg3301 <= ((|((forvar2947 == (8'hb5)) ^ $signed(forvar3081))) << reg3008);
                    end
                  else
                    begin
                      reg3301 <= (forvar3168 ?
                          forvar2922[(3'h6):(1'h0)] : ((!{forvar3007}) ?
                              reg2804 : reg3001));
                      reg3302 <= $signed(($unsigned($unsigned(reg3171)) ?
                          {(reg3193 ^ reg3250)} : reg2840));
                    end
                  for (forvar3303 = (1'h0); (forvar3303 < (2'h3)); forvar3303 = (forvar3303 + (1'h1)))
                    begin
                      reg3304 <= forvar3043;
                      reg3305 <= reg3304;
                      reg3306 <= forvar3070[(3'h4):(3'h4)];
                      reg3307 <= (!(^((~&reg3051) * reg2915)));
                    end
                  for (forvar3308 = (1'h0); (forvar3308 < (1'h1)); forvar3308 = (forvar3308 + (1'h1)))
                    begin
                      reg3309 <= {reg3283};
                      reg3310 <= {reg3117};
                    end
                end
              for (forvar3311 = (1'h0); (forvar3311 < (2'h3)); forvar3311 = (forvar3311 + (1'h1)))
                begin
                  for (forvar3312 = (1'h0); (forvar3312 < (2'h2)); forvar3312 = (forvar3312 + (1'h1)))
                    begin
                      reg3313 <= (^~reg2935[(3'h4):(3'h4)]);
                      reg3314 <= reg3232;
                      reg3315 <= reg3029;
                      reg3316 <= ($signed($signed(reg2790[(2'h3):(1'h0)])) & reg3147);
                    end
                  if ((8'hba))
                    begin
                      reg3317 <= reg3133;
                      reg3318 <= ($signed(reg3044[(1'h1):(1'h0)]) ?
                          $signed($signed({reg2837})) : forvar2868[(3'h6):(2'h3)]);
                      reg3319 <= $signed((-$unsigned($signed((8'h9c)))));
                      reg3320 <= reg3280[(4'hb):(3'h6)];
                    end
                  else
                    begin
                      reg3317 <= (~&(&$signed(reg3103[(4'hc):(3'h6)])));
                    end
                  for (forvar3321 = (1'h0); (forvar3321 < (2'h3)); forvar3321 = (forvar3321 + (1'h1)))
                    begin
                      reg3322 <= $unsigned(({$unsigned(reg3139)} != reg2911));
                      reg3323 <= $signed((+$signed(forvar2876[(4'hb):(4'ha)])));
                    end
                end
            end
          for (forvar3324 = (1'h0); (forvar3324 < (1'h1)); forvar3324 = (forvar3324 + (1'h1)))
            begin
              for (forvar3325 = (1'h0); (forvar3325 < (2'h3)); forvar3325 = (forvar3325 + (1'h1)))
                begin
                  reg3326 <= reg3026[(2'h2):(1'h0)];
                  for (forvar3327 = (1'h0); (forvar3327 < (2'h2)); forvar3327 = (forvar3327 + (1'h1)))
                    begin
                      reg3328 <= forvar3135[(3'h7):(1'h1)];
                      reg3329 <= $unsigned(reg2775);
                      reg3330 <= ((8'hb9) == ($unsigned((reg3233 ?
                              reg3274 : forvar2908)) ?
                          forvar2876[(4'ha):(3'h5)] : ($unsigned(forvar2764) != (forvar3110 > (8'hae)))));
                      reg3331 <= $unsigned(($unsigned((reg2898 * forvar3033)) | $signed((reg3140 ?
                          reg3036 : forvar3060))));
                    end
                end
              for (forvar3332 = (1'h0); (forvar3332 < (2'h2)); forvar3332 = (forvar3332 + (1'h1)))
                begin
                  if (reg2996[(1'h0):(1'h0)])
                    begin
                      reg3333 <= (~|$unsigned(reg2949));
                      reg3334 <= (reg3238[(2'h3):(1'h0)] ?
                          $signed((+$unsigned(reg2952))) : (^((reg3006 ?
                                  reg2798 : forvar3177) ?
                              wire2752 : (reg3136 >> forvar3122))));
                    end
                  else
                    begin
                      reg3333 <= $unsigned((&(|reg3072[(1'h1):(1'h1)])));
                    end
                  if (reg3034)
                    begin
                      reg3335 <= (~|($unsigned((!reg2994)) ?
                          (reg3174[(2'h3):(1'h0)] != (forvar2959 ?
                              forvar3296 : (8'hb8))) : $unsigned(reg2793)));
                      reg3336 <= forvar3255;
                      reg3337 <= (8'hb8);
                      reg3338 <= reg2946[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg3335 <= ($signed($signed(((8'hb8) != forvar3021))) ?
                          $signed(((forvar2808 ?
                              (8'haa) : forvar2891) < reg2963[(4'h9):(3'h7)])) : reg2820);
                    end
                  if (((reg3026 == reg2922) ?
                      $unsigned((8'hb3)) : (reg2781[(2'h2):(2'h2)] ?
                          ({forvar3091} ^~ $signed(forvar3228)) : ((forvar3210 ?
                                  (8'hb4) : reg2958) ?
                              $unsigned(reg2998) : reg3170[(3'h7):(3'h6)]))))
                    begin
                      reg3339 <= (~^((((8'ha2) ^~ reg3227) <= $signed(reg3193)) ?
                          (|(^reg3072)) : ($signed(reg2976) != (forvar2855 ?
                              reg2800 : forvar2821))));
                      reg3340 <= (-$signed((|reg3033[(2'h3):(1'h1)])));
                      reg3341 <= (((^reg3205) <<< ($signed(reg2860) >> (^~reg2771))) >>> (({reg2830} >>> (&forvar3122)) ?
                          reg2847 : {(forvar2775 ? reg3064 : forvar3285)}));
                      reg3342 <= $unsigned((~&$unsigned(forvar3091[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg3339 <= reg3306[(3'h7):(3'h4)];
                      reg3340 <= reg2935;
                    end
                end
              for (forvar3343 = (1'h0); (forvar3343 < (2'h2)); forvar3343 = (forvar3343 + (1'h1)))
                begin
                  for (forvar3344 = (1'h0); (forvar3344 < (2'h3)); forvar3344 = (forvar3344 + (1'h1)))
                    begin
                      reg3345 <= {(+reg3248[(1'h0):(1'h0)])};
                    end
                  for (forvar3346 = (1'h0); (forvar3346 < (1'h1)); forvar3346 = (forvar3346 + (1'h1)))
                    begin
                      reg3347 <= (reg2877[(4'he):(3'h4)] * (&reg3272));
                    end
                  for (forvar3348 = (1'h0); (forvar3348 < (2'h3)); forvar3348 = (forvar3348 + (1'h1)))
                    begin
                      reg3349 <= $signed(reg2853[(2'h3):(2'h2)]);
                    end
                end
              for (forvar3350 = (1'h0); (forvar3350 < (2'h2)); forvar3350 = (forvar3350 + (1'h1)))
                begin
                  if (($signed(((reg2805 >>> forvar2945) && (~reg2889))) ?
                      ((!reg3098) * ((forvar3292 >= reg3000) ?
                          $unsigned((8'ha9)) : $signed(forvar3052))) : reg2780[(3'h6):(3'h4)]))
                    begin
                      reg3351 <= $signed(reg3014[(3'h6):(1'h1)]);
                      reg3352 <= $signed(reg3098);
                      reg3353 <= $unsigned($signed($signed((reg3150 ?
                          reg2805 : reg2771))));
                    end
                  else
                    begin
                      reg3351 <= {reg2861[(1'h0):(1'h0)]};
                      reg3352 <= reg2843;
                      reg3353 <= (~^reg3329[(2'h3):(1'h0)]);
                    end
                  if (reg3298[(1'h0):(1'h0)])
                    begin
                      reg3354 <= reg3050;
                    end
                  else
                    begin
                      reg3354 <= ($signed($unsigned($signed(reg3085))) | (forvar3061 ?
                          (forvar3168 > reg2983) : (8'hb9)));
                      reg3355 <= (reg3188[(4'he):(2'h2)] + reg3098[(4'hb):(2'h2)]);
                    end
                  for (forvar3356 = (1'h0); (forvar3356 < (1'h0)); forvar3356 = (forvar3356 + (1'h1)))
                    begin
                      reg3357 <= (8'ha9);
                      reg3358 <= ({$unsigned(reg3322[(3'h4):(2'h3)])} <<< (((reg3206 <<< reg2877) ?
                          $signed((8'ha2)) : (reg2780 >= (8'ha9))) && $unsigned(((8'hb9) ?
                          reg3148 : reg3144))));
                    end
                end
            end
        end
      for (forvar3359 = (1'h0); (forvar3359 < (2'h2)); forvar3359 = (forvar3359 + (1'h1)))
        begin
          reg3360 <= (~&$signed(($signed(reg2947) && forvar3043[(3'h5):(1'h1)])));
          if ((((~$signed(reg3089)) | ((reg2946 ? reg2905 : (8'ha1)) ?
              $signed(reg3180) : $unsigned(reg3101))) + reg2823[(1'h1):(1'h1)]))
            begin
              reg3361 <= ($unsigned(reg3105[(4'hc):(4'hc)]) ?
                  $unsigned((^~(reg2834 <= forvar3210))) : (-($unsigned(reg2944) & (reg3333 * reg3156))));
              for (forvar3362 = (1'h0); (forvar3362 < (1'h0)); forvar3362 = (forvar3362 + (1'h1)))
                begin
                  for (forvar3363 = (1'h0); (forvar3363 < (2'h3)); forvar3363 = (forvar3363 + (1'h1)))
                    begin
                      reg3364 <= (-$unsigned($unsigned(reg2950[(2'h3):(1'h0)])));
                    end
                  for (forvar3365 = (1'h0); (forvar3365 < (1'h0)); forvar3365 = (forvar3365 + (1'h1)))
                    begin
                      reg3366 <= (^~(~&($signed(reg3276) == (forvar2774 ?
                          reg2862 : (8'hb8)))));
                      reg3367 <= ($signed($unsigned(reg3063)) ?
                          $signed((forvar3142[(2'h2):(1'h0)] ?
                              (reg2883 ? reg2828 : reg3273) : (reg2796 ?
                                  reg3137 : reg2945))) : $signed(forvar3102[(2'h3):(2'h3)]));
                    end
                  reg3368 <= $unsigned($unsigned($unsigned((reg2841 ~^ (8'hab)))));
                  if ($signed({$unsigned(reg2946)}))
                    begin
                      reg3369 <= reg2814[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg3369 <= {$signed(forvar2950)};
                    end
                end
              if ($signed($signed((&((8'haa) ? reg2772 : forvar2948)))))
                begin
                  reg3370 <= $signed((forvar2920[(1'h0):(1'h0)] > $unsigned(reg2925[(1'h0):(1'h0)])));
                  if (((&((~reg3086) ?
                      (!reg2766) : $unsigned(reg2811))) ^~ $signed(forvar2902)))
                    begin
                      reg3371 <= (reg2947[(3'h4):(3'h4)] ?
                          {$unsigned(reg3110[(2'h3):(2'h2)])} : ((reg3338 ?
                              (-reg3230) : (~forvar2829)) >> ((|(8'ha3)) && (&reg2853))));
                      reg3372 <= reg3171[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg3371 <= (^~$unsigned(($signed(reg2839) > reg3273)));
                      reg3372 <= (reg2999 <<< $signed((~|(~&(8'ha5)))));
                      reg3373 <= forvar3311;
                    end
                end
              else
                begin
                  if (reg2870)
                    begin
                      reg3370 <= (reg3062[(3'h6):(2'h3)] * $unsigned((reg2932 ?
                          {reg3227} : reg2994[(2'h3):(1'h0)])));
                      reg3371 <= (({reg3126} ?
                              forvar3311 : $unsigned(reg3298[(2'h2):(2'h2)])) ?
                          (($signed(reg3188) ?
                              $unsigned(reg2874) : (reg3304 >>> forvar2861)) & (^~reg3052)) : {$signed($unsigned(reg2893))});
                    end
                  else
                    begin
                      reg3370 <= (reg3111 >= $unsigned($unsigned(reg2769)));
                      reg3371 <= forvar2908[(2'h2):(2'h2)];
                    end
                  for (forvar3372 = (1'h0); (forvar3372 < (1'h1)); forvar3372 = (forvar3372 + (1'h1)))
                    begin
                      reg3373 <= ($unsigned(({reg3251} + $signed(forvar3012))) || ({(forvar3045 ?
                                  reg3020 : reg3112)} ?
                          (~|$unsigned(reg3349)) : ((reg2914 << reg3120) >= $signed(forvar3203))));
                      reg3374 <= $signed(($signed($signed(forvar2842)) == reg2946));
                      reg3375 <= {$signed($signed((~|reg2882)))};
                      reg3376 <= (($signed({reg3010}) ?
                          $signed(((8'ha6) ?
                              reg3329 : reg2759)) : (forvar3346[(3'h7):(1'h1)] - (reg3244 ?
                              (8'hb9) : reg2943))) & $unsigned(reg2943[(2'h2):(1'h0)]));
                    end
                  if (reg2939)
                    begin
                      reg3377 <= forvar3255;
                      reg3378 <= $unsigned($signed({reg3219}));
                    end
                  else
                    begin
                      reg3377 <= $unsigned($signed($signed($signed(reg3089))));
                    end
                  for (forvar3379 = (1'h0); (forvar3379 < (1'h0)); forvar3379 = (forvar3379 + (1'h1)))
                    begin
                      reg3380 <= (~^((&(reg2842 ~^ reg2882)) <<< reg3269[(2'h2):(2'h2)]));
                    end
                end
            end
          else
            begin
              for (forvar3361 = (1'h0); (forvar3361 < (1'h1)); forvar3361 = (forvar3361 + (1'h1)))
                begin
                  if ((reg2950[(3'h5):(2'h3)] | $unsigned((!reg3317))))
                    begin
                      reg3362 <= (|$unsigned(({reg2755} ?
                          (reg3199 ~^ forvar3157) : $signed(reg3009))));
                      reg3363 <= $unsigned(($unsigned(((8'hb1) ?
                          reg3295 : reg3091)) >= $signed($unsigned(forvar2968))));
                      reg3364 <= ((+{(~|forvar2764)}) ?
                          $signed({reg3208}) : ($signed(forvar3325[(3'h5):(1'h1)]) + (reg2788 ?
                              $unsigned(reg3225) : (forvar3321 || forvar3007))));
                      reg3365 <= forvar3091;
                    end
                  else
                    begin
                      reg3362 <= (reg2981[(2'h2):(1'h0)] | ((forvar3022[(1'h0):(1'h0)] * (reg3354 ?
                          reg2761 : reg2798)) >>> reg3143[(1'h1):(1'h0)]));
                    end
                end
              if ($unsigned(($signed(reg3352[(4'h9):(4'h8)]) ?
                  ((reg3349 ?
                      (8'hae) : reg2946) + (forvar3070 > reg2936)) : reg2924)))
                begin
                  reg3366 <= reg3219[(1'h1):(1'h0)];
                  if ($signed($signed(reg3250)))
                    begin
                      reg3367 <= ({$unsigned($unsigned(reg3252))} > reg3063[(1'h1):(1'h0)]);
                      reg3368 <= $unsigned(reg2977);
                    end
                  else
                    begin
                      reg3367 <= (({(reg3331 * reg3012)} & reg2959) ?
                          reg3147[(2'h2):(2'h2)] : $unsigned((~|$signed(forvar2842))));
                      reg3368 <= ($signed((forvar3007 ?
                              (8'hb6) : reg2959[(2'h3):(1'h0)])) ?
                          forvar2783 : {($unsigned(reg3096) > forvar2950)});
                      reg3369 <= reg2989;
                    end
                  if ((((^$unsigned(forvar3095)) ?
                          ($signed(reg2923) ?
                              ((8'hac) | reg3179) : $unsigned((8'hb3))) : (reg3208[(2'h3):(1'h1)] | $signed(reg3032))) ?
                      reg2989[(1'h0):(1'h0)] : $signed({$unsigned(reg2823)})))
                    begin
                      reg3370 <= $signed(reg3007[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg3370 <= reg3100[(3'h6):(1'h0)];
                    end
                  reg3371 <= ((~|($signed(reg2943) ?
                      reg3216[(1'h1):(1'h1)] : (reg2792 ?
                          reg2811 : reg3010))) <<< $unsigned(($signed((8'hb9)) ?
                      $signed(reg3233) : $signed(reg3107))));
                end
              else
                begin
                  if ($signed((8'h9c)))
                    begin
                      reg3366 <= reg3284[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3366 <= reg2801;
                    end
                  for (forvar3367 = (1'h0); (forvar3367 < (2'h2)); forvar3367 = (forvar3367 + (1'h1)))
                    begin
                      reg3368 <= $signed((+reg2866[(1'h0):(1'h0)]));
                    end
                  if ({reg3054[(3'h5):(3'h4)]})
                    begin
                      reg3369 <= (($signed((forvar2797 >>> (8'hb9))) ?
                          (!reg2813[(2'h2):(2'h2)]) : (8'hb4)) >= (8'hac));
                      reg3370 <= reg2883;
                      reg3371 <= (((8'hb8) ^ {forvar3237}) ?
                          (forvar2862[(4'hc):(4'h8)] >>> (8'hab)) : ($unsigned((8'h9c)) ?
                              (^((8'h9c) || reg2779)) : reg3038));
                    end
                  else
                    begin
                      reg3369 <= wire2752[(3'h5):(3'h4)];
                    end
                  for (forvar3372 = (1'h0); (forvar3372 < (1'h0)); forvar3372 = (forvar3372 + (1'h1)))
                    begin
                      reg3373 <= reg3047;
                      reg3374 <= (-reg2767);
                      reg3375 <= (((8'haf) <<< (~^{reg3096})) ~^ ((~&(~&(8'hb8))) ?
                          (~^$signed(forvar2826)) : reg3084[(2'h2):(2'h2)]));
                    end
                end
            end
          for (forvar3381 = (1'h0); (forvar3381 < (1'h0)); forvar3381 = (forvar3381 + (1'h1)))
            begin
              if ({reg3032})
                begin
                  if (({$unsigned({reg3024})} ?
                      reg2914 : {((reg3073 ?
                              (8'hb0) : forvar3187) ~^ reg2791)}))
                    begin
                      reg3382 <= reg3259;
                      reg3383 <= ((!(8'haf)) ^~ reg3025);
                      reg3384 <= (~reg3361);
                      reg3385 <= ((|(((8'hb0) * reg3047) ?
                              (reg3317 ? reg2932 : reg2860) : {(8'ha1)})) ?
                          $signed((|(reg2914 ?
                              reg3011 : reg2759))) : reg2869[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg3382 <= (~&$signed(reg3174));
                    end
                  if (((reg3137 ?
                      $unsigned((reg3261 ?
                          reg3203 : reg3145)) : {(~reg3316)}) | (((forvar2963 ?
                          reg3153 : reg3067) * forvar3109) ?
                      reg2922[(4'he):(3'h4)] : reg3233)))
                    begin
                      reg3386 <= reg2932[(3'h4):(2'h2)];
                      reg3387 <= (!reg3025);
                      reg3388 <= $signed(reg2926);
                      reg3389 <= forvar3344;
                    end
                  else
                    begin
                      reg3386 <= ((({reg3385} ?
                                  reg2777 : (forvar3186 ? reg2882 : (8'ha2))) ?
                              {reg3007[(1'h0):(1'h0)]} : reg3298[(1'h0):(1'h0)]) ?
                          reg3022[(2'h2):(1'h0)] : ($unsigned(((8'ha0) + reg3374)) ^ (reg3115[(2'h3):(1'h0)] ?
                              (^~(8'ha8)) : reg3159)));
                      reg3387 <= reg2869;
                      reg3388 <= reg3063;
                    end
                  for (forvar3390 = (1'h0); (forvar3390 < (1'h1)); forvar3390 = (forvar3390 + (1'h1)))
                    begin
                      reg3391 <= $signed($signed({(^reg3264)}));
                    end
                  reg3392 <= reg3229[(1'h1):(1'h1)];
                end
              else
                begin
                  for (forvar3382 = (1'h0); (forvar3382 < (1'h1)); forvar3382 = (forvar3382 + (1'h1)))
                    begin
                      reg3383 <= (8'hae);
                      reg3384 <= (~|reg2944[(1'h1):(1'h0)]);
                    end
                  reg3385 <= (($signed(reg2802) ?
                      reg2924 : (~^(forvar3200 < reg2788))) ~^ (reg2992 ?
                      {$signed(reg3012)} : reg2940));
                  reg3386 <= reg3256;
                end
            end
        end
      if ((~^reg2922))
        begin
          reg3393 <= (-$unsigned(($signed(forvar3061) <<< reg3366[(2'h2):(2'h2)])));
        end
      else
        begin
          reg3393 <= $signed({{$signed(reg2884)}});
          for (forvar3394 = (1'h0); (forvar3394 < (1'h0)); forvar3394 = (forvar3394 + (1'h1)))
            begin
              if ($unsigned(reg3010[(2'h2):(1'h1)]))
                begin
                  if ($signed($signed(reg2788[(3'h4):(1'h1)])))
                    begin
                      reg3395 <= $signed(({reg3144} && (~|(reg2938 ?
                          reg2816 : reg2825))));
                      reg3396 <= $unsigned({{reg2837}});
                    end
                  else
                    begin
                      reg3395 <= forvar2776[(3'h4):(2'h3)];
                      reg3396 <= forvar2876;
                    end
                  for (forvar3397 = (1'h0); (forvar3397 < (1'h1)); forvar3397 = (forvar3397 + (1'h1)))
                    begin
                      reg3398 <= $unsigned($signed((reg2811 - {reg2800})));
                      reg3399 <= $signed(($unsigned($signed(reg3264)) ~^ $signed(reg3110[(3'h5):(2'h3)])));
                      reg3400 <= $unsigned($unsigned(forvar2838[(2'h3):(2'h2)]));
                    end
                  for (forvar3401 = (1'h0); (forvar3401 < (2'h3)); forvar3401 = (forvar3401 + (1'h1)))
                    begin
                      reg3402 <= $unsigned(reg2833);
                      reg3403 <= {$unsigned((8'hb6))};
                    end
                  for (forvar3404 = (1'h0); (forvar3404 < (2'h2)); forvar3404 = (forvar3404 + (1'h1)))
                    begin
                      reg3405 <= ((8'ha0) ?
                          (!reg2846[(1'h0):(1'h0)]) : (reg3355[(2'h2):(1'h1)] << ($unsigned(reg2888) ^ (reg2875 || reg3039))));
                      reg3406 <= $signed($signed({(reg2853 <<< reg2773)}));
                    end
                end
              else
                begin
                  for (forvar3395 = (1'h0); (forvar3395 < (2'h3)); forvar3395 = (forvar3395 + (1'h1)))
                    begin
                      reg3396 <= $signed(((wire1763 ?
                          (reg2978 ?
                              (8'hb4) : forvar3016) : reg2755[(3'h5):(3'h4)]) <<< forvar2990[(1'h1):(1'h1)]));
                    end
                  for (forvar3397 = (1'h0); (forvar3397 < (1'h1)); forvar3397 = (forvar3397 + (1'h1)))
                    begin
                      reg3398 <= reg3228;
                      reg3399 <= reg3011[(3'h6):(2'h2)];
                      reg3400 <= $signed((8'hb1));
                      reg3401 <= $signed((((forvar2829 && (8'hb0)) && reg3015) ~^ ($unsigned(forvar2912) <= (forvar2770 * (8'hae)))));
                    end
                  for (forvar3402 = (1'h0); (forvar3402 < (1'h1)); forvar3402 = (forvar3402 + (1'h1)))
                    begin
                      reg3403 <= (^~$signed(({reg3236} ?
                          reg2977[(3'h7):(1'h0)] : ((8'ha1) ?
                              reg2841 : reg3196))));
                      reg3404 <= $unsigned(reg2807[(3'h4):(1'h0)]);
                      reg3405 <= ($signed((+$signed(reg3180))) ?
                          (reg3199[(4'he):(4'ha)] ?
                              $signed($unsigned(forvar3125)) : forvar3275[(4'h8):(3'h4)]) : $unsigned($unsigned($unsigned(reg2941))));
                    end
                end
              reg3407 <= ($signed($unsigned($signed((8'h9c)))) ?
                  ((^reg3221[(3'h7):(3'h6)]) > {{reg3101}}) : reg2920);
              if ($signed(((reg2989 ~^ {forvar3215}) == reg3405)))
                begin
                  if (reg3338[(2'h3):(1'h0)])
                    begin
                      reg3408 <= (^~($unsigned((~|wire1762)) | reg2967[(1'h1):(1'h0)]));
                      reg3409 <= ($signed(((forvar2925 ? reg2768 : reg2819) ?
                          $unsigned(forvar2865) : (~^reg3257))) == $signed((~^$signed(forvar3045))));
                      reg3410 <= {$signed(reg3396)};
                      reg3411 <= reg3257[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg3408 <= ($unsigned((+((8'ha1) ? (8'ha2) : reg2986))) ?
                          (reg2865[(4'hc):(3'h6)] - reg3319) : $unsigned(reg3192));
                    end
                  reg3412 <= {$signed($unsigned($signed(forvar2955)))};
                end
              else
                begin
                  for (forvar3408 = (1'h0); (forvar3408 < (2'h2)); forvar3408 = (forvar3408 + (1'h1)))
                    begin
                      reg3409 <= (8'hb8);
                    end
                  reg3410 <= forvar3205[(1'h1):(1'h1)];
                end
              for (forvar3413 = (1'h0); (forvar3413 < (1'h1)); forvar3413 = (forvar3413 + (1'h1)))
                begin
                  if (reg2935[(1'h0):(1'h0)])
                    begin
                      reg3414 <= $unsigned(reg2867);
                    end
                  else
                    begin
                      reg3414 <= reg2793[(1'h1):(1'h1)];
                      reg3415 <= $signed(($signed($signed(reg2915)) ?
                          (reg2995[(1'h1):(1'h0)] ?
                              (^reg2975) : {reg2853}) : ($unsigned(reg3314) ?
                              $unsigned((8'ha1)) : (reg2805 ?
                                  reg2864 : wire1760))));
                    end
                  for (forvar3416 = (1'h0); (forvar3416 < (2'h2)); forvar3416 = (forvar3416 + (1'h1)))
                    begin
                      reg3417 <= (({(reg3017 ^ reg3121)} << ((forvar3255 ?
                                  reg3141 : (8'h9f)) ?
                              {reg3039} : {(8'hb2)})) ?
                          ({reg3196[(2'h3):(1'h1)]} == ({reg3204} ?
                              (reg3300 ?
                                  reg2900 : reg3170) : reg3193[(2'h2):(1'h1)])) : (|reg3169[(4'h9):(4'h9)]));
                      reg3418 <= ((^(8'ha6)) + $signed(reg2957));
                      reg3419 <= (+$unsigned((reg2937[(4'hd):(1'h1)] >= (reg2881 - reg3082))));
                      reg3420 <= (!(($signed(reg3417) ?
                          (~|(8'ha4)) : (reg3044 >> reg3267)) < reg3316));
                    end
                  reg3421 <= ((^~(8'hae)) ?
                      {$signed($unsigned(reg2830))} : {({reg3270} - ((8'ha0) ?
                              forvar3394 : forvar2797))});
                  for (forvar3422 = (1'h0); (forvar3422 < (2'h2)); forvar3422 = (forvar3422 + (1'h1)))
                    begin
                      reg3423 <= ($signed($unsigned($signed(reg2927))) ?
                          wire2753[(4'h8):(3'h4)] : (!((^forvar3033) << $unsigned(reg2875))));
                    end
                end
            end
          for (forvar3424 = (1'h0); (forvar3424 < (2'h3)); forvar3424 = (forvar3424 + (1'h1)))
            begin
              reg3425 <= {((~|(reg3063 ? forvar3109 : (8'h9c))) ?
                      ($unsigned(reg3209) ?
                          (forvar3114 ?
                              reg3411 : reg3401) : (8'ha8)) : ($signed(forvar2958) ?
                          (^~forvar2797) : {reg3401}))};
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar3426 = (1'h0); (forvar3426 < (2'h3)); forvar3426 = (forvar3426 + (1'h1)))
        begin
          for (forvar3427 = (1'h0); (forvar3427 < (1'h0)); forvar3427 = (forvar3427 + (1'h1)))
            begin
              if ($unsigned(reg2883))
                begin
                  for (forvar3428 = (1'h0); (forvar3428 < (1'h1)); forvar3428 = (forvar3428 + (1'h1)))
                    begin
                      reg3429 <= (^(reg2756 <= (!reg3226[(2'h2):(1'h1)])));
                      reg3430 <= $signed($signed($signed((^forvar2920))));
                      reg3431 <= reg3185;
                      reg3432 <= reg3259[(3'h4):(2'h3)];
                    end
                  reg3433 <= (^(-(((8'hb8) >>> forvar3274) & reg3347[(1'h1):(1'h1)])));
                  if ($unsigned((($unsigned(forvar3130) != $signed((8'ha6))) ?
                      {$signed((8'haf))} : $signed({(8'ha2)}))))
                    begin
                      reg3434 <= $signed($unsigned((^~reg2995)));
                      reg3435 <= $unsigned((reg3367 >> (^~(forvar3350 >= reg2972))));
                      reg3436 <= $unsigned((~reg2848[(4'ha):(1'h1)]));
                    end
                  else
                    begin
                      reg3434 <= $signed($unsigned($signed(reg3217)));
                    end
                  for (forvar3437 = (1'h0); (forvar3437 < (2'h3)); forvar3437 = (forvar3437 + (1'h1)))
                    begin
                      reg3438 <= (&$signed(reg2884));
                      reg3439 <= ((8'ha5) ^~ (reg2939 ?
                          $unsigned(reg3287[(4'h9):(2'h3)]) : (~forvar2798[(2'h3):(1'h0)])));
                      reg3440 <= reg3073[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if (((((reg2941 ? reg2787 : forvar2855) ?
                          (forvar3283 ? reg2791 : reg2962) : (forvar2803 ?
                              reg2806 : forvar2808)) ?
                      ({(8'hac)} == {(8'h9c)}) : (+forvar2808[(3'h7):(2'h3)])) != ($signed(reg3009) && (-(~&reg3291)))))
                    begin
                      reg3428 <= reg3128[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg3428 <= forvar3297[(4'h8):(4'h8)];
                      reg3429 <= ({(&(reg2961 ?
                              (8'hab) : reg3162))} <<< reg2758[(1'h1):(1'h0)]);
                      reg3430 <= reg2876;
                      reg3431 <= reg2991[(4'ha):(2'h3)];
                    end
                end
              for (forvar3441 = (1'h0); (forvar3441 < (2'h2)); forvar3441 = (forvar3441 + (1'h1)))
                begin
                  reg3442 <= $unsigned(((reg3371 << ((8'h9d) + (8'hab))) ?
                      ($signed(reg2893) ?
                          $unsigned(reg3376) : (reg2898 << reg2780)) : reg3401[(2'h2):(2'h2)]));
                  if ((!(~^{wire1762})))
                    begin
                      reg3443 <= (forvar3011[(3'h7):(2'h2)] | reg3040);
                      reg3444 <= (8'hb3);
                      reg3445 <= {(|(~^(reg3171 ? reg3204 : forvar2865)))};
                    end
                  else
                    begin
                      reg3443 <= $signed($unsigned(reg3349));
                      reg3444 <= {$signed(((^reg3013) ? (8'hb4) : reg3064))};
                    end
                  reg3446 <= reg2828;
                  if ($signed(((((8'ha0) >> forvar3005) ^~ $unsigned(reg3189)) | ($unsigned(forvar3084) ?
                      (reg3243 ?
                          (8'hb9) : forvar3143) : (forvar3324 <= forvar3139)))))
                    begin
                      reg3447 <= $unsigned(((((8'ha7) >= reg3411) ?
                              (^~reg3403) : $unsigned(reg3001)) ?
                          ((-(8'h9f)) ? (|(8'ha0)) : (!(8'ha0))) : forvar3344));
                      reg3448 <= $unsigned({(^(reg2986 ? reg3393 : (8'hb2)))});
                      reg3449 <= forvar3350;
                    end
                  else
                    begin
                      reg3447 <= reg3282[(4'hd):(1'h1)];
                      reg3448 <= ((~((^~reg3047) ?
                              reg3104[(2'h3):(2'h2)] : (reg3024 ?
                                  reg3207 : reg2873))) ?
                          (+reg3100[(1'h0):(1'h0)]) : (^((forvar3428 == reg2852) ?
                              {(8'had)} : $signed(reg3349))));
                    end
                end
            end
        end
      for (forvar3450 = (1'h0); (forvar3450 < (2'h3)); forvar3450 = (forvar3450 + (1'h1)))
        begin
          for (forvar3451 = (1'h0); (forvar3451 < (2'h3)); forvar3451 = (forvar3451 + (1'h1)))
            begin
              reg3452 <= $unsigned($unsigned(forvar3164));
              for (forvar3453 = (1'h0); (forvar3453 < (1'h1)); forvar3453 = (forvar3453 + (1'h1)))
                begin
                  if ((~&($signed((!reg2915)) ^~ {$signed((8'hb9))})))
                    begin
                      reg3454 <= ($unsigned(($unsigned(reg3244) & {reg3391})) ?
                          reg2816[(2'h2):(2'h2)] : (~{$signed(reg2801)}));
                      reg3455 <= (+reg3195[(1'h1):(1'h0)]);
                      reg3456 <= {($signed($signed(reg2878)) ?
                              ($signed((8'hb3)) | (8'hb7)) : ($signed(reg2991) ?
                                  (reg3113 <= forvar2849) : {reg3353}))};
                    end
                  else
                    begin
                      reg3454 <= (+(+(reg3307[(3'h5):(1'h0)] != (forvar3437 ?
                          reg2914 : reg3096))));
                    end
                  for (forvar3457 = (1'h0); (forvar3457 < (1'h1)); forvar3457 = (forvar3457 + (1'h1)))
                    begin
                      reg3458 <= (!$unsigned((forvar3255[(1'h1):(1'h1)] | $signed(reg3226))));
                    end
                end
            end
        end
      reg3459 <= {$signed($signed((reg3329 ? reg3222 : (8'haa))))};
      for (forvar3460 = (1'h0); (forvar3460 < (2'h2)); forvar3460 = (forvar3460 + (1'h1)))
        begin
          if ($signed(reg2787))
            begin
              if (reg3338)
                begin
                  for (forvar3461 = (1'h0); (forvar3461 < (1'h0)); forvar3461 = (forvar3461 + (1'h1)))
                    begin
                      reg3462 <= {{reg2835}};
                      reg3463 <= $signed(reg2876[(1'h1):(1'h0)]);
                      reg3464 <= (8'ha7);
                      reg3465 <= (~&$unsigned($unsigned({reg2962})));
                    end
                  if ((forvar2968[(2'h3):(2'h2)] ~^ (reg3257[(1'h1):(1'h1)] ?
                      reg3268 : ($signed(forvar3016) != $signed((8'ha4))))))
                    begin
                      reg3466 <= {reg2879};
                      reg3467 <= $signed(($signed((+(8'haa))) * reg3155));
                      reg3468 <= (forvar3056 ?
                          reg3191 : $signed((!((8'hb8) ~^ reg3170))));
                    end
                  else
                    begin
                      reg3466 <= ((((~reg2922) ?
                                  reg2779 : (forvar3045 ? reg2998 : reg3029)) ?
                              (~|{reg3232}) : ((8'h9e) & $signed((8'ha2)))) ?
                          reg2876 : ($unsigned(reg2905[(3'h6):(3'h5)]) ?
                              (~&((8'hb7) ? reg3433 : reg2868)) : forvar2783));
                    end
                end
              else
                begin
                  if ((((reg3238[(3'h7):(3'h6)] ?
                          (reg3086 ?
                              reg2760 : reg3435) : forvar2945[(4'hc):(3'h7)]) ?
                      $signed((~&reg3391)) : $signed($signed(reg3105))) ^~ $signed(((reg3400 ?
                          (8'had) : forvar3395) ?
                      (~(8'hb7)) : reg3342[(3'h4):(3'h4)]))))
                    begin
                      reg3461 <= $signed((reg3006 ?
                          reg3120 : (reg2949[(4'hc):(4'ha)] ?
                              (forvar3183 >>> reg2982) : reg3364)));
                    end
                  else
                    begin
                      reg3461 <= reg3449;
                      reg3462 <= (forvar2917 ~^ reg2805);
                    end
                end
            end
          else
            begin
              for (forvar3461 = (1'h0); (forvar3461 < (1'h1)); forvar3461 = (forvar3461 + (1'h1)))
                begin
                  if ((reg3138[(3'h4):(1'h0)] >>> $signed(reg3374[(2'h3):(1'h0)])))
                    begin
                      reg3462 <= (~reg3035);
                    end
                  else
                    begin
                      reg3462 <= $signed(($unsigned(forvar3404[(3'h7):(1'h1)]) ?
                          (&(forvar2902 ?
                              reg3048 : reg3188)) : reg3073[(1'h0):(1'h0)]));
                      reg3463 <= reg3052[(3'h7):(3'h7)];
                    end
                  for (forvar3464 = (1'h0); (forvar3464 < (2'h3)); forvar3464 = (forvar3464 + (1'h1)))
                    begin
                      reg3465 <= ($unsigned(($signed(reg2978) ?
                              reg2823 : (forvar2822 ? reg2960 : (8'hb4)))) ?
                          forvar2801[(4'h9):(3'h6)] : $unsigned(($unsigned((8'ha4)) ?
                              {reg3137} : (~reg2813))));
                    end
                  for (forvar3466 = (1'h0); (forvar3466 < (2'h2)); forvar3466 = (forvar3466 + (1'h1)))
                    begin
                      reg3467 <= ($signed({reg3103[(4'hb):(3'h5)]}) ?
                          (&$signed((~&reg2761))) : forvar3325[(1'h1):(1'h1)]);
                      reg3468 <= ($unsigned(reg3257[(1'h1):(1'h0)]) & {((reg2810 ?
                              reg3057 : reg3176) ^ reg2834[(2'h3):(2'h2)])});
                    end
                  if ((!forvar2978[(2'h3):(2'h3)]))
                    begin
                      reg3469 <= ($unsigned((8'ha9)) ?
                          (8'ha4) : {{forvar2990}});
                      reg3470 <= reg3099;
                      reg3471 <= $unsigned($signed($unsigned($signed(forvar3441))));
                      reg3472 <= (~^($unsigned((~&forvar3223)) ?
                          reg2788[(2'h3):(2'h3)] : {$unsigned(forvar3297)}));
                    end
                  else
                    begin
                      reg3469 <= $signed(forvar3012);
                      reg3470 <= ($signed(($signed(reg2931) <<< reg2872[(1'h1):(1'h0)])) >= ((&(reg3106 ^ (8'haa))) ^~ (~|$signed(reg3431))));
                      reg3471 <= {reg3055};
                      reg3472 <= reg3391[(1'h1):(1'h1)];
                    end
                end
            end
          if (reg3180)
            begin
              if (forvar3242)
                begin
                  for (forvar3473 = (1'h0); (forvar3473 < (1'h1)); forvar3473 = (forvar3473 + (1'h1)))
                    begin
                      reg3474 <= {reg3304};
                      reg3475 <= reg3375;
                      reg3476 <= ($signed((&(~reg3108))) <<< (8'ha5));
                      reg3477 <= reg2925;
                    end
                  if ($signed($signed(reg3466)))
                    begin
                      reg3478 <= ($signed($unsigned(reg2939[(1'h0):(1'h0)])) ?
                          {(^$unsigned(reg3206))} : $signed($unsigned($signed(forvar3232))));
                    end
                  else
                    begin
                      reg3478 <= $signed(reg3270[(1'h1):(1'h0)]);
                      reg3479 <= $signed(forvar3461);
                      reg3480 <= ($unsigned(reg3243[(3'h5):(3'h5)]) == {(~&(reg3306 ?
                              reg3052 : reg3272))});
                    end
                  reg3481 <= $signed($signed({(forvar3297 ?
                          reg3367 : reg3231)}));
                end
              else
                begin
                  if (($signed(reg2773[(3'h7):(3'h5)]) ?
                      $signed($signed($unsigned(reg3222))) : $signed($signed(reg3015[(1'h1):(1'h1)]))))
                    begin
                      reg3473 <= reg3317;
                      reg3474 <= ({reg2784[(3'h7):(2'h3)]} ^~ $signed($signed(reg3005[(3'h6):(3'h5)])));
                      reg3475 <= reg2916[(3'h6):(3'h4)];
                      reg3476 <= ($signed(({reg2956} & (reg2880 != reg3373))) ^~ (~&(~|(forvar3210 ?
                          (8'ha2) : (8'hb3)))));
                    end
                  else
                    begin
                      reg3473 <= reg2995[(4'h8):(2'h2)];
                      reg3474 <= (~&reg3430[(3'h5):(3'h5)]);
                      reg3475 <= reg2952[(4'h9):(1'h1)];
                      reg3476 <= $unsigned((8'haa));
                    end
                  if (reg3097)
                    begin
                      reg3477 <= forvar3453[(1'h0):(1'h0)];
                      reg3478 <= {(($signed(reg3094) >> $unsigned(forvar3457)) ^ $unsigned((~^reg3144)))};
                    end
                  else
                    begin
                      reg3477 <= reg3339[(4'hb):(1'h1)];
                      reg3478 <= ((~((reg3078 ^ forvar3007) != (reg3033 ?
                          reg3202 : forvar2754))) && ((&(reg3473 ?
                          reg3289 : forvar3163)) ~^ (~^(reg3167 ?
                          forvar2783 : (8'hb6)))));
                      reg3479 <= reg2967[(1'h1):(1'h0)];
                    end
                end
              for (forvar3482 = (1'h0); (forvar3482 < (1'h1)); forvar3482 = (forvar3482 + (1'h1)))
                begin
                  if ({reg2813[(2'h3):(2'h3)]})
                    begin
                      reg3483 <= $signed(forvar3203[(4'h9):(2'h3)]);
                    end
                  else
                    begin
                      reg3483 <= reg2775;
                      reg3484 <= ({$signed(reg3211[(3'h7):(3'h5)])} >>> {$signed($unsigned(reg2928))});
                      reg3485 <= ($signed($signed($signed(forvar3292))) | ({reg3419} ~^ ({forvar3075} >> (8'ha3))));
                    end
                  reg3486 <= forvar3005[(3'h4):(2'h2)];
                  if ($unsigned($unsigned($signed(reg2999[(1'h0):(1'h0)]))))
                    begin
                      reg3487 <= reg2820[(4'ha):(1'h1)];
                    end
                  else
                    begin
                      reg3487 <= (!{(~forvar3095)});
                      reg3488 <= (({reg3077[(4'h8):(2'h2)]} ?
                          $unsigned($signed(reg3167)) : (|$unsigned(reg2878))) >> forvar2912);
                    end
                  for (forvar3489 = (1'h0); (forvar3489 < (2'h3)); forvar3489 = (forvar3489 + (1'h1)))
                    begin
                      reg3490 <= reg3333;
                      reg3491 <= $signed((($unsigned(reg3447) ?
                              (reg3026 ~^ reg3209) : (reg3072 ?
                                  reg2950 : reg3233)) ?
                          reg2819[(3'h5):(3'h4)] : (8'had)));
                    end
                end
              for (forvar3492 = (1'h0); (forvar3492 < (1'h0)); forvar3492 = (forvar3492 + (1'h1)))
                begin
                  for (forvar3493 = (1'h0); (forvar3493 < (2'h3)); forvar3493 = (forvar3493 + (1'h1)))
                    begin
                      reg3494 <= (|forvar3091);
                      reg3495 <= (reg3097 ?
                          $unsigned((&(reg3285 >> forvar3247))) : $unsigned((+forvar3112)));
                    end
                  if ($signed(((^reg3181) ?
                      (~((8'haa) & forvar3110)) : reg2957[(4'h9):(3'h6)])))
                    begin
                      reg3496 <= (reg2975[(2'h2):(2'h2)] || reg3225);
                      reg3497 <= $unsigned($unsigned(reg3341));
                      reg3498 <= forvar3090[(3'h4):(1'h0)];
                      reg3499 <= $signed(reg3369[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg3496 <= reg2758;
                      reg3497 <= reg3154[(3'h5):(2'h3)];
                      reg3498 <= $signed((|(~^reg3062[(4'hc):(2'h2)])));
                    end
                  for (forvar3500 = (1'h0); (forvar3500 < (1'h0)); forvar3500 = (forvar3500 + (1'h1)))
                    begin
                      reg3501 <= $unsigned(reg3341[(2'h3):(1'h0)]);
                    end
                end
            end
          else
            begin
              if (reg3233)
                begin
                  reg3473 <= ({forvar3451[(3'h4):(2'h2)]} <<< $signed($unsigned((reg3382 - reg3374))));
                end
              else
                begin
                  for (forvar3473 = (1'h0); (forvar3473 < (1'h1)); forvar3473 = (forvar3473 + (1'h1)))
                    begin
                      reg3474 <= reg2938;
                      reg3475 <= ((|$unsigned(reg3013)) - $signed(reg2945[(1'h0):(1'h0)]));
                    end
                end
              for (forvar3476 = (1'h0); (forvar3476 < (1'h0)); forvar3476 = (forvar3476 + (1'h1)))
                begin
                  for (forvar3477 = (1'h0); (forvar3477 < (2'h3)); forvar3477 = (forvar3477 + (1'h1)))
                    begin
                      reg3478 <= (($unsigned({reg2836}) ?
                          {(~^forvar3460)} : (~&(reg3410 ?
                              reg2927 : reg2794))) ^~ {reg3281[(1'h0):(1'h0)]});
                    end
                  if (((|((forvar3453 ? forvar3108 : reg3336) ?
                      (reg3018 ~^ reg3432) : reg3112)) || ($unsigned((!reg2968)) ?
                      (&reg3134) : $signed(reg2898))))
                    begin
                      reg3479 <= reg2789;
                      reg3480 <= reg2779;
                      reg3481 <= $signed($unsigned((+(^~reg2929))));
                    end
                  else
                    begin
                      reg3479 <= $unsigned({forvar2943});
                      reg3480 <= (($unsigned({reg3376}) <= $signed((forvar3288 - (8'hab)))) & {$unsigned($signed(reg3011))});
                    end
                end
              for (forvar3482 = (1'h0); (forvar3482 < (1'h1)); forvar3482 = (forvar3482 + (1'h1)))
                begin
                  for (forvar3483 = (1'h0); (forvar3483 < (1'h1)); forvar3483 = (forvar3483 + (1'h1)))
                    begin
                      reg3484 <= reg3317[(4'hc):(4'hb)];
                      reg3485 <= $unsigned((~^$signed($unsigned(forvar3344))));
                    end
                  for (forvar3486 = (1'h0); (forvar3486 < (2'h3)); forvar3486 = (forvar3486 + (1'h1)))
                    begin
                      reg3487 <= reg3372;
                      reg3488 <= {(reg2841[(1'h0):(1'h0)] ~^ forvar2919)};
                      reg3489 <= (^~(reg3360 ?
                          (^~reg3244[(1'h1):(1'h0)]) : (forvar3033[(2'h3):(2'h3)] ?
                              (reg2798 ? reg2983 : reg3309) : (|reg3231))));
                      reg3490 <= ($signed(reg2796) != $signed({forvar2892}));
                    end
                end
              for (forvar3491 = (1'h0); (forvar3491 < (2'h3)); forvar3491 = (forvar3491 + (1'h1)))
                begin
                  for (forvar3492 = (1'h0); (forvar3492 < (1'h1)); forvar3492 = (forvar3492 + (1'h1)))
                    begin
                      reg3493 <= (~|(^~$unsigned($signed(reg2939))));
                      reg3494 <= reg3365;
                    end
                end
            end
        end
    end
  module3502 modinst3602 (wire3601, clk, reg3205, reg3226, reg3095, reg3181, reg2868);
  module3603 modinst4018 (.wire3606(forvar3232), .clk(clk), .wire3604(reg3493), .wire3605(reg3229), .y(wire4017), .wire3608(reg2873), .wire3607(reg3363));
  assign wire4019 = forvar3186;
  always
    @(posedge clk) begin
      for (forvar4020 = (1'h0); (forvar4020 < (2'h3)); forvar4020 = (forvar4020 + (1'h1)))
        begin
          if ($unsigned((|reg3180[(3'h5):(1'h1)])))
            begin
              if ($unsigned(($unsigned((-reg2948)) ?
                  ($signed((8'hb8)) ?
                      {forvar3363} : $unsigned(forvar3492)) : {(forvar2993 ?
                          (8'ha9) : forvar3095)})))
                begin
                  for (forvar4021 = (1'h0); (forvar4021 < (1'h0)); forvar4021 = (forvar4021 + (1'h1)))
                    begin
                      reg4022 <= {{reg2769}};
                      reg4023 <= (^(reg3119 ?
                          forvar3152[(1'h0):(1'h0)] : (|reg3169[(3'h5):(1'h1)])));
                      reg4024 <= wire1760;
                      reg4025 <= forvar3343[(3'h5):(3'h4)];
                    end
                  for (forvar4026 = (1'h0); (forvar4026 < (1'h1)); forvar4026 = (forvar4026 + (1'h1)))
                    begin
                      reg4027 <= reg2894;
                    end
                end
              else
                begin
                  for (forvar4021 = (1'h0); (forvar4021 < (1'h0)); forvar4021 = (forvar4021 + (1'h1)))
                    begin
                      reg4022 <= (&$signed(reg3009[(1'h0):(1'h0)]));
                      reg4023 <= ((^forvar3010[(2'h2):(1'h1)]) + {$unsigned((~^reg3316))});
                      reg4024 <= $signed(reg3409[(1'h0):(1'h0)]);
                    end
                  reg4025 <= $unsigned($signed((~&{forvar3184})));
                end
            end
          else
            begin
              for (forvar4021 = (1'h0); (forvar4021 < (1'h1)); forvar4021 = (forvar4021 + (1'h1)))
                begin
                  if ((~^reg3200))
                    begin
                      reg4022 <= (($signed((~&reg2810)) ^~ wire1762[(1'h0):(1'h0)]) ^ (($signed(reg3124) ?
                          $unsigned(reg3377) : (forvar3232 ?
                              forvar3240 : reg2922)) * reg3444[(1'h0):(1'h0)]));
                      reg4023 <= reg3483[(3'h7):(3'h6)];
                      reg4024 <= {(8'hb3)};
                    end
                  else
                    begin
                      reg4022 <= (reg4024[(2'h2):(1'h1)] ?
                          ($unsigned((reg2827 ~^ reg3080)) | forvar3164[(3'h5):(3'h5)]) : $signed(forvar3095[(2'h3):(1'h0)]));
                      reg4023 <= ((~|{reg3009[(3'h5):(2'h2)]}) ?
                          reg3314[(3'h4):(3'h4)] : $unsigned(forvar2878[(2'h2):(2'h2)]));
                      reg4024 <= ((|$unsigned(reg2763)) ?
                          (($signed(reg2801) ?
                                  (forvar3265 - reg2895) : (reg2949 && reg2897)) ?
                              ($signed(forvar3491) ?
                                  (reg2869 ?
                                      reg2894 : reg3231) : {(8'hab)}) : forvar3365) : $signed(((forvar3045 ?
                                  forvar3348 : reg3073) ?
                              reg2755[(2'h3):(2'h2)] : (&forvar2754))));
                      reg4025 <= (^$signed(reg2988[(1'h0):(1'h0)]));
                    end
                end
              reg4026 <= (8'ha2);
              if ((-$unsigned($signed(reg3142))))
                begin
                  if (reg3412[(1'h0):(1'h0)])
                    begin
                      reg4027 <= (^~forvar3500);
                    end
                  else
                    begin
                      reg4027 <= forvar3275;
                      reg4028 <= (forvar2959 | forvar3457[(1'h0):(1'h0)]);
                    end
                  if ((reg3479[(1'h1):(1'h1)] ?
                      reg3478[(1'h1):(1'h1)] : reg2877))
                    begin
                      reg4029 <= forvar2799;
                      reg4030 <= ($signed(reg3109) * (($unsigned(forvar3285) ?
                              $unsigned(forvar3424) : (&(8'h9c))) ?
                          (reg3054 != (reg3188 ?
                              forvar3461 : (8'h9c))) : $signed($unsigned((8'hb1)))));
                      reg4031 <= reg2830[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg4029 <= forvar2944;
                      reg4030 <= reg3433;
                      reg4031 <= (!(reg3113[(2'h2):(1'h1)] ?
                          (^(reg3421 ?
                              (8'hb8) : reg2971)) : ($unsigned(reg3023) * (8'hb7))));
                    end
                  for (forvar4032 = (1'h0); (forvar4032 < (1'h1)); forvar4032 = (forvar4032 + (1'h1)))
                    begin
                      reg4033 <= reg3006;
                      reg4034 <= {reg3195[(1'h1):(1'h0)]};
                      reg4035 <= $signed(reg3021[(4'ha):(2'h3)]);
                      reg4036 <= $unsigned((($signed(reg2830) ?
                          (reg3333 == reg3097) : $signed(reg2888)) ~^ ((reg3342 ?
                          reg3404 : forvar3228) <= $unsigned((8'ha5)))));
                    end
                  for (forvar4037 = (1'h0); (forvar4037 < (2'h2)); forvar4037 = (forvar4037 + (1'h1)))
                    begin
                      reg4038 <= reg3433[(1'h1):(1'h1)];
                      reg4039 <= $signed(reg2860);
                    end
                end
              else
                begin
                  for (forvar4027 = (1'h0); (forvar4027 < (1'h1)); forvar4027 = (forvar4027 + (1'h1)))
                    begin
                      reg4028 <= (~&$unsigned(((^~reg3472) ?
                          $unsigned(reg2893) : $signed(forvar3492))));
                      reg4029 <= $unsigned((8'had));
                      reg4030 <= (~|reg2820[(3'h4):(1'h1)]);
                      reg4031 <= ($unsigned((((8'hb2) ? reg3373 : forvar3122) ?
                          (reg4035 >= reg3099) : reg2845[(2'h2):(1'h0)])) & $unsigned(($signed(reg3425) >> $signed(forvar3296))));
                    end
                  for (forvar4032 = (1'h0); (forvar4032 < (2'h3)); forvar4032 = (forvar4032 + (1'h1)))
                    begin
                      reg4033 <= reg4039;
                      reg4034 <= ((~&reg3092[(2'h2):(2'h2)]) ?
                          (~|(((8'ha8) ?
                              reg2854 : reg3338) | {forvar3344})) : ({reg3393[(3'h6):(1'h0)]} > $signed((~&reg2947))));
                      reg4035 <= reg3373;
                      reg4036 <= ({$signed($unsigned((8'h9c)))} >> ((+(~^reg2834)) >= (~^reg3487)));
                    end
                end
              reg4040 <= reg3372;
            end
          for (forvar4041 = (1'h0); (forvar4041 < (2'h2)); forvar4041 = (forvar4041 + (1'h1)))
            begin
              reg4042 <= (forvar3461[(2'h2):(1'h0)] - reg3418[(2'h2):(1'h1)]);
              reg4043 <= $unsigned((!reg3489));
              for (forvar4044 = (1'h0); (forvar4044 < (2'h3)); forvar4044 = (forvar4044 + (1'h1)))
                begin
                  for (forvar4045 = (1'h0); (forvar4045 < (1'h0)); forvar4045 = (forvar4045 + (1'h1)))
                    begin
                      reg4046 <= ($signed({forvar3274}) * $signed($unsigned(reg2888[(1'h1):(1'h1)])));
                      reg4047 <= $signed($signed(reg3338[(2'h3):(2'h3)]));
                      reg4048 <= ((reg3501[(1'h0):(1'h0)] & (~&$unsigned(reg2887))) << (((forvar3303 + (8'ha1)) ?
                              reg2840 : $unsigned(forvar2826)) ?
                          reg3083 : ((~^forvar3242) ? reg3038 : (8'hab))));
                      reg4049 <= (-$signed((^(reg3113 & (8'hb6)))));
                    end
                  reg4050 <= (^forvar3163[(4'h9):(1'h0)]);
                  reg4051 <= (((reg2884[(1'h1):(1'h0)] ?
                          (reg3204 ^ reg3055) : (8'ha0)) - ((~&reg3148) ?
                          (^forvar3365) : reg3386[(2'h2):(2'h2)])) ?
                      $signed(reg3018) : reg3298);
                end
            end
          for (forvar4052 = (1'h0); (forvar4052 < (1'h0)); forvar4052 = (forvar4052 + (1'h1)))
            begin
              for (forvar4053 = (1'h0); (forvar4053 < (2'h2)); forvar4053 = (forvar4053 + (1'h1)))
                begin
                  if ($signed($signed(($signed(forvar3240) >>> (~|forvar2931)))))
                    begin
                      reg4054 <= reg2967;
                      reg4055 <= reg3174;
                      reg4056 <= $signed($signed(reg3414[(2'h3):(1'h1)]));
                      reg4057 <= $signed($unsigned($unsigned((reg3252 >>> reg3423))));
                    end
                  else
                    begin
                      reg4054 <= reg2921;
                      reg4055 <= ((((reg2946 ? reg2955 : reg3499) ?
                                  (~&(8'haf)) : forvar3362) ?
                              forvar3009[(2'h2):(1'h0)] : (~^(reg3316 || reg4030))) ?
                          {$signed((~^reg2798))} : (-(~&$signed(reg3200))));
                      reg4056 <= {reg2915};
                    end
                end
              for (forvar4058 = (1'h0); (forvar4058 < (1'h1)); forvar4058 = (forvar4058 + (1'h1)))
                begin
                  if ({(reg3203[(2'h3):(2'h3)] ?
                          reg3160[(2'h2):(2'h2)] : {$signed(reg3442)})})
                    begin
                      reg4059 <= reg2988[(1'h1):(1'h0)];
                      reg4060 <= (forvar3187 ? forvar3254 : forvar3220);
                      reg4061 <= (^$signed(((reg3352 <= reg2961) == (reg2818 << reg2937))));
                    end
                  else
                    begin
                      reg4059 <= ($signed($unsigned($unsigned(reg3472))) ?
                          reg3473 : (((reg3251 ? (8'hb3) : forvar3011) ?
                                  (reg2806 ? reg2792 : forvar3139) : (reg3330 ?
                                      forvar2944 : forvar3271)) ?
                              (~|$unsigned(reg2906)) : (&(8'hb0))));
                      reg4060 <= (!reg3065[(1'h0):(1'h0)]);
                      reg4061 <= (~|reg2926[(1'h1):(1'h0)]);
                      reg4062 <= reg3244;
                    end
                  if ((($unsigned($unsigned((8'ha9))) << (forvar2797 ?
                          forvar3321[(1'h1):(1'h1)] : (reg3334 ?
                              forvar3350 : forvar2947))) ?
                      reg2845[(1'h0):(1'h0)] : ($signed(forvar3473) ?
                          $unsigned(forvar2899) : $signed((+reg3040)))))
                    begin
                      reg4063 <= ((&reg2758) <= $signed(reg3408[(1'h1):(1'h1)]));
                      reg4064 <= ((+(~&(reg2859 ?
                          reg3262 : reg2968))) >> (((forvar3275 != forvar3437) ?
                          (reg3319 ?
                              forvar2955 : reg2893) : forvar3087) < ((^(8'h9e)) | $unsigned(forvar3363))));
                      reg4065 <= reg3248;
                    end
                  else
                    begin
                      reg4063 <= $signed(reg3205[(3'h5):(3'h4)]);
                      reg4064 <= $signed(($unsigned((!forvar2955)) ?
                          (+$unsigned(reg3339)) : (~&{(8'ha5)})));
                      reg4065 <= $signed(reg3407[(1'h0):(1'h0)]);
                    end
                end
              if (forvar3404)
                begin
                  if ((reg3494 ?
                      (!{reg2922[(1'h1):(1'h0)]}) : forvar2959[(3'h7):(3'h4)]))
                    begin
                      reg4066 <= $unsigned((~^reg3291[(4'he):(4'he)]));
                      reg4067 <= (-reg2959[(1'h1):(1'h0)]);
                      reg4068 <= (~|{$unsigned($signed(reg3358))});
                      reg4069 <= $unsigned(((|reg2794) ?
                          {forvar3220} : $unsigned($signed(reg3181))));
                    end
                  else
                    begin
                      reg4066 <= ((^~reg3032) <= forvar3296[(3'h7):(1'h0)]);
                      reg4067 <= $unsigned(({$signed(forvar3007)} ?
                          (^~((8'haa) ~^ reg3377)) : $signed($signed(reg2766))));
                    end
                  if (reg3474)
                    begin
                      reg4070 <= (($signed($unsigned((8'haa))) ?
                          reg2784[(3'h6):(3'h6)] : ((+forvar2943) ?
                              (8'hb4) : (reg2862 ?
                                  reg2973 : forvar2968))) - reg3026[(4'h9):(1'h1)]);
                      reg4071 <= $unsigned(($unsigned({forvar3426}) ?
                          {(reg3368 ?
                                  (8'hba) : (8'hb3))} : reg3146[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg4070 <= ((^(reg2969[(1'h0):(1'h0)] << $signed((8'h9d)))) + ($unsigned((-(8'had))) ~^ (+$signed(reg3073))));
                      reg4071 <= (~&(forvar3255 >> reg4055));
                      reg4072 <= (!$signed($signed($signed(reg3307))));
                      reg4073 <= reg3287[(3'h6):(3'h5)];
                    end
                end
              else
                begin
                  if ($unsigned(((^~(~reg3391)) < $unsigned((&forvar4026)))))
                    begin
                      reg4066 <= reg2900[(3'h4):(3'h4)];
                      reg4067 <= ((^reg2802[(1'h1):(1'h1)]) ^ ((~|(reg3354 ?
                              reg2785 : reg2922)) ?
                          $unsigned((~^forvar3266)) : ($signed(reg3169) ?
                              (8'hab) : (reg3117 ? reg3225 : reg2824))));
                      reg4068 <= ($signed(forvar3006) ?
                          $signed(((8'hb3) ?
                              (~&reg2773) : $signed(reg3020))) : forvar4037);
                      reg4069 <= reg2803;
                    end
                  else
                    begin
                      reg4066 <= ($unsigned(((~|reg3238) || {reg3421})) > reg3370);
                      reg4067 <= forvar3151;
                    end
                  if ($signed((-$unsigned(reg4064))))
                    begin
                      reg4070 <= ((8'hb1) ?
                          $signed(forvar3165) : $signed(reg3401));
                    end
                  else
                    begin
                      reg4070 <= ((~^$signed($signed((8'hb2)))) <<< forvar4020);
                      reg4071 <= $unsigned($signed((-reg3173[(1'h0):(1'h0)])));
                    end
                  if ($signed({$signed(reg3269[(2'h2):(1'h1)])}))
                    begin
                      reg4072 <= (~($signed($signed(forvar3130)) ?
                          $signed($signed(reg4068)) : reg3408));
                      reg4073 <= $unsigned($signed((reg3132 <<< {(8'hb5)})));
                    end
                  else
                    begin
                      reg4072 <= (reg2851 & forvar3453);
                    end
                  for (forvar4074 = (1'h0); (forvar4074 < (2'h3)); forvar4074 = (forvar4074 + (1'h1)))
                    begin
                      reg4075 <= $unsigned(forvar2902);
                      reg4076 <= ((((~^reg3245) < (reg3435 >= (8'ha4))) && $unsigned($unsigned(reg4064))) ?
                          ((~|reg3173) ?
                              (^~reg3418[(2'h2):(1'h1)]) : ($signed(reg3415) ?
                                  (reg3129 ?
                                      reg2926 : (8'hb4)) : (reg3095 || forvar2964))) : $unsigned((reg3328[(2'h3):(2'h2)] - reg3320)));
                      reg4077 <= ((|$signed((&reg3360))) ?
                          $unsigned($signed(reg3071)) : $unsigned(reg3415[(3'h4):(2'h3)]));
                    end
                end
              if (reg2827[(1'h0):(1'h0)])
                begin
                  for (forvar4078 = (1'h0); (forvar4078 < (2'h3)); forvar4078 = (forvar4078 + (1'h1)))
                    begin
                      reg4079 <= (reg3309[(3'h5):(1'h1)] ?
                          $unsigned(reg3055[(2'h3):(1'h0)]) : (-$signed(reg3261[(1'h1):(1'h0)])));
                      reg4080 <= (^$signed(((forvar4045 >> reg3487) & $unsigned(forvar3095))));
                      reg4081 <= (~|(forvar3356[(1'h1):(1'h0)] ?
                          (|$unsigned(reg2973)) : (~|{reg3256})));
                    end
                  for (forvar4082 = (1'h0); (forvar4082 < (2'h3)); forvar4082 = (forvar4082 + (1'h1)))
                    begin
                      reg4083 <= (|$unsigned(reg3096));
                      reg4084 <= reg3020;
                    end
                  reg4085 <= (forvar3163 ^ forvar2969[(1'h0):(1'h0)]);
                  for (forvar4086 = (1'h0); (forvar4086 < (1'h1)); forvar4086 = (forvar4086 + (1'h1)))
                    begin
                      reg4087 <= reg2763;
                      reg4088 <= (forvar2826 ? {reg3444} : $signed(reg2948));
                      reg4089 <= $signed((~^$unsigned((!(8'ha6)))));
                    end
                end
              else
                begin
                  if (reg3420)
                    begin
                      reg4078 <= reg3211[(3'h4):(3'h4)];
                      reg4079 <= (~|((forvar3143 >>> {reg2904}) ^~ forvar3157[(3'h7):(2'h3)]));
                      reg4080 <= $unsigned({$signed((reg3169 ?
                              reg3020 : reg2991))});
                      reg4081 <= ((forvar3325 ?
                          $unsigned((reg3138 ?
                              (8'h9f) : forvar4021)) : $signed((~&(8'hb9)))) ~^ (|reg2906));
                    end
                  else
                    begin
                      reg4078 <= $unsigned($unsigned($unsigned((~|forvar3056))));
                      reg4079 <= (~|reg3131);
                      reg4080 <= reg3161[(2'h2):(2'h2)];
                    end
                  reg4082 <= reg3147[(2'h2):(1'h0)];
                  reg4083 <= (8'ha5);
                  for (forvar4084 = (1'h0); (forvar4084 < (1'h0)); forvar4084 = (forvar4084 + (1'h1)))
                    begin
                      reg4085 <= (reg4024 ?
                          ((8'ha7) || ((-forvar2920) ?
                              $unsigned(reg2792) : forvar3029[(1'h1):(1'h0)])) : $unsigned($unsigned(reg4078[(4'hb):(1'h1)])));
                      reg4086 <= {reg3120[(1'h1):(1'h0)]};
                      reg4087 <= ((+(forvar3007[(1'h1):(1'h0)] + $unsigned(reg2755))) << forvar3284);
                      reg4088 <= $unsigned(($unsigned({forvar3213}) ?
                          $signed(reg3277) : ({reg3452} * {reg2795})));
                    end
                end
            end
          if ((($unsigned((reg2863 ? reg4061 : forvar2862)) ?
              $signed(((8'ha5) ?
                  forvar3426 : reg2846)) : reg3355[(1'h0):(1'h0)]) ^ ((|(|reg3016)) >>> ($signed(reg4086) ?
              (reg3079 ? wire2753 : reg3149) : reg3176))))
            begin
              if ((8'hb1))
                begin
                  reg4090 <= $unsigned(reg3198);
                end
              else
                begin
                  if ((($unsigned((reg2966 ? reg3173 : forvar2866)) ?
                          forvar4021 : $signed({reg2951})) ?
                      $signed($unsigned(reg2980)) : reg2977))
                    begin
                      reg4090 <= reg2842[(1'h1):(1'h1)];
                      reg4091 <= $unsigned(($signed({reg3400}) == reg3366));
                      reg4092 <= reg3190;
                    end
                  else
                    begin
                      reg4090 <= (~$signed(reg3067));
                      reg4091 <= {$signed($signed(reg3459))};
                      reg4092 <= (reg3048 <<< (reg4047 ?
                          $unsigned($unsigned(reg2867)) : (|(-reg3185))));
                    end
                  for (forvar4093 = (1'h0); (forvar4093 < (2'h3)); forvar4093 = (forvar4093 + (1'h1)))
                    begin
                      reg4094 <= (^$unsigned($signed(forvar3215[(3'h7):(2'h3)])));
                      reg4095 <= $signed($signed({{forvar3203}}));
                      reg4096 <= reg4086;
                      reg4097 <= reg3147[(3'h4):(2'h2)];
                    end
                end
              for (forvar4098 = (1'h0); (forvar4098 < (1'h1)); forvar4098 = (forvar4098 + (1'h1)))
                begin
                  if (reg2973)
                    begin
                      reg4099 <= forvar3332[(3'h6):(1'h0)];
                      reg4100 <= (~&forvar2797[(3'h5):(2'h2)]);
                      reg4101 <= forvar3365;
                      reg4102 <= ($unsigned(({reg3185} ?
                              (!forvar3231) : $signed(reg3091))) ?
                          (8'ha8) : (~|($signed(reg3251) ?
                              forvar2944[(4'hc):(3'h5)] : (reg2865 ?
                                  forvar3426 : forvar3114))));
                    end
                  else
                    begin
                      reg4099 <= ((8'had) != $unsigned($signed((reg3368 > forvar3103))));
                      reg4100 <= (~&$signed(reg3208));
                      reg4101 <= (reg2889[(4'hb):(1'h1)] || reg3143);
                      reg4102 <= $signed($unsigned(({reg3403} ^ {reg4056})));
                    end
                end
              if (($unsigned(forvar2978) ?
                  {(~|reg2875[(2'h3):(1'h0)])} : ($signed(((8'hb0) ?
                      forvar3260 : reg3464)) != ({forvar2948} ?
                      (~^reg4100) : (reg3067 ? reg3443 : forvar3288)))))
                begin
                  for (forvar4103 = (1'h0); (forvar4103 < (2'h3)); forvar4103 = (forvar4103 + (1'h1)))
                    begin
                      reg4104 <= reg2904[(1'h0):(1'h0)];
                      reg4105 <= forvar2866;
                      reg4106 <= (reg3396 && (&(reg4033[(2'h3):(1'h1)] != $unsigned((8'hae)))));
                    end
                  for (forvar4107 = (1'h0); (forvar4107 < (2'h3)); forvar4107 = (forvar4107 + (1'h1)))
                    begin
                      reg4108 <= (reg4050[(3'h7):(3'h6)] ?
                          ({(reg3192 <= (8'ha5))} >>> $signed((reg2835 ?
                              reg2913 : reg2951))) : $unsigned((forvar3247 ?
                              $signed(reg4042) : (reg3485 ?
                                  reg3172 : forvar3346))));
                      reg4109 <= forvar2958;
                    end
                end
              else
                begin
                  reg4103 <= {(~|((^reg2860) ^ {reg3096}))};
                end
            end
          else
            begin
              for (forvar4090 = (1'h0); (forvar4090 < (2'h2)); forvar4090 = (forvar4090 + (1'h1)))
                begin
                  if ((reg4049 && reg2874[(3'h5):(1'h0)]))
                    begin
                      reg4091 <= reg2955[(3'h5):(1'h1)];
                      reg4092 <= reg3408[(1'h1):(1'h1)];
                      reg4093 <= (^~forvar2878);
                      reg4094 <= (~reg3412);
                    end
                  else
                    begin
                      reg4091 <= ((^({forvar3006} & (~^reg2976))) ?
                          {(^(^~reg4054))} : (~|(((8'hab) || reg2974) > reg2839[(2'h3):(2'h2)])));
                    end
                  if ((reg3228[(3'h6):(2'h3)] ?
                      (((forvar3151 & (8'h9f)) ?
                          ((8'hab) - reg3244) : $signed(reg2879)) <<< reg4069) : (-(!(~^reg3154)))))
                    begin
                      reg4095 <= forvar3453;
                      reg4096 <= (|{$unsigned({(8'hb5)})});
                      reg4097 <= (|reg3148);
                    end
                  else
                    begin
                      reg4095 <= reg3251;
                      reg4096 <= (forvar2993 ? forvar3441 : reg2947);
                      reg4097 <= $unsigned({(8'h9c)});
                      reg4098 <= $signed($unsigned(forvar3108[(4'hc):(4'hb)]));
                    end
                end
              reg4099 <= $signed(reg2913);
            end
        end
      for (forvar4110 = (1'h0); (forvar4110 < (1'h0)); forvar4110 = (forvar4110 + (1'h1)))
        begin
          for (forvar4111 = (1'h0); (forvar4111 < (1'h0)); forvar4111 = (forvar4111 + (1'h1)))
            begin
              reg4112 <= $signed($unsigned(((reg3110 ?
                  reg3338 : (8'haf)) ~^ (reg3084 >>> reg3430))));
              if ($signed(reg2872[(2'h2):(1'h1)]))
                begin
                  for (forvar4113 = (1'h0); (forvar4113 < (1'h0)); forvar4113 = (forvar4113 + (1'h1)))
                    begin
                      reg4114 <= {(reg3229[(2'h3):(1'h1)] ?
                              (~|$signed(reg3088)) : (-(forvar2919 ?
                                  reg2772 : reg2945)))};
                      reg4115 <= (forvar2776 ?
                          (forvar3427[(3'h5):(1'h0)] ?
                              (reg4102 ?
                                  (-reg2906) : $signed(reg3477)) : (forvar3394[(3'h5):(2'h2)] >= reg2798[(3'h5):(3'h5)])) : (~&$unsigned(forvar4110)));
                      reg4116 <= $unsigned((!(~forvar3367[(3'h6):(3'h4)])));
                    end
                end
              else
                begin
                  for (forvar4113 = (1'h0); (forvar4113 < (1'h1)); forvar4113 = (forvar4113 + (1'h1)))
                    begin
                      reg4114 <= ((($signed(reg3139) ?
                              reg4112[(2'h3):(1'h1)] : reg3358[(4'he):(4'h9)]) ?
                          reg3084 : {$unsigned(reg2860)}) && forvar4086);
                      reg4115 <= wire1761[(4'hc):(4'hc)];
                    end
                  for (forvar4116 = (1'h0); (forvar4116 < (1'h0)); forvar4116 = (forvar4116 + (1'h1)))
                    begin
                      reg4117 <= (8'hb9);
                      reg4118 <= (^~$unsigned($signed(forvar3408)));
                      reg4119 <= ((~&($unsigned(reg3209) && reg3142[(2'h3):(2'h3)])) ?
                          $unsigned(($signed(reg2847) ?
                              (~|reg3294) : forvar3143)) : forvar3007);
                      reg4120 <= $signed($signed(((reg4087 ?
                              forvar2849 : (8'hab)) ?
                          (reg3281 ? reg3236 : reg3216) : reg3499)));
                    end
                end
            end
          reg4121 <= reg3119;
          if (($unsigned(reg2852) ?
              {{(!reg2940)}} : $unsigned(reg3361[(1'h1):(1'h1)])))
            begin
              for (forvar4122 = (1'h0); (forvar4122 < (2'h3)); forvar4122 = (forvar4122 + (1'h1)))
                begin
                  for (forvar4123 = (1'h0); (forvar4123 < (2'h3)); forvar4123 = (forvar4123 + (1'h1)))
                    begin
                      reg4124 <= (^(8'hb7));
                      reg4125 <= ((reg2991[(4'hc):(4'hb)] <= $unsigned(reg3019[(3'h4):(3'h4)])) >>> {(~|(reg3405 ?
                              reg3158 : forvar3210))});
                      reg4126 <= (((^~reg3145) ?
                          $signed((&forvar3090)) : $signed((~&reg3044))) ^ reg3334);
                    end
                  reg4127 <= (reg4099[(4'h9):(1'h0)] ?
                      $signed(((|(8'hb9)) ?
                          {reg3438} : (~reg3380))) : $signed(((~|reg3273) - reg3463[(4'h9):(3'h7)])));
                end
              if (($unsigned($unsigned((reg2980 >>> reg3320))) == $unsigned(reg3487[(4'h9):(2'h2)])))
                begin
                  for (forvar4128 = (1'h0); (forvar4128 < (2'h3)); forvar4128 = (forvar4128 + (1'h1)))
                    begin
                      reg4129 <= reg3421;
                      reg4130 <= ((~&$signed((&(8'hb7)))) ^~ $unsigned($signed((reg2904 ?
                          (8'h9e) : reg4023))));
                    end
                end
              else
                begin
                  reg4128 <= (!{forvar3186[(1'h0):(1'h0)]});
                  if (wire4019[(3'h5):(3'h4)])
                    begin
                      reg4129 <= ($unsigned((~&(~|(8'haa)))) <= (reg3411[(2'h2):(1'h0)] * (wire4019 ?
                          forvar3047 : reg2959[(2'h2):(1'h0)])));
                      reg4130 <= reg3349[(2'h3):(2'h2)];
                      reg4131 <= reg3193[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4129 <= (&reg3407);
                    end
                end
              reg4132 <= reg3289;
            end
          else
            begin
              reg4122 <= {$unsigned(forvar3416[(3'h4):(1'h0)])};
            end
          for (forvar4133 = (1'h0); (forvar4133 < (1'h0)); forvar4133 = (forvar4133 + (1'h1)))
            begin
              for (forvar4134 = (1'h0); (forvar4134 < (2'h3)); forvar4134 = (forvar4134 + (1'h1)))
                begin
                  if ($unsigned(reg2851))
                    begin
                      reg4135 <= $unsigned(reg3161);
                      reg4136 <= $unsigned(reg3241[(1'h0):(1'h0)]);
                      reg4137 <= $signed($signed(reg3119));
                    end
                  else
                    begin
                      reg4135 <= {($signed((reg3376 ^ reg4137)) - ((forvar4111 ?
                              reg2965 : reg2787) < $signed(reg4083)))};
                    end
                  if ($unsigned((((reg3110 & forvar3139) ^ $signed(wire4019)) < $signed((+forvar2969)))))
                    begin
                      reg4138 <= ((~$signed((reg3176 ? wire1762 : reg3150))) ?
                          (reg4127 ?
                              reg2952[(3'h5):(3'h5)] : ((forvar2778 >> reg3387) ?
                                  (^reg3487) : (forvar2948 | (8'haf)))) : (&($unsigned(forvar3215) || $unsigned(reg4076))));
                      reg4139 <= $unsigned($unsigned(($unsigned(reg3170) ?
                          reg2962[(1'h0):(1'h0)] : $unsigned(reg3461))));
                      reg4140 <= $unsigned((~&$unsigned(wire3182[(3'h6):(2'h3)])));
                      reg4141 <= {$unsigned($signed($signed(reg3081)))};
                    end
                  else
                    begin
                      reg4138 <= $unsigned((-$signed($unsigned(reg3021))));
                      reg4139 <= forvar3453;
                      reg4140 <= ($unsigned($unsigned(reg2766)) ?
                          ((~^(reg2952 > (8'hb1))) ?
                              (8'haa) : (reg3104[(1'h1):(1'h0)] ?
                                  wire4019[(2'h3):(1'h0)] : $signed(reg3189))) : $unsigned($signed($unsigned(reg3063))));
                      reg4141 <= (reg3030[(2'h2):(1'h0)] <= $signed(((reg4025 ?
                          reg2831 : (8'hb7)) && $signed(forvar3265))));
                    end
                  if ((8'hb9))
                    begin
                      reg4142 <= reg2780;
                      reg4143 <= (($signed($unsigned(reg3214)) ?
                              forvar2777[(2'h3):(2'h3)] : reg2977) ?
                          ($unsigned(reg3446[(1'h0):(1'h0)]) || $signed($unsigned((8'hba)))) : (8'h9f));
                    end
                  else
                    begin
                      reg4142 <= (~|reg4049);
                    end
                end
              for (forvar4144 = (1'h0); (forvar4144 < (1'h1)); forvar4144 = (forvar4144 + (1'h1)))
                begin
                  if ($unsigned(($signed($unsigned((8'haf))) >= (reg3248 ?
                      reg3360 : forvar3426[(1'h1):(1'h1)]))))
                    begin
                      reg4145 <= {{((8'hb3) & {reg3433})}};
                      reg4146 <= $unsigned({forvar3365});
                    end
                  else
                    begin
                      reg4145 <= (($signed((forvar3473 ?
                          reg3068 : forvar3122)) * {(&reg3387)}) ^ {(^~((8'ha7) && reg2843))});
                      reg4146 <= $unsigned(reg3476[(1'h1):(1'h0)]);
                      reg4147 <= (({(reg2775 >>> reg3132)} ?
                          {reg2815[(4'hb):(3'h7)]} : (^$signed((8'hba)))) > (((reg2967 ?
                              reg3044 : (8'ha1)) != reg3362) ?
                          reg3023 : reg4097));
                    end
                  reg4148 <= (~&(~|reg4106[(4'h8):(4'h8)]));
                  for (forvar4149 = (1'h0); (forvar4149 < (1'h0)); forvar4149 = (forvar4149 + (1'h1)))
                    begin
                      reg4150 <= (^$signed(reg4056[(3'h6):(2'h2)]));
                      reg4151 <= ($signed(reg4112[(2'h2):(2'h2)]) ?
                          $unsigned((reg2841 ?
                              (8'hb0) : $signed((8'hb1)))) : (wire2749 ?
                              forvar3297 : reg3033[(2'h2):(2'h2)]));
                    end
                end
              if ((!(forvar3361 >>> reg3436)))
                begin
                  for (forvar4152 = (1'h0); (forvar4152 < (2'h2)); forvar4152 = (forvar4152 + (1'h1)))
                    begin
                      reg4153 <= (-(reg4073[(2'h2):(1'h0)] ?
                          (reg4085[(1'h0):(1'h0)] ?
                              reg2954[(1'h1):(1'h0)] : $unsigned(reg4129)) : ((8'haa) || $unsigned(reg3399))));
                      reg4154 <= forvar3491;
                      reg4155 <= $unsigned({(8'ha0)});
                    end
                  for (forvar4156 = (1'h0); (forvar4156 < (1'h1)); forvar4156 = (forvar4156 + (1'h1)))
                    begin
                      reg4157 <= (+((~reg2820) ?
                          reg3180 : {$unsigned(reg4137)}));
                    end
                  reg4158 <= $signed($signed(reg3053));
                  if ($unsigned($unsigned(reg2928[(2'h3):(2'h3)])))
                    begin
                      reg4159 <= forvar2931[(3'h5):(1'h0)];
                    end
                  else
                    begin
                      reg4159 <= $unsigned($signed(($signed(reg3338) ?
                          $unsigned(reg4114) : reg2938[(3'h5):(3'h4)])));
                      reg4160 <= (8'hb0);
                      reg4161 <= $signed({((reg3316 ?
                              forvar3453 : reg2970) & {(8'h9f)})});
                      reg4162 <= $signed($unsigned($signed((forvar3139 ?
                          reg2763 : forvar2963))));
                    end
                end
              else
                begin
                  if ($signed($signed($signed({reg3370}))))
                    begin
                      reg4152 <= (~&(8'hb7));
                      reg4153 <= $unsigned($signed({$unsigned(reg3009)}));
                    end
                  else
                    begin
                      reg4152 <= (^{$unsigned($unsigned(reg3385))});
                      reg4153 <= $unsigned(reg3239[(1'h1):(1'h0)]);
                    end
                  for (forvar4154 = (1'h0); (forvar4154 < (1'h0)); forvar4154 = (forvar4154 + (1'h1)))
                    begin
                      reg4155 <= reg4086[(3'h6):(3'h5)];
                      reg4156 <= $unsigned(($signed($signed(forvar4107)) ?
                          reg4031[(2'h3):(2'h3)] : $signed($unsigned(forvar2781))));
                      reg4157 <= (8'h9f);
                      reg4158 <= ($unsigned($signed((reg4061 == reg3294))) != reg3410[(1'h0):(1'h0)]);
                    end
                end
              reg4163 <= $signed((reg3263 && (((8'hb8) ~^ forvar2964) ?
                  $unsigned((8'had)) : (reg3218 > forvar2829))));
            end
        end
    end
  assign wire4164 = reg4073;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1219  (y, clk, wire1224, wire1223, wire1222, wire1221, wire1220);
  output wire [(32'h14c7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire1224;
  input wire [(4'hc):(1'h0)] wire1223;
  input wire signed [(3'h6):(1'h0)] wire1222;
  input wire signed [(4'he):(1'h0)] wire1221;
  input wire [(2'h3):(1'h0)] wire1220;
  wire [(3'h4):(1'h0)] wire1743;
  reg signed [(2'h2):(1'h0)] reg1742 = (1'h0);
  reg [(4'hf):(1'h0)] reg1720 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1717 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1716 = (1'h0);
  reg [(3'h5):(1'h0)] reg1715 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1741 = (1'h0);
  reg [(4'h9):(1'h0)] reg1739 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1738 = (1'h0);
  reg [(3'h7):(1'h0)] reg1734 = (1'h0);
  reg [(3'h6):(1'h0)] reg1740 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1739 = (1'h0);
  reg [(4'h8):(1'h0)] reg1738 = (1'h0);
  reg [(3'h7):(1'h0)] reg1737 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1736 = (1'h0);
  reg [(2'h2):(1'h0)] reg1735 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1734 = (1'h0);
  reg [(3'h4):(1'h0)] reg1731 = (1'h0);
  reg [(4'hf):(1'h0)] reg1728 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1724 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1733 = (1'h0);
  reg [(4'hd):(1'h0)] reg1732 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1731 = (1'h0);
  reg [(5'h10):(1'h0)] reg1730 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1729 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1728 = (1'h0);
  reg [(3'h7):(1'h0)] reg1727 = (1'h0);
  reg [(3'h6):(1'h0)] reg1726 = (1'h0);
  reg [(4'hc):(1'h0)] reg1725 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1724 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1723 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1722 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1721 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1720 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1719 = (1'h0);
  reg [(3'h7):(1'h0)] reg1718 = (1'h0);
  reg [(4'hc):(1'h0)] reg1717 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1716 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1715 = (1'h0);
  reg [(4'hb):(1'h0)] reg1714 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1713 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1712 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1711 = (1'h0);
  reg [(3'h7):(1'h0)] reg1710 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1709 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1708 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1707 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1706 = (1'h0);
  reg [(3'h4):(1'h0)] reg1705 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1704 = (1'h0);
  reg [(5'h10):(1'h0)] reg1703 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1702 = (1'h0);
  reg [(3'h5):(1'h0)] reg1701 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1700 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1699 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1697 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1698 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1697 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1696 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1695 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1694 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1693 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1692 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1691 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1690 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1689 = (1'h0);
  wire [(3'h6):(1'h0)] wire1688;
  reg signed [(3'h4):(1'h0)] reg1618 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1687 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1686 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1685 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1684 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1683 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1682 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1681 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1680 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1679 = (1'h0);
  reg [(4'ha):(1'h0)] reg1678 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1677 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1676 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1675 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1674 = (1'h0);
  reg [(4'he):(1'h0)] reg1673 = (1'h0);
  reg [(4'ha):(1'h0)] reg1672 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1671 = (1'h0);
  reg [(3'h6):(1'h0)] reg1670 = (1'h0);
  reg [(2'h2):(1'h0)] reg1657 = (1'h0);
  reg [(4'h8):(1'h0)] reg1669 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1668 = (1'h0);
  reg [(4'hd):(1'h0)] reg1667 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1666 = (1'h0);
  reg [(2'h2):(1'h0)] reg1665 = (1'h0);
  reg [(3'h5):(1'h0)] reg1664 = (1'h0);
  reg [(3'h6):(1'h0)] reg1663 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1662 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1661 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1660 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1659 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1658 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1657 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1656 = (1'h0);
  reg [(3'h7):(1'h0)] reg1655 = (1'h0);
  reg [(2'h3):(1'h0)] reg1654 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1653 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1652 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1651 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1650 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1649 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1648 = (1'h0);
  reg [(4'hd):(1'h0)] reg1647 = (1'h0);
  reg [(4'ha):(1'h0)] reg1646 = (1'h0);
  reg [(4'hb):(1'h0)] reg1645 = (1'h0);
  reg [(4'hb):(1'h0)] reg1644 = (1'h0);
  reg [(4'hb):(1'h0)] reg1643 = (1'h0);
  reg [(5'h10):(1'h0)] reg1642 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1641 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1640 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1639 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1637 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1638 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1637 = (1'h0);
  reg [(3'h7):(1'h0)] reg1636 = (1'h0);
  reg [(4'ha):(1'h0)] reg1635 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1634 = (1'h0);
  reg [(3'h4):(1'h0)] reg1633 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1632 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1631 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1630 = (1'h0);
  reg [(2'h3):(1'h0)] reg1629 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1628 = (1'h0);
  reg [(4'h8):(1'h0)] reg1627 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1626 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1625 = (1'h0);
  reg [(5'h10):(1'h0)] reg1624 = (1'h0);
  reg [(4'hc):(1'h0)] reg1623 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1622 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1621 = (1'h0);
  reg [(4'he):(1'h0)] forvar1620 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1619 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1618 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1601 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1599 = (1'h0);
  reg [(4'h9):(1'h0)] reg1617 = (1'h0);
  reg [(4'he):(1'h0)] reg1616 = (1'h0);
  reg [(2'h2):(1'h0)] reg1615 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1614 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1613 = (1'h0);
  reg [(2'h2):(1'h0)] reg1612 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1611 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1610 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1609 = (1'h0);
  reg [(3'h4):(1'h0)] reg1608 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1607 = (1'h0);
  reg [(2'h2):(1'h0)] reg1606 = (1'h0);
  reg [(4'hc):(1'h0)] reg1605 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1604 = (1'h0);
  reg [(5'h10):(1'h0)] reg1603 = (1'h0);
  reg [(2'h2):(1'h0)] reg1602 = (1'h0);
  reg [(4'he):(1'h0)] forvar1601 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1600 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1599 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1598 = (1'h0);
  reg [(3'h7):(1'h0)] reg1597 = (1'h0);
  wire [(4'h9):(1'h0)] wire1596;
  wire [(4'he):(1'h0)] wire1595;
  reg [(4'hc):(1'h0)] reg1594 = (1'h0);
  reg [(4'hf):(1'h0)] reg1593 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1592 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1591 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1590 = (1'h0);
  reg [(3'h4):(1'h0)] reg1589 = (1'h0);
  reg [(4'hc):(1'h0)] reg1588 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1587 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1586 = (1'h0);
  reg [(2'h2):(1'h0)] reg1585 = (1'h0);
  reg [(2'h2):(1'h0)] reg1584 = (1'h0);
  reg [(4'hd):(1'h0)] reg1583 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1582 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1581 = (1'h0);
  reg [(2'h2):(1'h0)] reg1580 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1579 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1578 = (1'h0);
  reg [(4'hc):(1'h0)] reg1577 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1576 = (1'h0);
  reg [(4'he):(1'h0)] reg1575 = (1'h0);
  reg [(4'hf):(1'h0)] reg1574 = (1'h0);
  reg [(4'hd):(1'h0)] reg1573 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1572 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1571 = (1'h0);
  reg [(4'ha):(1'h0)] reg1570 = (1'h0);
  reg [(4'ha):(1'h0)] reg1569 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1568 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1567 = (1'h0);
  reg [(4'hf):(1'h0)] reg1566 = (1'h0);
  reg [(4'hc):(1'h0)] reg1565 = (1'h0);
  reg [(4'ha):(1'h0)] reg1564 = (1'h0);
  reg [(4'hd):(1'h0)] reg1563 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1557 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1554 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1549 = (1'h0);
  reg [(4'hc):(1'h0)] reg1547 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1542 = (1'h0);
  reg [(4'h8):(1'h0)] reg1562 = (1'h0);
  reg [(2'h2):(1'h0)] reg1561 = (1'h0);
  reg [(4'ha):(1'h0)] reg1560 = (1'h0);
  reg [(3'h6):(1'h0)] reg1559 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1558 = (1'h0);
  reg [(3'h6):(1'h0)] reg1557 = (1'h0);
  reg [(3'h6):(1'h0)] reg1556 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1555 = (1'h0);
  reg [(3'h7):(1'h0)] reg1554 = (1'h0);
  reg [(4'h8):(1'h0)] reg1553 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1550 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1552 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1551 = (1'h0);
  reg [(4'h9):(1'h0)] reg1550 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1549 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1548 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1547 = (1'h0);
  reg [(2'h2):(1'h0)] reg1546 = (1'h0);
  reg [(3'h7):(1'h0)] reg1545 = (1'h0);
  reg [(5'h10):(1'h0)] reg1544 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1543 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1542 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1541 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1540 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1507 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1506 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1539 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1538 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1537 = (1'h0);
  reg [(4'hd):(1'h0)] reg1536 = (1'h0);
  reg [(3'h4):(1'h0)] reg1529 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1535 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1534 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1533 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1532 = (1'h0);
  reg [(3'h6):(1'h0)] reg1531 = (1'h0);
  reg [(3'h5):(1'h0)] reg1530 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1529 = (1'h0);
  reg [(3'h4):(1'h0)] reg1528 = (1'h0);
  reg [(3'h5):(1'h0)] reg1527 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1526 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1525 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1524 = (1'h0);
  reg [(3'h6):(1'h0)] reg1523 = (1'h0);
  reg [(3'h4):(1'h0)] reg1521 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1520 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1519 = (1'h0);
  reg [(3'h6):(1'h0)] reg1522 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1521 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1520 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1519 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1518 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1517 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1516 = (1'h0);
  reg [(3'h5):(1'h0)] reg1515 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1514 = (1'h0);
  reg [(4'hb):(1'h0)] reg1513 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1509 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1508 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1512 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1511 = (1'h0);
  reg [(4'hf):(1'h0)] reg1510 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1509 = (1'h0);
  reg [(4'h8):(1'h0)] reg1508 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1507 = (1'h0);
  reg [(3'h7):(1'h0)] reg1506 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1505 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1497 = (1'h0);
  reg [(3'h6):(1'h0)] reg1504 = (1'h0);
  reg [(4'he):(1'h0)] reg1503 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1502 = (1'h0);
  reg [(2'h3):(1'h0)] reg1501 = (1'h0);
  reg [(2'h3):(1'h0)] reg1500 = (1'h0);
  reg [(3'h6):(1'h0)] reg1496 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1493 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1489 = (1'h0);
  reg [(4'h8):(1'h0)] reg1490 = (1'h0);
  reg [(2'h2):(1'h0)] reg1499 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1498 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1497 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1496 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1495 = (1'h0);
  reg [(4'h8):(1'h0)] reg1494 = (1'h0);
  reg [(4'he):(1'h0)] reg1493 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1492 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1491 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1490 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1489 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1488 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1487 = (1'h0);
  reg [(4'hd):(1'h0)] reg1486 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1485 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1484 = (1'h0);
  reg [(4'he):(1'h0)] reg1483 = (1'h0);
  reg [(2'h2):(1'h0)] reg1482 = (1'h0);
  reg [(3'h6):(1'h0)] reg1481 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1480 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1479 = (1'h0);
  reg [(4'hc):(1'h0)] reg1478 = (1'h0);
  reg [(4'ha):(1'h0)] reg1477 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1476 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1475 = (1'h0);
  reg [(4'h9):(1'h0)] reg1474 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1473 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1472 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1471 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1470 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1469 = (1'h0);
  reg [(4'hd):(1'h0)] reg1468 = (1'h0);
  reg [(2'h2):(1'h0)] reg1467 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1466 = (1'h0);
  reg [(3'h7):(1'h0)] reg1465 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1464 = (1'h0);
  reg [(4'hb):(1'h0)] reg1463 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1462 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1461 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1460 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1459 = (1'h0);
  reg [(4'h9):(1'h0)] reg1458 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1453 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1457 = (1'h0);
  reg [(3'h6):(1'h0)] reg1456 = (1'h0);
  reg [(4'hf):(1'h0)] reg1455 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1454 = (1'h0);
  reg [(4'ha):(1'h0)] reg1453 = (1'h0);
  reg [(4'hd):(1'h0)] reg1444 = (1'h0);
  reg [(4'hb):(1'h0)] reg1452 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1451 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1450 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1449 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1448 = (1'h0);
  reg [(5'h10):(1'h0)] reg1447 = (1'h0);
  reg [(5'h10):(1'h0)] reg1446 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1445 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1444 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1443 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1442 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1441 = (1'h0);
  reg [(4'h8):(1'h0)] reg1440 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1439 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1408 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1411 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1394 = (1'h0);
  reg [(4'he):(1'h0)] forvar1391 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1414 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1410 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1409 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1405 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1404 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1397 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1402 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1401 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1398 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1395 = (1'h0);
  reg [(4'ha):(1'h0)] reg1392 = (1'h0);
  reg [(4'h9):(1'h0)] reg1383 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1436 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1434 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1438 = (1'h0);
  reg [(4'h8):(1'h0)] reg1437 = (1'h0);
  reg [(4'hb):(1'h0)] reg1436 = (1'h0);
  reg [(5'h10):(1'h0)] reg1435 = (1'h0);
  reg [(5'h10):(1'h0)] reg1434 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1433 = (1'h0);
  reg [(4'he):(1'h0)] reg1432 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1431 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1430 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1429 = (1'h0);
  reg [(3'h5):(1'h0)] reg1428 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1427 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1426 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1425 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1424 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1423 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1422 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1421 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1420 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1419 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1418 = (1'h0);
  reg [(2'h2):(1'h0)] reg1417 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1416 = (1'h0);
  reg [(4'ha):(1'h0)] reg1415 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1414 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1413 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1412 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1411 = (1'h0);
  reg [(3'h4):(1'h0)] reg1410 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1409 = (1'h0);
  reg [(4'hd):(1'h0)] reg1408 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1407 = (1'h0);
  reg [(4'hc):(1'h0)] reg1406 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1405 = (1'h0);
  reg [(2'h3):(1'h0)] reg1404 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1403 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1402 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1401 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1400 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1399 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1398 = (1'h0);
  reg [(2'h2):(1'h0)] reg1397 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1396 = (1'h0);
  reg [(5'h10):(1'h0)] reg1395 = (1'h0);
  reg [(2'h3):(1'h0)] reg1394 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1392 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1391 = (1'h0);
  reg [(4'he):(1'h0)] reg1390 = (1'h0);
  reg [(4'ha):(1'h0)] reg1389 = (1'h0);
  reg [(2'h2):(1'h0)] reg1388 = (1'h0);
  reg [(3'h6):(1'h0)] reg1387 = (1'h0);
  reg [(4'hb):(1'h0)] reg1386 = (1'h0);
  reg [(2'h3):(1'h0)] reg1385 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1384 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1383 = (1'h0);
  reg [(3'h6):(1'h0)] reg1382 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1381 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1380 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1378 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1376 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1372 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1379 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1378 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1377 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1376 = (1'h0);
  reg [(4'he):(1'h0)] reg1375 = (1'h0);
  reg [(4'he):(1'h0)] reg1374 = (1'h0);
  reg [(4'hd):(1'h0)] reg1373 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1372 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1371 = (1'h0);
  reg [(3'h4):(1'h0)] reg1370 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1369 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1367 = (1'h0);
  reg [(4'ha):(1'h0)] reg1366 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1364 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1363 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1358 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1353 = (1'h0);
  reg [(4'h8):(1'h0)] reg1347 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1344 = (1'h0);
  reg [(4'he):(1'h0)] forvar1343 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1338 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1355 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1368 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1367 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1366 = (1'h0);
  reg [(3'h4):(1'h0)] reg1365 = (1'h0);
  reg [(4'hc):(1'h0)] reg1364 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1363 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1362 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1361 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1360 = (1'h0);
  reg [(4'hb):(1'h0)] reg1359 = (1'h0);
  reg [(4'hb):(1'h0)] reg1358 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1357 = (1'h0);
  reg [(3'h7):(1'h0)] reg1356 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1355 = (1'h0);
  reg [(4'hc):(1'h0)] reg1354 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1353 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1352 = (1'h0);
  reg [(3'h5):(1'h0)] reg1351 = (1'h0);
  reg [(3'h4):(1'h0)] reg1350 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1349 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1348 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1347 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1346 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1345 = (1'h0);
  reg [(4'he):(1'h0)] reg1344 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1343 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1342 = (1'h0);
  reg [(3'h4):(1'h0)] reg1341 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1340 = (1'h0);
  reg [(2'h2):(1'h0)] reg1339 = (1'h0);
  reg [(2'h3):(1'h0)] reg1338 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1337 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1336 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1335 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1334 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1333 = (1'h0);
  reg [(3'h4):(1'h0)] reg1332 = (1'h0);
  reg [(5'h10):(1'h0)] reg1331 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1330 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1329 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1328 = (1'h0);
  reg [(2'h3):(1'h0)] reg1327 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1326 = (1'h0);
  reg [(4'he):(1'h0)] reg1325 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1324 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1320 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1319 = (1'h0);
  reg [(4'hd):(1'h0)] reg1311 = (1'h0);
  reg [(5'h10):(1'h0)] reg1317 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1315 = (1'h0);
  reg [(2'h3):(1'h0)] reg1312 = (1'h0);
  reg [(4'h8):(1'h0)] reg1323 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1322 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1321 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1320 = (1'h0);
  reg [(3'h5):(1'h0)] reg1319 = (1'h0);
  reg [(4'h9):(1'h0)] reg1318 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1317 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1316 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1315 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1314 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1313 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1312 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1311 = (1'h0);
  reg [(4'hf):(1'h0)] reg1310 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1309 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1308 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1307 = (1'h0);
  reg [(5'h10):(1'h0)] reg1306 = (1'h0);
  reg [(4'h9):(1'h0)] reg1305 = (1'h0);
  reg [(2'h2):(1'h0)] reg1304 = (1'h0);
  reg [(4'h8):(1'h0)] reg1303 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1302 = (1'h0);
  reg [(4'ha):(1'h0)] reg1301 = (1'h0);
  reg [(4'hf):(1'h0)] reg1300 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1299 = (1'h0);
  reg [(4'h9):(1'h0)] reg1298 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1297 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1296 = (1'h0);
  reg [(4'he):(1'h0)] reg1295 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1294 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1293 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1292 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1291 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1290 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1289 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1288 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1287 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1286 = (1'h0);
  wire [(3'h5):(1'h0)] wire1285;
  wire signed [(4'hc):(1'h0)] wire1284;
  reg [(4'ha):(1'h0)] reg1239 = (1'h0);
  reg [(3'h5):(1'h0)] reg1236 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1235 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1232 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1230 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1228 = (1'h0);
  reg [(4'ha):(1'h0)] reg1227 = (1'h0);
  reg [(4'h9):(1'h0)] reg1283 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1282 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1281 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1280 = (1'h0);
  reg [(2'h2):(1'h0)] reg1279 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1278 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1277 = (1'h0);
  reg [(4'h8):(1'h0)] reg1276 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1275 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1274 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1273 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1272 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1271 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1270 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1269 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1268 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1265 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1267 = (1'h0);
  reg [(4'hd):(1'h0)] reg1266 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1265 = (1'h0);
  reg [(2'h3):(1'h0)] reg1264 = (1'h0);
  reg [(4'ha):(1'h0)] reg1263 = (1'h0);
  reg [(2'h2):(1'h0)] reg1262 = (1'h0);
  reg [(4'hb):(1'h0)] reg1261 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1260 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1259 = (1'h0);
  reg [(4'hb):(1'h0)] reg1258 = (1'h0);
  reg [(4'hb):(1'h0)] reg1257 = (1'h0);
  reg [(4'ha):(1'h0)] reg1256 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1255 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1254 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1253 = (1'h0);
  reg [(3'h4):(1'h0)] reg1252 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1251 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1250 = (1'h0);
  reg [(3'h7):(1'h0)] reg1249 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1248 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1247 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1246 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1245 = (1'h0);
  reg [(4'h8):(1'h0)] reg1244 = (1'h0);
  reg [(4'he):(1'h0)] forvar1243 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1242 = (1'h0);
  reg [(4'hb):(1'h0)] reg1241 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1240 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1239 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1238 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1237 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1236 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1235 = (1'h0);
  reg [(3'h5):(1'h0)] reg1234 = (1'h0);
  reg [(2'h3):(1'h0)] reg1233 = (1'h0);
  reg [(2'h2):(1'h0)] reg1232 = (1'h0);
  reg [(3'h6):(1'h0)] reg1231 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1230 = (1'h0);
  reg [(4'he):(1'h0)] reg1229 = (1'h0);
  reg [(2'h3):(1'h0)] reg1228 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1227 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1226 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1225 = (1'h0);
  assign y = {wire1743,
                 reg1742,
                 reg1720,
                 forvar1717,
                 reg1716,
                 reg1715,
                 reg1741,
                 reg1739,
                 forvar1738,
                 reg1734,
                 reg1740,
                 forvar1739,
                 reg1738,
                 reg1737,
                 reg1736,
                 reg1735,
                 forvar1734,
                 reg1731,
                 reg1728,
                 forvar1724,
                 reg1733,
                 reg1732,
                 forvar1731,
                 reg1730,
                 reg1729,
                 forvar1728,
                 reg1727,
                 reg1726,
                 reg1725,
                 reg1724,
                 reg1723,
                 reg1722,
                 reg1721,
                 forvar1720,
                 reg1719,
                 reg1718,
                 reg1717,
                 forvar1716,
                 forvar1715,
                 reg1714,
                 reg1713,
                 reg1712,
                 reg1711,
                 reg1710,
                 forvar1709,
                 forvar1708,
                 reg1707,
                 reg1706,
                 reg1705,
                 forvar1704,
                 reg1703,
                 reg1702,
                 reg1701,
                 reg1700,
                 forvar1699,
                 forvar1697,
                 reg1698,
                 reg1697,
                 reg1696,
                 forvar1695,
                 forvar1694,
                 reg1693,
                 reg1692,
                 forvar1691,
                 forvar1690,
                 forvar1689,
                 wire1688,
                 reg1618,
                 reg1687,
                 reg1686,
                 reg1685,
                 reg1684,
                 forvar1683,
                 forvar1682,
                 reg1681,
                 reg1680,
                 reg1679,
                 reg1678,
                 forvar1677,
                 forvar1676,
                 forvar1675,
                 reg1674,
                 reg1673,
                 reg1672,
                 reg1671,
                 reg1670,
                 reg1657,
                 reg1669,
                 reg1668,
                 reg1667,
                 reg1666,
                 reg1665,
                 reg1664,
                 reg1663,
                 forvar1662,
                 reg1661,
                 reg1660,
                 reg1659,
                 reg1658,
                 forvar1657,
                 reg1656,
                 reg1655,
                 reg1654,
                 reg1653,
                 forvar1652,
                 reg1651,
                 forvar1650,
                 forvar1649,
                 forvar1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1640,
                 reg1639,
                 forvar1637,
                 reg1638,
                 reg1637,
                 reg1636,
                 reg1635,
                 forvar1634,
                 reg1633,
                 reg1632,
                 forvar1631,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1627,
                 forvar1626,
                 reg1625,
                 reg1624,
                 reg1623,
                 reg1622,
                 reg1621,
                 forvar1620,
                 reg1619,
                 forvar1618,
                 reg1601,
                 reg1599,
                 reg1617,
                 reg1616,
                 reg1615,
                 forvar1614,
                 forvar1613,
                 reg1612,
                 reg1611,
                 reg1610,
                 reg1609,
                 reg1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 reg1603,
                 reg1602,
                 forvar1601,
                 reg1600,
                 forvar1599,
                 forvar1598,
                 reg1597,
                 wire1596,
                 wire1595,
                 reg1594,
                 reg1593,
                 reg1592,
                 reg1591,
                 reg1590,
                 reg1589,
                 reg1588,
                 reg1587,
                 reg1586,
                 reg1585,
                 reg1584,
                 reg1583,
                 reg1582,
                 reg1581,
                 reg1580,
                 forvar1579,
                 forvar1578,
                 reg1577,
                 forvar1576,
                 reg1575,
                 reg1574,
                 reg1573,
                 forvar1572,
                 reg1571,
                 reg1570,
                 reg1569,
                 reg1568,
                 forvar1567,
                 reg1566,
                 reg1565,
                 reg1564,
                 reg1563,
                 forvar1557,
                 forvar1554,
                 forvar1549,
                 reg1547,
                 forvar1542,
                 reg1562,
                 reg1561,
                 reg1560,
                 reg1559,
                 reg1558,
                 reg1557,
                 reg1556,
                 reg1555,
                 reg1554,
                 reg1553,
                 forvar1550,
                 reg1552,
                 reg1551,
                 reg1550,
                 reg1549,
                 reg1548,
                 forvar1547,
                 reg1546,
                 reg1545,
                 reg1544,
                 forvar1543,
                 reg1542,
                 reg1541,
                 forvar1540,
                 reg1507,
                 forvar1506,
                 reg1539,
                 forvar1538,
                 reg1537,
                 reg1536,
                 reg1529,
                 reg1535,
                 reg1534,
                 reg1533,
                 reg1532,
                 reg1531,
                 reg1530,
                 forvar1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 reg1525,
                 forvar1524,
                 reg1523,
                 reg1521,
                 forvar1520,
                 reg1519,
                 reg1522,
                 forvar1521,
                 reg1520,
                 forvar1519,
                 reg1518,
                 reg1517,
                 reg1516,
                 reg1515,
                 reg1514,
                 reg1513,
                 reg1509,
                 forvar1508,
                 reg1512,
                 reg1511,
                 reg1510,
                 forvar1509,
                 reg1508,
                 forvar1507,
                 reg1506,
                 reg1505,
                 forvar1497,
                 reg1504,
                 reg1503,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1496,
                 forvar1493,
                 forvar1489,
                 reg1490,
                 reg1499,
                 reg1498,
                 reg1497,
                 forvar1496,
                 reg1495,
                 reg1494,
                 reg1493,
                 reg1492,
                 reg1491,
                 forvar1490,
                 reg1489,
                 forvar1488,
                 reg1487,
                 reg1486,
                 reg1485,
                 forvar1484,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1480,
                 forvar1479,
                 reg1478,
                 reg1477,
                 forvar1476,
                 reg1475,
                 reg1474,
                 forvar1473,
                 forvar1472,
                 reg1471,
                 reg1470,
                 forvar1469,
                 reg1468,
                 reg1467,
                 forvar1466,
                 reg1465,
                 forvar1464,
                 reg1463,
                 reg1462,
                 forvar1461,
                 forvar1460,
                 forvar1459,
                 reg1458,
                 forvar1453,
                 reg1457,
                 reg1456,
                 reg1455,
                 reg1454,
                 reg1453,
                 reg1444,
                 reg1452,
                 reg1451,
                 reg1450,
                 reg1449,
                 reg1448,
                 reg1447,
                 reg1446,
                 reg1445,
                 forvar1444,
                 reg1443,
                 reg1442,
                 forvar1441,
                 reg1440,
                 forvar1439,
                 forvar1408,
                 forvar1411,
                 forvar1394,
                 forvar1391,
                 reg1414,
                 forvar1410,
                 forvar1409,
                 reg1405,
                 forvar1404,
                 forvar1397,
                 reg1402,
                 reg1401,
                 forvar1398,
                 forvar1395,
                 reg1392,
                 reg1383,
                 forvar1436,
                 forvar1434,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1434,
                 forvar1433,
                 reg1432,
                 reg1431,
                 reg1430,
                 forvar1429,
                 reg1428,
                 reg1427,
                 forvar1426,
                 reg1425,
                 reg1424,
                 forvar1423,
                 reg1422,
                 reg1421,
                 reg1420,
                 forvar1419,
                 forvar1418,
                 reg1417,
                 reg1416,
                 reg1415,
                 forvar1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 reg1410,
                 reg1409,
                 reg1408,
                 reg1407,
                 reg1406,
                 forvar1405,
                 reg1404,
                 reg1403,
                 forvar1402,
                 forvar1401,
                 forvar1400,
                 reg1399,
                 reg1398,
                 reg1397,
                 reg1396,
                 reg1395,
                 reg1394,
                 reg1393,
                 forvar1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1386,
                 reg1385,
                 reg1384,
                 forvar1383,
                 reg1382,
                 reg1381,
                 reg1380,
                 forvar1378,
                 forvar1376,
                 reg1372,
                 reg1379,
                 reg1378,
                 reg1377,
                 reg1376,
                 reg1375,
                 reg1374,
                 reg1373,
                 forvar1372,
                 forvar1371,
                 reg1370,
                 reg1369,
                 forvar1367,
                 reg1366,
                 forvar1364,
                 forvar1363,
                 forvar1358,
                 forvar1353,
                 reg1347,
                 forvar1344,
                 forvar1343,
                 forvar1338,
                 reg1355,
                 reg1368,
                 reg1367,
                 forvar1366,
                 reg1365,
                 reg1364,
                 reg1363,
                 reg1362,
                 reg1361,
                 reg1360,
                 reg1359,
                 reg1358,
                 reg1357,
                 reg1356,
                 forvar1355,
                 reg1354,
                 reg1353,
                 reg1352,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 forvar1347,
                 reg1346,
                 reg1345,
                 reg1344,
                 reg1343,
                 reg1342,
                 reg1341,
                 reg1340,
                 reg1339,
                 reg1338,
                 forvar1337,
                 reg1336,
                 reg1335,
                 forvar1334,
                 reg1333,
                 reg1332,
                 reg1331,
                 reg1330,
                 forvar1329,
                 forvar1328,
                 reg1327,
                 reg1326,
                 reg1325,
                 forvar1324,
                 reg1320,
                 forvar1319,
                 reg1311,
                 reg1317,
                 forvar1315,
                 reg1312,
                 reg1323,
                 reg1322,
                 reg1321,
                 forvar1320,
                 reg1319,
                 reg1318,
                 forvar1317,
                 reg1316,
                 reg1315,
                 reg1314,
                 reg1313,
                 forvar1312,
                 forvar1311,
                 reg1310,
                 reg1309,
                 reg1308,
                 forvar1307,
                 reg1306,
                 reg1305,
                 reg1304,
                 reg1303,
                 forvar1302,
                 reg1301,
                 reg1300,
                 reg1299,
                 reg1298,
                 reg1297,
                 reg1296,
                 reg1295,
                 reg1294,
                 forvar1293,
                 reg1292,
                 reg1291,
                 reg1290,
                 reg1289,
                 forvar1288,
                 forvar1287,
                 forvar1286,
                 wire1285,
                 wire1284,
                 reg1239,
                 reg1236,
                 reg1235,
                 forvar1232,
                 reg1230,
                 forvar1228,
                 reg1227,
                 reg1283,
                 reg1282,
                 reg1281,
                 reg1280,
                 reg1279,
                 forvar1278,
                 forvar1277,
                 reg1276,
                 reg1275,
                 forvar1274,
                 forvar1273,
                 reg1272,
                 reg1271,
                 reg1270,
                 forvar1269,
                 reg1268,
                 forvar1265,
                 reg1267,
                 reg1266,
                 reg1265,
                 reg1264,
                 reg1263,
                 reg1262,
                 reg1261,
                 forvar1260,
                 reg1259,
                 reg1258,
                 reg1257,
                 reg1256,
                 forvar1255,
                 forvar1254,
                 reg1253,
                 reg1252,
                 reg1251,
                 reg1250,
                 reg1249,
                 forvar1248,
                 forvar1247,
                 reg1246,
                 reg1245,
                 reg1244,
                 forvar1243,
                 reg1242,
                 reg1241,
                 reg1240,
                 forvar1239,
                 reg1238,
                 reg1237,
                 forvar1236,
                 forvar1235,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1231,
                 forvar1230,
                 reg1229,
                 reg1228,
                 forvar1227,
                 forvar1226,
                 forvar1225,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($signed({$signed((~wire1223))}))
        begin
          for (forvar1225 = (1'h0); (forvar1225 < (1'h0)); forvar1225 = (forvar1225 + (1'h1)))
            begin
              for (forvar1226 = (1'h0); (forvar1226 < (2'h3)); forvar1226 = (forvar1226 + (1'h1)))
                begin
                  for (forvar1227 = (1'h0); (forvar1227 < (2'h2)); forvar1227 = (forvar1227 + (1'h1)))
                    begin
                      reg1228 <= ($signed($unsigned(((8'ha7) + wire1221))) ?
                          wire1224[(1'h0):(1'h0)] : wire1222[(1'h0):(1'h0)]);
                      reg1229 <= (-$signed((|(forvar1225 ?
                          forvar1226 : (8'hae)))));
                    end
                  for (forvar1230 = (1'h0); (forvar1230 < (1'h0)); forvar1230 = (forvar1230 + (1'h1)))
                    begin
                      reg1231 <= wire1222;
                      reg1232 <= reg1229[(4'hd):(4'hd)];
                      reg1233 <= (~$unsigned(wire1223));
                      reg1234 <= wire1220[(1'h1):(1'h0)];
                    end
                end
              for (forvar1235 = (1'h0); (forvar1235 < (1'h0)); forvar1235 = (forvar1235 + (1'h1)))
                begin
                  for (forvar1236 = (1'h0); (forvar1236 < (1'h0)); forvar1236 = (forvar1236 + (1'h1)))
                    begin
                      reg1237 <= $signed((((wire1222 ?
                              wire1221 : reg1229) && $unsigned(wire1223)) ?
                          $signed($unsigned(wire1222)) : (^~((8'hb5) ?
                              (8'h9c) : wire1224))));
                      reg1238 <= $signed({reg1231});
                    end
                  for (forvar1239 = (1'h0); (forvar1239 < (2'h3)); forvar1239 = (forvar1239 + (1'h1)))
                    begin
                      reg1240 <= forvar1226[(1'h0):(1'h0)];
                      reg1241 <= (-(forvar1235[(1'h1):(1'h0)] ?
                          reg1229 : $signed((~|wire1223))));
                      reg1242 <= ($signed($signed(wire1224)) ?
                          $signed((!(&forvar1226))) : reg1228);
                    end
                  for (forvar1243 = (1'h0); (forvar1243 < (2'h3)); forvar1243 = (forvar1243 + (1'h1)))
                    begin
                      reg1244 <= (wire1222 >>> ((((8'hb5) ?
                                  forvar1235 : reg1242) ?
                              reg1231 : $signed(forvar1225)) ?
                          forvar1235 : {$unsigned(forvar1225)}));
                      reg1245 <= $unsigned((^~($unsigned(forvar1235) ?
                          $unsigned(reg1244) : (reg1234 ?
                              reg1241 : forvar1236))));
                    end
                end
              reg1246 <= reg1228[(2'h2):(1'h1)];
              for (forvar1247 = (1'h0); (forvar1247 < (1'h0)); forvar1247 = (forvar1247 + (1'h1)))
                begin
                  for (forvar1248 = (1'h0); (forvar1248 < (2'h2)); forvar1248 = (forvar1248 + (1'h1)))
                    begin
                      reg1249 <= reg1233;
                    end
                  if (reg1240[(1'h0):(1'h0)])
                    begin
                      reg1250 <= reg1233;
                      reg1251 <= reg1238;
                      reg1252 <= (^{($signed(forvar1236) ?
                              (forvar1236 && wire1221) : (reg1231 ?
                                  reg1244 : reg1229))});
                      reg1253 <= ((~^(&$signed(forvar1248))) ^~ (($signed(reg1251) ?
                          {reg1242} : wire1222[(3'h4):(2'h3)]) * forvar1248));
                    end
                  else
                    begin
                      reg1250 <= forvar1230;
                      reg1251 <= ((8'h9d) ?
                          (~&$signed(forvar1243[(2'h2):(1'h1)])) : (^reg1244));
                    end
                end
            end
          for (forvar1254 = (1'h0); (forvar1254 < (2'h2)); forvar1254 = (forvar1254 + (1'h1)))
            begin
              for (forvar1255 = (1'h0); (forvar1255 < (2'h2)); forvar1255 = (forvar1255 + (1'h1)))
                begin
                  if ((~&$unsigned($unsigned($signed((8'h9f))))))
                    begin
                      reg1256 <= (reg1240 ?
                          ((~&$unsigned((8'haf))) | ($signed(forvar1225) ?
                              reg1242 : {wire1220})) : (~(!$signed(reg1241))));
                      reg1257 <= $unsigned($signed({$unsigned((8'h9d))}));
                      reg1258 <= {((reg1229[(4'hc):(1'h0)] ?
                              {reg1252} : (reg1228 == reg1232)) == (~|(~reg1231)))};
                    end
                  else
                    begin
                      reg1256 <= $unsigned((forvar1239[(4'ha):(3'h6)] <<< {forvar1235[(2'h2):(2'h2)]}));
                      reg1257 <= {((~$signed(wire1222)) ?
                              (&$signed(forvar1255)) : $signed(((8'hb9) || reg1241)))};
                    end
                  reg1259 <= forvar1255;
                  for (forvar1260 = (1'h0); (forvar1260 < (1'h0)); forvar1260 = (forvar1260 + (1'h1)))
                    begin
                      reg1261 <= (&$unsigned(((~&reg1250) ?
                          reg1228 : {reg1253})));
                      reg1262 <= ($signed(reg1246) ^ reg1252);
                      reg1263 <= forvar1235;
                      reg1264 <= $signed((!$signed(reg1241[(4'h8):(1'h0)])));
                    end
                end
              if (reg1241)
                begin
                  if ({(|forvar1248)})
                    begin
                      reg1265 <= (|(!forvar1235[(2'h3):(2'h2)]));
                      reg1266 <= wire1224[(2'h2):(1'h1)];
                      reg1267 <= reg1242;
                    end
                  else
                    begin
                      reg1265 <= ($unsigned(forvar1226[(3'h7):(3'h4)]) & $unsigned($unsigned(reg1267[(1'h1):(1'h0)])));
                      reg1266 <= reg1231;
                    end
                end
              else
                begin
                  for (forvar1265 = (1'h0); (forvar1265 < (1'h1)); forvar1265 = (forvar1265 + (1'h1)))
                    begin
                      reg1266 <= (~|$signed({(!reg1242)}));
                    end
                  reg1267 <= {forvar1225};
                  reg1268 <= $unsigned((^~(8'ha9)));
                  for (forvar1269 = (1'h0); (forvar1269 < (2'h3)); forvar1269 = (forvar1269 + (1'h1)))
                    begin
                      reg1270 <= reg1265;
                      reg1271 <= (8'had);
                      reg1272 <= $unsigned(reg1250[(2'h2):(1'h1)]);
                    end
                end
              for (forvar1273 = (1'h0); (forvar1273 < (2'h2)); forvar1273 = (forvar1273 + (1'h1)))
                begin
                  for (forvar1274 = (1'h0); (forvar1274 < (2'h2)); forvar1274 = (forvar1274 + (1'h1)))
                    begin
                      reg1275 <= {reg1258};
                      reg1276 <= $signed((~|reg1245[(3'h6):(3'h4)]));
                    end
                end
              for (forvar1277 = (1'h0); (forvar1277 < (1'h0)); forvar1277 = (forvar1277 + (1'h1)))
                begin
                  for (forvar1278 = (1'h0); (forvar1278 < (2'h2)); forvar1278 = (forvar1278 + (1'h1)))
                    begin
                      reg1279 <= (8'hb5);
                      reg1280 <= forvar1225[(3'h4):(1'h0)];
                      reg1281 <= $signed((($unsigned(reg1246) ?
                          $unsigned(reg1272) : {reg1272}) + (-(~reg1249))));
                    end
                  reg1282 <= (((^(reg1234 ? reg1264 : (8'hb4))) ?
                          (reg1234[(1'h1):(1'h1)] ^ (~&forvar1273)) : {{(8'ha3)}}) ?
                      $signed(reg1251[(4'h9):(1'h0)]) : $signed($unsigned(((8'hb6) == forvar1226))));
                end
            end
          reg1283 <= ({((^~reg1242) <<< {reg1266})} << (+$unsigned($unsigned(reg1270))));
        end
      else
        begin
          for (forvar1225 = (1'h0); (forvar1225 < (2'h2)); forvar1225 = (forvar1225 + (1'h1)))
            begin
              for (forvar1226 = (1'h0); (forvar1226 < (1'h0)); forvar1226 = (forvar1226 + (1'h1)))
                begin
                  reg1227 <= {{$signed({forvar1255})}};
                  for (forvar1228 = (1'h0); (forvar1228 < (1'h1)); forvar1228 = (forvar1228 + (1'h1)))
                    begin
                      reg1229 <= forvar1230[(3'h7):(1'h0)];
                      reg1230 <= reg1240[(2'h2):(2'h2)];
                      reg1231 <= $signed($signed((^$unsigned((8'ha1)))));
                    end
                  for (forvar1232 = (1'h0); (forvar1232 < (2'h3)); forvar1232 = (forvar1232 + (1'h1)))
                    begin
                      reg1233 <= $signed((8'hb1));
                      reg1234 <= (|(8'ha2));
                      reg1235 <= (~&reg1234[(1'h0):(1'h0)]);
                      reg1236 <= (($unsigned(forvar1228) >>> (&$unsigned(reg1231))) ^~ $signed(($signed(wire1221) ?
                          {forvar1225} : (reg1253 * reg1244))));
                    end
                  if ((+reg1242))
                    begin
                      reg1237 <= $signed($unsigned((|reg1227)));
                    end
                  else
                    begin
                      reg1237 <= {reg1227};
                      reg1238 <= (reg1270 ?
                          (reg1236 ?
                              forvar1248[(3'h7):(3'h7)] : {{forvar1236}}) : $signed(wire1222[(3'h5):(2'h3)]));
                      reg1239 <= $unsigned({$signed({reg1253})});
                    end
                end
            end
        end
    end
  assign wire1284 = $unsigned(forvar1232);
  assign wire1285 = $signed(reg1259);
  always
    @(posedge clk) begin
      for (forvar1286 = (1'h0); (forvar1286 < (2'h2)); forvar1286 = (forvar1286 + (1'h1)))
        begin
          for (forvar1287 = (1'h0); (forvar1287 < (2'h3)); forvar1287 = (forvar1287 + (1'h1)))
            begin
              if ($signed(($unsigned((|forvar1269)) ?
                  $signed(reg1253) : $signed(forvar1273))))
                begin
                  for (forvar1288 = (1'h0); (forvar1288 < (1'h1)); forvar1288 = (forvar1288 + (1'h1)))
                    begin
                      reg1289 <= ($signed(($unsigned(forvar1248) ?
                          forvar1236[(3'h7):(3'h5)] : (8'h9e))) + $signed($signed((reg1241 << reg1237))));
                    end
                end
              else
                begin
                  for (forvar1288 = (1'h0); (forvar1288 < (1'h0)); forvar1288 = (forvar1288 + (1'h1)))
                    begin
                      reg1289 <= reg1234;
                      reg1290 <= $signed($signed(forvar1278[(2'h3):(1'h1)]));
                      reg1291 <= $unsigned(reg1270[(3'h5):(2'h2)]);
                    end
                end
              if (wire1224)
                begin
                  reg1292 <= reg1272;
                  for (forvar1293 = (1'h0); (forvar1293 < (1'h0)); forvar1293 = (forvar1293 + (1'h1)))
                    begin
                      reg1294 <= (($signed((forvar1228 ? reg1283 : wire1220)) ?
                          ({(8'ha3)} - reg1271) : (!(wire1224 ?
                              reg1249 : reg1259))) >= forvar1239);
                      reg1295 <= $unsigned((^~(~&reg1230)));
                      reg1296 <= ((&$signed((wire1285 <= reg1271))) | reg1291);
                      reg1297 <= $unsigned(((reg1250 <= (+reg1263)) <<< ($unsigned(forvar1228) == (reg1251 < forvar1226))));
                    end
                  if ($signed($unsigned(reg1270)))
                    begin
                      reg1298 <= (~$unsigned(((8'ha3) + $unsigned(reg1295))));
                      reg1299 <= (($signed(reg1241) <<< forvar1287[(3'h5):(2'h3)]) || ((reg1238[(3'h5):(3'h4)] ?
                              $unsigned(reg1266) : {reg1242}) ?
                          reg1276 : ($unsigned(reg1227) >> (~|(8'haf)))));
                      reg1300 <= reg1281[(4'hf):(1'h1)];
                      reg1301 <= (~^(((reg1275 ? forvar1293 : reg1234) ?
                              (reg1296 && reg1246) : $unsigned(reg1296)) ?
                          reg1281 : reg1267[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg1298 <= ($signed(($unsigned(reg1265) & {reg1238})) & $unsigned($signed((reg1228 ?
                          (8'had) : (8'haf)))));
                    end
                end
              else
                begin
                  reg1292 <= $unsigned(reg1238[(1'h0):(1'h0)]);
                end
              for (forvar1302 = (1'h0); (forvar1302 < (2'h2)); forvar1302 = (forvar1302 + (1'h1)))
                begin
                  reg1303 <= $signed((~&({reg1238} ?
                      $unsigned(reg1263) : $unsigned(reg1300))));
                  if (reg1283)
                    begin
                      reg1304 <= $signed({{(forvar1288 ? reg1296 : reg1261)}});
                      reg1305 <= forvar1243;
                    end
                  else
                    begin
                      reg1304 <= $unsigned(reg1289[(1'h1):(1'h1)]);
                      reg1305 <= reg1271;
                      reg1306 <= $unsigned(forvar1288);
                    end
                end
              for (forvar1307 = (1'h0); (forvar1307 < (1'h0)); forvar1307 = (forvar1307 + (1'h1)))
                begin
                  reg1308 <= (({(reg1283 ? (8'ha5) : reg1230)} ?
                          $unsigned((8'hb4)) : reg1229[(2'h3):(2'h3)]) ?
                      (forvar1287[(3'h5):(2'h2)] & (|{(8'hb7)})) : reg1252);
                  reg1309 <= (($unsigned($unsigned(reg1234)) | {(reg1303 >> reg1233)}) ?
                      $unsigned($signed($unsigned(forvar1274))) : ($unsigned(forvar1248[(1'h1):(1'h0)]) <= {forvar1287}));
                end
            end
          if ((-reg1256))
            begin
              reg1310 <= forvar1278;
              for (forvar1311 = (1'h0); (forvar1311 < (1'h0)); forvar1311 = (forvar1311 + (1'h1)))
                begin
                  for (forvar1312 = (1'h0); (forvar1312 < (2'h3)); forvar1312 = (forvar1312 + (1'h1)))
                    begin
                      reg1313 <= {wire1223[(2'h2):(1'h1)]};
                      reg1314 <= $unsigned((|$unsigned(((8'ha5) ?
                          reg1275 : reg1276))));
                      reg1315 <= (~^reg1303);
                      reg1316 <= reg1258;
                    end
                  for (forvar1317 = (1'h0); (forvar1317 < (1'h0)); forvar1317 = (forvar1317 + (1'h1)))
                    begin
                      reg1318 <= (|((reg1295[(4'hd):(2'h3)] == (reg1251 + forvar1254)) >>> (forvar1243 ?
                          reg1251 : {(8'h9d)})));
                      reg1319 <= $signed((^~$unsigned(reg1227[(3'h4):(2'h2)])));
                    end
                  for (forvar1320 = (1'h0); (forvar1320 < (1'h1)); forvar1320 = (forvar1320 + (1'h1)))
                    begin
                      reg1321 <= wire1223[(4'hc):(4'hb)];
                      reg1322 <= ($signed(reg1253[(4'h8):(1'h1)]) - reg1270);
                      reg1323 <= reg1305;
                    end
                end
            end
          else
            begin
              reg1310 <= $unsigned((|((~|reg1321) & (reg1261 == forvar1235))));
              if ({$unsigned(((wire1222 || reg1261) <= forvar1288))})
                begin
                  for (forvar1311 = (1'h0); (forvar1311 < (2'h3)); forvar1311 = (forvar1311 + (1'h1)))
                    begin
                      reg1312 <= ($signed($signed((^~reg1263))) > $unsigned(reg1283));
                      reg1313 <= ((&reg1297) > ((!$unsigned(wire1222)) ?
                          reg1289 : $signed((wire1222 - reg1268))));
                      reg1314 <= (~&reg1257);
                    end
                  for (forvar1315 = (1'h0); (forvar1315 < (2'h2)); forvar1315 = (forvar1315 + (1'h1)))
                    begin
                      reg1316 <= $unsigned($signed((~&(wire1222 >>> reg1283))));
                      reg1317 <= (-reg1241);
                    end
                  reg1318 <= ((~&reg1297[(4'h8):(3'h6)]) << $unsigned(forvar1248[(4'h8):(3'h7)]));
                end
              else
                begin
                  reg1311 <= (~^$signed((((8'hab) ?
                      forvar1320 : reg1270) <= $signed(wire1221))));
                  for (forvar1312 = (1'h0); (forvar1312 < (1'h1)); forvar1312 = (forvar1312 + (1'h1)))
                    begin
                      reg1313 <= (~&$unsigned(((reg1311 ^~ reg1281) ?
                          reg1238 : $unsigned(reg1309))));
                      reg1314 <= forvar1278[(1'h1):(1'h0)];
                    end
                  if ($signed(({(^~reg1229)} ?
                      reg1267[(2'h2):(2'h2)] : $signed((forvar1315 <= reg1239)))))
                    begin
                      reg1315 <= $signed(forvar1293);
                      reg1316 <= $signed({$signed(forvar1286[(3'h4):(1'h1)])});
                      reg1317 <= (~&$unsigned((~^$signed(reg1304))));
                    end
                  else
                    begin
                      reg1315 <= {(reg1264[(1'h1):(1'h0)] << reg1317)};
                      reg1316 <= {forvar1287[(3'h5):(2'h3)]};
                    end
                end
              if ($unsigned(reg1231))
                begin
                  reg1319 <= (^((~^forvar1226[(2'h2):(2'h2)]) ?
                      ($unsigned(forvar1248) < {forvar1230}) : reg1241[(4'hb):(4'ha)]));
                  for (forvar1320 = (1'h0); (forvar1320 < (1'h1)); forvar1320 = (forvar1320 + (1'h1)))
                    begin
                      reg1321 <= reg1240[(1'h0):(1'h0)];
                    end
                  reg1322 <= $signed($signed(reg1296[(3'h7):(3'h6)]));
                end
              else
                begin
                  for (forvar1319 = (1'h0); (forvar1319 < (2'h3)); forvar1319 = (forvar1319 + (1'h1)))
                    begin
                      reg1320 <= $unsigned((reg1303[(3'h5):(2'h3)] >= reg1299[(4'ha):(4'h8)]));
                      reg1321 <= reg1282;
                      reg1322 <= ($signed((8'h9f)) * $unsigned(reg1279[(2'h2):(2'h2)]));
                      reg1323 <= forvar1307;
                    end
                  for (forvar1324 = (1'h0); (forvar1324 < (2'h3)); forvar1324 = (forvar1324 + (1'h1)))
                    begin
                      reg1325 <= reg1318;
                      reg1326 <= $signed((&$signed(reg1229)));
                      reg1327 <= {(reg1282[(2'h2):(1'h0)] * (reg1297[(1'h1):(1'h1)] < reg1250[(2'h3):(2'h3)]))};
                    end
                end
              for (forvar1328 = (1'h0); (forvar1328 < (2'h2)); forvar1328 = (forvar1328 + (1'h1)))
                begin
                  for (forvar1329 = (1'h0); (forvar1329 < (2'h2)); forvar1329 = (forvar1329 + (1'h1)))
                    begin
                      reg1330 <= (reg1319[(2'h3):(2'h3)] >> reg1233);
                      reg1331 <= (~reg1290[(1'h0):(1'h0)]);
                      reg1332 <= $unsigned(($signed($unsigned(reg1326)) + {(forvar1287 + reg1264)}));
                    end
                  reg1333 <= forvar1265;
                  for (forvar1334 = (1'h0); (forvar1334 < (2'h2)); forvar1334 = (forvar1334 + (1'h1)))
                    begin
                      reg1335 <= $unsigned((((reg1234 ?
                          forvar1227 : reg1296) <<< (~&reg1299)) - {(forvar1243 ?
                              reg1236 : forvar1329)}));
                    end
                  reg1336 <= ($unsigned(forvar1260) ?
                      (reg1229[(2'h2):(1'h0)] ?
                          ({(8'ha2)} ?
                              forvar1315 : $unsigned(reg1333)) : ((reg1311 ?
                              forvar1255 : forvar1317) & $unsigned(reg1240))) : (($unsigned(wire1220) ?
                          (reg1245 < (8'h9e)) : $unsigned(forvar1269)) | $signed(reg1261)));
                end
            end
          if (reg1300)
            begin
              if (reg1249)
                begin
                  for (forvar1337 = (1'h0); (forvar1337 < (1'h0)); forvar1337 = (forvar1337 + (1'h1)))
                    begin
                      reg1338 <= reg1310[(1'h0):(1'h0)];
                      reg1339 <= (~^$unsigned(reg1291));
                      reg1340 <= reg1305;
                      reg1341 <= (reg1316[(3'h7):(2'h3)] * (({reg1231} ?
                              (~^forvar1228) : reg1238[(3'h4):(1'h0)]) ?
                          reg1262[(1'h1):(1'h0)] : reg1322));
                    end
                end
              else
                begin
                  for (forvar1337 = (1'h0); (forvar1337 < (1'h0)); forvar1337 = (forvar1337 + (1'h1)))
                    begin
                      reg1338 <= $unsigned($unsigned((~&reg1252)));
                      reg1339 <= (reg1303[(2'h3):(1'h1)] >>> ($unsigned(reg1304) ?
                          (&(8'h9d)) : {{reg1251}}));
                      reg1340 <= {reg1228[(1'h1):(1'h0)]};
                      reg1341 <= (!$signed($signed({reg1291})));
                    end
                  reg1342 <= {$unsigned(reg1246[(2'h3):(1'h1)])};
                  if ((!$signed(forvar1254)))
                    begin
                      reg1343 <= ($signed(reg1317) ?
                          reg1272 : reg1257[(4'hb):(1'h0)]);
                      reg1344 <= (8'hb1);
                      reg1345 <= ((~$signed(reg1232)) >> (reg1261 >> {(8'hae)}));
                      reg1346 <= ($unsigned(((reg1343 ?
                          reg1342 : reg1316) + (reg1312 ?
                          reg1322 : forvar1286))) ^ $signed(reg1310[(4'ha):(3'h5)]));
                    end
                  else
                    begin
                      reg1343 <= (-((((8'hb9) > forvar1230) ?
                          $signed(wire1220) : (&reg1330)) >>> $unsigned($signed(wire1224))));
                      reg1344 <= ($unsigned(($unsigned(reg1316) <<< reg1233[(1'h0):(1'h0)])) ?
                          (wire1285[(1'h0):(1'h0)] ?
                              ((reg1310 ?
                                  reg1231 : reg1246) + $unsigned(forvar1312)) : reg1320[(1'h1):(1'h0)]) : {($signed((8'h9f)) ?
                                  (8'had) : {forvar1293})});
                      reg1345 <= ((^{forvar1307[(4'h9):(3'h5)]}) || (&reg1308[(2'h2):(1'h0)]));
                    end
                end
              for (forvar1347 = (1'h0); (forvar1347 < (1'h1)); forvar1347 = (forvar1347 + (1'h1)))
                begin
                  if ($unsigned($unsigned($signed(((8'hb3) ?
                      (8'haa) : reg1300)))))
                    begin
                      reg1348 <= $signed(reg1249);
                      reg1349 <= (forvar1255[(3'h4):(1'h0)] ?
                          ($signed(reg1309[(2'h2):(2'h2)]) ?
                              wire1220[(2'h2):(1'h0)] : (+(reg1276 ?
                                  reg1290 : reg1344))) : ($signed(forvar1311[(2'h3):(1'h0)]) ?
                              reg1256[(3'h5):(1'h1)] : {(reg1262 ?
                                      reg1267 : reg1316)}));
                      reg1350 <= reg1266[(3'h7):(1'h1)];
                    end
                  else
                    begin
                      reg1348 <= {$signed((8'had))};
                      reg1349 <= $unsigned((^($signed(reg1275) ?
                          forvar1317[(2'h3):(2'h3)] : (reg1257 ?
                              forvar1243 : reg1256))));
                      reg1350 <= ($signed((((8'haf) ?
                              forvar1243 : (8'had)) && (-reg1291))) ?
                          (~&((reg1236 <<< (8'ha0)) <<< (~^reg1263))) : (8'haa));
                      reg1351 <= $unsigned(((^(reg1301 ?
                          reg1237 : (8'h9d))) == ($unsigned((8'hb1)) ?
                          reg1272 : ((8'ha1) >>> (8'hb9)))));
                    end
                  if ((({$unsigned((8'hb6))} > ((forvar1288 == reg1350) * (reg1251 ?
                          reg1258 : reg1228))) ?
                      reg1294[(1'h1):(1'h1)] : ((reg1341[(1'h1):(1'h0)] ?
                          reg1265[(2'h3):(2'h3)] : reg1330[(4'hf):(4'hc)]) > (reg1320 ?
                          forvar1288 : forvar1260[(3'h5):(1'h0)]))))
                    begin
                      reg1352 <= (^$signed(((^forvar1324) && {forvar1287})));
                    end
                  else
                    begin
                      reg1352 <= (reg1245 >= (+reg1249[(1'h0):(1'h0)]));
                      reg1353 <= ($signed((^(reg1351 << reg1321))) ?
                          {forvar1227[(3'h6):(1'h0)]} : {(~(forvar1254 != forvar1317))});
                    end
                  reg1354 <= {(+reg1345)};
                end
              if (($signed($unsigned($unsigned((8'h9c)))) ?
                  {(~&(-reg1306))} : (-((&reg1322) ?
                      (8'hb1) : (reg1317 ? forvar1328 : forvar1273)))))
                begin
                  for (forvar1355 = (1'h0); (forvar1355 < (2'h3)); forvar1355 = (forvar1355 + (1'h1)))
                    begin
                      reg1356 <= $signed((forvar1255[(3'h4):(3'h4)] <= ((reg1349 ?
                              (8'h9e) : reg1280) ?
                          (&reg1301) : {forvar1278})));
                      reg1357 <= reg1267[(2'h3):(2'h2)];
                      reg1358 <= (reg1346[(3'h7):(1'h0)] ?
                          $signed($unsigned({forvar1302})) : {forvar1232[(4'h9):(1'h0)]});
                    end
                  if ($signed($unsigned(($unsigned(reg1276) <= $signed(reg1237)))))
                    begin
                      reg1359 <= reg1228;
                      reg1360 <= (~^$signed($unsigned(forvar1273[(1'h1):(1'h1)])));
                      reg1361 <= reg1352[(4'ha):(3'h5)];
                    end
                  else
                    begin
                      reg1359 <= (forvar1243[(4'ha):(4'ha)] ?
                          $unsigned((+$signed(forvar1347))) : $unsigned(reg1296[(4'hb):(2'h2)]));
                      reg1360 <= (($signed($unsigned(reg1229)) ?
                          (reg1335 && $signed(reg1246)) : (+reg1351)) & (|(reg1239[(3'h6):(1'h1)] ?
                          reg1271 : (8'hb5))));
                    end
                  if ({$signed({$unsigned(reg1304)})})
                    begin
                      reg1362 <= reg1283;
                      reg1363 <= reg1264;
                      reg1364 <= reg1230[(2'h2):(2'h2)];
                      reg1365 <= {{(forvar1287[(3'h5):(3'h4)] <<< $signed(reg1276))}};
                    end
                  else
                    begin
                      reg1362 <= $unsigned(reg1276);
                      reg1363 <= reg1297[(1'h1):(1'h0)];
                    end
                  for (forvar1366 = (1'h0); (forvar1366 < (2'h2)); forvar1366 = (forvar1366 + (1'h1)))
                    begin
                      reg1367 <= ((~^$unsigned((forvar1329 != reg1353))) - $unsigned($unsigned(reg1330)));
                      reg1368 <= ({{$signed(wire1284)}} ?
                          $unsigned((8'hb1)) : ($signed(forvar1225[(2'h3):(2'h3)]) ?
                              ($signed(forvar1337) ?
                                  $unsigned(forvar1248) : $unsigned((8'hb7))) : wire1221));
                    end
                end
              else
                begin
                  if ((reg1236 ?
                      ((^((8'hb1) ? (8'hae) : reg1252)) ?
                          forvar1324 : (~&$unsigned(reg1360))) : {(!{reg1339})}))
                    begin
                      reg1355 <= (!($signed(reg1241) ?
                          $unsigned(forvar1317[(3'h6):(3'h5)]) : $unsigned((reg1253 >= reg1331))));
                    end
                  else
                    begin
                      reg1355 <= $signed((8'ha9));
                    end
                  if ($unsigned($signed((&reg1300))))
                    begin
                      reg1356 <= $signed((8'hba));
                      reg1357 <= $signed(((((8'hb3) | (8'ha1)) ?
                          $unsigned(reg1300) : forvar1247[(4'ha):(4'h8)]) || (~&(~^forvar1324))));
                    end
                  else
                    begin
                      reg1356 <= reg1233;
                      reg1357 <= $unsigned(forvar1324[(1'h1):(1'h0)]);
                      reg1358 <= (~|reg1235);
                    end
                end
            end
          else
            begin
              for (forvar1337 = (1'h0); (forvar1337 < (2'h3)); forvar1337 = (forvar1337 + (1'h1)))
                begin
                  for (forvar1338 = (1'h0); (forvar1338 < (1'h0)); forvar1338 = (forvar1338 + (1'h1)))
                    begin
                      reg1339 <= $signed(($signed(forvar1324) ?
                          $signed($unsigned((8'hb8))) : ($signed(reg1314) >= (^(8'hb4)))));
                      reg1340 <= $signed(reg1290[(4'hc):(2'h3)]);
                      reg1341 <= reg1231[(1'h1):(1'h1)];
                      reg1342 <= (-forvar1315[(1'h1):(1'h1)]);
                    end
                end
              for (forvar1343 = (1'h0); (forvar1343 < (2'h2)); forvar1343 = (forvar1343 + (1'h1)))
                begin
                  for (forvar1344 = (1'h0); (forvar1344 < (1'h1)); forvar1344 = (forvar1344 + (1'h1)))
                    begin
                      reg1345 <= reg1345;
                      reg1346 <= $signed(($unsigned((-reg1348)) | $unsigned(reg1294)));
                      reg1347 <= forvar1337[(3'h4):(2'h2)];
                      reg1348 <= (-reg1320);
                    end
                  if ((~(~^reg1295)))
                    begin
                      reg1349 <= $signed((-((forvar1338 <<< reg1314) ?
                          $unsigned(wire1284) : (~|(8'h9d)))));
                      reg1350 <= $signed((reg1304 ?
                          forvar1324[(3'h4):(2'h3)] : {reg1340[(4'ha):(1'h1)]}));
                      reg1351 <= (((forvar1319[(2'h2):(1'h0)] >> (reg1348 ?
                              forvar1366 : wire1284)) | (8'hab)) ?
                          (((~&reg1265) ~^ (forvar1320 ?
                              reg1236 : reg1341)) - reg1363) : ((^forvar1329) ?
                              (!{forvar1226}) : ((reg1283 ?
                                  reg1297 : reg1264) & $unsigned(reg1306))));
                    end
                  else
                    begin
                      reg1349 <= $unsigned(forvar1307);
                      reg1350 <= reg1368;
                      reg1351 <= reg1326;
                      reg1352 <= ((reg1306 >= {forvar1319}) ?
                          $signed($signed((-forvar1343))) : reg1239);
                    end
                  for (forvar1353 = (1'h0); (forvar1353 < (2'h3)); forvar1353 = (forvar1353 + (1'h1)))
                    begin
                      reg1354 <= $signed(reg1363);
                      reg1355 <= ((|forvar1338[(2'h2):(2'h2)]) == (+reg1330));
                      reg1356 <= (~^reg1320[(3'h5):(3'h5)]);
                      reg1357 <= (|$unsigned(reg1244));
                    end
                  for (forvar1358 = (1'h0); (forvar1358 < (2'h2)); forvar1358 = (forvar1358 + (1'h1)))
                    begin
                      reg1359 <= $signed(reg1367);
                      reg1360 <= (|$signed((^~(+reg1271))));
                      reg1361 <= reg1305;
                      reg1362 <= forvar1260;
                    end
                end
              for (forvar1363 = (1'h0); (forvar1363 < (1'h1)); forvar1363 = (forvar1363 + (1'h1)))
                begin
                  for (forvar1364 = (1'h0); (forvar1364 < (1'h1)); forvar1364 = (forvar1364 + (1'h1)))
                    begin
                      reg1365 <= $signed(((~^(wire1220 ?
                              forvar1347 : reg1233)) ?
                          $signed(forvar1319) : ((&forvar1329) >= reg1343)));
                      reg1366 <= reg1332[(1'h0):(1'h0)];
                    end
                  for (forvar1367 = (1'h0); (forvar1367 < (2'h2)); forvar1367 = (forvar1367 + (1'h1)))
                    begin
                      reg1368 <= reg1351[(3'h4):(1'h0)];
                      reg1369 <= ((reg1340[(2'h2):(2'h2)] ?
                          {(~&forvar1347)} : (~|$unsigned(reg1365))) >= reg1250[(1'h1):(1'h0)]);
                    end
                end
            end
        end
      if ($unsigned((&reg1339[(2'h2):(2'h2)])))
        begin
          reg1370 <= $unsigned((+{forvar1255}));
          for (forvar1371 = (1'h0); (forvar1371 < (2'h3)); forvar1371 = (forvar1371 + (1'h1)))
            begin
              if ((^~$signed(((reg1252 ?
                  reg1358 : reg1292) ~^ $signed((8'haf))))))
                begin
                  for (forvar1372 = (1'h0); (forvar1372 < (1'h1)); forvar1372 = (forvar1372 + (1'h1)))
                    begin
                      reg1373 <= {{(reg1346 + forvar1265)}};
                      reg1374 <= {reg1268[(3'h4):(2'h3)]};
                      reg1375 <= forvar1248[(2'h2):(1'h0)];
                    end
                  reg1376 <= (reg1366 >> (!reg1341[(1'h1):(1'h1)]));
                  reg1377 <= {reg1303};
                  if (((~$unsigned($unsigned(reg1339))) - (+($unsigned(reg1353) * reg1335[(1'h0):(1'h0)]))))
                    begin
                      reg1378 <= $signed(reg1227);
                      reg1379 <= $unsigned((8'h9c));
                    end
                  else
                    begin
                      reg1378 <= ((forvar1288 | (^((8'hb8) ?
                          reg1272 : reg1310))) ^ reg1352);
                    end
                end
              else
                begin
                  if (((+(~(~&reg1332))) ?
                      {$signed(reg1242[(4'h8):(1'h0)])} : $unsigned(reg1235)))
                    begin
                      reg1372 <= {$signed($unsigned($signed(reg1300)))};
                      reg1373 <= (~^$signed($unsigned(((8'haa) ?
                          reg1341 : reg1316))));
                      reg1374 <= {{$signed((reg1327 ? reg1294 : forvar1329))}};
                      reg1375 <= (reg1305 ?
                          $signed($unsigned({reg1265})) : reg1332);
                    end
                  else
                    begin
                      reg1372 <= forvar1243[(2'h3):(1'h0)];
                      reg1373 <= (reg1340[(5'h10):(2'h3)] == $unsigned($signed($unsigned((8'hb2)))));
                      reg1374 <= reg1253;
                    end
                  for (forvar1376 = (1'h0); (forvar1376 < (2'h2)); forvar1376 = (forvar1376 + (1'h1)))
                    begin
                      reg1377 <= {$signed(($unsigned(forvar1288) * (~reg1266)))};
                    end
                  for (forvar1378 = (1'h0); (forvar1378 < (1'h1)); forvar1378 = (forvar1378 + (1'h1)))
                    begin
                      reg1379 <= reg1239;
                      reg1380 <= ((($unsigned(reg1327) > (reg1320 <= reg1240)) * forvar1329) ^~ {reg1230[(1'h0):(1'h0)]});
                      reg1381 <= $signed({$signed($unsigned(reg1232))});
                      reg1382 <= $signed(((!$signed(reg1352)) >>> $signed(((8'hb7) <= reg1358))));
                    end
                end
              for (forvar1383 = (1'h0); (forvar1383 < (1'h0)); forvar1383 = (forvar1383 + (1'h1)))
                begin
                  reg1384 <= (reg1292[(2'h2):(1'h1)] || $unsigned(((^~forvar1255) && reg1313[(3'h5):(1'h0)])));
                  if (((reg1321 ?
                      {forvar1302} : {(forvar1358 ?
                              reg1299 : reg1362)}) == ((~^reg1308) - forvar1358)))
                    begin
                      reg1385 <= $unsigned((+($signed(reg1283) ^~ reg1338)));
                      reg1386 <= reg1368;
                      reg1387 <= {forvar1328};
                      reg1388 <= $unsigned($signed(((|forvar1288) ?
                          (reg1279 ? wire1224 : (8'hb6)) : reg1318)));
                    end
                  else
                    begin
                      reg1385 <= $unsigned(($unsigned((forvar1307 && reg1236)) << forvar1254));
                      reg1386 <= ({{forvar1371[(3'h7):(3'h4)]}} << ((reg1331[(3'h7):(3'h7)] << reg1262) ?
                          ({reg1295} ?
                              reg1356[(1'h0):(1'h0)] : (|forvar1317)) : ((8'haa) ?
                              (^~reg1316) : $signed(reg1369))));
                    end
                  if ((reg1232 ?
                      $unsigned(reg1241[(2'h2):(1'h1)]) : $unsigned($unsigned({reg1351}))))
                    begin
                      reg1389 <= (((~((8'ha9) ?
                              reg1361 : reg1367)) == $unsigned(((8'h9f) << reg1311))) ?
                          (((-reg1298) | reg1289) >> reg1303[(3'h7):(1'h1)]) : reg1366[(4'ha):(4'ha)]);
                      reg1390 <= forvar1364[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1389 <= {$unsigned((-{forvar1302}))};
                      reg1390 <= forvar1324[(2'h2):(2'h2)];
                      reg1391 <= $signed((reg1342[(1'h1):(1'h0)] || forvar1355));
                    end
                  for (forvar1392 = (1'h0); (forvar1392 < (2'h3)); forvar1392 = (forvar1392 + (1'h1)))
                    begin
                      reg1393 <= forvar1343;
                      reg1394 <= $signed(reg1327[(1'h1):(1'h0)]);
                      reg1395 <= ($unsigned(forvar1319[(2'h2):(1'h1)]) && forvar1319[(1'h0):(1'h0)]);
                    end
                end
              if ((reg1306 ?
                  $signed(((forvar1312 != (8'ha2)) - forvar1383[(4'hb):(3'h7)])) : $signed(reg1230[(1'h1):(1'h0)])))
                begin
                  if (forvar1383)
                    begin
                      reg1396 <= {(reg1237[(3'h7):(3'h4)] ?
                              $unsigned((forvar1329 >>> forvar1302)) : {{forvar1227}})};
                    end
                  else
                    begin
                      reg1396 <= reg1227[(3'h5):(3'h4)];
                      reg1397 <= forvar1254[(3'h4):(1'h1)];
                      reg1398 <= forvar1364[(4'ha):(3'h4)];
                      reg1399 <= (((!(reg1262 ? (8'hb2) : reg1239)) ?
                              $unsigned((reg1339 ?
                                  reg1262 : reg1385)) : ((reg1241 ?
                                      reg1335 : (8'haa)) ?
                                  $unsigned(reg1344) : wire1285)) ?
                          (~(reg1389 ?
                              ((8'hb2) ?
                                  reg1386 : reg1333) : $unsigned(reg1295))) : ($signed((reg1257 ?
                              forvar1364 : forvar1338)) < forvar1307[(2'h3):(1'h0)]));
                    end
                end
              else
                begin
                  if (forvar1383[(4'h8):(1'h1)])
                    begin
                      reg1396 <= (8'hb8);
                      reg1397 <= (~^reg1361);
                      reg1398 <= (8'hac);
                    end
                  else
                    begin
                      reg1396 <= reg1297;
                      reg1397 <= ($signed($unsigned(forvar1328)) ?
                          {$signed((8'ha8))} : forvar1227);
                      reg1398 <= $signed(forvar1247);
                    end
                end
            end
          for (forvar1400 = (1'h0); (forvar1400 < (1'h1)); forvar1400 = (forvar1400 + (1'h1)))
            begin
              for (forvar1401 = (1'h0); (forvar1401 < (1'h1)); forvar1401 = (forvar1401 + (1'h1)))
                begin
                  for (forvar1402 = (1'h0); (forvar1402 < (1'h0)); forvar1402 = (forvar1402 + (1'h1)))
                    begin
                      reg1403 <= reg1353[(3'h5):(2'h3)];
                      reg1404 <= reg1362;
                    end
                  for (forvar1405 = (1'h0); (forvar1405 < (1'h1)); forvar1405 = (forvar1405 + (1'h1)))
                    begin
                      reg1406 <= (((+$unsigned(reg1282)) >> ((^~reg1394) != (~&reg1335))) <<< (+reg1352[(1'h1):(1'h1)]));
                      reg1407 <= (((+$signed(forvar1338)) ?
                              (+{reg1237}) : reg1240[(1'h0):(1'h0)]) ?
                          (-((forvar1277 < reg1296) ?
                              reg1241[(4'h9):(2'h3)] : reg1262)) : ((reg1326[(2'h3):(1'h0)] ?
                              (reg1282 ?
                                  (8'ha8) : (8'had)) : forvar1265[(3'h6):(2'h3)]) ^~ reg1301));
                      reg1408 <= {{forvar1293}};
                      reg1409 <= $unsigned($unsigned($signed($signed(reg1342))));
                    end
                  if ((($signed($signed(reg1268)) >= ($signed(wire1224) ?
                          (~reg1311) : $unsigned((8'ha0)))) ?
                      {{reg1313}} : (~&$unsigned({reg1393}))))
                    begin
                      reg1410 <= $signed(forvar1265);
                      reg1411 <= (~^(($unsigned(forvar1260) ?
                          reg1244[(2'h3):(1'h0)] : $signed(forvar1225)) < reg1236));
                      reg1412 <= $unsigned(forvar1254);
                      reg1413 <= $unsigned((8'ha0));
                    end
                  else
                    begin
                      reg1410 <= reg1348;
                      reg1411 <= {(^(~|(-reg1372)))};
                      reg1412 <= (|$signed($signed($unsigned(reg1253))));
                    end
                  for (forvar1414 = (1'h0); (forvar1414 < (1'h0)); forvar1414 = (forvar1414 + (1'h1)))
                    begin
                      reg1415 <= $unsigned($signed(reg1242[(4'ha):(2'h2)]));
                      reg1416 <= $signed($signed($unsigned(reg1407[(3'h4):(1'h0)])));
                    end
                end
              reg1417 <= (8'ha8);
              for (forvar1418 = (1'h0); (forvar1418 < (1'h1)); forvar1418 = (forvar1418 + (1'h1)))
                begin
                  for (forvar1419 = (1'h0); (forvar1419 < (1'h0)); forvar1419 = (forvar1419 + (1'h1)))
                    begin
                      reg1420 <= (+forvar1343[(2'h3):(1'h1)]);
                      reg1421 <= $unsigned({(reg1361 ?
                              (reg1410 || (8'hb1)) : {forvar1286})});
                      reg1422 <= reg1304;
                    end
                  for (forvar1423 = (1'h0); (forvar1423 < (2'h2)); forvar1423 = (forvar1423 + (1'h1)))
                    begin
                      reg1424 <= ($unsigned({reg1411[(2'h3):(2'h3)]}) ?
                          ($signed((reg1415 ?
                              (8'hba) : reg1407)) * $signed((reg1403 <= forvar1293))) : (8'hb9));
                      reg1425 <= (~^($signed((^reg1231)) ?
                          (^$unsigned(wire1220)) : ((reg1261 ?
                              (8'had) : reg1306) & $unsigned(forvar1419))));
                    end
                  for (forvar1426 = (1'h0); (forvar1426 < (2'h3)); forvar1426 = (forvar1426 + (1'h1)))
                    begin
                      reg1427 <= $signed(forvar1371);
                      reg1428 <= ($unsigned({$unsigned(reg1420)}) ?
                          $signed($signed($unsigned(reg1332))) : forvar1225);
                    end
                  for (forvar1429 = (1'h0); (forvar1429 < (1'h1)); forvar1429 = (forvar1429 + (1'h1)))
                    begin
                      reg1430 <= $unsigned(($unsigned((forvar1337 ?
                          reg1275 : reg1409)) || $unsigned($signed(reg1265))));
                      reg1431 <= $signed($signed($unsigned($unsigned(forvar1324))));
                      reg1432 <= $signed({({(8'h9e)} ^~ reg1378)});
                    end
                end
            end
          for (forvar1433 = (1'h0); (forvar1433 < (1'h1)); forvar1433 = (forvar1433 + (1'h1)))
            begin
              if (forvar1317)
                begin
                  reg1434 <= $signed(($unsigned((8'hb9)) ?
                      {(|reg1241)} : ((8'ha9) ? reg1326 : reg1363)));
                  if (reg1416)
                    begin
                      reg1435 <= ({$unsigned((reg1341 ~^ reg1327))} ?
                          reg1257 : reg1327);
                      reg1436 <= $unsigned($signed(($signed(reg1306) >> (forvar1372 ?
                          reg1289 : reg1409))));
                      reg1437 <= (~^(~^forvar1226[(1'h0):(1'h0)]));
                      reg1438 <= {($unsigned((reg1244 - reg1378)) > reg1358[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg1435 <= reg1380[(3'h6):(3'h4)];
                    end
                end
              else
                begin
                  for (forvar1434 = (1'h0); (forvar1434 < (2'h2)); forvar1434 = (forvar1434 + (1'h1)))
                    begin
                      reg1435 <= forvar1419[(2'h3):(1'h0)];
                    end
                  for (forvar1436 = (1'h0); (forvar1436 < (1'h0)); forvar1436 = (forvar1436 + (1'h1)))
                    begin
                      reg1437 <= $unsigned(((~$unsigned(reg1315)) ?
                          (reg1373 >= $signed(wire1224)) : forvar1307));
                      reg1438 <= ($unsigned($unsigned(reg1422)) == reg1367[(4'hd):(4'h8)]);
                    end
                end
            end
        end
      else
        begin
          reg1370 <= {(~^wire1224[(2'h2):(2'h2)])};
          for (forvar1371 = (1'h0); (forvar1371 < (2'h2)); forvar1371 = (forvar1371 + (1'h1)))
            begin
              for (forvar1372 = (1'h0); (forvar1372 < (2'h3)); forvar1372 = (forvar1372 + (1'h1)))
                begin
                  if ($signed((~&(~^(-(8'hb5))))))
                    begin
                      reg1373 <= (reg1411 >= {reg1399[(2'h2):(1'h1)]});
                      reg1374 <= ((&(~reg1266)) ?
                          {reg1437} : forvar1353[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1373 <= (reg1395[(4'hb):(1'h1)] ?
                          $signed({((8'ha5) - reg1347)}) : reg1359[(2'h2):(2'h2)]);
                    end
                  if ((({$unsigned(forvar1378)} ?
                          {$signed(wire1284)} : (reg1264 && reg1352[(4'h8):(3'h6)])) ?
                      {($unsigned((8'hae)) | reg1397)} : ((&(forvar1235 ?
                          reg1432 : (8'ha0))) <= (forvar1269[(2'h2):(2'h2)] ?
                          (~&reg1272) : (reg1364 ? reg1236 : reg1415)))))
                    begin
                      reg1375 <= (&$unsigned($signed(forvar1286)));
                      reg1376 <= (|$signed(reg1294));
                    end
                  else
                    begin
                      reg1375 <= ((((~|reg1279) << reg1264[(1'h1):(1'h0)]) - ($signed(reg1372) ?
                              (wire1285 != reg1309) : $signed(forvar1372))) ?
                          reg1327 : $unsigned((-(^~reg1394))));
                      reg1376 <= ({{(forvar1239 ?
                                  reg1336 : reg1389)}} ^ forvar1405[(3'h4):(2'h2)]);
                      reg1377 <= $signed(((((8'ha1) & (8'ha5)) ?
                          reg1420 : (~^(8'hb1))) && (~^forvar1228)));
                    end
                  for (forvar1378 = (1'h0); (forvar1378 < (2'h2)); forvar1378 = (forvar1378 + (1'h1)))
                    begin
                      reg1379 <= reg1388[(1'h1):(1'h1)];
                    end
                  if (((8'hac) ?
                      reg1417[(2'h2):(1'h1)] : (-(reg1408[(4'hd):(3'h7)] ?
                          $unsigned(reg1253) : {wire1223}))))
                    begin
                      reg1380 <= (((-((8'had) ?
                              reg1271 : reg1246)) >= {forvar1307}) ?
                          $signed(($signed(reg1436) ?
                              (forvar1426 & reg1397) : $signed(reg1267))) : $signed(reg1353));
                      reg1381 <= (~|reg1410);
                      reg1382 <= (reg1339 ?
                          reg1435[(3'h4):(3'h4)] : forvar1414);
                      reg1383 <= (reg1434 ?
                          $unsigned(($unsigned(reg1344) & {reg1317})) : (reg1351[(2'h3):(2'h2)] ?
                              {(~^reg1340)} : $unsigned((forvar1363 ?
                                  (8'ha0) : reg1415))));
                    end
                  else
                    begin
                      reg1380 <= $unsigned($signed({$signed(reg1416)}));
                    end
                end
              if ((($unsigned($unsigned(reg1398)) ?
                      $signed($signed(reg1437)) : {$signed(reg1353)}) ?
                  (&reg1330[(3'h7):(1'h0)]) : (~wire1224)))
                begin
                  reg1384 <= $signed(reg1430);
                end
              else
                begin
                  if ((8'hb4))
                    begin
                      reg1384 <= $signed(reg1425);
                      reg1385 <= ({reg1378[(1'h0):(1'h0)]} - $unsigned($unsigned($unsigned(wire1224))));
                      reg1386 <= (-$unsigned($unsigned((+forvar1347))));
                      reg1387 <= $signed(reg1280);
                    end
                  else
                    begin
                      reg1384 <= forvar1319;
                    end
                  if (reg1310[(3'h4):(1'h0)])
                    begin
                      reg1388 <= $signed(reg1435[(3'h6):(3'h6)]);
                      reg1389 <= (8'haf);
                    end
                  else
                    begin
                      reg1388 <= $unsigned($signed(reg1232[(1'h1):(1'h1)]));
                      reg1389 <= $signed($unsigned(reg1275));
                      reg1390 <= $unsigned((^$signed(reg1359)));
                    end
                end
            end
          if (reg1249[(1'h0):(1'h0)])
            begin
              reg1391 <= ((~^forvar1405) * reg1299[(4'hc):(4'hb)]);
              if (((-$signed((reg1242 << forvar1366))) ?
                  reg1398 : (^~reg1236[(1'h0):(1'h0)])))
                begin
                  if (((((8'hb9) * (~|reg1363)) ^ reg1239) >> ({forvar1247[(4'hb):(4'ha)]} > ((&reg1317) ?
                      reg1341 : ((8'hae) >> reg1425)))))
                    begin
                      reg1392 <= (8'haa);
                      reg1393 <= reg1364;
                      reg1394 <= forvar1247;
                    end
                  else
                    begin
                      reg1392 <= reg1349;
                      reg1393 <= (((+$signed(reg1299)) ?
                          {(8'hb7)} : ((!wire1224) ?
                              {reg1350} : $signed(forvar1225))) - (forvar1248[(3'h7):(3'h4)] < $signed((+(8'hab)))));
                    end
                  for (forvar1395 = (1'h0); (forvar1395 < (1'h1)); forvar1395 = (forvar1395 + (1'h1)))
                    begin
                      reg1396 <= (reg1245 > reg1421);
                      reg1397 <= (~^reg1340);
                    end
                  for (forvar1398 = (1'h0); (forvar1398 < (2'h3)); forvar1398 = (forvar1398 + (1'h1)))
                    begin
                      reg1399 <= reg1339[(2'h2):(1'h1)];
                    end
                  for (forvar1400 = (1'h0); (forvar1400 < (2'h2)); forvar1400 = (forvar1400 + (1'h1)))
                    begin
                      reg1401 <= reg1283;
                      reg1402 <= $unsigned((^{(forvar1319 <<< reg1410)}));
                      reg1403 <= ((-$unsigned((8'ha2))) == $unsigned((^reg1376)));
                    end
                end
              else
                begin
                  for (forvar1392 = (1'h0); (forvar1392 < (2'h3)); forvar1392 = (forvar1392 + (1'h1)))
                    begin
                      reg1393 <= (!forvar1315[(2'h3):(2'h3)]);
                      reg1394 <= (8'hac);
                      reg1395 <= (reg1338[(2'h2):(1'h0)] << $unsigned($unsigned((reg1406 || (8'hb5)))));
                    end
                  reg1396 <= {{wire1284[(2'h2):(2'h2)]}};
                  for (forvar1397 = (1'h0); (forvar1397 < (1'h0)); forvar1397 = (forvar1397 + (1'h1)))
                    begin
                      reg1398 <= (8'hb6);
                    end
                end
              for (forvar1404 = (1'h0); (forvar1404 < (2'h2)); forvar1404 = (forvar1404 + (1'h1)))
                begin
                  if (((8'hae) && {reg1320}))
                    begin
                      reg1405 <= ((~&((wire1284 ?
                          reg1251 : reg1339) & $signed(reg1347))) <<< ((!reg1290) && (~^(8'ha6))));
                    end
                  else
                    begin
                      reg1405 <= (&$unsigned($signed($signed(forvar1337))));
                    end
                  if ($unsigned(forvar1236))
                    begin
                      reg1406 <= reg1235[(4'he):(4'h9)];
                    end
                  else
                    begin
                      reg1406 <= ((~^$unsigned((reg1397 >>> reg1367))) <<< (^~reg1389));
                      reg1407 <= $signed(reg1356);
                      reg1408 <= $signed($unsigned($unsigned(reg1403[(1'h0):(1'h0)])));
                    end
                end
              for (forvar1409 = (1'h0); (forvar1409 < (1'h1)); forvar1409 = (forvar1409 + (1'h1)))
                begin
                  for (forvar1410 = (1'h0); (forvar1410 < (2'h2)); forvar1410 = (forvar1410 + (1'h1)))
                    begin
                      reg1411 <= {((&(~^forvar1227)) ?
                              reg1333 : $signed($unsigned(reg1341)))};
                      reg1412 <= $signed(reg1245[(3'h7):(3'h4)]);
                      reg1413 <= reg1310[(4'hd):(4'ha)];
                    end
                  if (((~$signed((reg1261 ?
                      reg1340 : reg1380))) ^ ($unsigned((reg1233 + forvar1429)) ?
                      reg1290 : {(^forvar1255)})))
                    begin
                      reg1414 <= reg1316;
                      reg1415 <= reg1246[(1'h1):(1'h0)];
                      reg1416 <= $unsigned((~&(^~$unsigned(reg1387))));
                      reg1417 <= $signed($signed(reg1332[(2'h3):(2'h2)]));
                    end
                  else
                    begin
                      reg1414 <= (8'ha5);
                      reg1415 <= $signed($unsigned($signed((reg1347 ~^ reg1338))));
                      reg1416 <= ($signed(reg1341[(2'h3):(1'h1)]) ?
                          forvar1225 : $signed($signed((reg1323 ?
                              reg1318 : (8'hb0)))));
                    end
                end
            end
          else
            begin
              for (forvar1391 = (1'h0); (forvar1391 < (1'h0)); forvar1391 = (forvar1391 + (1'h1)))
                begin
                  if ((~|(~&(|$signed(reg1236)))))
                    begin
                      reg1392 <= $signed($unsigned($unsigned(reg1253[(2'h3):(1'h1)])));
                    end
                  else
                    begin
                      reg1392 <= (reg1321 && $signed($signed(forvar1239)));
                      reg1393 <= reg1228;
                    end
                  for (forvar1394 = (1'h0); (forvar1394 < (2'h3)); forvar1394 = (forvar1394 + (1'h1)))
                    begin
                      reg1395 <= ($signed(reg1346[(2'h2):(2'h2)]) ?
                          reg1435 : reg1385[(1'h0):(1'h0)]);
                    end
                  if (reg1382)
                    begin
                      reg1396 <= (~reg1427[(3'h4):(2'h3)]);
                      reg1397 <= {forvar1287};
                      reg1398 <= ({$unsigned((reg1402 ?
                                  reg1244 : forvar1402))} ?
                          ((reg1353[(2'h2):(1'h0)] >> {(8'ha6)}) & ($unsigned(reg1262) > (forvar1230 ?
                              forvar1319 : reg1298))) : (|$unsigned(reg1380[(4'h9):(1'h1)])));
                      reg1399 <= forvar1401[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1396 <= (8'hb4);
                      reg1397 <= reg1229[(3'h5):(1'h1)];
                    end
                end
              for (forvar1400 = (1'h0); (forvar1400 < (2'h2)); forvar1400 = (forvar1400 + (1'h1)))
                begin
                  reg1401 <= $unsigned((forvar1392[(1'h0):(1'h0)] <= {$signed(reg1425)}));
                end
              reg1402 <= $signed(forvar1226[(3'h6):(2'h3)]);
              if (reg1360)
                begin
                  reg1403 <= $signed((~|$unsigned($signed(reg1230))));
                  for (forvar1404 = (1'h0); (forvar1404 < (2'h2)); forvar1404 = (forvar1404 + (1'h1)))
                    begin
                      reg1405 <= (!$unsigned($unsigned(forvar1293)));
                      reg1406 <= forvar1228[(1'h0):(1'h0)];
                      reg1407 <= (~|(reg1250 ?
                          $signed((reg1422 + reg1249)) : ({reg1375} >>> reg1356[(2'h3):(2'h2)])));
                      reg1408 <= ({(8'hb6)} <<< (($unsigned(forvar1419) >>> $unsigned((8'hac))) || ((~^forvar1358) != $unsigned(forvar1372))));
                    end
                  for (forvar1409 = (1'h0); (forvar1409 < (1'h0)); forvar1409 = (forvar1409 + (1'h1)))
                    begin
                      reg1410 <= $unsigned($signed(forvar1391[(1'h1):(1'h0)]));
                    end
                  for (forvar1411 = (1'h0); (forvar1411 < (1'h1)); forvar1411 = (forvar1411 + (1'h1)))
                    begin
                      reg1412 <= $signed(reg1310);
                      reg1413 <= ($signed(reg1374) ^ (~|((reg1354 >= forvar1410) <= $unsigned(reg1375))));
                    end
                end
              else
                begin
                  reg1403 <= ((|{$unsigned(forvar1293)}) - (&(forvar1273 ^~ reg1346)));
                  for (forvar1404 = (1'h0); (forvar1404 < (2'h3)); forvar1404 = (forvar1404 + (1'h1)))
                    begin
                      reg1405 <= $signed(forvar1254);
                      reg1406 <= (&reg1369[(2'h2):(2'h2)]);
                      reg1407 <= (8'hab);
                    end
                  for (forvar1408 = (1'h0); (forvar1408 < (2'h3)); forvar1408 = (forvar1408 + (1'h1)))
                    begin
                      reg1409 <= {$signed((-forvar1337[(2'h2):(1'h1)]))};
                      reg1410 <= forvar1397;
                      reg1411 <= {forvar1338};
                    end
                  if ($signed(forvar1334))
                    begin
                      reg1412 <= $unsigned($signed(($unsigned(reg1391) ?
                          (~&(8'hb4)) : forvar1367[(2'h3):(2'h3)])));
                      reg1413 <= reg1289;
                      reg1414 <= $signed($unsigned(reg1409[(4'h9):(2'h3)]));
                      reg1415 <= $signed((-$unsigned(forvar1293)));
                    end
                  else
                    begin
                      reg1412 <= ((~(forvar1236 + $unsigned(forvar1414))) <<< reg1236[(2'h3):(2'h3)]);
                      reg1413 <= forvar1408;
                      reg1414 <= {($signed((forvar1273 | reg1380)) | reg1347[(1'h1):(1'h1)])};
                      reg1415 <= $signed(reg1298[(1'h1):(1'h0)]);
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1439 = (1'h0); (forvar1439 < (1'h1)); forvar1439 = (forvar1439 + (1'h1)))
        begin
          reg1440 <= {forvar1226};
          if (reg1316[(3'h5):(2'h3)])
            begin
              if (reg1354)
                begin
                  for (forvar1441 = (1'h0); (forvar1441 < (1'h1)); forvar1441 = (forvar1441 + (1'h1)))
                    begin
                      reg1442 <= $unsigned(wire1284[(2'h3):(2'h2)]);
                      reg1443 <= ((forvar1344[(4'hc):(2'h2)] || $unsigned(forvar1278[(4'h8):(1'h1)])) && (+((reg1366 ?
                              reg1306 : reg1239) ?
                          {reg1407} : (!reg1386))));
                    end
                  for (forvar1444 = (1'h0); (forvar1444 < (2'h3)); forvar1444 = (forvar1444 + (1'h1)))
                    begin
                      reg1445 <= reg1432;
                      reg1446 <= ((($unsigned(reg1357) ?
                                  (reg1375 ?
                                      reg1438 : forvar1239) : $unsigned(forvar1225)) ?
                              $unsigned(reg1436[(4'ha):(2'h3)]) : reg1411) ?
                          (($unsigned(forvar1286) ?
                                  $unsigned(forvar1287) : (reg1276 - (8'hb1))) ?
                              ($signed(reg1238) ?
                                  (8'hb5) : (reg1313 ?
                                      wire1220 : reg1267)) : ({reg1295} ?
                                  {(8'hb3)} : $unsigned(reg1379))) : $unsigned($signed((reg1308 ~^ reg1270))));
                      reg1447 <= (+reg1432[(1'h1):(1'h1)]);
                    end
                  reg1448 <= reg1394[(2'h2):(2'h2)];
                  if (reg1422[(3'h5):(2'h3)])
                    begin
                      reg1449 <= ((-($unsigned(reg1345) ?
                              $signed(reg1321) : {reg1416})) ?
                          ($signed((forvar1232 ? (8'ha0) : forvar1255)) ?
                              (reg1232[(2'h2):(1'h1)] ?
                                  reg1346[(4'h8):(3'h7)] : forvar1311) : ($signed(reg1375) ^ (forvar1398 ?
                                  forvar1397 : reg1368))) : forvar1226[(3'h6):(3'h4)]);
                      reg1450 <= reg1398[(2'h3):(2'h3)];
                      reg1451 <= forvar1426;
                      reg1452 <= {$unsigned($unsigned(forvar1395))};
                    end
                  else
                    begin
                      reg1449 <= $signed($unsigned($unsigned((|reg1401))));
                      reg1450 <= $signed(($signed($signed(reg1327)) || reg1289));
                      reg1451 <= $unsigned((!((reg1438 ?
                          reg1370 : reg1357) ^~ reg1314)));
                      reg1452 <= {(~&((reg1436 ^ forvar1366) ?
                              (reg1396 ? reg1422 : reg1408) : {reg1346}))};
                    end
                end
              else
                begin
                  for (forvar1441 = (1'h0); (forvar1441 < (1'h1)); forvar1441 = (forvar1441 + (1'h1)))
                    begin
                      reg1442 <= {$unsigned($unsigned(reg1263))};
                      reg1443 <= $signed($signed({forvar1363[(3'h6):(1'h0)]}));
                      reg1444 <= (((reg1272[(1'h1):(1'h1)] >= reg1415[(3'h4):(2'h2)]) ?
                              (~^forvar1394[(4'h8):(1'h1)]) : (!((8'ha0) ?
                                  wire1222 : reg1358))) ?
                          $unsigned($unsigned(reg1372[(2'h3):(2'h2)])) : forvar1353[(1'h0):(1'h0)]);
                      reg1445 <= $signed($unsigned(reg1367));
                    end
                  if (reg1445)
                    begin
                      reg1446 <= reg1368[(1'h0):(1'h0)];
                      reg1447 <= ($unsigned(reg1305) > reg1232[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg1446 <= reg1351;
                    end
                  if ($signed((reg1308[(2'h3):(1'h0)] <<< reg1403[(3'h7):(3'h5)])))
                    begin
                      reg1448 <= ((~$unsigned((forvar1411 ?
                          reg1402 : wire1285))) ~^ (8'h9e));
                      reg1449 <= (forvar1371 <<< reg1431[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg1448 <= forvar1319[(1'h0):(1'h0)];
                      reg1449 <= (~^$unsigned($signed((~^reg1399))));
                      reg1450 <= $unsigned(forvar1371[(4'hc):(2'h3)]);
                    end
                end
              if ($unsigned(forvar1278))
                begin
                  if ($unsigned($signed(reg1306)))
                    begin
                      reg1453 <= (reg1422 | ((reg1408[(1'h1):(1'h0)] | (~|reg1375)) ?
                          reg1253 : ($signed(reg1359) > (forvar1391 ^~ reg1267))));
                      reg1454 <= ((wire1224[(1'h0):(1'h0)] ?
                          ({reg1351} != {forvar1441}) : $signed((reg1279 & reg1431))) & {($signed(forvar1286) ?
                              (reg1375 + reg1453) : (~&(8'h9c)))});
                      reg1455 <= (|(~|$unsigned((reg1259 ?
                          reg1388 : forvar1394))));
                    end
                  else
                    begin
                      reg1453 <= (~&($unsigned((8'hba)) ?
                          $signed({reg1241}) : ($unsigned(reg1454) ?
                              forvar1286 : {reg1266})));
                      reg1454 <= (reg1351 ?
                          ($signed({reg1257}) | (8'hae)) : {reg1323[(3'h4):(1'h1)]});
                      reg1455 <= ((reg1415 >= $unsigned($signed(forvar1319))) ?
                          $unsigned(forvar1273) : $signed(((reg1344 >>> forvar1243) ?
                              $unsigned(reg1244) : {forvar1225})));
                    end
                  reg1456 <= (8'hb5);
                  reg1457 <= reg1380;
                end
              else
                begin
                  for (forvar1453 = (1'h0); (forvar1453 < (1'h1)); forvar1453 = (forvar1453 + (1'h1)))
                    begin
                      reg1454 <= reg1338;
                    end
                end
              reg1458 <= $unsigned((reg1289 * {reg1395}));
            end
          else
            begin
              for (forvar1441 = (1'h0); (forvar1441 < (1'h1)); forvar1441 = (forvar1441 + (1'h1)))
                begin
                  if (((reg1420 || (~^$unsigned(forvar1344))) ^ (-forvar1366[(1'h0):(1'h0)])))
                    begin
                      reg1442 <= reg1416[(2'h3):(1'h1)];
                      reg1443 <= (~&((reg1239 ^ forvar1418[(3'h6):(3'h5)]) < (~|reg1428)));
                    end
                  else
                    begin
                      reg1442 <= (!((forvar1230 ?
                          $unsigned(reg1241) : {forvar1288}) && reg1392[(1'h0):(1'h0)]));
                      reg1443 <= $unsigned(($signed((~^reg1393)) ?
                          forvar1409 : reg1289[(2'h2):(1'h0)]));
                    end
                  for (forvar1444 = (1'h0); (forvar1444 < (1'h0)); forvar1444 = (forvar1444 + (1'h1)))
                    begin
                      reg1445 <= (reg1431 ?
                          (-reg1421[(1'h1):(1'h0)]) : forvar1311);
                      reg1446 <= (reg1336[(4'h8):(2'h3)] * ($signed($unsigned(reg1428)) ?
                          reg1364[(4'hb):(3'h4)] : (+reg1411)));
                    end
                  if ((-forvar1338[(4'h8):(3'h5)]))
                    begin
                      reg1447 <= reg1372[(3'h5):(2'h3)];
                      reg1448 <= reg1251[(4'hc):(3'h5)];
                      reg1449 <= (^reg1266[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1447 <= $signed(($unsigned((8'hb1)) ^~ (^reg1258)));
                      reg1448 <= $signed((8'hac));
                      reg1449 <= reg1290;
                    end
                  if (((((-reg1427) >= $unsigned(reg1271)) || reg1444) ~^ {$unsigned($unsigned(wire1285))}))
                    begin
                      reg1450 <= ({$signed($signed(forvar1311))} ?
                          $unsigned(forvar1409[(1'h0):(1'h0)]) : (~|({reg1437} >= (reg1249 ?
                              forvar1426 : (8'hb0)))));
                      reg1451 <= $unsigned(reg1385);
                      reg1452 <= (forvar1338 ?
                          reg1384[(1'h0):(1'h0)] : $unsigned($signed(reg1358)));
                    end
                  else
                    begin
                      reg1450 <= ((~(|(~|reg1279))) || (~^(reg1319 & $signed(forvar1429))));
                      reg1451 <= ((forvar1376[(4'hc):(3'h4)] ~^ forvar1419[(2'h3):(1'h0)]) ?
                          $unsigned((^~(8'hae))) : (({wire1222} ?
                                  $unsigned(reg1235) : reg1454) ?
                              ($signed(reg1244) < (forvar1433 ^ reg1349)) : $unsigned((reg1311 ?
                                  reg1264 : reg1310))));
                      reg1452 <= $unsigned(forvar1395);
                      reg1453 <= {$signed($unsigned(((8'hb7) ^ reg1411)))};
                    end
                end
              reg1454 <= $unsigned(($signed(reg1300) ?
                  $signed({reg1339}) : (~reg1259[(2'h3):(1'h0)])));
            end
          for (forvar1459 = (1'h0); (forvar1459 < (1'h1)); forvar1459 = (forvar1459 + (1'h1)))
            begin
              for (forvar1460 = (1'h0); (forvar1460 < (1'h0)); forvar1460 = (forvar1460 + (1'h1)))
                begin
                  for (forvar1461 = (1'h0); (forvar1461 < (1'h1)); forvar1461 = (forvar1461 + (1'h1)))
                    begin
                      reg1462 <= {{{{reg1413}}}};
                      reg1463 <= {(+$unsigned(reg1317[(4'hf):(4'h8)]))};
                    end
                end
              for (forvar1464 = (1'h0); (forvar1464 < (2'h2)); forvar1464 = (forvar1464 + (1'h1)))
                begin
                  reg1465 <= reg1437;
                  for (forvar1466 = (1'h0); (forvar1466 < (1'h1)); forvar1466 = (forvar1466 + (1'h1)))
                    begin
                      reg1467 <= $signed(((+(forvar1378 ? reg1290 : reg1251)) ?
                          {forvar1255} : forvar1239[(4'he):(3'h7)]));
                      reg1468 <= {(|reg1265)};
                    end
                  for (forvar1469 = (1'h0); (forvar1469 < (2'h2)); forvar1469 = (forvar1469 + (1'h1)))
                    begin
                      reg1470 <= $signed($unsigned($signed(reg1258)));
                      reg1471 <= $signed($signed(((^forvar1363) | $signed(forvar1434))));
                    end
                end
              for (forvar1472 = (1'h0); (forvar1472 < (1'h0)); forvar1472 = (forvar1472 + (1'h1)))
                begin
                  for (forvar1473 = (1'h0); (forvar1473 < (1'h0)); forvar1473 = (forvar1473 + (1'h1)))
                    begin
                      reg1474 <= (($unsigned(reg1445) ?
                          $unsigned((reg1282 ~^ (8'haf))) : ((|(8'hb3)) | ((8'ha2) || forvar1472))) != ((8'hb6) | $signed((reg1376 ?
                          reg1405 : reg1449))));
                      reg1475 <= reg1321[(2'h2):(1'h1)];
                    end
                  for (forvar1476 = (1'h0); (forvar1476 < (2'h3)); forvar1476 = (forvar1476 + (1'h1)))
                    begin
                      reg1477 <= $unsigned((reg1414[(1'h0):(1'h0)] ?
                          (~&(^reg1410)) : $signed((~reg1407))));
                    end
                  reg1478 <= reg1413;
                end
              if ((8'had))
                begin
                  for (forvar1479 = (1'h0); (forvar1479 < (2'h3)); forvar1479 = (forvar1479 + (1'h1)))
                    begin
                      reg1480 <= (~reg1290[(1'h1):(1'h0)]);
                      reg1481 <= $signed(reg1309);
                      reg1482 <= ($signed(((reg1405 >>> forvar1466) ?
                          {reg1386} : (forvar1405 ?
                              reg1463 : forvar1239))) || $unsigned($signed((!reg1290))));
                    end
                end
              else
                begin
                  for (forvar1479 = (1'h0); (forvar1479 < (2'h3)); forvar1479 = (forvar1479 + (1'h1)))
                    begin
                      reg1480 <= forvar1334[(3'h7):(3'h5)];
                      reg1481 <= ((~^$unsigned(reg1362[(2'h2):(1'h0)])) ?
                          (~|(((8'hba) * reg1427) | $signed(forvar1337))) : (-forvar1479));
                      reg1482 <= ((forvar1444[(3'h4):(2'h2)] - reg1405[(3'h4):(1'h0)]) ?
                          $unsigned((8'h9d)) : (~&reg1313));
                      reg1483 <= (forvar1236[(1'h0):(1'h0)] <= (((reg1343 >> reg1332) <= forvar1269) >>> reg1451));
                    end
                  for (forvar1484 = (1'h0); (forvar1484 < (1'h1)); forvar1484 = (forvar1484 + (1'h1)))
                    begin
                      reg1485 <= (~forvar1472);
                      reg1486 <= $signed(reg1303);
                      reg1487 <= $signed({(|(forvar1312 ?
                              forvar1228 : forvar1265))});
                    end
                end
            end
          if (reg1399[(3'h6):(3'h5)])
            begin
              if (forvar1401[(1'h0):(1'h0)])
                begin
                  for (forvar1488 = (1'h0); (forvar1488 < (1'h0)); forvar1488 = (forvar1488 + (1'h1)))
                    begin
                      reg1489 <= $unsigned({(reg1321 || reg1482[(1'h0):(1'h0)])});
                    end
                  for (forvar1490 = (1'h0); (forvar1490 < (1'h0)); forvar1490 = (forvar1490 + (1'h1)))
                    begin
                      reg1491 <= reg1463;
                      reg1492 <= reg1318;
                      reg1493 <= reg1384;
                      reg1494 <= wire1222[(3'h4):(3'h4)];
                    end
                  reg1495 <= ($unsigned(($unsigned(reg1405) < $signed(reg1428))) ?
                      $signed($unsigned($signed(reg1276))) : forvar1408);
                  for (forvar1496 = (1'h0); (forvar1496 < (2'h3)); forvar1496 = (forvar1496 + (1'h1)))
                    begin
                      reg1497 <= $unsigned(($signed((reg1250 ?
                          reg1443 : reg1372)) >= $signed(reg1414)));
                      reg1498 <= (|$unsigned(((forvar1255 ?
                          forvar1397 : reg1335) == $unsigned(reg1267))));
                      reg1499 <= reg1359[(3'h4):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar1488 = (1'h0); (forvar1488 < (1'h1)); forvar1488 = (forvar1488 + (1'h1)))
                    begin
                      reg1489 <= reg1438[(1'h0):(1'h0)];
                      reg1490 <= (8'hb1);
                    end
                end
            end
          else
            begin
              for (forvar1488 = (1'h0); (forvar1488 < (1'h0)); forvar1488 = (forvar1488 + (1'h1)))
                begin
                  for (forvar1489 = (1'h0); (forvar1489 < (2'h3)); forvar1489 = (forvar1489 + (1'h1)))
                    begin
                      reg1490 <= $unsigned($unsigned(($unsigned(reg1395) <<< forvar1278)));
                      reg1491 <= {(8'hb2)};
                      reg1492 <= $unsigned((8'hb5));
                    end
                  for (forvar1493 = (1'h0); (forvar1493 < (2'h3)); forvar1493 = (forvar1493 + (1'h1)))
                    begin
                      reg1494 <= {$unsigned(($signed(forvar1466) ?
                              (forvar1248 ? (8'ha6) : reg1491) : (~|reg1481)))};
                      reg1495 <= reg1396;
                      reg1496 <= reg1349[(3'h5):(1'h1)];
                    end
                end
              if ($signed((8'hb9)))
                begin
                  if ((8'ha9))
                    begin
                      reg1497 <= ($signed((~^$signed(wire1221))) <= reg1405[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg1497 <= (((&(forvar1398 ?
                              forvar1235 : reg1309)) | {(reg1270 == reg1227)}) ?
                          forvar1460[(3'h7):(1'h1)] : $signed(forvar1411));
                      reg1498 <= (&$unsigned(reg1410[(2'h2):(2'h2)]));
                      reg1499 <= (8'hb0);
                      reg1500 <= reg1436;
                    end
                  if (reg1500)
                    begin
                      reg1501 <= (((+(forvar1395 ?
                              reg1344 : reg1403)) && $signed(forvar1472[(4'h9):(2'h3)])) ?
                          $signed((^(^(8'ha9)))) : forvar1489[(1'h0):(1'h0)]);
                      reg1502 <= $unsigned(reg1335);
                      reg1503 <= forvar1312[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1501 <= {wire1284[(2'h2):(1'h0)]};
                      reg1502 <= ($unsigned((^~(~|forvar1444))) ?
                          $signed(((reg1462 < forvar1378) ?
                              $signed(forvar1409) : $unsigned((8'hab)))) : $unsigned(reg1244[(3'h7):(1'h0)]));
                      reg1503 <= $unsigned((reg1477 <= $signed(reg1326)));
                    end
                  reg1504 <= forvar1464[(4'h9):(3'h4)];
                end
              else
                begin
                  for (forvar1497 = (1'h0); (forvar1497 < (1'h1)); forvar1497 = (forvar1497 + (1'h1)))
                    begin
                      reg1498 <= (((!(+reg1391)) ?
                          {reg1391[(4'ha):(3'h7)]} : reg1322[(4'hf):(4'h9)]) <= $signed(((^~reg1321) ?
                          $signed(forvar1466) : (forvar1479 | (8'had)))));
                      reg1499 <= ({({reg1435} <<< (reg1482 & (8'hb3)))} << reg1344[(4'hb):(3'h5)]);
                      reg1500 <= $signed((~^$signed((forvar1273 ?
                          reg1463 : reg1342))));
                    end
                  reg1501 <= (!((!((8'ha4) ? reg1250 : reg1405)) ?
                      (((8'hb1) ? reg1232 : reg1420) ?
                          reg1283[(4'h8):(1'h1)] : $unsigned((8'ha2))) : (8'ha4)));
                end
            end
        end
      reg1505 <= $signed($unsigned($unsigned($unsigned((8'h9f)))));
      if ($unsigned(reg1454[(2'h3):(2'h3)]))
        begin
          reg1506 <= ({(reg1342[(3'h6):(3'h4)] ?
                  reg1395[(3'h4):(2'h3)] : (reg1325 >>> forvar1232))} >>> forvar1320);
          for (forvar1507 = (1'h0); (forvar1507 < (2'h2)); forvar1507 = (forvar1507 + (1'h1)))
            begin
              if (((({reg1230} ? (reg1422 + reg1338) : $signed(reg1238)) ?
                      forvar1489 : $unsigned((reg1309 ? reg1486 : reg1325))) ?
                  ({(reg1493 ?
                          reg1442 : reg1270)} <= (-$unsigned((8'ha9)))) : ((8'hb4) + $signed((reg1295 ?
                      forvar1419 : reg1283)))))
                begin
                  reg1508 <= $unsigned(reg1443);
                  for (forvar1509 = (1'h0); (forvar1509 < (1'h1)); forvar1509 = (forvar1509 + (1'h1)))
                    begin
                      reg1510 <= forvar1459[(1'h0):(1'h0)];
                      reg1511 <= $signed(((((8'h9e) ?
                              forvar1383 : forvar1337) ^~ (reg1332 * reg1483)) ?
                          ($signed(reg1380) ?
                              wire1223 : $signed(forvar1409)) : (((8'ha3) >>> reg1265) != reg1442)));
                      reg1512 <= $signed((($unsigned((8'ha0)) ?
                              {reg1333} : $unsigned(reg1417)) ?
                          ($signed(forvar1274) ?
                              (reg1399 >>> reg1239) : (reg1341 && reg1275)) : reg1297[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar1508 = (1'h0); (forvar1508 < (2'h3)); forvar1508 = (forvar1508 + (1'h1)))
                    begin
                      reg1509 <= reg1386;
                      reg1510 <= $signed($unsigned(reg1281[(3'h4):(3'h4)]));
                      reg1511 <= reg1271[(1'h0):(1'h0)];
                    end
                end
              if (reg1349)
                begin
                  if ((^~{$unsigned($unsigned((8'haa)))}))
                    begin
                      reg1513 <= reg1449;
                      reg1514 <= reg1364;
                      reg1515 <= reg1446;
                      reg1516 <= ($signed($unsigned((reg1270 ^ reg1347))) ?
                          $unsigned(reg1339[(2'h2):(2'h2)]) : (+wire1223[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg1513 <= reg1442;
                      reg1514 <= (-($signed((^reg1242)) < reg1493[(3'h4):(2'h3)]));
                    end
                  if ((8'ha5))
                    begin
                      reg1517 <= reg1451;
                    end
                  else
                    begin
                      reg1517 <= (~&(~&$unsigned(forvar1343)));
                      reg1518 <= $unsigned((reg1363 ?
                          {forvar1391[(3'h6):(3'h4)]} : forvar1288));
                    end
                  for (forvar1519 = (1'h0); (forvar1519 < (2'h3)); forvar1519 = (forvar1519 + (1'h1)))
                    begin
                      reg1520 <= forvar1358;
                    end
                  for (forvar1521 = (1'h0); (forvar1521 < (1'h1)); forvar1521 = (forvar1521 + (1'h1)))
                    begin
                      reg1522 <= (!(~|(8'hb8)));
                    end
                end
              else
                begin
                  if ((8'hb1))
                    begin
                      reg1513 <= forvar1235;
                      reg1514 <= {(^$unsigned($unsigned(reg1340)))};
                      reg1515 <= $signed({wire1220});
                      reg1516 <= reg1250;
                    end
                  else
                    begin
                      reg1513 <= {$unsigned(($signed(forvar1509) + $unsigned(reg1297)))};
                      reg1514 <= $signed(({(reg1490 ? (8'hb7) : (8'hab))} ?
                          ($unsigned(reg1304) == (reg1244 == reg1242)) : $signed(((8'hb2) <= reg1470))));
                    end
                  if ((|($signed((^~(8'hab))) ?
                      ($unsigned(forvar1419) ?
                          (reg1359 ?
                              (8'ha6) : (8'hb3)) : {reg1415}) : ((forvar1366 ?
                          reg1435 : forvar1302) >> $signed(reg1333)))))
                    begin
                      reg1517 <= $signed(((forvar1402 == (reg1463 ?
                          reg1401 : reg1504)) & reg1333));
                      reg1518 <= ((reg1358[(4'h8):(4'h8)] <<< reg1471[(4'ha):(1'h1)]) ?
                          (!reg1508) : $unsigned(($signed(forvar1401) > {(8'h9f)})));
                      reg1519 <= (^($signed({forvar1507}) ?
                          (|$signed(forvar1320)) : $signed($unsigned((8'h9f)))));
                    end
                  else
                    begin
                      reg1517 <= (|$unsigned($unsigned($unsigned(reg1289))));
                      reg1518 <= $signed(reg1474);
                    end
                  for (forvar1520 = (1'h0); (forvar1520 < (2'h2)); forvar1520 = (forvar1520 + (1'h1)))
                    begin
                      reg1521 <= (~^($unsigned(((8'h9d) && (8'hb2))) ?
                          $unsigned((reg1240 ?
                              reg1454 : forvar1410)) : reg1369[(4'h9):(3'h4)]));
                      reg1522 <= forvar1397;
                      reg1523 <= (reg1330 ?
                          ((8'hb0) || $signed((~&(8'had)))) : (($unsigned(reg1370) ?
                              ((8'hb3) ?
                                  forvar1243 : reg1336) : $unsigned(forvar1433)) <<< $signed(forvar1355[(3'h5):(1'h1)])));
                    end
                  for (forvar1524 = (1'h0); (forvar1524 < (2'h3)); forvar1524 = (forvar1524 + (1'h1)))
                    begin
                      reg1525 <= (^reg1497[(1'h1):(1'h0)]);
                      reg1526 <= (^{$signed($signed(reg1407))});
                      reg1527 <= ((~&(reg1275 ?
                          $signed(reg1495) : reg1392)) < (-(!((8'ha3) ?
                          reg1319 : reg1458))));
                    end
                end
              if (reg1465)
                begin
                  reg1528 <= (8'had);
                  for (forvar1529 = (1'h0); (forvar1529 < (2'h3)); forvar1529 = (forvar1529 + (1'h1)))
                    begin
                      reg1530 <= $signed(forvar1397);
                      reg1531 <= $unsigned($signed(($unsigned((8'ha5)) >> ((8'hba) ?
                          forvar1311 : (8'h9c)))));
                    end
                  if (forvar1488)
                    begin
                      reg1532 <= ($signed(forvar1439[(2'h2):(2'h2)]) ?
                          $unsigned($unsigned({reg1315})) : (((forvar1414 ?
                              reg1345 : reg1295) - (~forvar1320)) || reg1271));
                      reg1533 <= $unsigned(reg1390);
                      reg1534 <= {(($signed(forvar1423) ?
                              reg1501[(2'h3):(2'h3)] : $unsigned(reg1251)) * ((reg1445 ?
                              (8'hb9) : reg1457) <= $signed(reg1527)))};
                      reg1535 <= {(&$unsigned(reg1428))};
                    end
                  else
                    begin
                      reg1532 <= reg1387;
                      reg1533 <= (((reg1265 | $signed(reg1320)) <= forvar1324[(1'h0):(1'h0)]) ?
                          (8'hae) : $signed(reg1502[(1'h0):(1'h0)]));
                      reg1534 <= ((~^($signed((8'ha2)) ?
                              reg1404[(2'h3):(1'h0)] : reg1374)) ?
                          ((((8'ha5) ?
                              reg1316 : forvar1507) ^ (reg1275 || forvar1398)) != (~&$signed(forvar1311))) : (&((!reg1237) || $signed(reg1398))));
                      reg1535 <= $signed(reg1364);
                    end
                end
              else
                begin
                  if (((forvar1247 ~^ $signed(reg1297)) ?
                      $signed($unsigned((8'ha0))) : (forvar1311[(2'h2):(1'h0)] >>> $unsigned(((8'h9f) ?
                          wire1284 : reg1414)))))
                    begin
                      reg1528 <= (~|$unsigned($unsigned((!reg1365))));
                      reg1529 <= ({reg1335} ?
                          reg1261 : $signed($unsigned((reg1348 > forvar1444))));
                      reg1530 <= (~&{reg1386});
                      reg1531 <= reg1341[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg1528 <= (8'ha8);
                      reg1529 <= (8'haf);
                    end
                  if ((^$signed((^((8'h9d) && reg1528)))))
                    begin
                      reg1532 <= $unsigned((forvar1524[(3'h4):(2'h3)] + $unsigned($unsigned(reg1528))));
                    end
                  else
                    begin
                      reg1532 <= $unsigned((-reg1497));
                      reg1533 <= (^~reg1327[(1'h1):(1'h1)]);
                      reg1534 <= $unsigned($signed($unsigned((wire1221 ?
                          reg1359 : reg1335))));
                      reg1535 <= $signed(forvar1460[(4'hb):(3'h7)]);
                    end
                  if (forvar1466)
                    begin
                      reg1536 <= $unsigned(reg1521);
                    end
                  else
                    begin
                      reg1536 <= (&(reg1315 ?
                          reg1443[(3'h5):(1'h1)] : (reg1316 ?
                              (reg1380 << reg1515) : (8'hb2))));
                      reg1537 <= reg1251[(3'h6):(3'h6)];
                    end
                end
            end
          for (forvar1538 = (1'h0); (forvar1538 < (1'h0)); forvar1538 = (forvar1538 + (1'h1)))
            begin
              reg1539 <= {$signed($signed($signed(reg1509)))};
            end
        end
      else
        begin
          for (forvar1506 = (1'h0); (forvar1506 < (1'h0)); forvar1506 = (forvar1506 + (1'h1)))
            begin
              if (($signed({(^reg1505)}) ? reg1265[(1'h0):(1'h0)] : reg1402))
                begin
                  reg1507 <= ((!$unsigned(reg1405)) < forvar1488[(2'h3):(2'h2)]);
                  if (forvar1302[(1'h1):(1'h0)])
                    begin
                      reg1508 <= reg1504[(3'h5):(2'h2)];
                      reg1509 <= $signed((~(!$signed(reg1434))));
                    end
                  else
                    begin
                      reg1508 <= ((+{$signed(reg1282)}) ?
                          (forvar1239[(4'hf):(2'h3)] | (|(reg1413 ?
                              reg1492 : reg1402))) : $unsigned(reg1509));
                      reg1509 <= $unsigned($signed($signed((!reg1496))));
                    end
                end
              else
                begin
                  for (forvar1507 = (1'h0); (forvar1507 < (1'h1)); forvar1507 = (forvar1507 + (1'h1)))
                    begin
                      reg1508 <= ($signed((reg1325[(4'h9):(4'h8)] ?
                          {reg1414} : reg1249[(1'h0):(1'h0)])) + reg1445[(4'h8):(3'h6)]);
                      reg1509 <= (-(~reg1492));
                    end
                end
              reg1510 <= ((!reg1537) > forvar1461);
            end
        end
      for (forvar1540 = (1'h0); (forvar1540 < (1'h0)); forvar1540 = (forvar1540 + (1'h1)))
        begin
          reg1541 <= (reg1304 ?
              (!(forvar1444 ?
                  (+reg1354) : $signed(forvar1395))) : $unsigned((~|$unsigned(forvar1286))));
          if ($signed((({reg1240} & $unsigned(forvar1353)) ?
              reg1350 : (~&(-reg1414)))))
            begin
              reg1542 <= $unsigned((8'hb6));
              for (forvar1543 = (1'h0); (forvar1543 < (2'h2)); forvar1543 = (forvar1543 + (1'h1)))
                begin
                  if ($unsigned($unsigned(reg1236[(1'h1):(1'h1)])))
                    begin
                      reg1544 <= $signed(reg1386[(2'h3):(1'h0)]);
                      reg1545 <= ($signed((~|(&reg1425))) <= ($signed((~&(8'ha1))) && reg1318));
                      reg1546 <= forvar1473;
                    end
                  else
                    begin
                      reg1544 <= $unsigned(({$signed((8'hb4))} >= (|forvar1426[(1'h0):(1'h0)])));
                      reg1545 <= ((forvar1243 <= (^$unsigned(reg1539))) >> ({(reg1442 && reg1503)} || {(reg1409 ?
                              reg1482 : reg1344)}));
                      reg1546 <= $unsigned($signed($signed(reg1447)));
                    end
                  for (forvar1547 = (1'h0); (forvar1547 < (2'h2)); forvar1547 = (forvar1547 + (1'h1)))
                    begin
                      reg1548 <= (~&(|(|(reg1282 ~^ reg1521))));
                      reg1549 <= {$signed(((forvar1433 ?
                              forvar1524 : forvar1372) <<< (forvar1347 ^~ reg1416)))};
                    end
                end
              if (((((|reg1338) - (~&(8'ha0))) ? reg1375 : reg1427) ?
                  $unsigned($signed((reg1533 ?
                      reg1468 : reg1539))) : forvar1293[(1'h1):(1'h0)]))
                begin
                  if (reg1516)
                    begin
                      reg1550 <= (!{$unsigned(reg1279)});
                      reg1551 <= $unsigned(($unsigned((forvar1464 & reg1352)) <<< {(~&(8'h9f))}));
                    end
                  else
                    begin
                      reg1550 <= ((((reg1401 ?
                              (8'h9c) : reg1408) >> (~reg1312)) & reg1249[(1'h0):(1'h0)]) ?
                          (~(reg1448[(1'h0):(1'h0)] ?
                              (!wire1221) : (reg1509 ?
                                  reg1239 : (8'haf)))) : ($unsigned(forvar1419) >> $signed((|forvar1239))));
                    end
                  reg1552 <= reg1405;
                end
              else
                begin
                  for (forvar1550 = (1'h0); (forvar1550 < (1'h1)); forvar1550 = (forvar1550 + (1'h1)))
                    begin
                      reg1551 <= (((&(reg1390 ? (8'h9f) : reg1250)) ?
                          $unsigned(reg1364[(4'h8):(2'h2)]) : $signed((reg1306 ?
                              reg1527 : forvar1466))) ~^ (|reg1389[(2'h2):(2'h2)]));
                      reg1552 <= ($unsigned((reg1454 > (reg1548 ?
                          reg1450 : reg1369))) & reg1369[(1'h1):(1'h1)]);
                      reg1553 <= {(((forvar1493 ^~ (8'ha7)) ?
                                  $signed(forvar1466) : (forvar1488 ?
                                      reg1417 : reg1517)) ?
                              reg1414[(2'h3):(1'h0)] : $signed($unsigned(forvar1383)))};
                    end
                  if (($unsigned($signed((^~forvar1418))) ~^ reg1309[(3'h5):(3'h4)]))
                    begin
                      reg1554 <= $unsigned((!((8'ha4) ?
                          forvar1404[(1'h1):(1'h1)] : ((8'h9f) >>> (8'ha7)))));
                      reg1555 <= (!forvar1328[(4'ha):(3'h6)]);
                      reg1556 <= reg1233[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1554 <= (8'ha4);
                      reg1555 <= $signed({reg1492});
                      reg1556 <= (^$unsigned((reg1294 ?
                          $unsigned(reg1342) : $signed(reg1344))));
                    end
                  if ($unsigned($unsigned((forvar1343[(4'ha):(2'h2)] < reg1405[(3'h6):(3'h4)]))))
                    begin
                      reg1557 <= forvar1519[(4'ha):(2'h2)];
                      reg1558 <= $signed((~$unsigned($signed(forvar1459))));
                    end
                  else
                    begin
                      reg1557 <= $signed($unsigned((!$unsigned(reg1482))));
                      reg1558 <= reg1351[(2'h2):(2'h2)];
                      reg1559 <= (&$signed($unsigned($unsigned(reg1425))));
                      reg1560 <= reg1372;
                    end
                  if ((8'hb9))
                    begin
                      reg1561 <= (^($unsigned({reg1435}) >= reg1322[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg1561 <= reg1493;
                      reg1562 <= ($signed($signed($signed((8'h9e)))) ^ {(8'h9c)});
                    end
                end
            end
          else
            begin
              for (forvar1542 = (1'h0); (forvar1542 < (2'h3)); forvar1542 = (forvar1542 + (1'h1)))
                begin
                  for (forvar1543 = (1'h0); (forvar1543 < (1'h1)); forvar1543 = (forvar1543 + (1'h1)))
                    begin
                      reg1544 <= ((forvar1273[(1'h1):(1'h0)] ?
                          $signed((reg1396 ?
                              forvar1255 : reg1496)) : reg1514) | $unsigned(({forvar1311} ?
                          (reg1275 ?
                              reg1325 : reg1282) : $signed(forvar1235))));
                      reg1545 <= ($unsigned(reg1496) >= (~((+reg1401) ?
                          (+forvar1355) : $unsigned(forvar1269))));
                      reg1546 <= $unsigned((~|(forvar1286 ?
                          (-reg1407) : reg1309)));
                      reg1547 <= reg1438;
                    end
                  reg1548 <= $signed((~^(reg1263[(3'h6):(3'h5)] & $unsigned(forvar1479))));
                  for (forvar1549 = (1'h0); (forvar1549 < (2'h2)); forvar1549 = (forvar1549 + (1'h1)))
                    begin
                      reg1550 <= reg1440[(1'h0):(1'h0)];
                      reg1551 <= reg1369[(3'h6):(1'h0)];
                      reg1552 <= $unsigned($signed(forvar1277));
                      reg1553 <= $unsigned({$unsigned((reg1546 ?
                              forvar1243 : (8'hb0)))});
                    end
                  for (forvar1554 = (1'h0); (forvar1554 < (2'h3)); forvar1554 = (forvar1554 + (1'h1)))
                    begin
                      reg1555 <= (({reg1550[(3'h7):(3'h7)]} ^ ((forvar1255 >> forvar1367) && reg1308)) | reg1275[(1'h1):(1'h0)]);
                      reg1556 <= forvar1461;
                    end
                end
              for (forvar1557 = (1'h0); (forvar1557 < (2'h3)); forvar1557 = (forvar1557 + (1'h1)))
                begin
                  if (reg1319[(1'h0):(1'h0)])
                    begin
                      reg1558 <= {($signed(((8'ha9) ?
                              (8'hb9) : (8'haf))) >= ((~^reg1354) ?
                              (reg1407 >= reg1545) : (reg1458 == (8'hb5))))};
                      reg1559 <= $unsigned($signed(reg1389[(3'h6):(1'h0)]));
                      reg1560 <= reg1528;
                      reg1561 <= ((~^reg1357[(3'h6):(2'h2)]) >>> $unsigned((!(forvar1557 ?
                          reg1562 : forvar1410))));
                    end
                  else
                    begin
                      reg1558 <= (-forvar1248[(3'h4):(3'h4)]);
                      reg1559 <= (~^(forvar1378 ?
                          $unsigned(reg1493[(1'h0):(1'h0)]) : ($signed(forvar1344) || forvar1328)));
                      reg1560 <= $signed({$signed(reg1281[(4'ha):(1'h0)])});
                    end
                  if ({$unsigned(((^reg1233) >> $signed(reg1514)))})
                    begin
                      reg1562 <= (+($signed($signed(reg1552)) ?
                          {$unsigned(reg1251)} : reg1272));
                      reg1563 <= ((forvar1328 ?
                              (^{forvar1410}) : $signed($unsigned(reg1345))) ?
                          (reg1491[(3'h4):(2'h3)] == {(+forvar1506)}) : $signed(((forvar1414 | reg1232) <= $signed(reg1478))));
                      reg1564 <= $signed($signed($signed({forvar1286})));
                      reg1565 <= (^~($unsigned(((8'ha4) >= reg1498)) * ((forvar1320 >> forvar1429) > (reg1527 ?
                          forvar1411 : reg1397))));
                    end
                  else
                    begin
                      reg1562 <= reg1345[(1'h1):(1'h1)];
                      reg1563 <= (+(^forvar1433));
                      reg1564 <= ((~&(-{reg1366})) != ({$unsigned(reg1365)} ^ ((|forvar1235) != reg1508[(2'h2):(1'h0)])));
                      reg1565 <= $signed((^(reg1536[(3'h7):(3'h4)] ?
                          (reg1315 - forvar1398) : $signed(reg1507))));
                    end
                end
              reg1566 <= reg1562[(4'h8):(2'h2)];
              for (forvar1567 = (1'h0); (forvar1567 < (2'h3)); forvar1567 = (forvar1567 + (1'h1)))
                begin
                  if ($unsigned(reg1389[(3'h5):(2'h2)]))
                    begin
                      reg1568 <= ((+((wire1223 | reg1539) ?
                              (reg1242 ? reg1299 : reg1364) : reg1229)) ?
                          (forvar1293 ?
                              reg1447[(5'h10):(4'hf)] : {(reg1526 ?
                                      reg1258 : (8'ha8))}) : reg1557[(3'h6):(2'h3)]);
                      reg1569 <= (($unsigned($unsigned(reg1281)) ~^ (~|(~&forvar1243))) ^ forvar1554[(1'h0):(1'h0)]);
                      reg1570 <= reg1486;
                      reg1571 <= (^((8'h9e) ?
                          ({reg1449} ?
                              reg1381[(3'h5):(3'h5)] : (8'ha0)) : forvar1265));
                    end
                  else
                    begin
                      reg1568 <= (8'ha7);
                      reg1569 <= (+$unsigned((reg1381[(1'h1):(1'h0)] >>> (reg1359 - reg1520))));
                      reg1570 <= ($unsigned($signed($signed(reg1509))) ?
                          forvar1395 : (reg1410 << (reg1465[(3'h7):(3'h7)] && (~^reg1427))));
                    end
                  for (forvar1572 = (1'h0); (forvar1572 < (2'h2)); forvar1572 = (forvar1572 + (1'h1)))
                    begin
                      reg1573 <= reg1406[(2'h3):(1'h0)];
                      reg1574 <= ((^~$unsigned((~(8'ha6)))) ?
                          {$unsigned({reg1317})} : reg1343[(4'h9):(4'h9)]);
                      reg1575 <= reg1494[(3'h6):(1'h0)];
                    end
                end
            end
          for (forvar1576 = (1'h0); (forvar1576 < (1'h1)); forvar1576 = (forvar1576 + (1'h1)))
            begin
              reg1577 <= reg1467[(1'h1):(1'h1)];
              for (forvar1578 = (1'h0); (forvar1578 < (2'h2)); forvar1578 = (forvar1578 + (1'h1)))
                begin
                  for (forvar1579 = (1'h0); (forvar1579 < (2'h3)); forvar1579 = (forvar1579 + (1'h1)))
                    begin
                      reg1580 <= $unsigned($signed(reg1490[(3'h6):(3'h4)]));
                    end
                  reg1581 <= $unsigned($signed(reg1517));
                  if ((reg1505[(3'h4):(1'h0)] ?
                      (&($unsigned(reg1507) < (reg1241 ^ reg1566))) : $signed($unsigned((reg1368 ?
                          reg1417 : (8'hb5))))))
                    begin
                      reg1582 <= (reg1393 ?
                          $unsigned(((~(8'ha8)) <= (wire1223 & reg1250))) : $signed({(~reg1458)}));
                      reg1583 <= $signed(reg1361);
                    end
                  else
                    begin
                      reg1582 <= (((((8'h9c) - forvar1423) ~^ $signed(forvar1472)) <= {$signed(reg1580)}) ?
                          wire1222[(3'h4):(2'h2)] : {(reg1455 == reg1485[(1'h0):(1'h0)])});
                    end
                  if (reg1449[(3'h5):(1'h1)])
                    begin
                      reg1584 <= ($signed($signed(forvar1312[(3'h6):(1'h0)])) || $signed((^~$signed(forvar1243))));
                      reg1585 <= $signed($signed(((~&reg1384) + (reg1420 >= reg1407))));
                      reg1586 <= $signed((reg1397[(1'h0):(1'h0)] ?
                          $unsigned((-forvar1542)) : {((8'ha9) & (8'hba))}));
                      reg1587 <= (~|reg1348[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1584 <= (((!{reg1504}) & (reg1388 != $unsigned((8'hb9)))) ?
                          $unsigned(forvar1317) : {reg1474[(2'h3):(1'h0)]});
                      reg1585 <= (-$signed(reg1390[(1'h0):(1'h0)]));
                      reg1586 <= forvar1433[(2'h3):(2'h3)];
                    end
                end
              if (((((reg1303 ? forvar1414 : (8'hac)) ?
                          ((8'ha2) != forvar1274) : ((8'haf) ?
                              forvar1479 : reg1305)) ?
                      $signed((&wire1223)) : ((&reg1322) ?
                          reg1550 : $unsigned(reg1529))) ?
                  (((forvar1434 ^ forvar1459) & {forvar1353}) ?
                      $signed((reg1373 == forvar1260)) : (~(-forvar1434))) : (((reg1236 ^ reg1415) ?
                      reg1271[(3'h6):(3'h6)] : reg1509[(3'h6):(1'h1)]) > reg1394[(1'h0):(1'h0)])))
                begin
                  reg1588 <= (($signed((^~(8'ha5))) - (!(8'h9f))) ?
                      {reg1539} : reg1447[(3'h4):(2'h3)]);
                  reg1589 <= forvar1434[(1'h1):(1'h1)];
                end
              else
                begin
                  reg1588 <= (($unsigned({(8'h9c)}) <= (reg1381[(3'h4):(3'h4)] + (reg1453 ?
                      reg1406 : forvar1337))) ^~ reg1532);
                  if ((^~$signed(reg1422)))
                    begin
                      reg1589 <= $unsigned($signed($unsigned((reg1559 * reg1431))));
                    end
                  else
                    begin
                      reg1589 <= ((forvar1255[(1'h0):(1'h0)] - (~|(reg1263 > forvar1260))) ?
                          $signed(forvar1255[(1'h1):(1'h0)]) : $unsigned($signed((reg1319 == forvar1461))));
                      reg1590 <= (($signed(reg1502) ?
                          (forvar1543 ?
                              $signed(forvar1461) : (reg1580 ^ reg1309)) : $unsigned((forvar1265 * reg1387))) - (!wire1285[(1'h1):(1'h0)]));
                    end
                  if (($unsigned((|$signed((8'hb6)))) ?
                      ($signed({reg1263}) ?
                          $signed(reg1504[(1'h1):(1'h0)]) : (reg1397 ?
                              $unsigned(reg1507) : $unsigned((8'ha5)))) : reg1520))
                    begin
                      reg1591 <= reg1237[(4'hb):(4'h9)];
                      reg1592 <= reg1279;
                      reg1593 <= forvar1524[(1'h0):(1'h0)];
                      reg1594 <= (($signed($unsigned(reg1443)) ?
                              forvar1391 : (!(reg1502 ^ reg1574))) ?
                          ($unsigned((8'hb3)) == wire1284) : ($unsigned($unsigned((8'haa))) || (reg1408[(3'h6):(1'h0)] ?
                              $unsigned((8'hac)) : reg1397)));
                    end
                  else
                    begin
                      reg1591 <= (8'h9f);
                      reg1592 <= forvar1497[(4'hb):(1'h1)];
                    end
                end
            end
        end
    end
  assign wire1595 = ($signed(($unsigned((8'h9c)) ?
                        $unsigned(forvar1473) : $signed((8'ha6)))) < {(reg1239 ?
                            reg1525 : (forvar1423 ? reg1586 : reg1502))});
  assign wire1596 = ($unsigned(forvar1235[(2'h2):(2'h2)]) ?
                        forvar1547[(2'h3):(2'h2)] : reg1467);
  always
    @(posedge clk) begin
      reg1597 <= (-reg1299[(4'hb):(3'h6)]);
      for (forvar1598 = (1'h0); (forvar1598 < (1'h1)); forvar1598 = (forvar1598 + (1'h1)))
        begin
          if (reg1375)
            begin
              for (forvar1599 = (1'h0); (forvar1599 < (1'h0)); forvar1599 = (forvar1599 + (1'h1)))
                begin
                  reg1600 <= $signed((reg1330 ?
                      reg1377 : (^~((8'hab) << forvar1509))));
                  for (forvar1601 = (1'h0); (forvar1601 < (1'h0)); forvar1601 = (forvar1601 + (1'h1)))
                    begin
                      reg1602 <= {$signed(((forvar1601 ^ reg1556) ?
                              $unsigned((8'hb4)) : (+reg1522)))};
                      reg1603 <= (!reg1241);
                      reg1604 <= reg1545[(1'h0):(1'h0)];
                    end
                  if ($signed($signed(forvar1286)))
                    begin
                      reg1605 <= ((reg1244[(3'h6):(3'h6)] ?
                              forvar1543 : ((|(8'ha8)) | (8'ha1))) ?
                          (~|$signed((-reg1434))) : (reg1457[(4'hc):(4'ha)] << reg1428[(1'h1):(1'h1)]));
                      reg1606 <= reg1317;
                      reg1607 <= (~&$unsigned(reg1410));
                      reg1608 <= (reg1501[(1'h1):(1'h1)] ?
                          $signed(((reg1519 && reg1355) | ((8'hb6) < reg1363))) : $signed($signed(forvar1429)));
                    end
                  else
                    begin
                      reg1605 <= reg1438;
                      reg1606 <= {({reg1394} | reg1290[(3'h5):(3'h4)])};
                      reg1607 <= $unsigned($unsigned(($unsigned((8'hb5)) ?
                          (forvar1521 ^ reg1290) : ((8'hb0) ?
                              (8'ha2) : reg1345))));
                    end
                  if ((~&(reg1550 ?
                      (reg1315[(3'h4):(1'h0)] >>> $signed((8'hb0))) : ((forvar1353 <<< (8'h9d)) ?
                          reg1382 : forvar1225[(3'h4):(2'h3)]))))
                    begin
                      reg1609 <= (reg1421 >>> ((reg1453[(3'h6):(3'h5)] || (^reg1374)) != (^((8'ha7) ?
                          reg1493 : forvar1317))));
                      reg1610 <= (-(|reg1447));
                      reg1611 <= $unsigned($signed($signed($signed(reg1384))));
                    end
                  else
                    begin
                      reg1609 <= forvar1461;
                    end
                end
              reg1612 <= forvar1429;
              for (forvar1613 = (1'h0); (forvar1613 < (1'h0)); forvar1613 = (forvar1613 + (1'h1)))
                begin
                  for (forvar1614 = (1'h0); (forvar1614 < (2'h3)); forvar1614 = (forvar1614 + (1'h1)))
                    begin
                      reg1615 <= (($signed((reg1404 ?
                              forvar1265 : forvar1255)) ?
                          forvar1418 : ($signed(reg1513) <= (reg1443 ?
                              reg1556 : reg1462))) == {(~^$signed(forvar1436))});
                      reg1616 <= $signed(wire1595[(3'h6):(3'h6)]);
                      reg1617 <= reg1296[(4'ha):(3'h7)];
                    end
                end
            end
          else
            begin
              if (((8'hac) <= reg1573[(3'h4):(2'h2)]))
                begin
                  for (forvar1599 = (1'h0); (forvar1599 < (1'h1)); forvar1599 = (forvar1599 + (1'h1)))
                    begin
                      reg1600 <= $unsigned({$signed(forvar1355[(2'h2):(1'h0)])});
                    end
                  for (forvar1601 = (1'h0); (forvar1601 < (2'h3)); forvar1601 = (forvar1601 + (1'h1)))
                    begin
                      reg1602 <= (~^$unsigned($signed($signed((8'hb2)))));
                      reg1603 <= reg1246;
                      reg1604 <= (+reg1458[(2'h3):(1'h0)]);
                      reg1605 <= (~reg1377[(2'h3):(1'h1)]);
                    end
                end
              else
                begin
                  if ($unsigned((~^(&(reg1516 ? forvar1398 : (8'ha9))))))
                    begin
                      reg1599 <= ($signed($signed((forvar1410 ?
                          reg1317 : forvar1247))) ^ (((forvar1423 ?
                                  forvar1433 : reg1264) ?
                              reg1318[(4'h8):(3'h4)] : $unsigned(reg1507)) ?
                          {wire1220[(2'h3):(2'h2)]} : {$signed(forvar1433)}));
                      reg1600 <= (8'hb1);
                      reg1601 <= reg1505[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1599 <= (~reg1447[(2'h2):(1'h0)]);
                      reg1600 <= $signed(reg1266);
                      reg1601 <= $unsigned($unsigned(reg1275[(1'h0):(1'h0)]));
                    end
                end
            end
        end
      if (forvar1337)
        begin
          for (forvar1618 = (1'h0); (forvar1618 < (2'h2)); forvar1618 = (forvar1618 + (1'h1)))
            begin
              reg1619 <= ($unsigned(reg1383) >> reg1583);
              for (forvar1620 = (1'h0); (forvar1620 < (2'h2)); forvar1620 = (forvar1620 + (1'h1)))
                begin
                  reg1621 <= (-(8'ha1));
                  if ($signed(($signed(reg1403) | $signed((!reg1611)))))
                    begin
                      reg1622 <= $unsigned({$unsigned((forvar1496 ?
                              reg1446 : forvar1408))});
                    end
                  else
                    begin
                      reg1622 <= (reg1551[(2'h2):(1'h0)] ?
                          $unsigned({(^forvar1288)}) : reg1506);
                      reg1623 <= $signed(($signed((reg1443 ~^ reg1428)) ?
                          (8'hb8) : forvar1599));
                      reg1624 <= {$signed(reg1395)};
                      reg1625 <= $signed(({reg1309} ?
                          $unsigned($signed(forvar1343)) : ($signed(reg1407) ?
                              reg1612 : (reg1471 ^~ reg1511))));
                    end
                  for (forvar1626 = (1'h0); (forvar1626 < (2'h2)); forvar1626 = (forvar1626 + (1'h1)))
                    begin
                      reg1627 <= ($unsigned($signed((forvar1371 != reg1298))) ^ reg1388);
                      reg1628 <= (~^(~forvar1414[(2'h2):(2'h2)]));
                      reg1629 <= $unsigned((&reg1477));
                      reg1630 <= $unsigned($unsigned(reg1500[(1'h0):(1'h0)]));
                    end
                  for (forvar1631 = (1'h0); (forvar1631 < (1'h1)); forvar1631 = (forvar1631 + (1'h1)))
                    begin
                      reg1632 <= (forvar1436[(4'he):(4'hd)] >> reg1395);
                      reg1633 <= (8'ha2);
                    end
                end
              if ($signed($unsigned(reg1404)))
                begin
                  for (forvar1634 = (1'h0); (forvar1634 < (2'h2)); forvar1634 = (forvar1634 + (1'h1)))
                    begin
                      reg1635 <= (&reg1491);
                    end
                  if (forvar1320)
                    begin
                      reg1636 <= {(!$signed((reg1485 ? reg1404 : (8'hab))))};
                    end
                  else
                    begin
                      reg1636 <= ($signed($signed((reg1629 ?
                              reg1304 : wire1596))) ?
                          $signed($signed(reg1262)) : (((forvar1618 ?
                                  reg1386 : forvar1260) ?
                              {(8'hb2)} : $unsigned(reg1605)) == forvar1614));
                      reg1637 <= $signed($unsigned(($unsigned(forvar1567) >>> (|reg1610))));
                      reg1638 <= (forvar1439[(1'h1):(1'h1)] == (((forvar1598 << forvar1540) > reg1477) ?
                          ((forvar1464 | reg1413) >>> (forvar1459 && reg1340)) : reg1534[(4'hb):(4'hb)]));
                    end
                end
              else
                begin
                  for (forvar1634 = (1'h0); (forvar1634 < (1'h1)); forvar1634 = (forvar1634 + (1'h1)))
                    begin
                      reg1635 <= (forvar1529 ?
                          ($unsigned($unsigned(reg1315)) ?
                              ((-forvar1402) ?
                                  $unsigned(forvar1460) : (8'hac)) : (reg1570 != reg1521[(1'h1):(1'h1)])) : forvar1613);
                      reg1636 <= ($signed((&$unsigned(reg1393))) ?
                          reg1311[(4'h9):(1'h1)] : reg1360[(1'h1):(1'h1)]);
                    end
                  for (forvar1637 = (1'h0); (forvar1637 < (2'h3)); forvar1637 = (forvar1637 + (1'h1)))
                    begin
                      reg1638 <= $unsigned($signed($unsigned($signed((8'hb7)))));
                      reg1639 <= ($signed(({forvar1312} ?
                          $signed((8'ha5)) : $unsigned(reg1364))) - (($unsigned(forvar1543) > (reg1444 ?
                              reg1504 : reg1315)) ?
                          (~&(forvar1334 ?
                              reg1427 : reg1388)) : $unsigned(reg1448[(1'h1):(1'h0)])));
                      reg1640 <= reg1447;
                      reg1641 <= (~^{reg1279[(2'h2):(2'h2)]});
                    end
                  reg1642 <= $signed(($signed((~&reg1496)) ?
                      reg1605 : $signed($signed((8'had)))));
                  if ($unsigned({{reg1465[(2'h3):(1'h1)]}}))
                    begin
                      reg1643 <= reg1521;
                      reg1644 <= (reg1493 & $unsigned({((8'hb9) ^~ forvar1599)}));
                      reg1645 <= reg1310;
                      reg1646 <= (^(reg1639 ? reg1396 : $unsigned(reg1327)));
                    end
                  else
                    begin
                      reg1643 <= $signed((+{reg1386[(4'ha):(4'h8)]}));
                    end
                end
            end
          reg1647 <= (forvar1476[(4'hf):(2'h2)] ~^ (reg1249 & ((reg1281 != reg1237) ?
              $unsigned(reg1446) : forvar1254[(3'h6):(1'h0)])));
          for (forvar1648 = (1'h0); (forvar1648 < (2'h3)); forvar1648 = (forvar1648 + (1'h1)))
            begin
              for (forvar1649 = (1'h0); (forvar1649 < (1'h1)); forvar1649 = (forvar1649 + (1'h1)))
                begin
                  for (forvar1650 = (1'h0); (forvar1650 < (2'h3)); forvar1650 = (forvar1650 + (1'h1)))
                    begin
                      reg1651 <= (~^reg1553[(2'h3):(1'h1)]);
                    end
                  for (forvar1652 = (1'h0); (forvar1652 < (2'h2)); forvar1652 = (forvar1652 + (1'h1)))
                    begin
                      reg1653 <= $unsigned(($unsigned($signed(reg1408)) + (8'ha8)));
                      reg1654 <= ((^~reg1428) >= ((~forvar1519) ?
                          (8'hba) : reg1586[(4'h8):(3'h6)]));
                      reg1655 <= (^~(^~(~&reg1318[(3'h6):(3'h4)])));
                    end
                end
              reg1656 <= (!(((forvar1232 ?
                  forvar1400 : reg1373) <= (^reg1391)) ^ forvar1439[(1'h0):(1'h0)]));
              if (forvar1634[(3'h6):(1'h0)])
                begin
                  for (forvar1657 = (1'h0); (forvar1657 < (1'h0)); forvar1657 = (forvar1657 + (1'h1)))
                    begin
                      reg1658 <= ((^~((8'ha8) ?
                              (forvar1273 ?
                                  forvar1334 : reg1344) : reg1394[(1'h1):(1'h0)])) ?
                          $signed($unsigned(reg1625[(3'h5):(3'h4)])) : ($signed((8'hb6)) >> (((8'hb0) ?
                              reg1573 : reg1491) || $signed(forvar1489))));
                      reg1659 <= forvar1579[(3'h4):(1'h0)];
                      reg1660 <= $unsigned((8'ha5));
                      reg1661 <= reg1356[(2'h2):(1'h0)];
                    end
                  for (forvar1662 = (1'h0); (forvar1662 < (2'h3)); forvar1662 = (forvar1662 + (1'h1)))
                    begin
                      reg1663 <= (reg1585 ?
                          ((8'hab) ?
                              $unsigned($signed(forvar1293)) : $signed((~reg1581))) : (reg1645[(1'h0):(1'h0)] > reg1465[(1'h1):(1'h1)]));
                      reg1664 <= (8'hac);
                      reg1665 <= (&$unsigned($unsigned((reg1604 && forvar1423))));
                    end
                  if ({((((8'hb0) == (8'hab)) >>> (reg1369 ?
                              reg1251 : forvar1497)) ?
                          reg1647 : $unsigned($unsigned(forvar1411)))})
                    begin
                      reg1666 <= reg1518;
                      reg1667 <= (forvar1626[(3'h4):(2'h3)] ^ $unsigned((|reg1377)));
                      reg1668 <= $unsigned($unsigned(reg1615));
                      reg1669 <= (&reg1606[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg1666 <= reg1259[(4'hb):(4'h9)];
                      reg1667 <= $unsigned(reg1659);
                      reg1668 <= forvar1273[(1'h0):(1'h0)];
                      reg1669 <= reg1356;
                    end
                end
              else
                begin
                  reg1657 <= (~^($unsigned((+reg1351)) ?
                      {(!reg1604)} : reg1321[(3'h5):(3'h5)]));
                end
              if ($unsigned((((8'ha8) ?
                      (reg1639 ? reg1667 : reg1227) : (reg1494 ?
                          wire1595 : reg1546)) ?
                  ((|reg1410) <<< $signed((8'hb4))) : ((forvar1347 >> forvar1519) * reg1610))))
                begin
                  reg1670 <= {(^reg1633[(1'h0):(1'h0)])};
                  if (($unsigned(reg1597) ?
                      {$unsigned(reg1453[(1'h0):(1'h0)])} : reg1644))
                    begin
                      reg1671 <= (reg1502[(1'h1):(1'h1)] ~^ ($unsigned(reg1520) < reg1600[(1'h1):(1'h1)]));
                      reg1672 <= (~&$signed({$unsigned(reg1369)}));
                      reg1673 <= ({reg1320[(2'h3):(1'h1)]} ?
                          $signed(($signed(reg1409) ?
                              (reg1340 ?
                                  reg1671 : reg1642) : $unsigned(reg1319))) : $signed(((~reg1438) << reg1544)));
                      reg1674 <= $signed(reg1325[(4'h8):(2'h2)]);
                    end
                  else
                    begin
                      reg1671 <= ($unsigned(((reg1531 ? reg1368 : (8'hb4)) ?
                          $unsigned(reg1364) : reg1335[(2'h2):(1'h1)])) ~^ reg1304[(1'h0):(1'h0)]);
                      reg1672 <= {($signed((reg1353 < reg1647)) ?
                              (-reg1363[(2'h2):(1'h0)]) : $unsigned($unsigned(reg1554)))};
                      reg1673 <= ($unsigned(reg1387[(1'h0):(1'h0)]) ?
                          reg1415[(3'h5):(3'h5)] : ((8'h9c) ?
                              (8'ha8) : (reg1270[(1'h0):(1'h0)] >= (reg1296 ?
                                  (8'hab) : reg1369))));
                    end
                end
              else
                begin
                  if ($unsigned(reg1497[(1'h1):(1'h0)]))
                    begin
                      reg1670 <= forvar1436;
                    end
                  else
                    begin
                      reg1670 <= (((~^$unsigned(forvar1626)) == $signed((reg1558 && forvar1226))) ?
                          (~&$signed((&reg1296))) : ((~|(reg1450 ?
                              (8'ha8) : reg1395)) > ((reg1554 ?
                              forvar1404 : reg1446) >> (&forvar1493))));
                    end
                end
            end
          for (forvar1675 = (1'h0); (forvar1675 < (1'h0)); forvar1675 = (forvar1675 + (1'h1)))
            begin
              for (forvar1676 = (1'h0); (forvar1676 < (2'h2)); forvar1676 = (forvar1676 + (1'h1)))
                begin
                  for (forvar1677 = (1'h0); (forvar1677 < (2'h2)); forvar1677 = (forvar1677 + (1'h1)))
                    begin
                      reg1678 <= (reg1392[(3'h4):(1'h0)] >= ((reg1420[(4'h8):(4'h8)] + (+forvar1255)) < (8'hb3)));
                      reg1679 <= reg1635;
                    end
                  if ($signed($signed(($signed(reg1589) ?
                      (forvar1634 ?
                          reg1511 : forvar1235) : $unsigned(reg1417)))))
                    begin
                      reg1680 <= $unsigned($unsigned(forvar1543));
                    end
                  else
                    begin
                      reg1680 <= ((({reg1659} <<< $unsigned(forvar1614)) ?
                              $signed((^forvar1254)) : $signed((&forvar1278))) ?
                          $unsigned(reg1612[(2'h2):(1'h0)]) : (8'haa));
                      reg1681 <= $signed(((^$signed(reg1672)) >>> reg1347));
                    end
                end
              for (forvar1682 = (1'h0); (forvar1682 < (2'h2)); forvar1682 = (forvar1682 + (1'h1)))
                begin
                  for (forvar1683 = (1'h0); (forvar1683 < (2'h3)); forvar1683 = (forvar1683 + (1'h1)))
                    begin
                      reg1684 <= reg1669;
                      reg1685 <= $signed($signed((-(reg1536 - reg1679))));
                    end
                  if (reg1268)
                    begin
                      reg1686 <= ($unsigned((((8'h9d) ^~ reg1657) && reg1294[(3'h4):(3'h4)])) ?
                          (~&reg1355) : $signed(forvar1273[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg1686 <= $signed(reg1421[(1'h1):(1'h1)]);
                      reg1687 <= (~|(($signed(reg1372) ?
                              (forvar1439 <<< forvar1567) : $signed(reg1349)) ?
                          $unsigned((forvar1287 ?
                              (8'hb1) : reg1424)) : $signed((8'hac))));
                    end
                end
            end
        end
      else
        begin
          reg1618 <= (((~&(reg1332 | forvar1307)) ?
                  $unsigned((~&reg1562)) : ((reg1323 ? reg1594 : forvar1614) ?
                      $unsigned(reg1504) : reg1632)) ?
              ((-(forvar1543 ?
                  forvar1353 : (8'hb3))) != $signed($unsigned(reg1564))) : $signed(((~reg1398) * $unsigned(reg1638))));
        end
    end
  assign wire1688 = (-reg1518);
  always
    @(posedge clk) begin
      for (forvar1689 = (1'h0); (forvar1689 < (2'h3)); forvar1689 = (forvar1689 + (1'h1)))
        begin
          for (forvar1690 = (1'h0); (forvar1690 < (2'h3)); forvar1690 = (forvar1690 + (1'h1)))
            begin
              for (forvar1691 = (1'h0); (forvar1691 < (2'h3)); forvar1691 = (forvar1691 + (1'h1)))
                begin
                  if (((|$unsigned($signed(reg1424))) == reg1317[(4'hd):(2'h3)]))
                    begin
                      reg1692 <= reg1295[(2'h2):(1'h0)];
                      reg1693 <= ($unsigned($signed(reg1259)) ?
                          (forvar1328 ~^ reg1599[(3'h5):(1'h0)]) : $signed($unsigned((+forvar1328))));
                    end
                  else
                    begin
                      reg1692 <= ((-$unsigned($signed(reg1402))) && reg1432[(4'h9):(3'h7)]);
                      reg1693 <= (reg1581 - $signed({$signed((8'hb5))}));
                    end
                end
            end
          if ((~|reg1684[(2'h3):(2'h3)]))
            begin
              for (forvar1694 = (1'h0); (forvar1694 < (1'h0)); forvar1694 = (forvar1694 + (1'h1)))
                begin
                  for (forvar1695 = (1'h0); (forvar1695 < (2'h2)); forvar1695 = (forvar1695 + (1'h1)))
                    begin
                      reg1696 <= (!$unsigned(forvar1401));
                    end
                end
              reg1697 <= reg1231[(1'h0):(1'h0)];
              reg1698 <= (+$signed(forvar1372));
            end
          else
            begin
              for (forvar1694 = (1'h0); (forvar1694 < (2'h2)); forvar1694 = (forvar1694 + (1'h1)))
                begin
                  for (forvar1695 = (1'h0); (forvar1695 < (1'h1)); forvar1695 = (forvar1695 + (1'h1)))
                    begin
                      reg1696 <= (8'hb2);
                    end
                  for (forvar1697 = (1'h0); (forvar1697 < (2'h2)); forvar1697 = (forvar1697 + (1'h1)))
                    begin
                      reg1698 <= $unsigned($unsigned(forvar1598));
                    end
                  for (forvar1699 = (1'h0); (forvar1699 < (1'h1)); forvar1699 = (forvar1699 + (1'h1)))
                    begin
                      reg1700 <= (reg1412 - ($signed(reg1674) ?
                          $unsigned((reg1305 ^ (8'hb4))) : reg1551[(1'h0):(1'h0)]));
                      reg1701 <= {reg1406};
                      reg1702 <= ((-reg1532) > reg1355);
                      reg1703 <= forvar1378[(2'h2):(1'h1)];
                    end
                  for (forvar1704 = (1'h0); (forvar1704 < (2'h2)); forvar1704 = (forvar1704 + (1'h1)))
                    begin
                      reg1705 <= reg1551[(1'h0):(1'h0)];
                      reg1706 <= $signed($signed((~^(~|reg1556))));
                      reg1707 <= reg1416[(3'h4):(1'h1)];
                    end
                end
              for (forvar1708 = (1'h0); (forvar1708 < (2'h2)); forvar1708 = (forvar1708 + (1'h1)))
                begin
                  for (forvar1709 = (1'h0); (forvar1709 < (2'h3)); forvar1709 = (forvar1709 + (1'h1)))
                    begin
                      reg1710 <= $unsigned($signed(($signed(reg1545) - {reg1582})));
                      reg1711 <= {$signed(((reg1594 ? forvar1363 : reg1693) ?
                              forvar1255 : {reg1415}))};
                      reg1712 <= (reg1702 ?
                          (~&(~|$signed(forvar1579))) : $unsigned(forvar1508));
                    end
                  if ($signed((reg1448 ?
                      {$signed(forvar1441)} : reg1305[(3'h5):(3'h5)])))
                    begin
                      reg1713 <= reg1449[(4'hd):(2'h3)];
                      reg1714 <= forvar1411[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg1713 <= $unsigned((^~forvar1371[(3'h7):(3'h5)]));
                    end
                end
            end
          if (((~&reg1432) + $unsigned(forvar1488[(4'hb):(4'h8)])))
            begin
              for (forvar1715 = (1'h0); (forvar1715 < (1'h0)); forvar1715 = (forvar1715 + (1'h1)))
                begin
                  for (forvar1716 = (1'h0); (forvar1716 < (2'h3)); forvar1716 = (forvar1716 + (1'h1)))
                    begin
                      reg1717 <= forvar1334[(3'h7):(2'h3)];
                      reg1718 <= reg1549;
                      reg1719 <= (((reg1687 ?
                              $unsigned((8'ha8)) : (forvar1493 ?
                                  reg1422 : forvar1690)) ?
                          reg1696 : {(8'hb9)}) <= reg1671);
                    end
                  for (forvar1720 = (1'h0); (forvar1720 < (1'h0)); forvar1720 = (forvar1720 + (1'h1)))
                    begin
                      reg1721 <= forvar1520[(4'hc):(3'h7)];
                      reg1722 <= (((|{reg1354}) ~^ reg1692) ?
                          forvar1691[(2'h3):(2'h3)] : $unsigned((8'hae)));
                    end
                end
              if (forvar1400[(4'h9):(1'h0)])
                begin
                  if ($signed(($unsigned(reg1351[(2'h3):(1'h0)]) + reg1571[(3'h7):(2'h2)])))
                    begin
                      reg1723 <= reg1552[(3'h5):(2'h2)];
                      reg1724 <= forvar1408[(1'h1):(1'h0)];
                      reg1725 <= ($unsigned(forvar1695) ?
                          forvar1243 : $signed(forvar1695));
                      reg1726 <= $signed(((-reg1568) ?
                          {(reg1477 - (8'hac))} : ((reg1492 ?
                              reg1657 : reg1635) >>> $signed(forvar1459))));
                    end
                  else
                    begin
                      reg1723 <= (|$signed(((+(8'hb2)) ?
                          reg1644[(4'ha):(4'h8)] : $unsigned(reg1497))));
                    end
                  reg1727 <= $unsigned(forvar1550[(1'h1):(1'h1)]);
                  for (forvar1728 = (1'h0); (forvar1728 < (1'h0)); forvar1728 = (forvar1728 + (1'h1)))
                    begin
                      reg1729 <= forvar1278[(3'h4):(3'h4)];
                      reg1730 <= {forvar1320};
                    end
                  for (forvar1731 = (1'h0); (forvar1731 < (1'h0)); forvar1731 = (forvar1731 + (1'h1)))
                    begin
                      reg1732 <= $signed((+reg1360[(2'h3):(1'h0)]));
                      reg1733 <= $signed((8'ha5));
                    end
                end
              else
                begin
                  reg1723 <= reg1665[(1'h1):(1'h0)];
                  for (forvar1724 = (1'h0); (forvar1724 < (2'h2)); forvar1724 = (forvar1724 + (1'h1)))
                    begin
                      reg1725 <= ((reg1499[(2'h2):(2'h2)] & $unsigned($signed((8'h9f)))) << forvar1410);
                    end
                  if (reg1601[(2'h3):(1'h0)])
                    begin
                      reg1726 <= reg1406;
                      reg1727 <= (~&{reg1443});
                      reg1728 <= ($signed($signed(reg1617[(2'h2):(1'h0)])) ?
                          (((8'haa) ? $unsigned(forvar1613) : reg1571) ?
                              $unsigned($signed(reg1235)) : {$unsigned(reg1585)}) : $unsigned(({forvar1614} <<< $signed(reg1447))));
                      reg1729 <= reg1374[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg1726 <= $signed((8'hb7));
                      reg1727 <= reg1581;
                      reg1728 <= (forvar1648 < $signed(($unsigned(forvar1572) ?
                          $unsigned(reg1465) : (forvar1364 ?
                              reg1421 : forvar1549))));
                      reg1729 <= (($signed(((8'hb9) ~^ reg1387)) ?
                              reg1249 : reg1664) ?
                          ($signed((forvar1473 + reg1592)) >= (reg1526 ?
                              ((8'ha7) ^~ forvar1230) : ((8'h9e) >> forvar1367))) : reg1432[(1'h0):(1'h0)]);
                    end
                  if ({reg1559})
                    begin
                      reg1730 <= (reg1333 ?
                          (8'haf) : {$signed((~^forvar1572))});
                      reg1731 <= $unsigned((reg1710[(3'h6):(3'h4)] >> $unsigned(reg1229)));
                      reg1732 <= reg1495;
                    end
                  else
                    begin
                      reg1730 <= $unsigned($unsigned(reg1549[(3'h5):(2'h2)]));
                      reg1731 <= $signed($signed(reg1359[(3'h6):(2'h2)]));
                    end
                end
              if (reg1486[(2'h3):(1'h1)])
                begin
                  for (forvar1734 = (1'h0); (forvar1734 < (2'h2)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= reg1296;
                      reg1736 <= $signed($signed((forvar1433 ?
                          (-reg1367) : {reg1581})));
                      reg1737 <= $signed(reg1263);
                    end
                  reg1738 <= forvar1634[(3'h6):(1'h0)];
                  for (forvar1739 = (1'h0); (forvar1739 < (1'h0)); forvar1739 = (forvar1739 + (1'h1)))
                    begin
                      reg1740 <= reg1280;
                    end
                end
              else
                begin
                  if (((^~$unsigned((reg1295 && reg1685))) - reg1693))
                    begin
                      reg1734 <= (~^(({reg1244} ?
                              $unsigned(reg1592) : $signed(reg1310)) ?
                          $signed((+reg1575)) : reg1706[(1'h0):(1'h0)]));
                      reg1735 <= $signed($signed($unsigned($unsigned(reg1673))));
                      reg1736 <= $unsigned($signed({(reg1309 ?
                              reg1463 : reg1251)}));
                      reg1737 <= reg1729;
                    end
                  else
                    begin
                      reg1734 <= $signed(reg1227);
                      reg1735 <= reg1587[(1'h0):(1'h0)];
                      reg1736 <= (~^$signed(((forvar1433 <<< reg1308) == reg1396[(2'h2):(2'h2)])));
                    end
                  for (forvar1738 = (1'h0); (forvar1738 < (2'h2)); forvar1738 = (forvar1738 + (1'h1)))
                    begin
                      reg1739 <= (~&{((reg1267 ? (8'had) : forvar1613) ?
                              $signed(reg1701) : (wire1223 ?
                                  reg1313 : forvar1434))});
                      reg1740 <= reg1534[(2'h2):(2'h2)];
                    end
                end
              reg1741 <= (((&(reg1229 ?
                  reg1301 : reg1320)) != reg1435[(1'h1):(1'h1)]) ~^ ($unsigned($signed(forvar1488)) || ((~|reg1256) & reg1591[(3'h7):(1'h0)])));
            end
          else
            begin
              if ($unsigned($unsigned($signed($unsigned((8'had))))))
                begin
                  reg1715 <= (~^forvar1460);
                  reg1716 <= $signed($signed(forvar1709));
                  for (forvar1717 = (1'h0); (forvar1717 < (2'h3)); forvar1717 = (forvar1717 + (1'h1)))
                    begin
                      reg1718 <= {$unsigned(({reg1698} + (8'ha7)))};
                      reg1719 <= forvar1507;
                      reg1720 <= reg1258;
                    end
                end
              else
                begin
                  if ($signed((reg1311 == $signed((~&(8'hb4))))))
                    begin
                      reg1715 <= (-$signed((reg1453[(4'h8):(1'h0)] ?
                          {forvar1426} : (reg1527 ^~ forvar1410))));
                      reg1716 <= $signed((reg1684[(3'h5):(2'h3)] ?
                          $unsigned($signed(reg1391)) : $signed($unsigned(forvar1506))));
                    end
                  else
                    begin
                      reg1715 <= $unsigned(forvar1542);
                    end
                end
              reg1721 <= (8'hb0);
            end
        end
      reg1742 <= reg1564;
    end
  assign wire1743 = (forvar1479 ^~ ((-$signed(reg1450)) ?
                        ((-reg1370) > $unsigned(reg1728)) : (reg1272[(3'h4):(2'h3)] >>> {reg1263})));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1001  (y, clk, wire1005, wire1004, wire1003, wire1002);
  output wire [(32'h6c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire1005;
  input wire [(3'h5):(1'h0)] wire1004;
  input wire [(4'h9):(1'h0)] wire1003;
  input wire [(3'h6):(1'h0)] wire1002;
  wire signed [(4'h8):(1'h0)] wire1017;
  reg signed [(4'ha):(1'h0)] reg1016 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire1015;
  wire [(4'h8):(1'h0)] wire1014;
  wire signed [(5'h10):(1'h0)] wire1013;
  wire [(4'hd):(1'h0)] wire1012;
  wire [(3'h6):(1'h0)] wire1011;
  wire [(4'h8):(1'h0)] wire1010;
  wire [(5'h10):(1'h0)] wire1009;
  wire [(2'h3):(1'h0)] wire1008;
  wire signed [(2'h3):(1'h0)] wire1007;
  wire signed [(2'h3):(1'h0)] wire1006;
  assign y = {wire1017,
                 reg1016,
                 wire1015,
                 wire1014,
                 wire1013,
                 wire1012,
                 wire1011,
                 wire1010,
                 wire1009,
                 wire1008,
                 wire1007,
                 wire1006,
                 (1'h0)};
  assign wire1006 = ($unsigned(wire1002[(3'h4):(1'h0)]) & ($unsigned((~|wire1003)) ?
                        wire1005 : $signed({wire1004})));
  assign wire1007 = {(wire1006 <= $unsigned($unsigned(wire1006)))};
  assign wire1008 = (wire1005[(3'h5):(2'h2)] ? wire1003 : wire1004);
  assign wire1009 = $unsigned(wire1005[(2'h2):(2'h2)]);
  assign wire1010 = wire1005[(3'h7):(3'h5)];
  assign wire1011 = wire1009;
  assign wire1012 = (8'ha0);
  assign wire1013 = wire1002[(3'h5):(2'h2)];
  assign wire1014 = wire1003[(1'h1):(1'h1)];
  assign wire1015 = $signed(wire1003[(3'h7):(2'h3)]);
  always
    @(posedge clk) begin
      reg1016 <= $signed((-$signed({wire1010})));
    end
  assign wire1017 = ({((wire1009 ? (8'ha2) : wire1005) ?
                                ((8'hb6) ?
                                    (8'ha7) : wire1003) : $unsigned(wire1012))} ?
                        (wire1014[(3'h7):(2'h2)] - wire1014) : ((wire1013 ?
                            (^~(8'had)) : wire1004) ^~ $signed((wire1006 > wire1002))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3603
#( parameter param4016 = {(((^(8'hab)) == ((8'ha1) ? (8'hac) : (8'h9f))) + (|((8'ha6) ? (8'ha2) : (8'hb0))))} )
(y, clk, wire3608, wire3607, wire3606, wire3605, wire3604);
  output wire [(32'h1142):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire3608;
  input wire signed [(4'ha):(1'h0)] wire3607;
  input wire [(4'hc):(1'h0)] wire3606;
  input wire [(4'ha):(1'h0)] wire3605;
  input wire [(4'hb):(1'h0)] wire3604;
  wire [(4'he):(1'h0)] wire4015;
  reg signed [(4'ha):(1'h0)] reg4014 = (1'h0);
  reg [(4'hd):(1'h0)] reg4004 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4000 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3999 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3998 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3993 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3989 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3988 = (1'h0);
  reg [(4'ha):(1'h0)] reg3986 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3981 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3975 = (1'h0);
  reg [(4'ha):(1'h0)] reg3974 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3971 = (1'h0);
  reg [(4'ha):(1'h0)] reg4013 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4012 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4011 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4010 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4009 = (1'h0);
  reg [(2'h3):(1'h0)] reg4008 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4007 = (1'h0);
  reg [(3'h4):(1'h0)] reg4006 = (1'h0);
  reg [(3'h5):(1'h0)] reg4005 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4004 = (1'h0);
  reg [(4'h9):(1'h0)] reg4003 = (1'h0);
  reg [(3'h7):(1'h0)] reg4002 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4001 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4000 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3999 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3998 = (1'h0);
  reg [(2'h3):(1'h0)] reg3997 = (1'h0);
  reg [(5'h10):(1'h0)] reg3996 = (1'h0);
  reg [(4'hc):(1'h0)] reg3995 = (1'h0);
  reg [(3'h5):(1'h0)] reg3990 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3994 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3993 = (1'h0);
  reg [(4'he):(1'h0)] reg3992 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3991 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3990 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3989 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3988 = (1'h0);
  reg [(4'hc):(1'h0)] reg3970 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3969 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3966 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3964 = (1'h0);
  reg [(4'hd):(1'h0)] reg3984 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3980 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3976 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3987 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3986 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3985 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3984 = (1'h0);
  reg [(2'h2):(1'h0)] reg3983 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3982 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3981 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3980 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3979 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3978 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3977 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3976 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3963 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3975 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3974 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3973 = (1'h0);
  reg [(2'h3):(1'h0)] reg3972 = (1'h0);
  reg [(3'h5):(1'h0)] reg3971 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3970 = (1'h0);
  reg [(3'h5):(1'h0)] reg3969 = (1'h0);
  reg [(4'he):(1'h0)] reg3968 = (1'h0);
  reg [(4'hb):(1'h0)] reg3967 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3966 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3965 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3964 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3963 = (1'h0);
  wire [(4'h9):(1'h0)] wire3962;
  wire signed [(3'h7):(1'h0)] wire3961;
  reg [(3'h5):(1'h0)] reg3960 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3959 = (1'h0);
  reg [(4'hb):(1'h0)] reg3958 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3957 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3956 = (1'h0);
  reg [(3'h7):(1'h0)] reg3955 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3954 = (1'h0);
  reg [(4'ha):(1'h0)] reg3953 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3952 = (1'h0);
  reg [(4'he):(1'h0)] forvar3951 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3950 = (1'h0);
  reg [(5'h10):(1'h0)] reg3949 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3948 = (1'h0);
  reg [(3'h7):(1'h0)] reg3947 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3946 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3945 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3944 = (1'h0);
  reg [(4'hd):(1'h0)] reg3943 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3942 = (1'h0);
  reg [(5'h10):(1'h0)] reg3941 = (1'h0);
  reg [(4'hf):(1'h0)] reg3940 = (1'h0);
  reg [(3'h7):(1'h0)] reg3939 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3938 = (1'h0);
  reg [(4'hf):(1'h0)] reg3937 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3936 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3935 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3934 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3933 = (1'h0);
  reg [(3'h5):(1'h0)] reg3932 = (1'h0);
  reg [(4'hb):(1'h0)] reg3931 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3930 = (1'h0);
  reg [(4'ha):(1'h0)] reg3929 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3928 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3927 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3926 = (1'h0);
  reg [(4'hd):(1'h0)] reg3925 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3924 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3923 = (1'h0);
  reg [(3'h7):(1'h0)] reg3922 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3921 = (1'h0);
  reg [(4'he):(1'h0)] forvar3920 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3919 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3915 = (1'h0);
  reg [(4'hb):(1'h0)] reg3920 = (1'h0);
  reg [(2'h2):(1'h0)] reg3919 = (1'h0);
  reg [(4'hd):(1'h0)] reg3918 = (1'h0);
  reg [(4'h9):(1'h0)] reg3917 = (1'h0);
  reg [(4'hc):(1'h0)] reg3916 = (1'h0);
  reg [(3'h7):(1'h0)] reg3915 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3914 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3913 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3912 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3911 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3910 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3909 = (1'h0);
  reg [(4'h8):(1'h0)] reg3908 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3907 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3906 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3905 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3904 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3903 = (1'h0);
  reg [(3'h4):(1'h0)] reg3902 = (1'h0);
  reg [(2'h3):(1'h0)] reg3901 = (1'h0);
  reg [(5'h10):(1'h0)] reg3900 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3899 = (1'h0);
  reg [(4'hb):(1'h0)] reg3899 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3892 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3898 = (1'h0);
  reg [(4'h9):(1'h0)] reg3897 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3894 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3885 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3878 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3877 = (1'h0);
  reg [(3'h5):(1'h0)] reg3875 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3869 = (1'h0);
  reg [(4'ha):(1'h0)] reg3870 = (1'h0);
  reg [(4'hc):(1'h0)] reg3867 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3896 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3889 = (1'h0);
  reg [(4'ha):(1'h0)] reg3895 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3894 = (1'h0);
  reg [(4'hb):(1'h0)] reg3893 = (1'h0);
  reg [(3'h5):(1'h0)] reg3892 = (1'h0);
  reg [(3'h5):(1'h0)] reg3891 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3890 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3889 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3888 = (1'h0);
  reg [(2'h3):(1'h0)] reg3887 = (1'h0);
  reg [(4'he):(1'h0)] reg3886 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3885 = (1'h0);
  reg [(4'hf):(1'h0)] reg3884 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3883 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3882 = (1'h0);
  reg [(4'hf):(1'h0)] reg3881 = (1'h0);
  reg [(4'he):(1'h0)] reg3880 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3879 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3878 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3877 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3876 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar3875 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3874 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3873 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3872 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3871 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3870 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3869 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3868 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3867 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3866 = (1'h0);
  reg [(4'ha):(1'h0)] reg3858 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3855 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3854 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3865 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3864 = (1'h0);
  reg [(4'h8):(1'h0)] reg3863 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3862 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3861 = (1'h0);
  reg [(4'hb):(1'h0)] reg3860 = (1'h0);
  reg [(3'h6):(1'h0)] reg3859 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3858 = (1'h0);
  reg [(4'hc):(1'h0)] reg3857 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3856 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3855 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3854 = (1'h0);
  reg [(4'hc):(1'h0)] reg3853 = (1'h0);
  reg [(3'h7):(1'h0)] reg3852 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3851 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3850 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3849 = (1'h0);
  reg [(4'ha):(1'h0)] reg3848 = (1'h0);
  reg [(2'h2):(1'h0)] reg3847 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3846 = (1'h0);
  reg [(4'hf):(1'h0)] reg3845 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3844 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3843 = (1'h0);
  reg [(4'hd):(1'h0)] reg3842 = (1'h0);
  reg [(2'h3):(1'h0)] reg3841 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3840 = (1'h0);
  reg [(3'h5):(1'h0)] reg3839 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3838 = (1'h0);
  reg [(4'hc):(1'h0)] reg3837 = (1'h0);
  reg [(4'hc):(1'h0)] reg3836 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3835 = (1'h0);
  reg [(3'h4):(1'h0)] reg3834 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3833 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3832 = (1'h0);
  reg [(3'h7):(1'h0)] reg3831 = (1'h0);
  reg [(5'h10):(1'h0)] reg3830 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3829 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3828 = (1'h0);
  reg [(4'ha):(1'h0)] reg3827 = (1'h0);
  reg [(4'hc):(1'h0)] reg3826 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3825 = (1'h0);
  reg [(3'h7):(1'h0)] reg3824 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3823 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3820 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3822 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3821 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3820 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar3819 = (1'h0);
  reg [(3'h5):(1'h0)] reg3818 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3817 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3816 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3815 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3814 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3812 = (1'h0);
  reg [(4'hf):(1'h0)] reg3811 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3810 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3813 = (1'h0);
  reg [(4'hb):(1'h0)] reg3812 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3811 = (1'h0);
  reg [(4'hd):(1'h0)] reg3810 = (1'h0);
  reg [(4'hd):(1'h0)] reg3809 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3808 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3807 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3806 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3805 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3804 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3803 = (1'h0);
  reg [(4'he):(1'h0)] reg3802 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3801 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3800 = (1'h0);
  reg [(4'hf):(1'h0)] reg3799 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3798 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3797 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3796 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3795 = (1'h0);
  reg [(4'hc):(1'h0)] reg3785 = (1'h0);
  reg [(3'h6):(1'h0)] reg3794 = (1'h0);
  reg [(3'h5):(1'h0)] reg3793 = (1'h0);
  reg [(3'h4):(1'h0)] reg3792 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3791 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3790 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3789 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3788 = (1'h0);
  reg [(3'h5):(1'h0)] reg3787 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3786 = (1'h0);
  reg [(4'hf):(1'h0)] forvar3785 = (1'h0);
  reg [(4'hb):(1'h0)] reg3784 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3783 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3782 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3781 = (1'h0);
  reg [(4'hf):(1'h0)] reg3780 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3779 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3778 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3777 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3776 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3775 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3774 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3773 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3772 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3771 = (1'h0);
  reg [(4'h9):(1'h0)] reg3770 = (1'h0);
  reg [(5'h10):(1'h0)] reg3769 = (1'h0);
  reg [(4'hb):(1'h0)] reg3768 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3767 = (1'h0);
  reg [(2'h3):(1'h0)] reg3766 = (1'h0);
  reg [(3'h6):(1'h0)] reg3765 = (1'h0);
  reg [(3'h6):(1'h0)] reg3764 = (1'h0);
  reg [(5'h10):(1'h0)] reg3763 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3762 = (1'h0);
  reg [(4'hf):(1'h0)] reg3761 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3760 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3759 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3758 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3757 = (1'h0);
  reg [(4'hc):(1'h0)] reg3756 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3755 = (1'h0);
  reg [(3'h4):(1'h0)] reg3754 = (1'h0);
  reg [(4'hc):(1'h0)] reg3753 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3752 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3751 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3750 = (1'h0);
  reg [(5'h10):(1'h0)] reg3749 = (1'h0);
  reg [(3'h4):(1'h0)] reg3748 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3747 = (1'h0);
  reg [(4'hc):(1'h0)] reg3746 = (1'h0);
  reg [(2'h2):(1'h0)] reg3745 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3744 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3743 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3742 = (1'h0);
  reg [(4'he):(1'h0)] reg3741 = (1'h0);
  reg [(4'h9):(1'h0)] reg3740 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3739 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3738 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3737 = (1'h0);
  reg [(3'h5):(1'h0)] reg3736 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3735 = (1'h0);
  reg [(4'hf):(1'h0)] reg3734 = (1'h0);
  reg [(5'h10):(1'h0)] reg3733 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3732 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3731 = (1'h0);
  reg [(5'h10):(1'h0)] reg3730 = (1'h0);
  reg [(4'hd):(1'h0)] reg3729 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3728 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar3727 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3726 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3725 = (1'h0);
  reg [(4'hc):(1'h0)] reg3724 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3723 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3722 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg3721 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3720 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3719 = (1'h0);
  reg [(4'he):(1'h0)] forvar3716 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar3714 = (1'h0);
  reg [(2'h3):(1'h0)] reg3711 = (1'h0);
  reg [(3'h5):(1'h0)] reg3718 = (1'h0);
  reg [(4'he):(1'h0)] reg3717 = (1'h0);
  reg [(4'h9):(1'h0)] reg3716 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3715 = (1'h0);
  reg [(4'hc):(1'h0)] reg3714 = (1'h0);
  reg [(3'h7):(1'h0)] reg3713 = (1'h0);
  reg [(4'ha):(1'h0)] reg3712 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3711 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3710 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3709 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3708 = (1'h0);
  reg [(4'h8):(1'h0)] reg3707 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3706 = (1'h0);
  reg [(3'h7):(1'h0)] reg3705 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3704 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3703 = (1'h0);
  reg [(4'he):(1'h0)] reg3702 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3701 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3700 = (1'h0);
  reg [(4'ha):(1'h0)] forvar3699 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3698 = (1'h0);
  reg [(4'ha):(1'h0)] reg3697 = (1'h0);
  reg [(3'h7):(1'h0)] reg3696 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3695 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3694 = (1'h0);
  reg [(4'hd):(1'h0)] reg3693 = (1'h0);
  reg [(4'ha):(1'h0)] reg3692 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3691 = (1'h0);
  reg [(4'ha):(1'h0)] reg3690 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3689 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3688 = (1'h0);
  reg [(5'h10):(1'h0)] reg3687 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar3686 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3685 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3684 = (1'h0);
  reg [(4'hc):(1'h0)] reg3683 = (1'h0);
  reg [(4'hd):(1'h0)] reg3682 = (1'h0);
  reg [(4'hd):(1'h0)] reg3681 = (1'h0);
  reg [(4'ha):(1'h0)] reg3680 = (1'h0);
  reg [(4'hf):(1'h0)] reg3679 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3678 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3678 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3677 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3676 = (1'h0);
  reg [(4'he):(1'h0)] reg3675 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3674 = (1'h0);
  reg [(4'hc):(1'h0)] reg3673 = (1'h0);
  reg [(4'hf):(1'h0)] reg3672 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3671 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3670 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3669 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3668 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3667 = (1'h0);
  reg [(5'h10):(1'h0)] reg3666 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3644 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3642 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3645 = (1'h0);
  reg [(4'hc):(1'h0)] reg3640 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3638 = (1'h0);
  reg [(4'hd):(1'h0)] reg3665 = (1'h0);
  reg [(4'hb):(1'h0)] reg3664 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3663 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3662 = (1'h0);
  reg [(3'h4):(1'h0)] reg3661 = (1'h0);
  reg [(3'h7):(1'h0)] reg3660 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3659 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3659 = (1'h0);
  reg [(3'h6):(1'h0)] reg3658 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3657 = (1'h0);
  reg [(4'hf):(1'h0)] reg3656 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3655 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3654 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3653 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3652 = (1'h0);
  reg [(4'he):(1'h0)] forvar3648 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3647 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3651 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3650 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg3649 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3648 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3647 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3634 = (1'h0);
  reg [(3'h5):(1'h0)] reg3646 = (1'h0);
  reg [(2'h3):(1'h0)] reg3645 = (1'h0);
  reg [(4'hd):(1'h0)] reg3644 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3643 = (1'h0);
  reg [(4'hb):(1'h0)] reg3642 = (1'h0);
  reg [(4'hd):(1'h0)] reg3641 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3640 = (1'h0);
  reg [(3'h7):(1'h0)] reg3639 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3638 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3637 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3636 = (1'h0);
  reg [(2'h2):(1'h0)] reg3635 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3634 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3633 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3632 = (1'h0);
  reg [(3'h5):(1'h0)] reg3631 = (1'h0);
  reg [(2'h3):(1'h0)] forvar3622 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3618 = (1'h0);
  reg [(4'hd):(1'h0)] reg3630 = (1'h0);
  reg [(3'h7):(1'h0)] forvar3627 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3626 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3628 = (1'h0);
  reg [(5'h10):(1'h0)] reg3627 = (1'h0);
  reg [(4'hc):(1'h0)] forvar3626 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3625 = (1'h0);
  reg [(3'h6):(1'h0)] reg3624 = (1'h0);
  reg [(3'h4):(1'h0)] reg3623 = (1'h0);
  reg [(3'h4):(1'h0)] reg3622 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3621 = (1'h0);
  reg [(4'hb):(1'h0)] reg3620 = (1'h0);
  reg [(3'h7):(1'h0)] reg3619 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3618 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg3617 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3616 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3615 = (1'h0);
  reg [(4'hc):(1'h0)] reg3614 = (1'h0);
  reg [(4'hd):(1'h0)] reg3613 = (1'h0);
  reg [(4'ha):(1'h0)] reg3612 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar3611 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3610 = (1'h0);
  wire [(2'h3):(1'h0)] wire3609;
  assign y = {wire4015,
                 reg4014,
                 reg4004,
                 forvar4000,
                 reg3999,
                 reg3998,
                 forvar3993,
                 forvar3989,
                 reg3988,
                 reg3986,
                 forvar3981,
                 forvar3975,
                 reg3974,
                 forvar3971,
                 reg4013,
                 reg4012,
                 reg4011,
                 reg4010,
                 forvar4009,
                 reg4008,
                 reg4007,
                 reg4006,
                 reg4005,
                 forvar4004,
                 reg4003,
                 reg4002,
                 reg4001,
                 reg4000,
                 forvar3999,
                 forvar3998,
                 reg3997,
                 reg3996,
                 reg3995,
                 reg3990,
                 reg3994,
                 reg3993,
                 reg3992,
                 reg3991,
                 forvar3990,
                 reg3989,
                 forvar3988,
                 reg3970,
                 forvar3969,
                 reg3966,
                 forvar3964,
                 reg3984,
                 forvar3980,
                 forvar3976,
                 reg3987,
                 forvar3986,
                 reg3985,
                 forvar3984,
                 reg3983,
                 reg3982,
                 reg3981,
                 reg3980,
                 reg3979,
                 reg3978,
                 reg3977,
                 reg3976,
                 reg3963,
                 reg3975,
                 forvar3974,
                 reg3973,
                 reg3972,
                 reg3971,
                 forvar3970,
                 reg3969,
                 reg3968,
                 reg3967,
                 forvar3966,
                 reg3965,
                 reg3964,
                 forvar3963,
                 wire3962,
                 wire3961,
                 reg3960,
                 reg3959,
                 reg3958,
                 reg3957,
                 forvar3956,
                 reg3955,
                 forvar3954,
                 reg3953,
                 reg3952,
                 forvar3951,
                 reg3950,
                 reg3949,
                 forvar3948,
                 reg3947,
                 reg3946,
                 forvar3945,
                 forvar3944,
                 reg3943,
                 reg3942,
                 reg3941,
                 reg3940,
                 reg3939,
                 forvar3938,
                 reg3937,
                 forvar3936,
                 forvar3935,
                 reg3934,
                 reg3933,
                 reg3932,
                 reg3931,
                 forvar3930,
                 reg3929,
                 forvar3928,
                 reg3927,
                 forvar3926,
                 reg3925,
                 reg3924,
                 forvar3923,
                 reg3922,
                 reg3921,
                 forvar3920,
                 forvar3919,
                 forvar3915,
                 reg3920,
                 reg3919,
                 reg3918,
                 reg3917,
                 reg3916,
                 reg3915,
                 forvar3914,
                 reg3913,
                 reg3912,
                 reg3911,
                 reg3910,
                 forvar3909,
                 reg3908,
                 reg3907,
                 reg3906,
                 reg3905,
                 forvar3904,
                 reg3903,
                 reg3902,
                 reg3901,
                 reg3900,
                 forvar3899,
                 reg3899,
                 forvar3892,
                 reg3898,
                 reg3897,
                 forvar3894,
                 reg3885,
                 reg3878,
                 forvar3877,
                 reg3875,
                 forvar3869,
                 reg3870,
                 reg3867,
                 reg3896,
                 reg3889,
                 reg3895,
                 reg3894,
                 reg3893,
                 reg3892,
                 reg3891,
                 reg3890,
                 forvar3889,
                 reg3888,
                 reg3887,
                 reg3886,
                 forvar3885,
                 reg3884,
                 forvar3883,
                 reg3882,
                 reg3881,
                 reg3880,
                 reg3879,
                 forvar3878,
                 reg3877,
                 reg3876,
                 forvar3875,
                 reg3874,
                 reg3873,
                 reg3872,
                 reg3871,
                 forvar3870,
                 reg3869,
                 reg3868,
                 forvar3867,
                 forvar3866,
                 reg3858,
                 reg3855,
                 forvar3854,
                 reg3865,
                 reg3864,
                 reg3863,
                 forvar3862,
                 reg3861,
                 reg3860,
                 reg3859,
                 forvar3858,
                 reg3857,
                 reg3856,
                 forvar3855,
                 reg3854,
                 reg3853,
                 reg3852,
                 reg3851,
                 forvar3850,
                 reg3849,
                 reg3848,
                 reg3847,
                 reg3846,
                 reg3845,
                 forvar3844,
                 reg3843,
                 reg3842,
                 reg3841,
                 forvar3840,
                 reg3839,
                 reg3838,
                 reg3837,
                 reg3836,
                 reg3835,
                 reg3834,
                 reg3833,
                 reg3832,
                 reg3831,
                 reg3830,
                 forvar3829,
                 reg3828,
                 reg3827,
                 reg3826,
                 reg3825,
                 reg3824,
                 forvar3823,
                 forvar3820,
                 reg3822,
                 forvar3821,
                 reg3820,
                 forvar3819,
                 reg3818,
                 reg3817,
                 reg3816,
                 reg3815,
                 forvar3814,
                 forvar3812,
                 reg3811,
                 forvar3810,
                 reg3813,
                 reg3812,
                 forvar3811,
                 reg3810,
                 reg3809,
                 forvar3808,
                 forvar3807,
                 reg3806,
                 forvar3805,
                 forvar3804,
                 reg3803,
                 reg3802,
                 reg3801,
                 reg3800,
                 reg3799,
                 forvar3798,
                 forvar3797,
                 forvar3796,
                 reg3795,
                 reg3785,
                 reg3794,
                 reg3793,
                 reg3792,
                 reg3791,
                 reg3790,
                 reg3789,
                 reg3788,
                 reg3787,
                 reg3786,
                 forvar3785,
                 reg3784,
                 reg3783,
                 reg3782,
                 forvar3781,
                 reg3780,
                 reg3779,
                 reg3778,
                 reg3777,
                 forvar3776,
                 reg3775,
                 forvar3774,
                 reg3773,
                 reg3772,
                 reg3771,
                 reg3770,
                 reg3769,
                 reg3768,
                 reg3767,
                 reg3766,
                 reg3765,
                 reg3764,
                 reg3763,
                 reg3762,
                 reg3761,
                 forvar3760,
                 forvar3759,
                 forvar3758,
                 reg3757,
                 reg3756,
                 forvar3755,
                 reg3754,
                 reg3753,
                 reg3752,
                 reg3751,
                 forvar3750,
                 reg3749,
                 reg3748,
                 reg3747,
                 reg3746,
                 reg3745,
                 reg3744,
                 forvar3743,
                 forvar3742,
                 reg3741,
                 reg3740,
                 reg3739,
                 reg3738,
                 forvar3737,
                 reg3736,
                 reg3735,
                 reg3734,
                 reg3733,
                 forvar3732,
                 reg3731,
                 reg3730,
                 reg3729,
                 forvar3728,
                 forvar3727,
                 reg3726,
                 forvar3725,
                 reg3724,
                 reg3723,
                 reg3722,
                 reg3721,
                 forvar3720,
                 reg3719,
                 forvar3716,
                 forvar3714,
                 reg3711,
                 reg3718,
                 reg3717,
                 reg3716,
                 reg3715,
                 reg3714,
                 reg3713,
                 reg3712,
                 forvar3711,
                 reg3710,
                 reg3709,
                 reg3708,
                 reg3707,
                 reg3706,
                 reg3705,
                 forvar3704,
                 reg3703,
                 reg3702,
                 forvar3701,
                 reg3700,
                 forvar3699,
                 reg3698,
                 reg3697,
                 reg3696,
                 forvar3695,
                 forvar3694,
                 reg3693,
                 reg3692,
                 reg3691,
                 reg3690,
                 forvar3689,
                 forvar3688,
                 reg3687,
                 forvar3686,
                 reg3685,
                 reg3684,
                 reg3683,
                 reg3682,
                 reg3681,
                 reg3680,
                 reg3679,
                 forvar3678,
                 reg3678,
                 reg3677,
                 reg3676,
                 reg3675,
                 reg3674,
                 reg3673,
                 reg3672,
                 reg3671,
                 forvar3670,
                 reg3669,
                 forvar3668,
                 forvar3667,
                 reg3666,
                 forvar3644,
                 forvar3642,
                 forvar3645,
                 reg3640,
                 forvar3638,
                 reg3665,
                 reg3664,
                 forvar3663,
                 reg3662,
                 reg3661,
                 reg3660,
                 forvar3659,
                 reg3659,
                 reg3658,
                 reg3657,
                 reg3656,
                 reg3655,
                 forvar3654,
                 reg3653,
                 reg3652,
                 forvar3648,
                 reg3647,
                 reg3651,
                 reg3650,
                 reg3649,
                 reg3648,
                 forvar3647,
                 reg3634,
                 reg3646,
                 reg3645,
                 reg3644,
                 reg3643,
                 reg3642,
                 reg3641,
                 forvar3640,
                 reg3639,
                 reg3638,
                 reg3637,
                 reg3636,
                 reg3635,
                 forvar3634,
                 reg3633,
                 reg3632,
                 reg3631,
                 forvar3622,
                 forvar3618,
                 reg3630,
                 forvar3627,
                 reg3626,
                 reg3629,
                 reg3628,
                 reg3627,
                 forvar3626,
                 reg3625,
                 reg3624,
                 reg3623,
                 reg3622,
                 reg3621,
                 reg3620,
                 reg3619,
                 reg3618,
                 reg3617,
                 forvar3616,
                 reg3615,
                 reg3614,
                 reg3613,
                 reg3612,
                 forvar3611,
                 forvar3610,
                 wire3609,
                 (1'h0)};
  assign wire3609 = (wire3608[(5'h10):(4'hf)] & {((8'ha5) ?
                            $unsigned(wire3605) : $signed(wire3605))});
  always
    @(posedge clk) begin
      for (forvar3610 = (1'h0); (forvar3610 < (1'h0)); forvar3610 = (forvar3610 + (1'h1)))
        begin
          if ((-wire3609[(2'h2):(1'h1)]))
            begin
              for (forvar3611 = (1'h0); (forvar3611 < (2'h3)); forvar3611 = (forvar3611 + (1'h1)))
                begin
                  if (wire3606[(3'h6):(2'h3)])
                    begin
                      reg3612 <= wire3606[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg3612 <= ((~&forvar3610[(2'h2):(1'h1)]) ?
                          (wire3604 >= ($signed(wire3607) < $signed(reg3612))) : ({$signed(wire3604)} != {(~|wire3608)}));
                      reg3613 <= (+$signed((|wire3606)));
                      reg3614 <= ((+($signed(forvar3611) >>> {reg3613})) ?
                          wire3608 : forvar3610[(2'h3):(2'h3)]);
                      reg3615 <= $unsigned($signed(reg3612));
                    end
                  for (forvar3616 = (1'h0); (forvar3616 < (2'h3)); forvar3616 = (forvar3616 + (1'h1)))
                    begin
                      reg3617 <= $unsigned((~|forvar3616));
                      reg3618 <= $signed(reg3615);
                      reg3619 <= $unsigned(wire3608[(4'h9):(4'h8)]);
                      reg3620 <= ((((reg3617 ? reg3613 : (8'hb6)) ?
                          (-(8'ha8)) : $signed(reg3617)) & ((reg3612 ?
                          (8'hba) : forvar3616) || (forvar3611 ?
                          reg3614 : reg3617))) >> ((((8'h9e) ?
                                  reg3613 : forvar3611) ?
                              wire3607[(2'h3):(2'h3)] : wire3606[(4'hb):(4'h9)]) ?
                          reg3618 : ($unsigned(reg3614) ?
                              (&reg3614) : wire3606[(3'h4):(1'h1)])));
                    end
                  reg3621 <= reg3615;
                  if ($signed((wire3608[(4'hd):(4'hd)] ^~ {$signed(reg3614)})))
                    begin
                      reg3622 <= (^~$signed($signed((8'h9d))));
                      reg3623 <= ($unsigned(((~^reg3619) != $signed(reg3614))) ?
                          forvar3616 : (($unsigned(reg3621) <= $unsigned(reg3621)) ~^ $unsigned((reg3614 ?
                              reg3619 : wire3605))));
                    end
                  else
                    begin
                      reg3622 <= ((~|(^((8'hb8) <<< forvar3610))) ?
                          wire3607 : wire3608);
                      reg3623 <= ($unsigned(wire3604) ?
                          (^forvar3610) : reg3620);
                      reg3624 <= forvar3611;
                      reg3625 <= $unsigned($unsigned((8'hae)));
                    end
                end
              if ($signed($signed(reg3617)))
                begin
                  for (forvar3626 = (1'h0); (forvar3626 < (2'h3)); forvar3626 = (forvar3626 + (1'h1)))
                    begin
                      reg3627 <= (((((8'hb0) ? (8'hb6) : reg3617) ?
                              reg3612 : $unsigned(reg3620)) <= {(!reg3618)}) ?
                          $signed($signed($signed(reg3613))) : (|{$unsigned((8'ha7))}));
                      reg3628 <= (reg3621[(3'h7):(1'h1)] ?
                          {(~reg3620)} : (reg3612 ?
                              ((^reg3621) >= (reg3612 ?
                                  reg3614 : (8'ha0))) : ((~|reg3615) ?
                                  reg3623 : (wire3607 | reg3627))));
                      reg3629 <= {(8'hac)};
                    end
                end
              else
                begin
                  reg3626 <= (~|reg3623[(1'h0):(1'h0)]);
                  for (forvar3627 = (1'h0); (forvar3627 < (2'h2)); forvar3627 = (forvar3627 + (1'h1)))
                    begin
                      reg3628 <= forvar3626;
                      reg3629 <= (~&(|{reg3627[(4'h8):(4'h8)]}));
                    end
                  reg3630 <= (~^((!(wire3609 << forvar3610)) * $unsigned($signed(wire3607))));
                end
            end
          else
            begin
              for (forvar3611 = (1'h0); (forvar3611 < (1'h1)); forvar3611 = (forvar3611 + (1'h1)))
                begin
                  if ($unsigned((^~(8'ha5))))
                    begin
                      reg3612 <= (8'ha2);
                      reg3613 <= wire3606;
                      reg3614 <= $signed({reg3626[(3'h5):(3'h5)]});
                      reg3615 <= {{$unsigned(wire3605)}};
                    end
                  else
                    begin
                      reg3612 <= {(-reg3623)};
                      reg3613 <= ($unsigned(($signed(reg3623) <<< reg3612)) ?
                          (+reg3625) : forvar3610[(3'h4):(3'h4)]);
                      reg3614 <= reg3630[(3'h7):(3'h7)];
                      reg3615 <= $signed((-(~&$signed(reg3623))));
                    end
                  for (forvar3616 = (1'h0); (forvar3616 < (1'h0)); forvar3616 = (forvar3616 + (1'h1)))
                    begin
                      reg3617 <= ((^(8'had)) >>> ((~|(~(8'hb7))) >= $unsigned((^reg3615))));
                    end
                  for (forvar3618 = (1'h0); (forvar3618 < (1'h1)); forvar3618 = (forvar3618 + (1'h1)))
                    begin
                      reg3619 <= ($signed(forvar3626[(4'ha):(4'h9)]) ?
                          wire3608 : $unsigned(forvar3610[(3'h5):(2'h3)]));
                      reg3620 <= wire3605;
                    end
                end
              if ($signed(((&reg3621[(2'h3):(2'h3)]) ?
                  $unsigned({reg3628}) : (reg3617 >= (&reg3617)))))
                begin
                  reg3621 <= $signed(forvar3626[(2'h2):(1'h0)]);
                  for (forvar3622 = (1'h0); (forvar3622 < (2'h3)); forvar3622 = (forvar3622 + (1'h1)))
                    begin
                      reg3623 <= reg3621;
                      reg3624 <= {($signed(reg3613) ?
                              ((~^reg3613) >> (forvar3610 + forvar3622)) : reg3613[(4'hd):(3'h6)])};
                      reg3625 <= ((|wire3606[(2'h3):(1'h0)]) ?
                          $unsigned($unsigned(((8'hb7) ?
                              reg3617 : reg3612))) : $unsigned(reg3625[(5'h10):(5'h10)]));
                      reg3626 <= $signed({reg3613});
                    end
                end
              else
                begin
                  if ({reg3628[(1'h1):(1'h0)]})
                    begin
                      reg3621 <= $unsigned($unsigned(((reg3612 + reg3615) ?
                          $signed((8'ha5)) : reg3618[(2'h3):(2'h2)])));
                      reg3622 <= reg3623[(1'h0):(1'h0)];
                      reg3623 <= $signed((^{forvar3610[(2'h3):(2'h2)]}));
                    end
                  else
                    begin
                      reg3621 <= (($unsigned((^~reg3627)) >>> $unsigned($unsigned(reg3620))) && $unsigned((^~(8'ha5))));
                      reg3622 <= reg3622[(2'h2):(1'h0)];
                    end
                  if ((~^$unsigned((((8'hb0) ? reg3629 : wire3607) ?
                      (&forvar3616) : (&forvar3626)))))
                    begin
                      reg3624 <= $signed(wire3606);
                      reg3625 <= wire3609;
                      reg3626 <= reg3614;
                    end
                  else
                    begin
                      reg3624 <= reg3617;
                    end
                  if (forvar3626[(4'hb):(3'h6)])
                    begin
                      reg3627 <= {(8'ha4)};
                      reg3628 <= {$signed(({reg3612} ?
                              reg3614[(3'h7):(3'h5)] : (forvar3610 ?
                                  (8'hba) : forvar3616)))};
                      reg3629 <= $signed((^reg3624[(2'h2):(2'h2)]));
                    end
                  else
                    begin
                      reg3627 <= {forvar3622[(2'h2):(1'h1)]};
                      reg3628 <= (forvar3611[(1'h1):(1'h1)] | (8'ha1));
                      reg3629 <= (^(((reg3613 ? reg3624 : (8'hb2)) ?
                          (^~forvar3611) : reg3621) <<< {{reg3622}}));
                    end
                  if (reg3618[(1'h1):(1'h0)])
                    begin
                      reg3630 <= (|$signed(reg3614));
                      reg3631 <= $signed(reg3623);
                    end
                  else
                    begin
                      reg3630 <= $unsigned((~&(|{wire3604})));
                      reg3631 <= forvar3616[(2'h3):(1'h0)];
                      reg3632 <= {(reg3614 ^~ $unsigned((-wire3606)))};
                    end
                end
              reg3633 <= {$signed(reg3617[(4'hb):(3'h6)])};
            end
          if ((8'h9e))
            begin
              if ($unsigned(reg3627))
                begin
                  for (forvar3634 = (1'h0); (forvar3634 < (2'h3)); forvar3634 = (forvar3634 + (1'h1)))
                    begin
                      reg3635 <= (wire3606[(4'hb):(1'h1)] < wire3604);
                    end
                  if (reg3618)
                    begin
                      reg3636 <= $unsigned(reg3618);
                      reg3637 <= (forvar3626 & $signed((~|$unsigned(forvar3626))));
                      reg3638 <= (({{reg3612}} != ({reg3627} ?
                          (reg3623 << (8'hb3)) : $signed(forvar3616))) <<< $signed(((&(8'hb2)) ^~ reg3623)));
                      reg3639 <= reg3627[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg3636 <= reg3637[(4'hc):(4'h8)];
                      reg3637 <= ((wire3606[(1'h0):(1'h0)] ?
                          ($signed(reg3612) ^~ reg3629[(3'h4):(2'h3)]) : (8'h9d)) < reg3639[(2'h2):(2'h2)]);
                      reg3638 <= ((-$signed((forvar3610 ?
                          wire3606 : wire3607))) - ((~(reg3623 ?
                              (8'hb1) : forvar3618)) ?
                          ((&forvar3627) ?
                              $unsigned(reg3639) : (~|reg3626)) : reg3624[(1'h0):(1'h0)]));
                    end
                  for (forvar3640 = (1'h0); (forvar3640 < (2'h3)); forvar3640 = (forvar3640 + (1'h1)))
                    begin
                      reg3641 <= ((($signed(reg3620) >> $signed(forvar3626)) ?
                          (forvar3618[(4'hc):(3'h6)] != $unsigned((8'hba))) : forvar3610[(1'h1):(1'h1)]) || ($unsigned(((8'hb8) ?
                              reg3635 : (8'hac))) ?
                          (forvar3618 ?
                              (wire3609 <<< forvar3640) : $unsigned(reg3636)) : $unsigned(reg3623)));
                      reg3642 <= {{(^reg3641)}};
                    end
                  if (({(forvar3610[(3'h5):(2'h2)] ?
                              {reg3626} : $signed(reg3635))} ?
                      wire3606[(4'h8):(3'h6)] : forvar3618))
                    begin
                      reg3643 <= (forvar3618[(1'h0):(1'h0)] ?
                          (reg3637[(3'h4):(1'h1)] | ($unsigned(reg3625) ?
                              (-(8'hb8)) : $signed(wire3606))) : (~reg3641));
                      reg3644 <= ((({(8'ha5)} <<< reg3622) ?
                          (|(~wire3606)) : $unsigned((~^reg3612))) == $signed((~&$unsigned((8'hb7)))));
                      reg3645 <= $signed($signed($signed({wire3604})));
                      reg3646 <= ((!$unsigned(reg3627[(2'h2):(1'h0)])) <<< ($signed($unsigned(reg3635)) ?
                          $signed(((8'ha0) ?
                              forvar3634 : reg3613)) : ($unsigned(reg3622) < $signed((8'ha7)))));
                    end
                  else
                    begin
                      reg3643 <= $signed(wire3607[(4'h8):(3'h5)]);
                      reg3644 <= (^~((reg3645[(1'h1):(1'h1)] ?
                          (forvar3618 ?
                              reg3613 : reg3639) : (8'hb6)) >= forvar3611));
                      reg3645 <= reg3643[(2'h3):(2'h3)];
                    end
                end
              else
                begin
                  reg3634 <= $signed($signed(wire3604[(2'h2):(2'h2)]));
                  if (wire3606)
                    begin
                      reg3635 <= (+$unsigned((|{wire3606})));
                    end
                  else
                    begin
                      reg3635 <= (reg3612 < $signed(((reg3617 ?
                          reg3630 : forvar3616) >> $signed(reg3643))));
                      reg3636 <= reg3613[(2'h2):(1'h0)];
                      reg3637 <= (reg3642[(4'h8):(4'h8)] ^ ((^$unsigned(reg3626)) ?
                          ($signed((8'haf)) << wire3604) : reg3645[(1'h0):(1'h0)]));
                      reg3638 <= $signed(reg3614[(4'h8):(3'h4)]);
                    end
                end
              if (forvar3618)
                begin
                  for (forvar3647 = (1'h0); (forvar3647 < (2'h2)); forvar3647 = (forvar3647 + (1'h1)))
                    begin
                      reg3648 <= reg3645[(2'h3):(1'h0)];
                      reg3649 <= $unsigned($unsigned(reg3612));
                      reg3650 <= ((-($signed(reg3628) ?
                              $signed(wire3606) : reg3619)) ?
                          $signed(reg3634[(3'h7):(1'h0)]) : forvar3627[(3'h6):(1'h1)]);
                      reg3651 <= ($signed(reg3636) ?
                          reg3615 : reg3624[(3'h6):(2'h2)]);
                    end
                end
              else
                begin
                  reg3647 <= wire3607[(4'h9):(3'h7)];
                  for (forvar3648 = (1'h0); (forvar3648 < (2'h2)); forvar3648 = (forvar3648 + (1'h1)))
                    begin
                      reg3649 <= reg3625;
                      reg3650 <= ({$unsigned((reg3650 & reg3634))} ?
                          forvar3627 : {reg3651[(3'h6):(3'h4)]});
                      reg3651 <= {($signed(reg3636) ?
                              $signed((reg3620 ?
                                  reg3632 : (8'haf))) : $unsigned((~&reg3623)))};
                      reg3652 <= (($signed(forvar3618) & $signed(((8'hab) ?
                              reg3642 : reg3648))) ?
                          (8'hb3) : reg3651[(4'hb):(3'h5)]);
                    end
                  reg3653 <= $unsigned((^$signed(forvar3640[(4'ha):(3'h7)])));
                  for (forvar3654 = (1'h0); (forvar3654 < (1'h0)); forvar3654 = (forvar3654 + (1'h1)))
                    begin
                      reg3655 <= (((-{reg3631}) ?
                          forvar3626[(4'ha):(1'h1)] : forvar3640) * reg3623);
                    end
                end
              if ((((^(forvar3611 ? reg3650 : reg3621)) ?
                  wire3609 : (^(reg3650 ? (8'hab) : reg3620))) >>> (8'ha4)))
                begin
                  if ($unsigned(reg3637[(2'h2):(2'h2)]))
                    begin
                      reg3656 <= wire3605;
                      reg3657 <= $signed((~$signed($signed(reg3626))));
                      reg3658 <= $unsigned((+(reg3652[(4'hc):(3'h5)] ?
                          reg3620[(4'hb):(3'h4)] : reg3628[(2'h2):(2'h2)])));
                      reg3659 <= ((~^(^((8'hb3) ? reg3657 : reg3615))) ?
                          (({reg3634} ?
                              (forvar3616 != reg3621) : (reg3653 + reg3612)) & ((8'ha9) ^~ $signed(reg3648))) : {(8'hba)});
                    end
                  else
                    begin
                      reg3656 <= (~{(~^{forvar3647})});
                      reg3657 <= $unsigned($signed($signed({reg3647})));
                      reg3658 <= {$signed(forvar3654)};
                      reg3659 <= reg3613[(3'h6):(3'h5)];
                    end
                end
              else
                begin
                  if (($unsigned(($signed(reg3626) ?
                          (reg3643 ? reg3630 : reg3650) : $signed(reg3647))) ?
                      (forvar3648[(1'h1):(1'h1)] ?
                          {(^forvar3626)} : {(^~reg3628)}) : (-reg3634)))
                    begin
                      reg3656 <= $signed((~&reg3636[(1'h0):(1'h0)]));
                      reg3657 <= (reg3613 ?
                          $unsigned(reg3653) : ({$signed(reg3627)} ?
                              $signed($signed(reg3613)) : $signed((reg3627 ?
                                  reg3612 : wire3604))));
                    end
                  else
                    begin
                      reg3656 <= ({(8'hb1)} ?
                          ((wire3608 << (forvar3610 ? reg3627 : wire3607)) ?
                              reg3643 : ((reg3635 ?
                                  reg3628 : reg3637) & (~reg3636))) : forvar3626[(3'h7):(3'h6)]);
                      reg3657 <= $unsigned((reg3620 + reg3625[(2'h2):(1'h0)]));
                      reg3658 <= ($signed(forvar3622[(1'h0):(1'h0)]) <= (~^((~|reg3613) >= forvar3634[(1'h0):(1'h0)])));
                    end
                  for (forvar3659 = (1'h0); (forvar3659 < (1'h0)); forvar3659 = (forvar3659 + (1'h1)))
                    begin
                      reg3660 <= (($unsigned((~^reg3636)) ?
                          reg3647 : reg3634) != reg3652[(3'h7):(3'h6)]);
                      reg3661 <= (8'hb1);
                      reg3662 <= ({reg3644[(1'h0):(1'h0)]} ?
                          $signed($signed(forvar3610[(1'h0):(1'h0)])) : reg3618);
                    end
                  for (forvar3663 = (1'h0); (forvar3663 < (2'h3)); forvar3663 = (forvar3663 + (1'h1)))
                    begin
                      reg3664 <= {(((forvar3640 < (8'hab)) - ((8'ha6) - forvar3634)) ?
                              $unsigned((reg3661 >> reg3628)) : ((wire3604 ?
                                      reg3649 : forvar3654) ?
                                  (reg3653 || (8'ha3)) : (+reg3660)))};
                      reg3665 <= (8'hba);
                    end
                end
            end
          else
            begin
              reg3634 <= $signed((8'ha4));
              if (((forvar3654[(3'h7):(3'h7)] << (((8'hac) * (8'ha2)) >> $signed(reg3643))) ?
                  (((reg3625 ? reg3623 : forvar3616) ~^ reg3653) ?
                      $unsigned($signed(reg3659)) : reg3637) : (~^$unsigned($signed(reg3647)))))
                begin
                  if (((reg3639 >> {$unsigned(reg3612)}) ?
                      (forvar3626[(3'h5):(2'h2)] ?
                          $signed((reg3620 ?
                              (8'hab) : reg3628)) : (8'hb1)) : (~&reg3657[(1'h1):(1'h0)])))
                    begin
                      reg3635 <= reg3652;
                      reg3636 <= $unsigned(reg3658);
                    end
                  else
                    begin
                      reg3635 <= (!$signed((-reg3652[(3'h4):(2'h2)])));
                      reg3636 <= (~|$signed($signed((~&reg3644))));
                      reg3637 <= reg3619;
                      reg3638 <= $signed(wire3604);
                    end
                  reg3639 <= reg3652;
                end
              else
                begin
                  reg3635 <= {({reg3631[(1'h0):(1'h0)]} >> ((8'ha9) ?
                          (reg3647 ? reg3624 : forvar3626) : (reg3619 ?
                              forvar3622 : reg3626)))};
                  if ($unsigned(($unsigned((reg3644 <<< wire3607)) ?
                      (!{reg3658}) : {(~^reg3635)})))
                    begin
                      reg3636 <= reg3647[(4'hf):(3'h4)];
                      reg3637 <= $signed($signed((|(reg3656 >> reg3625))));
                    end
                  else
                    begin
                      reg3636 <= ({(&((8'ha7) ?
                              reg3643 : reg3632))} >> reg3661[(3'h4):(1'h1)]);
                      reg3637 <= ((-{$signed((8'hb9))}) >> {($unsigned(forvar3618) ?
                              forvar3647[(1'h1):(1'h0)] : (reg3612 < reg3649))});
                    end
                  for (forvar3638 = (1'h0); (forvar3638 < (2'h3)); forvar3638 = (forvar3638 + (1'h1)))
                    begin
                      reg3639 <= $signed($unsigned((wire3609[(2'h3):(2'h3)] | reg3664[(2'h2):(2'h2)])));
                      reg3640 <= reg3657[(4'hc):(2'h2)];
                      reg3641 <= (-$signed($signed($signed(reg3636))));
                    end
                end
              if ({((-$unsigned(forvar3611)) ?
                      reg3631[(1'h1):(1'h1)] : (&$signed((8'ha1))))})
                begin
                  if ($signed({reg3635[(1'h1):(1'h1)]}))
                    begin
                      reg3642 <= (-(8'ha2));
                      reg3643 <= reg3650[(4'hb):(3'h4)];
                      reg3644 <= $unsigned({reg3659[(4'hd):(3'h5)]});
                    end
                  else
                    begin
                      reg3642 <= reg3642[(4'h8):(3'h6)];
                      reg3643 <= ((reg3665 ?
                              $unsigned((|forvar3616)) : (8'ha8)) ?
                          $signed(reg3625[(3'h6):(1'h1)]) : (reg3641 ?
                              $signed(wire3607[(2'h3):(2'h2)]) : ((reg3631 << reg3630) ?
                                  (8'hb1) : $signed(wire3606))));
                      reg3644 <= reg3652;
                    end
                  for (forvar3645 = (1'h0); (forvar3645 < (2'h3)); forvar3645 = (forvar3645 + (1'h1)))
                    begin
                      reg3646 <= $signed(forvar3634);
                      reg3647 <= reg3647;
                      reg3648 <= reg3628[(1'h1):(1'h0)];
                      reg3649 <= ($unsigned((reg3648[(1'h1):(1'h0)] ^~ $signed(forvar3627))) ^~ $signed((~^(+reg3641))));
                    end
                  if ($unsigned(reg3644))
                    begin
                      reg3650 <= (-(&$unsigned((+reg3632))));
                      reg3651 <= reg3642[(1'h1):(1'h0)];
                      reg3652 <= (^reg3658);
                    end
                  else
                    begin
                      reg3650 <= $unsigned($unsigned(reg3619));
                      reg3651 <= (^~$unsigned((!$signed(reg3619))));
                    end
                  reg3653 <= $signed($unsigned(((wire3608 ?
                      (8'hac) : reg3615) == $unsigned((8'haa)))));
                end
              else
                begin
                  for (forvar3642 = (1'h0); (forvar3642 < (2'h2)); forvar3642 = (forvar3642 + (1'h1)))
                    begin
                      reg3643 <= reg3624;
                    end
                  for (forvar3644 = (1'h0); (forvar3644 < (1'h0)); forvar3644 = (forvar3644 + (1'h1)))
                    begin
                      reg3645 <= $unsigned(forvar3638[(3'h6):(3'h6)]);
                      reg3646 <= $unsigned($signed($unsigned((^~(8'ha2)))));
                      reg3647 <= {($unsigned((reg3614 ^~ reg3653)) ?
                              forvar3642 : reg3619[(3'h5):(3'h5)])};
                    end
                end
              for (forvar3654 = (1'h0); (forvar3654 < (2'h3)); forvar3654 = (forvar3654 + (1'h1)))
                begin
                  if ((&((reg3615[(2'h2):(2'h2)] == ((8'haa) ?
                          reg3636 : forvar3659)) ?
                      ($signed(reg3642) ?
                          ((8'ha8) ?
                              (8'h9f) : (8'hba)) : reg3646[(3'h5):(3'h4)]) : (forvar3645[(3'h4):(2'h2)] <= (~^forvar3648)))))
                    begin
                      reg3655 <= $unsigned(($signed({(8'hb7)}) ?
                          {wire3607[(2'h2):(2'h2)]} : $signed($unsigned(reg3626))));
                    end
                  else
                    begin
                      reg3655 <= wire3604[(3'h4):(1'h1)];
                      reg3656 <= reg3642;
                      reg3657 <= $unsigned(((reg3625[(3'h5):(3'h4)] ?
                          $signed(reg3627) : $signed(reg3633)) != wire3609));
                      reg3658 <= reg3638;
                    end
                end
            end
        end
      reg3666 <= $unsigned($signed(reg3657[(1'h0):(1'h0)]));
      for (forvar3667 = (1'h0); (forvar3667 < (2'h2)); forvar3667 = (forvar3667 + (1'h1)))
        begin
          for (forvar3668 = (1'h0); (forvar3668 < (2'h2)); forvar3668 = (forvar3668 + (1'h1)))
            begin
              reg3669 <= (&$unsigned((~reg3620)));
              for (forvar3670 = (1'h0); (forvar3670 < (2'h2)); forvar3670 = (forvar3670 + (1'h1)))
                begin
                  reg3671 <= $unsigned((~($unsigned(wire3605) ?
                      $unsigned((8'hb6)) : $unsigned((8'ha7)))));
                  reg3672 <= $unsigned($signed($unsigned($signed((8'ha1)))));
                  reg3673 <= (((reg3660 ?
                          (reg3652 ^ reg3666) : (reg3661 ?
                              reg3662 : reg3651)) || {(|wire3608)}) ?
                      (wire3609[(1'h0):(1'h0)] ~^ $unsigned($signed(forvar3654))) : ((reg3653[(3'h6):(3'h6)] ?
                          (reg3653 <<< forvar3644) : $unsigned(reg3643)) <= $signed($unsigned(wire3606))));
                  reg3674 <= ($signed(reg3626) << (^{reg3645[(1'h0):(1'h0)]}));
                end
              reg3675 <= ({reg3646} << (($unsigned(forvar3634) ?
                  reg3614 : reg3672) >>> ({(8'hb3)} ?
                  reg3662[(3'h4):(2'h2)] : (reg3629 ? reg3641 : reg3656))));
              reg3676 <= $unsigned((~^(forvar3611 ?
                  reg3619 : (reg3664 >> forvar3627))));
            end
          reg3677 <= {((+$unsigned((8'hb3))) >>> $unsigned(wire3609))};
        end
      if ((forvar3622 >= $unsigned($unsigned(forvar3622))))
        begin
          reg3678 <= reg3671;
        end
      else
        begin
          for (forvar3678 = (1'h0); (forvar3678 < (2'h2)); forvar3678 = (forvar3678 + (1'h1)))
            begin
              if ({(^(wire3604 ? reg3623 : $signed(reg3647)))})
                begin
                  if ((|(-$signed((reg3613 & forvar3626)))))
                    begin
                      reg3679 <= reg3623;
                      reg3680 <= reg3671[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg3679 <= reg3679[(2'h2):(1'h0)];
                    end
                  if ((reg3661[(3'h4):(2'h2)] && reg3613))
                    begin
                      reg3681 <= reg3625[(3'h5):(2'h2)];
                      reg3682 <= $signed(({(+reg3657)} * (reg3639[(1'h0):(1'h0)] & reg3645[(1'h1):(1'h1)])));
                      reg3683 <= reg3679;
                      reg3684 <= ((^reg3638[(4'ha):(4'ha)]) ?
                          (($unsigned((8'hb6)) ?
                                  $unsigned(forvar3616) : $signed(reg3618)) ?
                              $unsigned((reg3632 > reg3676)) : ({forvar3663} ?
                                  (8'hac) : reg3656)) : ((!forvar3638[(3'h5):(1'h1)]) ?
                              $signed(((8'hb5) ?
                                  wire3604 : reg3623)) : $signed(reg3673[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg3681 <= reg3624;
                      reg3682 <= reg3671;
                      reg3683 <= (~^(({reg3621} >= (reg3655 ?
                          (8'ha2) : reg3666)) <<< (forvar3618[(3'h5):(2'h2)] ?
                          ((8'hab) <<< (8'ha8)) : {forvar3668})));
                      reg3684 <= $unsigned(reg3656);
                    end
                end
              else
                begin
                  if ((reg3664[(4'hb):(4'h8)] ?
                      (~^(^reg3648)) : reg3637[(3'h7):(3'h6)]))
                    begin
                      reg3679 <= ((reg3648[(1'h1):(1'h1)] << ($unsigned(forvar3663) ?
                          (+reg3641) : (^~forvar3640))) ^~ (~|(^~((8'haa) ?
                          reg3620 : forvar3616))));
                      reg3680 <= $unsigned(({(reg3650 >>> reg3638)} ?
                          ($unsigned(forvar3642) > wire3609) : $signed($signed(reg3684))));
                    end
                  else
                    begin
                      reg3679 <= (reg3656[(4'ha):(4'h9)] & ($signed($signed(reg3649)) ?
                          ((&(8'hb5)) ?
                              $signed(forvar3678) : $unsigned(forvar3648)) : $signed(reg3678)));
                    end
                  reg3681 <= (reg3679[(2'h3):(1'h0)] ?
                      ($signed($signed(forvar3634)) <<< {(&(8'hac))}) : wire3606);
                  if ($unsigned(forvar3638))
                    begin
                      reg3682 <= $signed((-forvar3654));
                      reg3683 <= ($signed(reg3624[(3'h5):(2'h2)]) ?
                          {{wire3609[(2'h2):(2'h2)]}} : forvar3667);
                      reg3684 <= $signed(reg3613);
                      reg3685 <= reg3627[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg3682 <= $unsigned(reg3680[(4'h8):(1'h0)]);
                      reg3683 <= reg3634[(1'h0):(1'h0)];
                      reg3684 <= reg3636;
                    end
                  for (forvar3686 = (1'h0); (forvar3686 < (2'h2)); forvar3686 = (forvar3686 + (1'h1)))
                    begin
                      reg3687 <= ((wire3607[(2'h2):(1'h1)] ?
                          reg3644 : reg3646[(2'h2):(2'h2)]) - {forvar3622[(1'h0):(1'h0)]});
                    end
                end
              for (forvar3688 = (1'h0); (forvar3688 < (2'h2)); forvar3688 = (forvar3688 + (1'h1)))
                begin
                  for (forvar3689 = (1'h0); (forvar3689 < (2'h3)); forvar3689 = (forvar3689 + (1'h1)))
                    begin
                      reg3690 <= {$signed((8'hb0))};
                      reg3691 <= (-(((reg3644 == reg3631) != wire3609) ?
                          $signed((reg3633 ?
                              reg3641 : reg3612)) : $unsigned((|forvar3648))));
                      reg3692 <= (forvar3668 ?
                          reg3621 : ($unsigned(reg3671) ?
                              (forvar3668 && {forvar3686}) : ($signed(reg3622) ~^ $unsigned(forvar3642))));
                      reg3693 <= forvar3616;
                    end
                end
            end
          for (forvar3694 = (1'h0); (forvar3694 < (2'h3)); forvar3694 = (forvar3694 + (1'h1)))
            begin
              for (forvar3695 = (1'h0); (forvar3695 < (2'h2)); forvar3695 = (forvar3695 + (1'h1)))
                begin
                  if ($signed((^~{reg3646[(3'h5):(3'h5)]})))
                    begin
                      reg3696 <= $signed((($signed(reg3678) ?
                              (+reg3642) : {forvar3645}) ?
                          ((&reg3632) ^ (reg3628 != reg3662)) : $unsigned($signed(reg3684))));
                    end
                  else
                    begin
                      reg3696 <= $signed(reg3657[(2'h3):(2'h2)]);
                      reg3697 <= reg3687[(4'hc):(2'h3)];
                      reg3698 <= {$unsigned((reg3647[(4'ha):(4'ha)] <<< forvar3611))};
                    end
                  for (forvar3699 = (1'h0); (forvar3699 < (1'h0)); forvar3699 = (forvar3699 + (1'h1)))
                    begin
                      reg3700 <= {wire3605[(3'h5):(1'h0)]};
                    end
                  for (forvar3701 = (1'h0); (forvar3701 < (1'h0)); forvar3701 = (forvar3701 + (1'h1)))
                    begin
                      reg3702 <= ((({forvar3659} ?
                              reg3652[(4'he):(3'h7)] : reg3649[(3'h5):(3'h4)]) != $unsigned((~^reg3636))) ?
                          $signed((reg3673 ?
                              forvar3663 : forvar3688)) : reg3669);
                      reg3703 <= ($unsigned($unsigned((^~forvar3659))) <= $unsigned(wire3605[(3'h5):(1'h0)]));
                    end
                  for (forvar3704 = (1'h0); (forvar3704 < (1'h1)); forvar3704 = (forvar3704 + (1'h1)))
                    begin
                      reg3705 <= $unsigned($unsigned(reg3678));
                      reg3706 <= (^reg3700[(4'h9):(2'h3)]);
                      reg3707 <= {reg3639};
                      reg3708 <= (8'hb8);
                    end
                end
              reg3709 <= $signed(((^(forvar3688 >>> reg3632)) <= $signed($signed(reg3656))));
              if ((~$unsigned({{reg3647}})))
                begin
                  reg3710 <= $unsigned($signed($signed({reg3623})));
                  for (forvar3711 = (1'h0); (forvar3711 < (2'h3)); forvar3711 = (forvar3711 + (1'h1)))
                    begin
                      reg3712 <= $signed(reg3710[(4'h9):(3'h4)]);
                      reg3713 <= {forvar3689[(3'h7):(1'h1)]};
                      reg3714 <= $unsigned(forvar3688);
                    end
                  if ($unsigned(reg3690[(3'h7):(2'h3)]))
                    begin
                      reg3715 <= (-(reg3634 ?
                          (~|(8'ha7)) : (~^$unsigned(reg3650))));
                      reg3716 <= $signed(reg3637[(4'hf):(2'h2)]);
                      reg3717 <= wire3607[(2'h3):(1'h0)];
                      reg3718 <= {((|(reg3659 ? forvar3634 : reg3623)) ?
                              $unsigned(reg3645) : reg3626[(1'h1):(1'h1)])};
                    end
                  else
                    begin
                      reg3715 <= reg3622;
                      reg3716 <= wire3604[(4'h9):(2'h3)];
                    end
                end
              else
                begin
                  if ($unsigned(wire3609))
                    begin
                      reg3710 <= {$signed(((~&reg3693) ?
                              forvar3648 : (reg3633 != reg3682)))};
                      reg3711 <= $signed(($signed((reg3634 | reg3645)) ?
                          ((reg3707 ? wire3606 : forvar3616) ?
                              reg3700 : $unsigned(reg3621)) : (forvar3711 ^ (^(8'ha7)))));
                    end
                  else
                    begin
                      reg3710 <= (reg3641 ?
                          ($unsigned((^reg3644)) || $unsigned((^(8'had)))) : (forvar3711 ?
                              forvar3668 : (!reg3629[(2'h3):(2'h3)])));
                      reg3711 <= (($unsigned($unsigned(reg3712)) ?
                          ($unsigned(reg3693) ?
                              $signed(reg3615) : reg3632[(1'h1):(1'h0)]) : $unsigned($signed(forvar3695))) < (reg3690[(4'ha):(4'h8)] ?
                          $unsigned((~^reg3669)) : {(~|reg3666)}));
                      reg3712 <= forvar3670[(3'h5):(3'h4)];
                      reg3713 <= (({(reg3630 ? reg3623 : (8'hb3))} ?
                          (~((8'ha0) && (8'hb4))) : (~|$unsigned(wire3606))) <<< $signed($unsigned(reg3660)));
                    end
                  for (forvar3714 = (1'h0); (forvar3714 < (1'h0)); forvar3714 = (forvar3714 + (1'h1)))
                    begin
                      reg3715 <= reg3671;
                    end
                  for (forvar3716 = (1'h0); (forvar3716 < (2'h3)); forvar3716 = (forvar3716 + (1'h1)))
                    begin
                      reg3717 <= ((~|$unsigned((^forvar3678))) ?
                          $signed(($unsigned(reg3669) ?
                              (wire3607 ?
                                  reg3714 : forvar3699) : $unsigned(forvar3688))) : $signed(reg3692[(4'h9):(3'h7)]));
                      reg3718 <= $signed($signed(forvar3670));
                      reg3719 <= (reg3716[(3'h7):(3'h5)] && ({$unsigned(forvar3695)} ?
                          (&$signed(forvar3704)) : $signed({reg3682})));
                    end
                  for (forvar3720 = (1'h0); (forvar3720 < (2'h2)); forvar3720 = (forvar3720 + (1'h1)))
                    begin
                      reg3721 <= (&$unsigned(reg3692));
                      reg3722 <= ((-(8'had)) ?
                          (((forvar3668 == (8'h9f)) >= $unsigned(forvar3659)) & reg3614) : (8'ha1));
                      reg3723 <= $signed(({(|reg3651)} ?
                          forvar3667 : (forvar3688[(1'h1):(1'h0)] << $signed((8'ha8)))));
                      reg3724 <= $signed((((~&(8'hb5)) ?
                              (reg3698 <<< (8'ha3)) : (reg3622 * reg3641)) ?
                          reg3697[(4'h9):(1'h1)] : forvar3616));
                    end
                end
              for (forvar3725 = (1'h0); (forvar3725 < (1'h0)); forvar3725 = (forvar3725 + (1'h1)))
                begin
                  reg3726 <= $unsigned({{$unsigned(reg3649)}});
                end
            end
          for (forvar3727 = (1'h0); (forvar3727 < (2'h3)); forvar3727 = (forvar3727 + (1'h1)))
            begin
              for (forvar3728 = (1'h0); (forvar3728 < (2'h2)); forvar3728 = (forvar3728 + (1'h1)))
                begin
                  if (reg3705)
                    begin
                      reg3729 <= {reg3637[(3'h7):(3'h4)]};
                      reg3730 <= $unsigned((+reg3692[(4'ha):(3'h4)]));
                      reg3731 <= ({$signed((forvar3727 ? reg3626 : reg3645))} ?
                          (^($unsigned(forvar3689) == {forvar3654})) : ((8'haf) != $unsigned((wire3607 != reg3678))));
                    end
                  else
                    begin
                      reg3729 <= reg3685[(1'h0):(1'h0)];
                    end
                  for (forvar3732 = (1'h0); (forvar3732 < (1'h0)); forvar3732 = (forvar3732 + (1'h1)))
                    begin
                      reg3733 <= reg3666;
                      reg3734 <= $signed($unsigned(reg3675));
                      reg3735 <= (reg3626 ?
                          (&($unsigned(wire3606) + (-forvar3654))) : (~($signed(forvar3616) ?
                              $signed(reg3626) : (reg3633 >>> reg3617))));
                      reg3736 <= ((8'haa) < reg3659);
                    end
                  for (forvar3737 = (1'h0); (forvar3737 < (1'h1)); forvar3737 = (forvar3737 + (1'h1)))
                    begin
                      reg3738 <= (~^(wire3607[(4'h9):(3'h6)] ?
                          $signed($unsigned(reg3714)) : {reg3624}));
                      reg3739 <= $signed(forvar3634);
                      reg3740 <= (~^(!$unsigned((&reg3612))));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      reg3741 <= $unsigned({(^~(8'ha6))});
      for (forvar3742 = (1'h0); (forvar3742 < (1'h1)); forvar3742 = (forvar3742 + (1'h1)))
        begin
          if (reg3617)
            begin
              for (forvar3743 = (1'h0); (forvar3743 < (1'h0)); forvar3743 = (forvar3743 + (1'h1)))
                begin
                  if ((8'ha6))
                    begin
                      reg3744 <= ({reg3723} ?
                          $unsigned(forvar3714[(3'h5):(3'h4)]) : reg3622[(1'h1):(1'h1)]);
                      reg3745 <= {{$signed(reg3693)}};
                      reg3746 <= $signed($signed($signed(reg3660[(3'h6):(1'h0)])));
                    end
                  else
                    begin
                      reg3744 <= $unsigned({$unsigned($signed(wire3608))});
                      reg3745 <= reg3653;
                    end
                  if ($unsigned(reg3684[(3'h5):(3'h4)]))
                    begin
                      reg3747 <= $signed($unsigned($signed({(8'hb4)})));
                      reg3748 <= forvar3728;
                      reg3749 <= reg3693[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3747 <= ($unsigned(($signed((8'hb9)) ?
                              (!reg3665) : $signed((8'hb4)))) ?
                          reg3713[(1'h1):(1'h1)] : forvar3732);
                    end
                  for (forvar3750 = (1'h0); (forvar3750 < (1'h0)); forvar3750 = (forvar3750 + (1'h1)))
                    begin
                      reg3751 <= reg3639[(2'h2):(1'h1)];
                      reg3752 <= $unsigned(reg3702);
                      reg3753 <= (forvar3638[(4'ha):(4'h9)] + $signed({(+reg3690)}));
                      reg3754 <= reg3641[(4'hd):(4'h9)];
                    end
                  for (forvar3755 = (1'h0); (forvar3755 < (1'h0)); forvar3755 = (forvar3755 + (1'h1)))
                    begin
                      reg3756 <= $unsigned($unsigned($signed(((8'ha4) ?
                          (8'ha2) : (8'haf)))));
                      reg3757 <= $unsigned((^(~&((8'hb9) ?
                          reg3674 : reg3692))));
                    end
                end
            end
          else
            begin
              for (forvar3743 = (1'h0); (forvar3743 < (1'h1)); forvar3743 = (forvar3743 + (1'h1)))
                begin
                  if ($unsigned(reg3709))
                    begin
                      reg3744 <= {((&(reg3678 ?
                              reg3634 : forvar3663)) < {((8'hab) ?
                                  (8'hb7) : reg3702)})};
                    end
                  else
                    begin
                      reg3744 <= {((~&$signed(reg3628)) < $signed((~(8'hb0))))};
                      reg3745 <= reg3715[(4'hd):(4'hd)];
                      reg3746 <= $unsigned(((8'haf) >= (~^$unsigned(forvar3670))));
                    end
                end
            end
          for (forvar3758 = (1'h0); (forvar3758 < (1'h1)); forvar3758 = (forvar3758 + (1'h1)))
            begin
              for (forvar3759 = (1'h0); (forvar3759 < (2'h2)); forvar3759 = (forvar3759 + (1'h1)))
                begin
                  for (forvar3760 = (1'h0); (forvar3760 < (2'h2)); forvar3760 = (forvar3760 + (1'h1)))
                    begin
                      reg3761 <= (($unsigned(((8'ha9) ?
                              (8'h9f) : reg3629)) || ((forvar3760 ?
                              (8'ha6) : (8'hb8)) == $unsigned((8'hb9)))) ?
                          $signed(((forvar3670 ~^ reg3680) ?
                              $unsigned(reg3741) : {reg3687})) : $unsigned((|(reg3684 ?
                              reg3629 : reg3665))));
                      reg3762 <= {(((reg3617 + reg3678) ^ $signed(wire3607)) * reg3621[(3'h4):(1'h1)])};
                      reg3763 <= (^reg3748);
                      reg3764 <= ($unsigned($unsigned((reg3669 >>> reg3671))) ?
                          ((reg3745 < ((8'haf) ? (8'hb7) : reg3627)) ?
                              $signed((forvar3647 ?
                                  reg3690 : forvar3742)) : $signed($signed(reg3624))) : (~|$signed((&reg3763))));
                    end
                end
              if ((reg3744 ?
                  {$signed(reg3632)} : $signed(((reg3749 ?
                      reg3620 : reg3748) ^ $signed(reg3661)))))
                begin
                  if ($signed(reg3753))
                    begin
                      reg3765 <= reg3666[(1'h1):(1'h1)];
                      reg3766 <= $signed($signed({(~|forvar3704)}));
                    end
                  else
                    begin
                      reg3765 <= forvar3758;
                      reg3766 <= (((reg3745 ?
                          (reg3684 ?
                              reg3716 : reg3630) : reg3729[(3'h5):(2'h2)]) && {(^reg3647)}) ^ (!(forvar3699 ?
                          forvar3720[(3'h4):(2'h3)] : $unsigned((8'ha1)))));
                    end
                  if ($signed(((-reg3639) <= forvar3654)))
                    begin
                      reg3767 <= reg3676[(1'h0):(1'h0)];
                      reg3768 <= reg3705[(1'h1):(1'h1)];
                      reg3769 <= (~((&$signed((8'ha1))) && (-{reg3680})));
                      reg3770 <= $unsigned(reg3751);
                    end
                  else
                    begin
                      reg3767 <= $unsigned($unsigned((-$signed(forvar3714))));
                      reg3768 <= (($unsigned(((8'ha2) ? (8'h9c) : reg3617)) ?
                              ((reg3702 >> (8'ha9)) | (reg3639 > (8'hac))) : ((reg3718 + reg3627) - reg3618[(3'h5):(1'h0)])) ?
                          {wire3605} : ($signed($unsigned(reg3631)) ^ forvar3611));
                      reg3769 <= reg3765[(3'h6):(1'h0)];
                    end
                  if (reg3715[(3'h4):(2'h3)])
                    begin
                      reg3771 <= ($unsigned($unsigned($unsigned((8'hb2)))) >= $signed((!forvar3663[(4'ha):(4'h8)])));
                    end
                  else
                    begin
                      reg3771 <= forvar3714;
                    end
                  if ($signed(forvar3654[(4'h8):(1'h0)]))
                    begin
                      reg3772 <= (|reg3617[(2'h2):(2'h2)]);
                      reg3773 <= $unsigned($unsigned($signed(forvar3720[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg3772 <= (reg3634 ?
                          $signed(($unsigned(reg3731) ^~ (reg3674 || reg3716))) : reg3678[(2'h2):(2'h2)]);
                    end
                end
              else
                begin
                  reg3765 <= reg3700;
                end
              for (forvar3774 = (1'h0); (forvar3774 < (2'h3)); forvar3774 = (forvar3774 + (1'h1)))
                begin
                  reg3775 <= $signed(($signed((~reg3666)) >>> forvar3750[(2'h2):(2'h2)]));
                  for (forvar3776 = (1'h0); (forvar3776 < (1'h0)); forvar3776 = (forvar3776 + (1'h1)))
                    begin
                      reg3777 <= forvar3618[(1'h1):(1'h1)];
                      reg3778 <= ($unsigned((wire3609[(1'h1):(1'h1)] ?
                          forvar3668 : (reg3710 ?
                              reg3773 : reg3733))) >> ($unsigned((-reg3625)) ?
                          forvar3645[(2'h2):(1'h1)] : $signed($signed(reg3715))));
                      reg3779 <= $signed(((~&{reg3762}) >> {$signed(wire3606)}));
                      reg3780 <= $unsigned({(~(reg3696 ? reg3744 : reg3739))});
                    end
                  for (forvar3781 = (1'h0); (forvar3781 < (1'h1)); forvar3781 = (forvar3781 + (1'h1)))
                    begin
                      reg3782 <= reg3684[(2'h3):(1'h1)];
                      reg3783 <= reg3733;
                    end
                end
              if (((reg3698 <<< (|(reg3740 ?
                  forvar3701 : reg3779))) >> $signed({(reg3625 != (8'hb2))})))
                begin
                  reg3784 <= (reg3665[(3'h7):(3'h5)] ?
                      reg3614[(4'hc):(2'h3)] : ((reg3735[(3'h6):(3'h4)] != (forvar3699 + forvar3627)) ?
                          reg3647 : forvar3616));
                  for (forvar3785 = (1'h0); (forvar3785 < (2'h3)); forvar3785 = (forvar3785 + (1'h1)))
                    begin
                      reg3786 <= ((((forvar3688 >> reg3672) <<< forvar3785[(4'h9):(3'h4)]) ?
                          reg3628[(1'h1):(1'h0)] : $signed((reg3629 > reg3733))) << $unsigned((reg3696[(2'h3):(1'h0)] ?
                          forvar3647[(2'h3):(2'h3)] : $unsigned(reg3756))));
                      reg3787 <= reg3719;
                      reg3788 <= wire3605;
                      reg3789 <= $signed($signed((~&(reg3767 ?
                          reg3710 : reg3746))));
                    end
                  reg3790 <= (~&reg3784);
                  if ($signed(reg3698[(1'h1):(1'h0)]))
                    begin
                      reg3791 <= ($signed($signed((reg3643 ~^ (8'ha2)))) ?
                          $unsigned($unsigned((reg3707 >> reg3770))) : $signed(((^~forvar3727) || $unsigned((8'hb4)))));
                      reg3792 <= forvar3640;
                      reg3793 <= forvar3781[(4'h9):(3'h5)];
                      reg3794 <= reg3793[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg3791 <= (-($unsigned((^reg3655)) ?
                          reg3683 : ({reg3659} == (+forvar3688))));
                      reg3792 <= ((|{forvar3695[(3'h7):(3'h5)]}) & $unsigned((~|reg3719)));
                    end
                end
              else
                begin
                  reg3784 <= ((^~(reg3634[(2'h2):(2'h2)] & ((8'hb8) ?
                      reg3731 : forvar3774))) ~^ (reg3696[(1'h1):(1'h0)] & (reg3664[(2'h2):(2'h2)] ?
                      (~&forvar3755) : forvar3647[(3'h6):(3'h6)])));
                  if ((~^($unsigned($unsigned(reg3678)) >= {reg3714[(4'h8):(3'h4)]})))
                    begin
                      reg3785 <= ($unsigned($signed((reg3787 ?
                              wire3606 : reg3747))) ?
                          (reg3613[(3'h6):(2'h3)] ?
                              ($unsigned(reg3770) ?
                                  (reg3751 ?
                                      reg3635 : forvar3645) : (~&(8'ha6))) : $signed($signed((8'hab)))) : $signed($signed(((8'hab) ?
                              reg3648 : reg3731))));
                      reg3786 <= $unsigned((forvar3785[(2'h3):(2'h3)] ?
                          reg3690[(4'ha):(2'h3)] : reg3650));
                      reg3787 <= forvar3668;
                      reg3788 <= reg3714;
                    end
                  else
                    begin
                      reg3785 <= ((&$signed(forvar3699)) >= reg3716);
                      reg3786 <= $signed($unsigned((8'ha1)));
                    end
                end
            end
          reg3795 <= reg3631;
          for (forvar3796 = (1'h0); (forvar3796 < (2'h2)); forvar3796 = (forvar3796 + (1'h1)))
            begin
              for (forvar3797 = (1'h0); (forvar3797 < (1'h0)); forvar3797 = (forvar3797 + (1'h1)))
                begin
                  for (forvar3798 = (1'h0); (forvar3798 < (2'h2)); forvar3798 = (forvar3798 + (1'h1)))
                    begin
                      reg3799 <= (forvar3796 ? reg3679 : reg3751);
                      reg3800 <= (~^$signed($signed(reg3626[(4'hb):(3'h6)])));
                      reg3801 <= $unsigned({$signed($unsigned(reg3752))});
                      reg3802 <= $signed(reg3703[(1'h1):(1'h0)]);
                    end
                  reg3803 <= $unsigned((((^~reg3716) - (reg3660 ^ (8'haa))) == (-reg3676[(2'h2):(1'h0)])));
                end
              for (forvar3804 = (1'h0); (forvar3804 < (2'h3)); forvar3804 = (forvar3804 + (1'h1)))
                begin
                  for (forvar3805 = (1'h0); (forvar3805 < (1'h0)); forvar3805 = (forvar3805 + (1'h1)))
                    begin
                      reg3806 <= (~|{reg3733});
                    end
                end
              for (forvar3807 = (1'h0); (forvar3807 < (1'h0)); forvar3807 = (forvar3807 + (1'h1)))
                begin
                  for (forvar3808 = (1'h0); (forvar3808 < (2'h3)); forvar3808 = (forvar3808 + (1'h1)))
                    begin
                      reg3809 <= ($signed(reg3621[(1'h0):(1'h0)]) * (((reg3719 ?
                                  forvar3804 : reg3638) ?
                              (reg3631 ?
                                  forvar3781 : (8'ha4)) : ((8'ha2) + reg3791)) ?
                          (~(reg3772 + reg3752)) : forvar3688[(3'h6):(2'h3)]));
                    end
                end
              if ($unsigned(forvar3699))
                begin
                  reg3810 <= $unsigned($unsigned(((8'ha9) + {reg3643})));
                  for (forvar3811 = (1'h0); (forvar3811 < (1'h1)); forvar3811 = (forvar3811 + (1'h1)))
                    begin
                      reg3812 <= $signed({(8'hac)});
                      reg3813 <= ($signed(forvar3807[(3'h4):(2'h2)]) ?
                          forvar3759[(1'h1):(1'h1)] : {{$signed(forvar3618)}});
                    end
                end
              else
                begin
                  for (forvar3810 = (1'h0); (forvar3810 < (1'h1)); forvar3810 = (forvar3810 + (1'h1)))
                    begin
                      reg3811 <= $unsigned(((~&{(8'haa)}) ?
                          forvar3647 : (8'ha8)));
                    end
                  for (forvar3812 = (1'h0); (forvar3812 < (2'h2)); forvar3812 = (forvar3812 + (1'h1)))
                    begin
                      reg3813 <= $unsigned($unsigned({(8'hb1)}));
                    end
                  for (forvar3814 = (1'h0); (forvar3814 < (1'h1)); forvar3814 = (forvar3814 + (1'h1)))
                    begin
                      reg3815 <= $unsigned((((forvar3699 ?
                              reg3793 : reg3762) > wire3606) ?
                          reg3696[(3'h7):(3'h4)] : $unsigned(wire3607[(1'h0):(1'h0)])));
                      reg3816 <= (+$signed({(~|forvar3634)}));
                      reg3817 <= (~^((^~$signed(forvar3711)) ^~ $signed((forvar3704 >>> reg3681))));
                      reg3818 <= ((((forvar3742 ? reg3653 : forvar3725) ?
                              wire3609[(1'h1):(1'h0)] : reg3627) ?
                          ($signed(reg3719) ?
                              forvar3622 : (reg3679 ?
                                  (8'hb7) : (8'hb0))) : $signed($signed(wire3604))) * forvar3699[(3'h5):(2'h2)]);
                    end
                end
            end
        end
      for (forvar3819 = (1'h0); (forvar3819 < (1'h0)); forvar3819 = (forvar3819 + (1'h1)))
        begin
          if ((+forvar3807))
            begin
              reg3820 <= ({forvar3670} >>> $unsigned((8'ha0)));
              for (forvar3821 = (1'h0); (forvar3821 < (2'h3)); forvar3821 = (forvar3821 + (1'h1)))
                begin
                  reg3822 <= (~&($signed($signed(reg3649)) << reg3779));
                end
            end
          else
            begin
              for (forvar3820 = (1'h0); (forvar3820 < (1'h0)); forvar3820 = (forvar3820 + (1'h1)))
                begin
                  for (forvar3821 = (1'h0); (forvar3821 < (1'h1)); forvar3821 = (forvar3821 + (1'h1)))
                    begin
                      reg3822 <= (8'ha0);
                    end
                  for (forvar3823 = (1'h0); (forvar3823 < (2'h2)); forvar3823 = (forvar3823 + (1'h1)))
                    begin
                      reg3824 <= reg3664;
                      reg3825 <= (^~{forvar3678[(2'h2):(1'h1)]});
                      reg3826 <= $signed((reg3696 <= (^~$unsigned(forvar3737))));
                      reg3827 <= $signed((8'ha3));
                    end
                end
            end
          reg3828 <= (($signed((forvar3695 == reg3747)) && ((8'h9f) && (~&reg3642))) * (reg3698[(2'h2):(1'h1)] < $signed((forvar3626 < (8'hb9)))));
          for (forvar3829 = (1'h0); (forvar3829 < (2'h3)); forvar3829 = (forvar3829 + (1'h1)))
            begin
              if (($signed({((8'haa) ? reg3676 : (8'hb0))}) ?
                  $signed(reg3678[(4'h9):(2'h2)]) : (((-reg3630) * forvar3694) ~^ ((^reg3799) - $signed(reg3810)))))
                begin
                  if (($unsigned({(reg3736 || (8'ha6))}) ?
                      (~^$unsigned($signed((8'hb9)))) : reg3801))
                    begin
                      reg3830 <= {(reg3816[(3'h6):(3'h6)] ?
                              (&forvar3727) : forvar3808[(2'h2):(1'h1)])};
                      reg3831 <= (reg3801 ?
                          $signed($unsigned($unsigned(reg3775))) : (($signed(reg3638) ?
                                  wire3609[(2'h2):(1'h1)] : reg3772) ?
                              $unsigned(forvar3627[(2'h2):(1'h0)]) : {(reg3795 ^ forvar3804)}));
                      reg3832 <= forvar3701;
                      reg3833 <= $unsigned({reg3749});
                    end
                  else
                    begin
                      reg3830 <= (+$unsigned(($signed(reg3741) << $unsigned(reg3726))));
                      reg3831 <= {($signed(forvar3699[(4'h9):(1'h1)]) ?
                              (^(&reg3617)) : $unsigned(reg3827[(2'h2):(1'h1)]))};
                      reg3832 <= {reg3632[(1'h0):(1'h0)]};
                      reg3833 <= {reg3692[(4'ha):(4'h9)]};
                    end
                  if ($unsigned(reg3717))
                    begin
                      reg3834 <= $signed((8'hb0));
                      reg3835 <= (forvar3667 ?
                          reg3734[(1'h0):(1'h0)] : ((^(forvar3796 && (8'ha1))) ?
                              reg3666[(4'hc):(4'hb)] : (reg3711 ?
                                  (~^reg3711) : (~^forvar3647))));
                      reg3836 <= reg3675;
                      reg3837 <= (($signed(reg3673) ?
                              (!forvar3634) : {(forvar3694 ?
                                      reg3751 : (8'ha2))}) ?
                          reg3647 : $signed($signed($signed(reg3627))));
                    end
                  else
                    begin
                      reg3834 <= $signed((|({(8'hab)} | (&reg3657))));
                      reg3835 <= ((reg3799 ?
                          reg3719[(1'h0):(1'h0)] : (forvar3711[(2'h3):(2'h3)] ?
                              (forvar3807 ?
                                  reg3822 : (8'hb8)) : forvar3798[(4'h9):(4'h9)])) == $signed($unsigned($unsigned(reg3816))));
                      reg3836 <= (!(reg3791[(3'h4):(3'h4)] ?
                          reg3775 : (~&$unsigned(forvar3743))));
                    end
                  if ($signed(($unsigned((~&forvar3760)) ?
                      ((forvar3634 >>> wire3608) << {forvar3640}) : {reg3684})))
                    begin
                      reg3838 <= (forvar3759 & reg3800[(3'h7):(2'h2)]);
                    end
                  else
                    begin
                      reg3838 <= (^~$signed($unsigned($unsigned((8'hb0)))));
                      reg3839 <= {$unsigned($signed($unsigned((8'haf))))};
                    end
                end
              else
                begin
                  if ($unsigned(reg3652[(1'h1):(1'h1)]))
                    begin
                      reg3830 <= $signed((^((reg3625 ?
                          forvar3627 : (8'ha5)) + (+(8'hb0)))));
                      reg3831 <= reg3835[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg3830 <= (($unsigned((8'hb6)) ?
                              $signed(reg3715) : $signed((reg3631 | reg3752))) ?
                          $unsigned((reg3754 || (reg3802 ?
                              reg3792 : reg3650))) : (forvar3720 == {(reg3620 ?
                                  forvar3743 : forvar3759)}));
                      reg3831 <= ((^$unsigned({reg3791})) ^ reg3633);
                      reg3832 <= $signed({$signed((reg3800 ?
                              forvar3616 : (8'hb7)))});
                    end
                end
              for (forvar3840 = (1'h0); (forvar3840 < (1'h0)); forvar3840 = (forvar3840 + (1'h1)))
                begin
                  if (forvar3622[(2'h3):(1'h1)])
                    begin
                      reg3841 <= $unsigned(((8'hb3) ?
                          reg3637 : reg3786[(1'h0):(1'h0)]));
                      reg3842 <= $signed((reg3625[(2'h3):(2'h3)] > $signed({reg3640})));
                      reg3843 <= reg3660;
                    end
                  else
                    begin
                      reg3841 <= {(forvar3616[(4'ha):(3'h7)] ?
                              ($unsigned(reg3660) * (|(8'hb2))) : (forvar3654 >> (forvar3774 != reg3618)))};
                    end
                  for (forvar3844 = (1'h0); (forvar3844 < (2'h2)); forvar3844 = (forvar3844 + (1'h1)))
                    begin
                      reg3845 <= $signed(forvar3796);
                    end
                  if ($unsigned(forvar3640))
                    begin
                      reg3846 <= ((-((~&(8'hac)) ^ (~|reg3645))) != reg3628);
                      reg3847 <= (-(~$unsigned(((8'hae) ? reg3615 : reg3676))));
                      reg3848 <= ((8'hb0) ?
                          (((~|reg3721) && reg3733) ?
                              (forvar3638 ?
                                  reg3669 : ((8'h9e) ?
                                      (8'ha9) : wire3605)) : reg3837) : (^~(reg3627 ?
                              (forvar3820 + reg3778) : (reg3639 ?
                                  reg3723 : reg3735))));
                      reg3849 <= ((($signed((8'ha3)) != (!forvar3688)) ?
                          $signed($signed((8'ha6))) : forvar3647[(3'h6):(2'h3)]) ~^ ((^~reg3775) ?
                          {(forvar3640 < reg3791)} : ((forvar3797 && forvar3829) ?
                              forvar3626[(4'hb):(1'h1)] : $unsigned((8'hb8)))));
                    end
                  else
                    begin
                      reg3846 <= reg3623;
                      reg3847 <= reg3839;
                      reg3848 <= forvar3626;
                      reg3849 <= (^forvar3688[(1'h1):(1'h0)]);
                    end
                end
              if (({(-(reg3680 + reg3792))} >>> $unsigned((forvar3667 ?
                  reg3666 : (-(8'hb9))))))
                begin
                  for (forvar3850 = (1'h0); (forvar3850 < (1'h1)); forvar3850 = (forvar3850 + (1'h1)))
                    begin
                      reg3851 <= (({forvar3728[(1'h1):(1'h0)]} ?
                              $unsigned((~^reg3618)) : (|forvar3797[(2'h2):(1'h1)])) ?
                          $signed(reg3812[(4'h8):(3'h4)]) : ($unsigned((forvar3785 ?
                              forvar3850 : reg3710)) ^~ reg3782[(3'h7):(3'h5)]));
                      reg3852 <= reg3822[(3'h6):(3'h6)];
                      reg3853 <= reg3655[(1'h1):(1'h0)];
                      reg3854 <= forvar3610[(1'h1):(1'h1)];
                    end
                  for (forvar3855 = (1'h0); (forvar3855 < (1'h0)); forvar3855 = (forvar3855 + (1'h1)))
                    begin
                      reg3856 <= (!(~|$unsigned($signed(reg3839))));
                      reg3857 <= {$signed((^~$unsigned((8'h9d))))};
                    end
                  for (forvar3858 = (1'h0); (forvar3858 < (1'h1)); forvar3858 = (forvar3858 + (1'h1)))
                    begin
                      reg3859 <= reg3638[(5'h10):(2'h2)];
                      reg3860 <= ($unsigned(((reg3835 != reg3788) * {reg3769})) * ($unsigned($signed(reg3617)) | $signed((^(8'h9e)))));
                      reg3861 <= $signed((forvar3855 ^ (^~(reg3825 ?
                          (8'ha6) : forvar3699))));
                    end
                  for (forvar3862 = (1'h0); (forvar3862 < (2'h2)); forvar3862 = (forvar3862 + (1'h1)))
                    begin
                      reg3863 <= (|reg3740);
                      reg3864 <= forvar3670[(3'h4):(3'h4)];
                      reg3865 <= reg3713;
                    end
                end
              else
                begin
                  for (forvar3850 = (1'h0); (forvar3850 < (1'h1)); forvar3850 = (forvar3850 + (1'h1)))
                    begin
                      reg3851 <= $unsigned($signed(({(8'hac)} ~^ $signed(reg3740))));
                      reg3852 <= ((reg3786[(1'h1):(1'h0)] ?
                              ((wire3606 | (8'hb8)) ?
                                  reg3749[(3'h4):(3'h4)] : reg3693[(3'h6):(3'h4)]) : (reg3708[(4'hb):(3'h5)] ?
                                  (forvar3648 && (8'h9f)) : reg3665[(2'h2):(2'h2)])) ?
                          reg3731[(3'h5):(1'h1)] : reg3785[(3'h5):(1'h1)]);
                      reg3853 <= (reg3665 ?
                          $unsigned($unsigned(reg3845[(1'h1):(1'h0)])) : reg3659[(4'hf):(4'hd)]);
                    end
                  for (forvar3854 = (1'h0); (forvar3854 < (1'h1)); forvar3854 = (forvar3854 + (1'h1)))
                    begin
                      reg3855 <= reg3643;
                      reg3856 <= $signed((|($unsigned(reg3786) ?
                          ((8'ha1) ^ reg3788) : (reg3780 ?
                              reg3809 : forvar3668))));
                      reg3857 <= {($signed(reg3834[(1'h1):(1'h1)]) <= $unsigned((-reg3863)))};
                    end
                  if ($signed((((reg3813 >= reg3863) - (reg3658 ?
                          reg3612 : reg3834)) ?
                      (reg3706 < forvar3796[(3'h5):(1'h0)]) : forvar3742)))
                    begin
                      reg3858 <= reg3682;
                      reg3859 <= $unsigned((~^($unsigned((8'ha0)) * ((8'hba) ?
                          forvar3820 : forvar3670))));
                      reg3860 <= ((&$signed((reg3707 ? reg3767 : reg3849))) ?
                          (~|$unsigned(reg3724[(4'h8):(3'h7)])) : (((reg3864 ?
                                  reg3691 : reg3749) <= (~&reg3800)) ?
                              reg3859 : reg3673[(3'h6):(1'h1)]));
                      reg3861 <= forvar3618[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg3858 <= (reg3649 ?
                          reg3671 : ($signed(reg3711) ^ $signed(reg3832)));
                      reg3859 <= ($unsigned($unsigned(reg3762)) ^~ $signed((^~forvar3814)));
                    end
                  for (forvar3862 = (1'h0); (forvar3862 < (2'h2)); forvar3862 = (forvar3862 + (1'h1)))
                    begin
                      reg3863 <= {$unsigned((~^reg3736))};
                      reg3864 <= (|{$signed((reg3816 << reg3708))});
                      reg3865 <= ($unsigned((~^$signed(reg3857))) < wire3607[(3'h7):(3'h6)]);
                    end
                end
            end
        end
      if (reg3731[(3'h4):(2'h2)])
        begin
          for (forvar3866 = (1'h0); (forvar3866 < (2'h2)); forvar3866 = (forvar3866 + (1'h1)))
            begin
              for (forvar3867 = (1'h0); (forvar3867 < (1'h1)); forvar3867 = (forvar3867 + (1'h1)))
                begin
                  reg3868 <= $unsigned((~|(reg3630 & ((8'h9d) ?
                      reg3712 : reg3735))));
                  reg3869 <= forvar3622[(1'h0):(1'h0)];
                  for (forvar3870 = (1'h0); (forvar3870 < (1'h1)); forvar3870 = (forvar3870 + (1'h1)))
                    begin
                      reg3871 <= {{{reg3652[(3'h5):(3'h4)]}}};
                    end
                  if ((8'ha2))
                    begin
                      reg3872 <= ((reg3835 != wire3604) ?
                          (-(+reg3647[(4'hd):(4'hd)])) : ($unsigned($signed(forvar3812)) ^ (forvar3634[(1'h1):(1'h0)] ?
                              (~|reg3641) : (reg3673 || forvar3759))));
                    end
                  else
                    begin
                      reg3872 <= ($unsigned(({forvar3704} ?
                              (reg3740 && reg3812) : $unsigned(reg3626))) ?
                          ((^{reg3700}) <<< reg3855[(4'h9):(3'h7)]) : {(~(!(8'hae)))});
                      reg3873 <= forvar3686;
                      reg3874 <= wire3604;
                    end
                end
              for (forvar3875 = (1'h0); (forvar3875 < (1'h1)); forvar3875 = (forvar3875 + (1'h1)))
                begin
                  reg3876 <= (!reg3734[(2'h2):(1'h1)]);
                  reg3877 <= (reg3656[(4'h9):(4'h8)] ?
                      (reg3687 ?
                          ($signed(reg3745) ?
                              $unsigned(reg3770) : {(8'haa)}) : ($signed(reg3629) != (reg3693 ?
                              reg3785 : reg3691))) : (|{(reg3872 ?
                              (8'had) : forvar3711)}));
                end
              for (forvar3878 = (1'h0); (forvar3878 < (2'h3)); forvar3878 = (forvar3878 + (1'h1)))
                begin
                  if ({(!$signed((reg3696 || reg3703)))})
                    begin
                      reg3879 <= forvar3668;
                      reg3880 <= ((((reg3810 + reg3643) | {(8'hb3)}) ?
                              reg3691[(1'h0):(1'h0)] : ($signed(reg3757) || (^~forvar3878))) ?
                          (forvar3844 ?
                              ({forvar3814} ?
                                  $unsigned((8'hb8)) : $signed(reg3752)) : reg3864[(1'h0):(1'h0)]) : $unsigned($unsigned(((8'hba) ?
                              reg3853 : forvar3659))));
                      reg3881 <= forvar3627[(1'h1):(1'h0)];
                      reg3882 <= $unsigned(reg3682);
                    end
                  else
                    begin
                      reg3879 <= ($signed($signed(forvar3858[(4'hf):(3'h6)])) & reg3751);
                      reg3880 <= forvar3610[(1'h1):(1'h0)];
                      reg3881 <= {(8'h9c)};
                    end
                  for (forvar3883 = (1'h0); (forvar3883 < (2'h3)); forvar3883 = (forvar3883 + (1'h1)))
                    begin
                      reg3884 <= $signed(forvar3742[(2'h3):(1'h1)]);
                    end
                end
              if ($unsigned(reg3625[(2'h3):(2'h3)]))
                begin
                  for (forvar3885 = (1'h0); (forvar3885 < (1'h0)); forvar3885 = (forvar3885 + (1'h1)))
                    begin
                      reg3886 <= reg3780;
                      reg3887 <= ((~&($signed(reg3651) ?
                          reg3749[(1'h0):(1'h0)] : (reg3739 > reg3723))) || $unsigned(reg3765));
                      reg3888 <= ($unsigned($signed({reg3702})) ?
                          reg3806[(1'h0):(1'h0)] : $unsigned(reg3749[(4'ha):(2'h2)]));
                    end
                  for (forvar3889 = (1'h0); (forvar3889 < (2'h2)); forvar3889 = (forvar3889 + (1'h1)))
                    begin
                      reg3890 <= $unsigned((reg3801[(1'h1):(1'h0)] ?
                          $signed({reg3656}) : $signed($signed(reg3627))));
                      reg3891 <= {($signed((wire3608 ? forvar3781 : reg3812)) ?
                              ((forvar3694 ^~ reg3633) ?
                                  {reg3747} : reg3745) : (+$signed(forvar3889)))};
                    end
                  if ($signed(forvar3805[(3'h5):(2'h2)]))
                    begin
                      reg3892 <= (reg3669 ?
                          ((&((8'hae) ^~ reg3802)) || reg3852[(3'h4):(1'h0)]) : reg3710[(4'hc):(3'h7)]);
                      reg3893 <= $unsigned($signed(((!(8'h9f)) ?
                          (~^reg3636) : reg3884)));
                      reg3894 <= ($unsigned({(reg3833 + reg3880)}) >> (~(+$unsigned(forvar3808))));
                      reg3895 <= $unsigned($unsigned(reg3831));
                    end
                  else
                    begin
                      reg3892 <= (~^(^((&(8'ha5)) || (reg3810 << reg3891))));
                    end
                end
              else
                begin
                  for (forvar3885 = (1'h0); (forvar3885 < (1'h0)); forvar3885 = (forvar3885 + (1'h1)))
                    begin
                      reg3886 <= reg3872[(1'h0):(1'h0)];
                      reg3887 <= ((^~$unsigned((forvar3737 == reg3621))) ?
                          ((&{reg3748}) ?
                              $unsigned(forvar3728) : {(reg3693 * reg3852)}) : ($unsigned(((8'h9f) * reg3786)) <= reg3680));
                    end
                  if (reg3738)
                    begin
                      reg3888 <= $signed(((~&reg3793[(2'h2):(1'h1)]) >>> ((^~forvar3695) && (8'h9c))));
                      reg3889 <= (+{(~^(~&reg3851))});
                    end
                  else
                    begin
                      reg3888 <= reg3873;
                      reg3889 <= (reg3669 >>> reg3817);
                    end
                end
            end
          reg3896 <= $unsigned((~$signed((-reg3835))));
        end
      else
        begin
          for (forvar3866 = (1'h0); (forvar3866 < (1'h1)); forvar3866 = (forvar3866 + (1'h1)))
            begin
              reg3867 <= ((^~$unsigned(forvar3668[(2'h2):(1'h0)])) ?
                  (($unsigned(reg3806) ?
                      {forvar3814} : $signed(reg3702)) ^~ forvar3885[(1'h0):(1'h0)]) : ($signed((+reg3624)) < ((+reg3612) || reg3882[(3'h6):(3'h4)])));
              reg3868 <= ($unsigned($signed($unsigned(reg3757))) ?
                  reg3795 : (((!forvar3688) ?
                          (forvar3840 | reg3834) : (8'ha8)) ?
                      (^~$signed(forvar3699)) : $unsigned($unsigned(reg3886))));
              if ((-$signed({reg3620[(4'h9):(1'h1)]})))
                begin
                  if ({((-$signed(forvar3805)) && ((^~reg3677) < reg3703[(1'h1):(1'h1)]))})
                    begin
                      reg3869 <= (~&(((reg3855 ?
                              forvar3862 : (8'hb0)) == {reg3873}) ?
                          (8'hb1) : (~^(reg3818 ? reg3799 : forvar3634))));
                      reg3870 <= $unsigned(reg3832);
                      reg3871 <= $unsigned({((+reg3864) ^ {reg3642})});
                    end
                  else
                    begin
                      reg3869 <= $unsigned(((-{reg3641}) ~^ reg3801));
                    end
                end
              else
                begin
                  for (forvar3869 = (1'h0); (forvar3869 < (2'h3)); forvar3869 = (forvar3869 + (1'h1)))
                    begin
                      reg3870 <= (reg3827[(1'h0):(1'h0)] + reg3665);
                    end
                  reg3871 <= reg3830[(3'h5):(3'h4)];
                  if ((forvar3820[(2'h3):(1'h1)] ?
                      $unsigned(((forvar3820 ~^ reg3863) != wire3609[(2'h3):(2'h2)])) : reg3655[(3'h4):(1'h1)]))
                    begin
                      reg3872 <= (forvar3678 ?
                          reg3822[(4'ha):(4'ha)] : $unsigned(((reg3822 ?
                                  reg3806 : (8'ha0)) ?
                              $signed(reg3711) : (8'hb2))));
                      reg3873 <= $unsigned(reg3869[(3'h6):(3'h6)]);
                      reg3874 <= $signed($signed((!$signed(forvar3699))));
                      reg3875 <= (-({((8'ha3) ?
                              reg3770 : (8'hb8))} <= $signed((reg3753 > reg3769))));
                    end
                  else
                    begin
                      reg3872 <= (forvar3867[(4'ha):(2'h3)] <<< reg3757[(4'ha):(1'h1)]);
                      reg3873 <= $signed((($signed(reg3872) + reg3801[(1'h0):(1'h0)]) + {reg3773[(5'h10):(4'hc)]}));
                      reg3874 <= $unsigned(reg3859);
                    end
                  reg3876 <= (~|reg3709[(2'h3):(2'h2)]);
                end
              for (forvar3877 = (1'h0); (forvar3877 < (1'h1)); forvar3877 = (forvar3877 + (1'h1)))
                begin
                  if (reg3726[(1'h0):(1'h0)])
                    begin
                      reg3878 <= ((reg3687[(4'hc):(4'hc)] ?
                              (!(+reg3793)) : reg3656) ?
                          (forvar3808[(3'h6):(2'h3)] >>> (reg3791 <= forvar3850)) : ($unsigned(reg3868) ?
                              reg3655 : {$unsigned(forvar3659)}));
                    end
                  else
                    begin
                      reg3878 <= (-(!($signed(reg3746) ~^ {reg3623})));
                    end
                  if ($unsigned(reg3642[(1'h0):(1'h0)]))
                    begin
                      reg3879 <= reg3891[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg3879 <= reg3733[(3'h7):(3'h6)];
                      reg3880 <= $unsigned($signed({reg3827}));
                      reg3881 <= (reg3803 - $signed((forvar3711 <<< reg3722[(3'h4):(2'h2)])));
                      reg3882 <= $signed((((+forvar3634) ^ $unsigned(reg3716)) <<< $unsigned(reg3864[(1'h0):(1'h0)])));
                    end
                  for (forvar3883 = (1'h0); (forvar3883 < (2'h2)); forvar3883 = (forvar3883 + (1'h1)))
                    begin
                      reg3884 <= (reg3873 ^~ $unsigned($signed($signed(reg3661))));
                      reg3885 <= reg3835;
                    end
                  if (reg3811[(4'h9):(2'h3)])
                    begin
                      reg3886 <= $unsigned($unsigned((^forvar3720)));
                      reg3887 <= forvar3829;
                    end
                  else
                    begin
                      reg3886 <= ({((forvar3750 ?
                                  reg3752 : forvar3634) ^~ $unsigned(reg3764))} ?
                          $signed($signed($unsigned(reg3658))) : forvar3648);
                      reg3887 <= {$unsigned($unsigned((reg3678 + (8'had))))};
                      reg3888 <= ($unsigned(((reg3873 || forvar3670) + (reg3856 << reg3838))) ?
                          ((+(^~reg3868)) == (~^(forvar3627 ?
                              (8'hb8) : reg3627))) : reg3707[(4'h8):(4'h8)]);
                    end
                end
            end
          for (forvar3889 = (1'h0); (forvar3889 < (1'h1)); forvar3889 = (forvar3889 + (1'h1)))
            begin
              if ($unsigned((forvar3644[(2'h3):(1'h1)] ?
                  (~^reg3641) : ({reg3816} ? forvar3858 : (^~(8'ha3))))))
                begin
                  if (reg3765[(1'h1):(1'h1)])
                    begin
                      reg3890 <= (reg3876[(2'h2):(1'h1)] ?
                          $signed(reg3680) : reg3644[(4'h9):(3'h4)]);
                      reg3891 <= forvar3758;
                      reg3892 <= (forvar3867[(3'h4):(1'h1)] ?
                          $signed(($unsigned(reg3692) ?
                              $unsigned((8'hb3)) : (~forvar3807))) : {reg3809});
                    end
                  else
                    begin
                      reg3890 <= ($signed(reg3846) ?
                          (^((reg3831 << forvar3688) ?
                              $unsigned(reg3873) : $unsigned(forvar3670))) : (~(+(&reg3800))));
                      reg3891 <= reg3838;
                      reg3892 <= (reg3834 ?
                          ($signed($unsigned(forvar3678)) ?
                              ((reg3681 ?
                                  (8'hab) : (8'ha4)) <= $unsigned(forvar3737)) : ((reg3890 | (8'hb3)) <= $unsigned(reg3726))) : (~^$unsigned($signed(reg3707))));
                      reg3893 <= ({$signed((reg3700 > reg3715))} - (((8'h9c) ^ (&reg3718)) << (|(|reg3658))));
                    end
                  for (forvar3894 = (1'h0); (forvar3894 < (1'h0)); forvar3894 = (forvar3894 + (1'h1)))
                    begin
                      reg3895 <= ($unsigned(forvar3638[(2'h2):(2'h2)]) ?
                          (&{(~&reg3864)}) : ({reg3730} - reg3756));
                      reg3896 <= reg3614[(2'h3):(1'h0)];
                      reg3897 <= {$unsigned($signed(forvar3804[(3'h4):(1'h1)]))};
                      reg3898 <= $signed((~reg3836[(4'hb):(1'h1)]));
                    end
                end
              else
                begin
                  reg3890 <= (-{{forvar3654}});
                  reg3891 <= wire3606[(4'ha):(4'h9)];
                  for (forvar3892 = (1'h0); (forvar3892 < (1'h0)); forvar3892 = (forvar3892 + (1'h1)))
                    begin
                      reg3893 <= (reg3780[(4'ha):(1'h0)] ?
                          $unsigned(($signed(reg3718) ?
                              (forvar3648 ?
                                  forvar3798 : forvar3869) : {reg3754})) : ((-(8'hb2)) >>> ($unsigned(forvar3642) < (reg3638 != reg3842))));
                      reg3894 <= forvar3688[(2'h2):(1'h1)];
                    end
                end
              if ((~|reg3892[(2'h3):(1'h1)]))
                begin
                  reg3899 <= reg3838[(3'h7):(3'h4)];
                end
              else
                begin
                  for (forvar3899 = (1'h0); (forvar3899 < (2'h2)); forvar3899 = (forvar3899 + (1'h1)))
                    begin
                      reg3900 <= (reg3800 && {forvar3610});
                      reg3901 <= $signed(((~|$unsigned((8'ha5))) ?
                          wire3607[(1'h0):(1'h0)] : $signed($unsigned(forvar3694))));
                      reg3902 <= $unsigned(reg3612[(4'h8):(3'h7)]);
                      reg3903 <= ($signed($unsigned({reg3712})) ?
                          $unsigned($unsigned((~|reg3665))) : $signed($unsigned(reg3747)));
                    end
                  for (forvar3904 = (1'h0); (forvar3904 < (1'h1)); forvar3904 = (forvar3904 + (1'h1)))
                    begin
                      reg3905 <= (reg3879 ?
                          forvar3622 : ({forvar3760[(2'h2):(2'h2)]} ?
                              $unsigned(reg3651[(4'hf):(1'h1)]) : $signed((reg3843 ?
                                  forvar3875 : (8'hb7)))));
                      reg3906 <= reg3735;
                      reg3907 <= {$unsigned((reg3905[(4'h9):(1'h0)] ?
                              forvar3688 : forvar3634[(3'h7):(3'h4)]))};
                      reg3908 <= $signed((~|(~reg3879)));
                    end
                  for (forvar3909 = (1'h0); (forvar3909 < (2'h2)); forvar3909 = (forvar3909 + (1'h1)))
                    begin
                      reg3910 <= $unsigned((reg3856[(3'h4):(2'h3)] ?
                          reg3894 : $unsigned($unsigned(forvar3616))));
                      reg3911 <= (+(reg3899 ?
                          (+(forvar3611 >> reg3896)) : reg3713));
                      reg3912 <= forvar3878;
                      reg3913 <= forvar3737;
                    end
                end
            end
          if ($unsigned(reg3835[(3'h5):(2'h3)]))
            begin
              if ($unsigned($unsigned(reg3693)))
                begin
                  for (forvar3914 = (1'h0); (forvar3914 < (1'h1)); forvar3914 = (forvar3914 + (1'h1)))
                    begin
                      reg3915 <= $unsigned(reg3665[(1'h0):(1'h0)]);
                      reg3916 <= $signed((($signed(reg3753) >> reg3729[(4'hc):(4'h8)]) || (~forvar3688)));
                      reg3917 <= $unsigned($unsigned($unsigned(forvar3695[(2'h2):(1'h1)])));
                      reg3918 <= ($signed({$signed(reg3885)}) ?
                          ({{reg3895}} > {{forvar3701}}) : ((8'h9d) ?
                              {forvar3805} : $unsigned($unsigned(reg3880))));
                    end
                  if (forvar3728[(3'h4):(3'h4)])
                    begin
                      reg3919 <= $unsigned($unsigned({forvar3878[(2'h3):(1'h0)]}));
                    end
                  else
                    begin
                      reg3919 <= ($unsigned({reg3745}) != forvar3909);
                      reg3920 <= forvar3759[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar3914 = (1'h0); (forvar3914 < (1'h0)); forvar3914 = (forvar3914 + (1'h1)))
                    begin
                      reg3915 <= forvar3867[(3'h5):(1'h1)];
                      reg3916 <= $unsigned({((forvar3634 ? reg3849 : (8'h9d)) ?
                              $signed(reg3620) : (~&reg3865))});
                      reg3917 <= (~^$signed(({reg3614} ?
                          $unsigned((8'hab)) : (reg3753 <= reg3865))));
                    end
                  reg3918 <= (+{reg3700[(2'h3):(2'h2)]});
                  reg3919 <= $unsigned((reg3747 & (~&$unsigned(forvar3737))));
                end
            end
          else
            begin
              for (forvar3914 = (1'h0); (forvar3914 < (1'h0)); forvar3914 = (forvar3914 + (1'h1)))
                begin
                  for (forvar3915 = (1'h0); (forvar3915 < (2'h3)); forvar3915 = (forvar3915 + (1'h1)))
                    begin
                      reg3916 <= $signed((((~reg3815) ?
                              ((8'ha9) | forvar3883) : (reg3771 ?
                                  forvar3909 : reg3788)) ?
                          $unsigned(reg3912[(1'h1):(1'h0)]) : $unsigned((8'hae))));
                      reg3917 <= (((!$signed((8'ha9))) ?
                              $signed($signed(forvar3611)) : ($unsigned(reg3635) ?
                                  $unsigned(reg3620) : $signed(forvar3742))) ?
                          $signed((&forvar3855[(3'h5):(1'h0)])) : $signed((~$signed(reg3633))));
                      reg3918 <= reg3768;
                    end
                end
              for (forvar3919 = (1'h0); (forvar3919 < (1'h1)); forvar3919 = (forvar3919 + (1'h1)))
                begin
                  for (forvar3920 = (1'h0); (forvar3920 < (2'h2)); forvar3920 = (forvar3920 + (1'h1)))
                    begin
                      reg3921 <= ((reg3787[(2'h3):(2'h3)] ?
                          (~$unsigned(forvar3686)) : $signed($signed(forvar3840))) >= {$unsigned(forvar3885)});
                      reg3922 <= (+(-$unsigned(reg3711[(2'h3):(2'h3)])));
                    end
                  for (forvar3923 = (1'h0); (forvar3923 < (2'h2)); forvar3923 = (forvar3923 + (1'h1)))
                    begin
                      reg3924 <= (forvar3855 && $signed((-{(8'hac)})));
                      reg3925 <= (forvar3870[(2'h2):(1'h1)] >= (forvar3750[(1'h1):(1'h0)] ?
                          forvar3866[(1'h0):(1'h0)] : $unsigned((reg3621 ?
                              forvar3622 : reg3792))));
                    end
                end
              for (forvar3926 = (1'h0); (forvar3926 < (1'h0)); forvar3926 = (forvar3926 + (1'h1)))
                begin
                  reg3927 <= reg3816[(5'h10):(5'h10)];
                  for (forvar3928 = (1'h0); (forvar3928 < (1'h0)); forvar3928 = (forvar3928 + (1'h1)))
                    begin
                      reg3929 <= (reg3885[(2'h2):(1'h0)] <<< (reg3748 <= ($signed(forvar3699) != reg3658)));
                    end
                  for (forvar3930 = (1'h0); (forvar3930 < (2'h2)); forvar3930 = (forvar3930 + (1'h1)))
                    begin
                      reg3931 <= ((^~(forvar3659[(3'h7):(3'h4)] + reg3851[(3'h4):(1'h0)])) || reg3815[(4'hc):(3'h5)]);
                      reg3932 <= reg3818[(3'h4):(3'h4)];
                      reg3933 <= ((reg3856 ?
                          $unsigned($unsigned((8'h9e))) : ((reg3918 ?
                                  (8'ha5) : reg3625) ?
                              reg3873[(2'h2):(1'h0)] : (&reg3783))) <<< ((~|(reg3801 ?
                              reg3836 : reg3646)) ?
                          ((reg3693 && reg3656) ?
                              ((8'hab) ?
                                  reg3640 : reg3872) : forvar3688[(2'h3):(1'h1)]) : reg3632[(2'h2):(1'h0)]));
                      reg3934 <= $signed((($unsigned(reg3629) == (~^reg3775)) ?
                          ((&forvar3611) ?
                              reg3782[(1'h0):(1'h0)] : $signed((8'h9d))) : (forvar3727 ?
                              $signed(forvar3870) : (8'ha0))));
                    end
                end
            end
          for (forvar3935 = (1'h0); (forvar3935 < (1'h0)); forvar3935 = (forvar3935 + (1'h1)))
            begin
              for (forvar3936 = (1'h0); (forvar3936 < (1'h0)); forvar3936 = (forvar3936 + (1'h1)))
                begin
                  reg3937 <= ((reg3719[(1'h0):(1'h0)] * reg3867[(4'h9):(2'h3)]) ?
                      reg3788 : $unsigned((^(+reg3852))));
                  for (forvar3938 = (1'h0); (forvar3938 < (1'h0)); forvar3938 = (forvar3938 + (1'h1)))
                    begin
                      reg3939 <= (reg3724 || reg3849);
                      reg3940 <= $signed((reg3848 ?
                          $signed($signed(reg3729)) : reg3741));
                    end
                  if ((((!$unsigned(reg3636)) ?
                      $unsigned(reg3718) : (+(reg3785 ?
                          (8'hab) : reg3656))) <<< reg3705))
                    begin
                      reg3941 <= $unsigned($signed($signed((|reg3630))));
                      reg3942 <= {(^~((&reg3902) >>> reg3633))};
                    end
                  else
                    begin
                      reg3941 <= (^~((+(~forvar3814)) ?
                          forvar3716 : (~(forvar3899 ? reg3853 : reg3822))));
                    end
                end
              reg3943 <= (|$signed(reg3757[(4'h9):(2'h2)]));
              for (forvar3944 = (1'h0); (forvar3944 < (1'h0)); forvar3944 = (forvar3944 + (1'h1)))
                begin
                  for (forvar3945 = (1'h0); (forvar3945 < (1'h1)); forvar3945 = (forvar3945 + (1'h1)))
                    begin
                      reg3946 <= ((|$unsigned({reg3896})) ?
                          (~&$signed(reg3726[(3'h5):(3'h4)])) : ($signed(reg3739) - $signed((reg3671 << reg3838))));
                      reg3947 <= {($signed($signed(reg3856)) ?
                              $unsigned(reg3810) : {((8'haf) ?
                                      forvar3701 : forvar3877)})};
                    end
                  for (forvar3948 = (1'h0); (forvar3948 < (2'h3)); forvar3948 = (forvar3948 + (1'h1)))
                    begin
                      reg3949 <= $signed(forvar3919);
                      reg3950 <= {{(reg3690 >>> wire3605)}};
                    end
                end
              for (forvar3951 = (1'h0); (forvar3951 < (2'h2)); forvar3951 = (forvar3951 + (1'h1)))
                begin
                  if (reg3922)
                    begin
                      reg3952 <= reg3692[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg3952 <= (&((^~reg3941) ^ reg3751[(2'h3):(2'h3)]));
                      reg3953 <= $unsigned((~^(^(forvar3760 ^ reg3841))));
                    end
                  for (forvar3954 = (1'h0); (forvar3954 < (1'h0)); forvar3954 = (forvar3954 + (1'h1)))
                    begin
                      reg3955 <= reg3792[(2'h3):(1'h1)];
                    end
                  for (forvar3956 = (1'h0); (forvar3956 < (2'h3)); forvar3956 = (forvar3956 + (1'h1)))
                    begin
                      reg3957 <= $unsigned(reg3855[(4'h9):(3'h4)]);
                      reg3958 <= $unsigned(reg3865);
                      reg3959 <= (($signed($signed(reg3873)) ?
                          reg3950 : reg3621[(2'h3):(1'h1)]) << $signed($unsigned($signed(reg3828))));
                      reg3960 <= (-($unsigned(((8'ha0) - reg3644)) != (|(reg3626 ?
                          reg3890 : forvar3667))));
                    end
                end
            end
        end
    end
  assign wire3961 = ($unsigned((^~reg3940)) - (($unsigned(reg3878) ?
                            (!reg3719) : (reg3911 ? reg3754 : reg3794)) ?
                        forvar3728 : $signed(reg3959[(1'h0):(1'h0)])));
  assign wire3962 = (($unsigned((reg3642 == reg3722)) ^ forvar3954) ?
                        reg3723[(2'h3):(2'h2)] : (~|$unsigned(reg3733[(4'hf):(4'he)])));
  always
    @(posedge clk) begin
      if ((+$signed($unsigned((~|forvar3936)))))
        begin
          if (($unsigned(reg3915[(3'h7):(2'h3)]) ?
              ($unsigned($unsigned((8'hb8))) >= (forvar3855[(2'h3):(1'h0)] >>> {reg3878})) : ((^$signed(reg3893)) & $signed({reg3729}))))
            begin
              if ((($unsigned(forvar3935) >= (-(reg3733 ? reg3693 : (8'hb5)))) ?
                  ($unsigned(reg3960[(1'h1):(1'h0)]) ^ forvar3678[(1'h0):(1'h0)]) : ((&reg3793[(3'h5):(1'h1)]) << $signed({reg3631}))))
                begin
                  for (forvar3963 = (1'h0); (forvar3963 < (1'h1)); forvar3963 = (forvar3963 + (1'h1)))
                    begin
                      reg3964 <= ((reg3841 ?
                          forvar3866[(1'h1):(1'h0)] : $unsigned((forvar3923 >> (8'ha2)))) >>> $unsigned(reg3952[(3'h4):(2'h3)]));
                      reg3965 <= {$unsigned(((~|forvar3870) ?
                              {forvar3774} : reg3767))};
                    end
                  for (forvar3966 = (1'h0); (forvar3966 < (1'h1)); forvar3966 = (forvar3966 + (1'h1)))
                    begin
                      reg3967 <= reg3769[(4'hc):(3'h6)];
                      reg3968 <= ((|reg3630[(4'h9):(1'h0)]) ?
                          {$unsigned((~|reg3784))} : ((reg3726 ?
                              $unsigned(forvar3699) : (reg3687 ?
                                  reg3625 : forvar3616)) || ($unsigned(reg3892) ?
                              (reg3683 && reg3784) : (forvar3701 ?
                                  reg3780 : reg3624))));
                      reg3969 <= $unsigned((($unsigned(reg3848) ~^ reg3910[(4'h8):(2'h3)]) == forvar3956[(3'h6):(3'h4)]));
                    end
                  for (forvar3970 = (1'h0); (forvar3970 < (1'h1)); forvar3970 = (forvar3970 + (1'h1)))
                    begin
                      reg3971 <= (($unsigned($signed(reg3790)) & reg3888[(1'h0):(1'h0)]) ?
                          forvar3923[(1'h0):(1'h0)] : (($unsigned(reg3710) ^ reg3634[(4'hb):(4'h8)]) ?
                              ((forvar3797 + reg3847) ?
                                  $unsigned(reg3669) : (reg3644 ?
                                      (8'hb8) : reg3946)) : reg3846[(1'h1):(1'h1)]));
                      reg3972 <= $unsigned((8'ha5));
                      reg3973 <= $unsigned($unsigned(reg3752[(1'h0):(1'h0)]));
                    end
                  for (forvar3974 = (1'h0); (forvar3974 < (1'h0)); forvar3974 = (forvar3974 + (1'h1)))
                    begin
                      reg3975 <= reg3706;
                    end
                end
              else
                begin
                  if (reg3631[(2'h3):(1'h0)])
                    begin
                      reg3963 <= reg3855[(1'h1):(1'h1)];
                      reg3964 <= $unsigned($unsigned((forvar3611[(3'h7):(2'h2)] || reg3630)));
                    end
                  else
                    begin
                      reg3963 <= $signed({forvar3854});
                      reg3964 <= (reg3833 + reg3789[(1'h0):(1'h0)]);
                      reg3965 <= (8'ha5);
                    end
                end
              if (reg3871[(3'h6):(1'h1)])
                begin
                  if ($signed((^~$signed(reg3632))))
                    begin
                      reg3976 <= reg3738;
                      reg3977 <= (-($unsigned(reg3705) ^ ((forvar3742 ?
                          (8'ha3) : forvar3634) ^ reg3820[(3'h7):(1'h1)])));
                      reg3978 <= reg3964[(3'h4):(1'h0)];
                      reg3979 <= (8'hb9);
                    end
                  else
                    begin
                      reg3976 <= reg3718[(2'h2):(1'h1)];
                      reg3977 <= {$unsigned($signed(reg3665[(2'h2):(2'h2)]))};
                    end
                  if ($signed((~&$signed($signed(reg3863)))))
                    begin
                      reg3980 <= ((+reg3769[(3'h4):(1'h1)]) ?
                          $signed((+(+reg3817))) : $unsigned($unsigned(reg3957[(1'h1):(1'h1)])));
                      reg3981 <= reg3773;
                      reg3982 <= {(|$signed((reg3870 ? reg3903 : (8'ha2))))};
                    end
                  else
                    begin
                      reg3980 <= reg3714[(4'h9):(3'h4)];
                      reg3981 <= (|(^~$unsigned($signed((8'hab)))));
                      reg3982 <= reg3901;
                      reg3983 <= $unsigned((((reg3809 ? reg3953 : (8'hb5)) ?
                          ((8'hb4) ?
                              forvar3645 : (8'h9c)) : (8'hb3)) ~^ reg3722[(3'h5):(1'h0)]));
                    end
                  for (forvar3984 = (1'h0); (forvar3984 < (2'h2)); forvar3984 = (forvar3984 + (1'h1)))
                    begin
                      reg3985 <= forvar3935[(4'hf):(2'h2)];
                    end
                  for (forvar3986 = (1'h0); (forvar3986 < (1'h0)); forvar3986 = (forvar3986 + (1'h1)))
                    begin
                      reg3987 <= wire3962[(2'h2):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar3976 = (1'h0); (forvar3976 < (1'h1)); forvar3976 = (forvar3976 + (1'h1)))
                    begin
                      reg3977 <= $unsigned($unsigned(reg3898[(4'h9):(1'h1)]));
                      reg3978 <= ((~&$unsigned({reg3978})) * reg3794);
                    end
                  reg3979 <= $unsigned({((forvar3695 ? forvar3855 : reg3690) ?
                          (forvar3814 ?
                              (8'hb9) : forvar3805) : $unsigned(reg3625))});
                  for (forvar3980 = (1'h0); (forvar3980 < (1'h1)); forvar3980 = (forvar3980 + (1'h1)))
                    begin
                      reg3981 <= {((reg3893[(2'h3):(2'h3)] ?
                                  (reg3784 ?
                                      forvar3956 : (8'hac)) : (^(8'hb0))) ?
                              {((8'ha7) ?
                                      reg3708 : forvar3808)} : ($signed(reg3841) && (^reg3978)))};
                      reg3982 <= reg3847;
                      reg3983 <= forvar3920;
                      reg3984 <= ((^$signed((~reg3825))) < ($signed((~&forvar3963)) < ($signed(reg3717) >= (^(8'ha5)))));
                    end
                end
            end
          else
            begin
              for (forvar3963 = (1'h0); (forvar3963 < (1'h0)); forvar3963 = (forvar3963 + (1'h1)))
                begin
                  for (forvar3964 = (1'h0); (forvar3964 < (2'h3)); forvar3964 = (forvar3964 + (1'h1)))
                    begin
                      reg3965 <= {$signed(((reg3703 ^~ reg3771) ?
                              reg3900 : reg3724))};
                      reg3966 <= ((~forvar3877) ?
                          (8'hae) : (reg3943 || reg3888[(1'h0):(1'h0)]));
                      reg3967 <= reg3845;
                      reg3968 <= (forvar3743 ?
                          (((reg3782 > reg3751) ^ (reg3739 && reg3910)) ?
                              (~^$signed(forvar3704)) : {reg3761}) : $signed($signed((8'ha7))));
                    end
                end
              for (forvar3969 = (1'h0); (forvar3969 < (1'h1)); forvar3969 = (forvar3969 + (1'h1)))
                begin
                  reg3970 <= reg3752[(1'h1):(1'h1)];
                  reg3971 <= forvar3711[(2'h3):(2'h2)];
                end
            end
          for (forvar3988 = (1'h0); (forvar3988 < (1'h0)); forvar3988 = (forvar3988 + (1'h1)))
            begin
              reg3989 <= reg3888;
              if ($signed((reg3848 ?
                  forvar3951[(4'h8):(2'h3)] : (reg3643 >> {reg3884}))))
                begin
                  for (forvar3990 = (1'h0); (forvar3990 < (1'h0)); forvar3990 = (forvar3990 + (1'h1)))
                    begin
                      reg3991 <= {reg3964[(2'h2):(1'h1)]};
                      reg3992 <= $signed((|($unsigned(forvar3899) | (8'hb9))));
                      reg3993 <= $signed(forvar3694[(4'h9):(2'h2)]);
                      reg3994 <= ((-$unsigned((~&(8'hae)))) ?
                          $unsigned(reg3981) : reg3772[(4'hb):(2'h2)]);
                    end
                end
              else
                begin
                  reg3990 <= {$unsigned((forvar3796 >= ((8'haf) ?
                          reg3677 : reg3771)))};
                  if ((~$unsigned(reg3745[(2'h2):(1'h1)])))
                    begin
                      reg3991 <= (&forvar3808[(3'h5):(1'h1)]);
                    end
                  else
                    begin
                      reg3991 <= reg3615[(2'h3):(2'h3)];
                      reg3992 <= ((reg3761 > (forvar3727[(2'h3):(2'h3)] <<< (reg3717 > (8'hba)))) ?
                          (($signed(reg3851) * (reg3872 <<< reg3958)) <= $unsigned($signed(reg3941))) : $signed({(reg3884 >= (8'hac))}));
                      reg3993 <= reg3640;
                    end
                  if (reg3685[(1'h0):(1'h0)])
                    begin
                      reg3994 <= (~&($unsigned($signed((8'ha3))) <<< ((~^reg3775) ^ (~reg3979))));
                      reg3995 <= reg3868[(3'h7):(1'h0)];
                      reg3996 <= (^forvar3948[(2'h2):(1'h0)]);
                      reg3997 <= reg3877[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3994 <= (reg3771[(2'h3):(1'h1)] || $unsigned($signed($signed(reg3925))));
                    end
                end
              for (forvar3998 = (1'h0); (forvar3998 < (2'h3)); forvar3998 = (forvar3998 + (1'h1)))
                begin
                  for (forvar3999 = (1'h0); (forvar3999 < (2'h2)); forvar3999 = (forvar3999 + (1'h1)))
                    begin
                      reg4000 <= $unsigned((^(|$unsigned(reg3965))));
                      reg4001 <= (-$unsigned(({reg3803} ?
                          reg3977[(1'h0):(1'h0)] : reg3919)));
                      reg4002 <= ($unsigned(reg3647[(4'hf):(2'h3)]) << {$unsigned($signed((8'hb8)))});
                      reg4003 <= $unsigned({(~^reg3752)});
                    end
                  for (forvar4004 = (1'h0); (forvar4004 < (1'h0)); forvar4004 = (forvar4004 + (1'h1)))
                    begin
                      reg4005 <= ($signed((&reg3786)) ?
                          (forvar3670[(3'h5):(1'h0)] & reg3711[(1'h1):(1'h1)]) : (~$signed($signed(reg3978))));
                      reg4006 <= {{(reg3768[(4'hb):(4'ha)] <= (reg3984 ?
                                  (8'had) : reg3924))}};
                      reg4007 <= forvar3969[(3'h4):(2'h2)];
                    end
                  reg4008 <= (~^(8'ha3));
                  for (forvar4009 = (1'h0); (forvar4009 < (2'h2)); forvar4009 = (forvar4009 + (1'h1)))
                    begin
                      reg4010 <= $signed(forvar3954);
                      reg4011 <= $signed($unsigned($unsigned({reg3910})));
                      reg4012 <= (reg3619[(1'h1):(1'h0)] | $signed((8'ha8)));
                      reg4013 <= $unsigned(reg3959);
                    end
                end
            end
        end
      else
        begin
          for (forvar3963 = (1'h0); (forvar3963 < (2'h2)); forvar3963 = (forvar3963 + (1'h1)))
            begin
              if (reg3649)
                begin
                  if (($signed($signed(reg3659[(4'h9):(1'h0)])) ?
                      reg3786 : $signed(forvar3743[(1'h0):(1'h0)])))
                    begin
                      reg3964 <= $unsigned(reg3882);
                      reg3965 <= {$unsigned($signed(reg4005))};
                    end
                  else
                    begin
                      reg3964 <= ($unsigned($unsigned($unsigned(forvar3823))) - $signed(reg3627[(1'h0):(1'h0)]));
                    end
                  for (forvar3966 = (1'h0); (forvar3966 < (1'h0)); forvar3966 = (forvar3966 + (1'h1)))
                    begin
                      reg3967 <= reg3816;
                      reg3968 <= {(reg3656 >>> forvar3805[(4'he):(4'h8)])};
                      reg3969 <= ((((+reg3749) ^ {reg3680}) ?
                              ($signed(reg3673) >= reg3765[(3'h4):(2'h3)]) : ((reg3615 <<< reg3678) ?
                                  (reg3708 && forvar3878) : reg3651)) ?
                          (+(~&$signed(reg3918))) : (~|($unsigned(forvar3980) ?
                              reg3726 : reg3993)));
                      reg3970 <= forvar3892;
                    end
                end
              else
                begin
                  if (((reg3931 ?
                          (|$unsigned(forvar3678)) : ((+reg3731) ?
                              reg3920 : $signed(reg3624))) ?
                      (~^($signed(reg3987) & reg4003[(4'h8):(2'h3)])) : $unsigned(reg3846)))
                    begin
                      reg3964 <= $signed({(reg3861 >> $signed(reg3918))});
                      reg3965 <= forvar3820[(4'h9):(3'h6)];
                    end
                  else
                    begin
                      reg3964 <= reg3795[(3'h6):(3'h4)];
                    end
                  for (forvar3966 = (1'h0); (forvar3966 < (2'h2)); forvar3966 = (forvar3966 + (1'h1)))
                    begin
                      reg3967 <= (~^((forvar3889 ?
                          {forvar3951} : (forvar3695 ?
                              reg3790 : (8'hb6))) - $signed({reg3791})));
                      reg3968 <= $signed($signed(reg3649));
                      reg3969 <= {$signed({(reg3882 ? wire3962 : (8'hab))})};
                      reg3970 <= reg3997;
                    end
                  for (forvar3971 = (1'h0); (forvar3971 < (2'h2)); forvar3971 = (forvar3971 + (1'h1)))
                    begin
                      reg3972 <= (reg4003[(2'h2):(1'h1)] ?
                          forvar3701[(1'h0):(1'h0)] : forvar3862[(3'h4):(2'h3)]);
                      reg3973 <= $unsigned($signed({(forvar3935 ?
                              reg3669 : reg3982)}));
                      reg3974 <= (reg3994[(4'hd):(4'h9)] ?
                          (reg3751[(1'h1):(1'h0)] - ((forvar3704 + reg3832) >= {forvar3894})) : ((((8'hb7) ?
                                  reg3973 : forvar3648) ?
                              $signed(reg3772) : $unsigned((8'haf))) || $signed({reg3893})));
                    end
                end
              for (forvar3975 = (1'h0); (forvar3975 < (1'h1)); forvar3975 = (forvar3975 + (1'h1)))
                begin
                  if ((((forvar3807 && reg3683) + ((reg3612 > reg3801) >= reg3976)) || $signed({{(8'hac)}})))
                    begin
                      reg3976 <= ($signed((reg3820[(2'h3):(2'h2)] ?
                              ((8'ha2) ?
                                  (8'ha8) : (8'h9e)) : $signed(reg3963))) ?
                          reg3685 : reg3678[(2'h2):(1'h0)]);
                      reg3977 <= reg3646;
                      reg3978 <= reg3716;
                      reg3979 <= $unsigned((^~(~|(reg3637 <= reg3846))));
                    end
                  else
                    begin
                      reg3976 <= {(($unsigned(reg3643) << (reg3800 & forvar3986)) << $signed($unsigned(forvar3711)))};
                      reg3977 <= (~&((&$signed(reg3894)) ?
                          $unsigned($signed(reg4003)) : (reg3979 <<< {(8'hab)})));
                    end
                end
              for (forvar3980 = (1'h0); (forvar3980 < (1'h0)); forvar3980 = (forvar3980 + (1'h1)))
                begin
                  for (forvar3981 = (1'h0); (forvar3981 < (2'h3)); forvar3981 = (forvar3981 + (1'h1)))
                    begin
                      reg3982 <= {$unsigned({(forvar3945 <<< forvar3878)})};
                      reg3983 <= ((((reg3723 & (8'haf)) >>> (reg3614 ?
                              reg3816 : forvar3798)) * forvar3875[(4'h8):(3'h6)]) ?
                          $signed($signed((reg3662 ?
                              reg3757 : (8'hac)))) : {forvar3948});
                      reg3984 <= $unsigned(reg3974);
                      reg3985 <= ((-({reg3786} > (~forvar3909))) ?
                          $unsigned((+{forvar3858})) : $unsigned((~&{reg3697})));
                    end
                  reg3986 <= {$signed($unsigned((forvar3999 ?
                          reg3648 : reg3679)))};
                  if ((reg3678[(4'h9):(3'h5)] << (&(8'hb3))))
                    begin
                      reg3987 <= ((~&reg3922[(2'h3):(1'h1)]) ?
                          $unsigned(($signed(reg3651) <<< reg3990[(2'h2):(2'h2)])) : ((+(forvar3755 ?
                                  forvar3964 : reg3903)) ?
                              reg3783 : $signed((^~reg3693))));
                    end
                  else
                    begin
                      reg3987 <= reg3666[(4'ha):(4'h8)];
                      reg3988 <= (reg3713[(3'h4):(3'h4)] - {{$signed(reg3783)}});
                    end
                  for (forvar3989 = (1'h0); (forvar3989 < (2'h3)); forvar3989 = (forvar3989 + (1'h1)))
                    begin
                      reg3990 <= forvar3850;
                      reg3991 <= (~&$unsigned({$unsigned(reg3715)}));
                      reg3992 <= ($signed((forvar3670 > reg3965[(4'h8):(3'h5)])) ?
                          reg3624 : $unsigned({(~^reg3614)}));
                    end
                end
              if (reg3779)
                begin
                  for (forvar3993 = (1'h0); (forvar3993 < (1'h0)); forvar3993 = (forvar3993 + (1'h1)))
                    begin
                      reg3994 <= {($unsigned((^reg3761)) ?
                              $signed(reg3889[(3'h7):(2'h2)]) : $unsigned(reg3775))};
                      reg3995 <= {reg3900};
                      reg3996 <= {$unsigned(reg3721)};
                    end
                end
              else
                begin
                  for (forvar3993 = (1'h0); (forvar3993 < (2'h2)); forvar3993 = (forvar3993 + (1'h1)))
                    begin
                      reg3994 <= (reg3888 << reg4011[(4'hb):(4'h8)]);
                      reg3995 <= (((^~(reg3853 < (8'hb1))) ?
                          (wire3962 * (8'ha4)) : $unsigned($unsigned(forvar3776))) <<< $signed(((|reg3679) <<< (~|reg3639))));
                    end
                  reg3996 <= (reg3795 <<< $signed($signed(reg3713[(2'h3):(1'h1)])));
                  if (reg3684)
                    begin
                      reg3997 <= (reg3946 ?
                          $signed(reg3864) : (forvar3970 | ((8'h9f) ?
                              $unsigned(forvar3819) : $unsigned((8'haf)))));
                      reg3998 <= $unsigned(forvar3870);
                      reg3999 <= (forvar3638[(3'h4):(1'h1)] ~^ $unsigned(($unsigned((8'h9c)) - (^~reg3939))));
                    end
                  else
                    begin
                      reg3997 <= reg3785[(3'h4):(3'h4)];
                      reg3998 <= (^$unsigned((8'h9c)));
                    end
                  for (forvar4000 = (1'h0); (forvar4000 < (2'h3)); forvar4000 = (forvar4000 + (1'h1)))
                    begin
                      reg4001 <= $signed(forvar3686);
                      reg4002 <= ({reg3756[(4'h9):(3'h7)]} ^~ ($signed(reg3942) || $unsigned(forvar3725)));
                      reg4003 <= ($unsigned(($unsigned(forvar3986) ?
                          $signed(reg3785) : (reg3952 ?
                              forvar3688 : (8'had)))) <= reg3993[(3'h6):(1'h0)]);
                    end
                end
            end
          reg4004 <= $unsigned($unsigned((+forvar3971[(2'h3):(2'h2)])));
        end
      reg4014 <= $signed((&$unsigned($unsigned(reg3626))));
    end
  assign wire4015 = $unsigned(($signed(((8'haf) <<< forvar3776)) ?
                        $signed($unsigned(reg3690)) : forvar3951[(4'ha):(2'h2)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module3502
#( parameter param3600 = ((~^((~(8'h9f)) == ((8'h9f) ? (8'h9e) : (8'hb1)))) > {((~^(8'hac)) << ((8'ha5) ? (8'hab) : (8'ha2)))}) )
(y, clk, wire3507, wire3506, wire3505, wire3504, wire3503);
  output wire [(32'h482):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire3507;
  input wire signed [(3'h4):(1'h0)] wire3506;
  input wire signed [(2'h2):(1'h0)] wire3505;
  input wire signed [(3'h6):(1'h0)] wire3504;
  input wire [(3'h5):(1'h0)] wire3503;
  wire [(3'h6):(1'h0)] wire3599;
  wire [(2'h3):(1'h0)] wire3598;
  wire [(4'hb):(1'h0)] wire3597;
  wire signed [(3'h4):(1'h0)] wire3596;
  wire signed [(4'hf):(1'h0)] wire3595;
  reg signed [(4'hf):(1'h0)] reg3594 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3562 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3561 = (1'h0);
  reg [(4'hb):(1'h0)] reg3560 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3559 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3557 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3556 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3554 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3551 = (1'h0);
  reg [(3'h5):(1'h0)] forvar3546 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3539 = (1'h0);
  reg [(3'h7):(1'h0)] reg3548 = (1'h0);
  reg [(3'h7):(1'h0)] reg3547 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3543 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3542 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar3530 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3525 = (1'h0);
  reg [(3'h6):(1'h0)] reg3524 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3520 = (1'h0);
  reg [(4'h9):(1'h0)] forvar3514 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3512 = (1'h0);
  reg [(4'hf):(1'h0)] reg3593 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3592 = (1'h0);
  reg [(3'h4):(1'h0)] reg3591 = (1'h0);
  reg [(2'h2):(1'h0)] reg3590 = (1'h0);
  reg [(3'h4):(1'h0)] reg3589 = (1'h0);
  reg [(5'h10):(1'h0)] reg3588 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg3587 = (1'h0);
  reg [(4'h8):(1'h0)] reg3586 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3585 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3584 = (1'h0);
  reg [(4'h8):(1'h0)] reg3583 = (1'h0);
  reg [(4'he):(1'h0)] reg3582 = (1'h0);
  reg [(3'h6):(1'h0)] forvar3581 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3580 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3579 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3578 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3577 = (1'h0);
  reg [(4'hf):(1'h0)] reg3576 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3575 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3574 = (1'h0);
  reg [(4'hd):(1'h0)] reg3573 = (1'h0);
  reg [(3'h5):(1'h0)] reg3571 = (1'h0);
  reg [(4'hb):(1'h0)] forvar3570 = (1'h0);
  reg [(3'h7):(1'h0)] reg3572 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar3571 = (1'h0);
  reg [(4'h8):(1'h0)] reg3570 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3569 = (1'h0);
  reg [(3'h4):(1'h0)] reg3568 = (1'h0);
  reg [(5'h10):(1'h0)] reg3567 = (1'h0);
  reg [(4'hb):(1'h0)] reg3566 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3565 = (1'h0);
  reg [(4'hd):(1'h0)] reg3564 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3563 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar3562 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3561 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3560 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3559 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar3550 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3558 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg3557 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3556 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3555 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3554 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3553 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3552 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg3551 = (1'h0);
  reg [(4'hf):(1'h0)] reg3550 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3549 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3548 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar3547 = (1'h0);
  reg [(5'h10):(1'h0)] forvar3544 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3546 = (1'h0);
  reg [(2'h3):(1'h0)] reg3545 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3544 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg3543 = (1'h0);
  reg [(4'h8):(1'h0)] forvar3542 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3541 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg3540 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3539 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3538 = (1'h0);
  reg [(4'hb):(1'h0)] reg3537 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg3536 = (1'h0);
  reg [(5'h10):(1'h0)] reg3535 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3534 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3533 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3532 = (1'h0);
  reg [(4'hc):(1'h0)] reg3533 = (1'h0);
  reg [(2'h2):(1'h0)] forvar3532 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg3531 = (1'h0);
  reg [(4'h8):(1'h0)] reg3530 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3529 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar3517 = (1'h0);
  reg [(3'h4):(1'h0)] reg3515 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3528 = (1'h0);
  reg [(4'hb):(1'h0)] reg3527 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg3526 = (1'h0);
  reg [(2'h3):(1'h0)] reg3525 = (1'h0);
  reg [(3'h4):(1'h0)] forvar3524 = (1'h0);
  reg [(2'h2):(1'h0)] reg3523 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3522 = (1'h0);
  reg [(5'h10):(1'h0)] reg3521 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg3520 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar3519 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg3518 = (1'h0);
  reg [(2'h2):(1'h0)] reg3517 = (1'h0);
  reg [(2'h2):(1'h0)] reg3516 = (1'h0);
  reg [(4'he):(1'h0)] forvar3515 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar3511 = (1'h0);
  reg signed [(4'he):(1'h0)] reg3510 = (1'h0);
  reg [(4'hb):(1'h0)] reg3514 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg3513 = (1'h0);
  reg [(2'h2):(1'h0)] reg3512 = (1'h0);
  reg [(2'h3):(1'h0)] reg3511 = (1'h0);
  reg [(4'hd):(1'h0)] forvar3510 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar3509 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire3508;
  assign y = {wire3599,
                 wire3598,
                 wire3597,
                 wire3596,
                 wire3595,
                 reg3594,
                 reg3562,
                 forvar3561,
                 reg3560,
                 reg3559,
                 forvar3557,
                 forvar3556,
                 reg3554,
                 forvar3551,
                 forvar3546,
                 forvar3539,
                 reg3548,
                 reg3547,
                 forvar3543,
                 reg3542,
                 forvar3530,
                 forvar3525,
                 reg3524,
                 forvar3520,
                 forvar3514,
                 forvar3512,
                 reg3593,
                 reg3592,
                 reg3591,
                 reg3590,
                 reg3589,
                 reg3588,
                 reg3587,
                 reg3586,
                 reg3585,
                 forvar3584,
                 reg3583,
                 reg3582,
                 forvar3581,
                 reg3580,
                 forvar3579,
                 forvar3578,
                 reg3577,
                 reg3576,
                 forvar3575,
                 reg3574,
                 reg3573,
                 reg3571,
                 forvar3570,
                 reg3572,
                 forvar3571,
                 reg3570,
                 reg3569,
                 reg3568,
                 reg3567,
                 reg3566,
                 reg3565,
                 reg3564,
                 reg3563,
                 forvar3562,
                 reg3561,
                 forvar3560,
                 forvar3559,
                 forvar3550,
                 reg3558,
                 reg3557,
                 reg3556,
                 reg3555,
                 forvar3554,
                 reg3553,
                 reg3552,
                 reg3551,
                 reg3550,
                 reg3549,
                 forvar3548,
                 forvar3547,
                 forvar3544,
                 reg3546,
                 reg3545,
                 reg3544,
                 reg3543,
                 forvar3542,
                 reg3541,
                 reg3540,
                 reg3539,
                 reg3538,
                 reg3537,
                 reg3536,
                 reg3535,
                 reg3534,
                 forvar3533,
                 reg3532,
                 reg3533,
                 forvar3532,
                 reg3531,
                 reg3530,
                 reg3529,
                 forvar3517,
                 reg3515,
                 reg3528,
                 reg3527,
                 reg3526,
                 reg3525,
                 forvar3524,
                 reg3523,
                 reg3522,
                 reg3521,
                 reg3520,
                 forvar3519,
                 reg3518,
                 reg3517,
                 reg3516,
                 forvar3515,
                 forvar3511,
                 reg3510,
                 reg3514,
                 reg3513,
                 reg3512,
                 reg3511,
                 forvar3510,
                 forvar3509,
                 wire3508,
                 (1'h0)};
  assign wire3508 = $signed($unsigned((+{(8'ha4)})));
  always
    @(posedge clk) begin
      if (wire3506[(3'h4):(2'h3)])
        begin
          for (forvar3509 = (1'h0); (forvar3509 < (1'h1)); forvar3509 = (forvar3509 + (1'h1)))
            begin
              if ($signed(wire3505))
                begin
                  for (forvar3510 = (1'h0); (forvar3510 < (2'h3)); forvar3510 = (forvar3510 + (1'h1)))
                    begin
                      reg3511 <= ((forvar3510 != $unsigned($unsigned(wire3508))) * ($unsigned((^(8'ha7))) == (~{wire3508})));
                      reg3512 <= forvar3509[(4'hd):(4'hc)];
                    end
                  reg3513 <= $signed(forvar3510[(4'h9):(3'h4)]);
                  reg3514 <= (wire3504[(1'h1):(1'h0)] ? wire3503 : wire3508);
                end
              else
                begin
                  reg3510 <= reg3514[(4'hb):(4'h8)];
                  for (forvar3511 = (1'h0); (forvar3511 < (1'h0)); forvar3511 = (forvar3511 + (1'h1)))
                    begin
                      reg3512 <= $signed((((~|wire3504) ?
                          (forvar3511 ?
                              (8'hb1) : (8'ha1)) : $signed(wire3505)) >> ((reg3513 ?
                          wire3508 : wire3507) | $signed(reg3513))));
                      reg3513 <= wire3504;
                      reg3514 <= ((^~$unsigned({reg3514})) > (($signed(wire3505) & $signed(reg3510)) > (~{reg3511})));
                    end
                end
              if (({$unsigned({reg3514})} ?
                  {reg3514[(3'h6):(2'h2)]} : ($signed($signed(forvar3510)) ?
                      (^$signed(wire3506)) : $unsigned({forvar3510}))))
                begin
                  for (forvar3515 = (1'h0); (forvar3515 < (1'h0)); forvar3515 = (forvar3515 + (1'h1)))
                    begin
                      reg3516 <= reg3512[(2'h2):(1'h0)];
                      reg3517 <= ((8'hba) << $unsigned((reg3512 != $unsigned((8'hb8)))));
                      reg3518 <= wire3506[(1'h1):(1'h1)];
                    end
                  for (forvar3519 = (1'h0); (forvar3519 < (1'h0)); forvar3519 = (forvar3519 + (1'h1)))
                    begin
                      reg3520 <= (wire3505[(1'h0):(1'h0)] ?
                          forvar3509 : (+((forvar3509 ?
                              wire3503 : wire3507) ~^ (+reg3516))));
                    end
                  if ($signed(((&reg3510[(4'ha):(3'h7)]) ^~ reg3518)))
                    begin
                      reg3521 <= wire3507;
                      reg3522 <= forvar3510[(3'h5):(3'h5)];
                      reg3523 <= (8'hb6);
                    end
                  else
                    begin
                      reg3521 <= $signed(reg3512);
                      reg3522 <= {(reg3522 || (|$signed(wire3505)))};
                    end
                  for (forvar3524 = (1'h0); (forvar3524 < (2'h3)); forvar3524 = (forvar3524 + (1'h1)))
                    begin
                      reg3525 <= (^~(|((reg3510 ~^ wire3505) ^ (reg3518 ?
                          wire3505 : (8'hb4)))));
                      reg3526 <= {((8'haf) != (8'hb2))};
                      reg3527 <= (|$unsigned((reg3517 ?
                          (~&reg3510) : {(8'hb2)})));
                      reg3528 <= ({$signed((forvar3515 ?
                              (8'hba) : forvar3511))} >>> $unsigned($signed($unsigned(forvar3511))));
                    end
                end
              else
                begin
                  if ($unsigned($signed($signed($unsigned((8'hb3))))))
                    begin
                      reg3515 <= (&(8'h9f));
                      reg3516 <= reg3520;
                    end
                  else
                    begin
                      reg3515 <= (($unsigned((reg3526 << reg3514)) ?
                              {(+reg3528)} : $unsigned((reg3526 ?
                                  reg3517 : forvar3510))) ?
                          (!(~&(wire3508 ?
                              reg3513 : wire3506))) : ({$signed(reg3527)} & wire3504[(3'h4):(3'h4)]));
                    end
                  for (forvar3517 = (1'h0); (forvar3517 < (2'h3)); forvar3517 = (forvar3517 + (1'h1)))
                    begin
                      reg3518 <= $signed($signed($signed((^(8'hac)))));
                    end
                  for (forvar3519 = (1'h0); (forvar3519 < (1'h0)); forvar3519 = (forvar3519 + (1'h1)))
                    begin
                      reg3520 <= $unsigned(reg3515);
                    end
                end
              if ((($unsigned($signed(forvar3515)) ?
                  (reg3526[(4'h9):(1'h0)] >= wire3507[(3'h7):(3'h4)]) : $signed(wire3506)) != (({reg3520} >>> {reg3517}) ?
                  ((wire3508 ?
                      reg3522 : (8'hb7)) | wire3504) : (~|(reg3517 && forvar3511)))))
                begin
                  if (reg3523)
                    begin
                      reg3529 <= $signed(reg3525);
                    end
                  else
                    begin
                      reg3529 <= $unsigned(({reg3513} > (^$unsigned(wire3507))));
                      reg3530 <= $unsigned($signed(forvar3524[(1'h1):(1'h0)]));
                      reg3531 <= (~|$unsigned(reg3528[(3'h5):(3'h5)]));
                    end
                  for (forvar3532 = (1'h0); (forvar3532 < (1'h0)); forvar3532 = (forvar3532 + (1'h1)))
                    begin
                      reg3533 <= (($unsigned($signed(reg3525)) ?
                          ($signed(reg3510) ^ (reg3513 && (8'h9f))) : ((reg3513 ?
                                  forvar3509 : wire3506) ?
                              $signed((8'h9d)) : (reg3510 ?
                                  reg3516 : reg3529))) ^~ $signed($signed(reg3527)));
                    end
                end
              else
                begin
                  reg3529 <= (forvar3517 ?
                      (forvar3519[(2'h3):(1'h1)] < {(forvar3510 ?
                              reg3530 : reg3512)}) : wire3507[(3'h5):(1'h0)]);
                  if (wire3508)
                    begin
                      reg3530 <= $unsigned((($unsigned(reg3514) ?
                          forvar3519 : (&reg3520)) && ({reg3516} ?
                          reg3529[(2'h2):(1'h0)] : (!reg3527))));
                      reg3531 <= (($signed($signed(reg3517)) ?
                          (8'ha5) : reg3515[(3'h4):(3'h4)]) >> ($unsigned(reg3513) ?
                          ((!wire3505) || reg3513) : (~&(reg3525 ?
                              (8'ha0) : wire3508))));
                      reg3532 <= ($signed(({(8'hb7)} * forvar3519)) ?
                          {((wire3507 ?
                                  reg3525 : reg3522) | forvar3511)} : forvar3524[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg3530 <= (forvar3519 ?
                          reg3516[(1'h1):(1'h1)] : (~^((~&reg3514) ?
                              $signed(forvar3532) : (8'haa))));
                    end
                  for (forvar3533 = (1'h0); (forvar3533 < (2'h3)); forvar3533 = (forvar3533 + (1'h1)))
                    begin
                      reg3534 <= (!reg3512[(1'h1):(1'h0)]);
                      reg3535 <= reg3533[(3'h4):(1'h0)];
                      reg3536 <= $unsigned($unsigned(forvar3533));
                    end
                  if ((^((~&reg3529) < (&(reg3529 & reg3529)))))
                    begin
                      reg3537 <= $unsigned($unsigned(($unsigned(reg3515) ?
                          $unsigned((8'hb1)) : (wire3503 ?
                              reg3531 : wire3508))));
                    end
                  else
                    begin
                      reg3537 <= (8'hb2);
                      reg3538 <= (|$signed(reg3531));
                      reg3539 <= reg3523;
                      reg3540 <= {($unsigned(reg3511[(1'h1):(1'h1)]) ~^ ($signed(reg3527) ?
                              reg3525 : ((8'h9c) >>> reg3510)))};
                    end
                end
              reg3541 <= reg3527[(3'h7):(1'h1)];
            end
          for (forvar3542 = (1'h0); (forvar3542 < (1'h1)); forvar3542 = (forvar3542 + (1'h1)))
            begin
              reg3543 <= ($unsigned(($signed(reg3515) ? {reg3536} : reg3515)) ?
                  $signed({{reg3525}}) : (reg3535 ~^ forvar3511[(2'h3):(2'h3)]));
              if (reg3513)
                begin
                  if ({$signed(({reg3537} ^~ (~|(8'hb8))))})
                    begin
                      reg3544 <= (reg3528[(3'h6):(3'h5)] ^ {$signed((reg3531 ?
                              reg3510 : reg3538))});
                    end
                  else
                    begin
                      reg3544 <= $signed((~^({wire3505} ?
                          (reg3513 | forvar3509) : $signed(reg3536))));
                      reg3545 <= forvar3532;
                    end
                  reg3546 <= $unsigned(forvar3542[(4'h8):(1'h1)]);
                end
              else
                begin
                  for (forvar3544 = (1'h0); (forvar3544 < (1'h1)); forvar3544 = (forvar3544 + (1'h1)))
                    begin
                      reg3545 <= $unsigned((wire3507 ?
                          $unsigned((wire3504 ^~ reg3535)) : $unsigned(reg3522)));
                      reg3546 <= reg3525[(2'h2):(1'h1)];
                    end
                end
            end
          for (forvar3547 = (1'h0); (forvar3547 < (1'h0)); forvar3547 = (forvar3547 + (1'h1)))
            begin
              for (forvar3548 = (1'h0); (forvar3548 < (1'h0)); forvar3548 = (forvar3548 + (1'h1)))
                begin
                  reg3549 <= ({$unsigned((&forvar3533))} | {forvar3544[(3'h6):(3'h4)]});
                end
              if ($signed(reg3543[(3'h7):(2'h3)]))
                begin
                  if (reg3531)
                    begin
                      reg3550 <= (8'hac);
                    end
                  else
                    begin
                      reg3550 <= $signed(reg3529[(3'h5):(2'h2)]);
                      reg3551 <= (((reg3526 + (8'hba)) >= $signed($signed(reg3541))) ?
                          (reg3536[(3'h5):(1'h0)] >= {(reg3513 ?
                                  forvar3548 : (8'hb8))}) : $signed((~^(reg3522 * reg3516))));
                      reg3552 <= forvar3519;
                      reg3553 <= reg3521;
                    end
                  for (forvar3554 = (1'h0); (forvar3554 < (1'h1)); forvar3554 = (forvar3554 + (1'h1)))
                    begin
                      reg3555 <= $signed(reg3521[(4'h8):(2'h2)]);
                      reg3556 <= $unsigned(wire3506[(1'h1):(1'h1)]);
                      reg3557 <= {reg3521[(4'hc):(4'h9)]};
                      reg3558 <= reg3523;
                    end
                end
              else
                begin
                  for (forvar3550 = (1'h0); (forvar3550 < (1'h1)); forvar3550 = (forvar3550 + (1'h1)))
                    begin
                      reg3551 <= (((-reg3557) > $unsigned((~|reg3541))) || $unsigned((!$signed(forvar3517))));
                      reg3552 <= forvar3517;
                    end
                end
              for (forvar3559 = (1'h0); (forvar3559 < (2'h2)); forvar3559 = (forvar3559 + (1'h1)))
                begin
                  for (forvar3560 = (1'h0); (forvar3560 < (1'h0)); forvar3560 = (forvar3560 + (1'h1)))
                    begin
                      reg3561 <= $signed($signed(reg3536));
                    end
                  for (forvar3562 = (1'h0); (forvar3562 < (2'h2)); forvar3562 = (forvar3562 + (1'h1)))
                    begin
                      reg3563 <= (($unsigned({wire3507}) ?
                          ((~wire3507) >> (forvar3532 ?
                              reg3539 : forvar3554)) : ((-(8'ha8)) ?
                              (reg3539 && reg3512) : (forvar3559 > reg3528))) >> $signed(forvar3562[(2'h3):(1'h0)]));
                      reg3564 <= $unsigned(reg3539);
                    end
                  if (reg3513[(1'h0):(1'h0)])
                    begin
                      reg3565 <= $signed(reg3515);
                      reg3566 <= $unsigned((reg3510[(4'he):(4'h9)] ?
                          reg3520 : (reg3515 ?
                              $signed(reg3561) : forvar3559[(2'h2):(1'h0)])));
                      reg3567 <= reg3557[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg3565 <= (~(forvar3511[(3'h4):(1'h0)] << $unsigned($signed(reg3511))));
                      reg3566 <= reg3513[(3'h5):(2'h2)];
                      reg3567 <= {(reg3540[(1'h0):(1'h0)] ?
                              $unsigned((reg3553 ?
                                  reg3515 : reg3540)) : (^(!reg3515)))};
                      reg3568 <= $unsigned(forvar3559[(1'h1):(1'h0)]);
                    end
                  reg3569 <= $unsigned(((&$unsigned(reg3511)) ?
                      reg3527[(2'h2):(2'h2)] : reg3561));
                end
              if ($unsigned(((~&{forvar3532}) & $unsigned({forvar3562}))))
                begin
                  reg3570 <= ((reg3544[(3'h6):(3'h6)] && $signed(reg3530)) & forvar3547[(2'h2):(2'h2)]);
                  for (forvar3571 = (1'h0); (forvar3571 < (1'h1)); forvar3571 = (forvar3571 + (1'h1)))
                    begin
                      reg3572 <= (~|$signed($signed((~&reg3516))));
                    end
                end
              else
                begin
                  for (forvar3570 = (1'h0); (forvar3570 < (2'h3)); forvar3570 = (forvar3570 + (1'h1)))
                    begin
                      reg3571 <= (-wire3508);
                      reg3572 <= $signed((($signed((8'h9f)) == (reg3536 + reg3511)) ?
                          $signed((|(8'hb4))) : (~(reg3536 <= reg3557))));
                    end
                  if ((wire3507[(2'h3):(1'h1)] <<< $unsigned($unsigned($signed(reg3543)))))
                    begin
                      reg3573 <= {$unsigned(reg3552)};
                    end
                  else
                    begin
                      reg3573 <= {(-forvar3562[(3'h7):(2'h3)])};
                      reg3574 <= reg3516;
                    end
                  for (forvar3575 = (1'h0); (forvar3575 < (2'h2)); forvar3575 = (forvar3575 + (1'h1)))
                    begin
                      reg3576 <= $signed({forvar3547});
                      reg3577 <= ({(~^$signed(reg3572))} - reg3511[(2'h2):(2'h2)]);
                    end
                end
            end
          for (forvar3578 = (1'h0); (forvar3578 < (2'h2)); forvar3578 = (forvar3578 + (1'h1)))
            begin
              for (forvar3579 = (1'h0); (forvar3579 < (2'h2)); forvar3579 = (forvar3579 + (1'h1)))
                begin
                  reg3580 <= reg3558;
                  for (forvar3581 = (1'h0); (forvar3581 < (2'h3)); forvar3581 = (forvar3581 + (1'h1)))
                    begin
                      reg3582 <= reg3551;
                      reg3583 <= {$unsigned(wire3508[(3'h5):(1'h1)])};
                    end
                  for (forvar3584 = (1'h0); (forvar3584 < (2'h3)); forvar3584 = (forvar3584 + (1'h1)))
                    begin
                      reg3585 <= $unsigned($signed((!(~^forvar3510))));
                      reg3586 <= $signed($signed((8'h9f)));
                      reg3587 <= ($signed((wire3503[(1'h1):(1'h1)] == (8'ha2))) < ({$unsigned(reg3565)} ?
                          $unsigned(reg3532[(3'h4):(1'h0)]) : reg3534));
                      reg3588 <= ($signed(($signed((8'ha8)) >>> reg3531)) || (~|(((8'ha2) <= reg3510) > (+wire3503))));
                    end
                  if ({$signed($unsigned($unsigned(reg3531)))})
                    begin
                      reg3589 <= (8'hac);
                      reg3590 <= {{reg3564}};
                      reg3591 <= (~$signed($signed($unsigned(reg3546))));
                      reg3592 <= {(forvar3519 ?
                              $unsigned(forvar3550[(1'h1):(1'h1)]) : reg3537[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg3589 <= reg3589[(3'h4):(1'h0)];
                      reg3590 <= $signed(reg3553);
                      reg3591 <= $signed({(8'h9f)});
                    end
                end
              reg3593 <= reg3564;
            end
        end
      else
        begin
          for (forvar3509 = (1'h0); (forvar3509 < (1'h1)); forvar3509 = (forvar3509 + (1'h1)))
            begin
              reg3510 <= ((reg3561 <<< (&reg3523[(1'h0):(1'h0)])) ?
                  forvar3510[(3'h6):(3'h6)] : reg3523[(1'h0):(1'h0)]);
              for (forvar3511 = (1'h0); (forvar3511 < (2'h2)); forvar3511 = (forvar3511 + (1'h1)))
                begin
                  for (forvar3512 = (1'h0); (forvar3512 < (2'h3)); forvar3512 = (forvar3512 + (1'h1)))
                    begin
                      reg3513 <= reg3589[(2'h3):(1'h1)];
                    end
                  for (forvar3514 = (1'h0); (forvar3514 < (2'h3)); forvar3514 = (forvar3514 + (1'h1)))
                    begin
                      reg3515 <= reg3532;
                      reg3516 <= $signed(({forvar3571} ?
                          (reg3573[(3'h4):(3'h4)] ?
                              $signed((8'hab)) : reg3543) : (((8'haf) ?
                                  forvar3514 : (8'ha2)) ?
                              $unsigned(reg3543) : (reg3536 ?
                                  wire3504 : reg3553))));
                      reg3517 <= $signed(($signed($unsigned(forvar3581)) ?
                          ($signed(reg3586) ?
                              reg3582[(4'hd):(1'h1)] : $unsigned(reg3530)) : forvar3550[(1'h1):(1'h1)]));
                      reg3518 <= $unsigned($signed(($signed(reg3534) ^~ $signed(forvar3514))));
                    end
                end
            end
          for (forvar3519 = (1'h0); (forvar3519 < (1'h0)); forvar3519 = (forvar3519 + (1'h1)))
            begin
              if (reg3593)
                begin
                  for (forvar3520 = (1'h0); (forvar3520 < (2'h3)); forvar3520 = (forvar3520 + (1'h1)))
                    begin
                      reg3521 <= reg3555;
                      reg3522 <= $signed(({(reg3518 << reg3539)} ?
                          (~^$unsigned(forvar3533)) : (^(reg3588 ?
                              reg3536 : reg3530))));
                      reg3523 <= {forvar3550[(3'h4):(1'h1)]};
                      reg3524 <= $unsigned($signed(($unsigned((8'h9f)) ?
                          {forvar3515} : $unsigned(forvar3548))));
                    end
                end
              else
                begin
                  if ({($unsigned((reg3524 ?
                          (8'h9c) : forvar3511)) || $signed(forvar3533))})
                    begin
                      reg3520 <= reg3566;
                      reg3521 <= $signed(($unsigned((~&(8'hb8))) ?
                          $signed((^forvar3560)) : ((~wire3507) || $unsigned((8'hb8)))));
                      reg3522 <= reg3526;
                      reg3523 <= (+(8'ha2));
                    end
                  else
                    begin
                      reg3520 <= (^($unsigned($signed(forvar3509)) ?
                          (&reg3546) : $signed((8'ha8))));
                      reg3521 <= (-forvar3542[(3'h4):(2'h2)]);
                    end
                  reg3524 <= reg3530;
                  for (forvar3525 = (1'h0); (forvar3525 < (2'h2)); forvar3525 = (forvar3525 + (1'h1)))
                    begin
                      reg3526 <= $signed(reg3550);
                      reg3527 <= (reg3586 - reg3564);
                      reg3528 <= (~&(8'had));
                      reg3529 <= reg3568;
                    end
                end
              for (forvar3530 = (1'h0); (forvar3530 < (2'h3)); forvar3530 = (forvar3530 + (1'h1)))
                begin
                  if ($signed($signed({(~&reg3520)})))
                    begin
                      reg3531 <= reg3537[(3'h4):(2'h3)];
                      reg3532 <= {($unsigned((reg3526 ?
                              reg3589 : (8'hae))) <= ((wire3505 ~^ forvar3571) ?
                              ((8'haa) ? reg3580 : forvar3510) : (reg3521 ?
                                  reg3561 : (8'hb0))))};
                      reg3533 <= reg3549;
                    end
                  else
                    begin
                      reg3531 <= (8'ha6);
                      reg3532 <= forvar3510[(2'h3):(1'h1)];
                      reg3533 <= reg3561[(1'h1):(1'h1)];
                      reg3534 <= $unsigned(((8'had) ?
                          (forvar3550 & (-forvar3525)) : $unsigned(reg3552)));
                    end
                  if ($unsigned(($unsigned((-reg3557)) ?
                      {(^reg3568)} : reg3520)))
                    begin
                      reg3535 <= ((({reg3516} >= $signed(reg3553)) ?
                          forvar3578[(1'h0):(1'h0)] : {(~&reg3521)}) ~^ $unsigned($unsigned($signed(reg3586))));
                      reg3536 <= reg3540[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg3535 <= $unsigned($unsigned((|$unsigned(reg3530))));
                      reg3536 <= ((~^(~^{forvar3524})) ?
                          $signed(reg3511[(2'h3):(2'h3)]) : $unsigned(reg3520));
                      reg3537 <= reg3520[(1'h0):(1'h0)];
                    end
                end
              reg3538 <= (!$unsigned((reg3540[(3'h4):(1'h1)] > $unsigned(reg3528))));
            end
          if ((8'hae))
            begin
              if ((reg3540[(3'h4):(1'h1)] <= $signed(forvar3514[(3'h7):(2'h3)])))
                begin
                  reg3539 <= $unsigned($signed(($unsigned((8'ha3)) ?
                      {reg3550} : (&forvar3544))));
                  if (($unsigned(reg3590) ? reg3591 : (~^reg3551)))
                    begin
                      reg3540 <= (~(($unsigned((8'hb8)) != ((8'ha5) ?
                              forvar3584 : reg3511)) ?
                          {(forvar3509 ? reg3535 : reg3585)} : (forvar3581 ?
                              reg3514[(4'ha):(4'ha)] : forvar3509)));
                    end
                  else
                    begin
                      reg3540 <= (^~$signed(((reg3524 ?
                          reg3510 : reg3524) & (!reg3557))));
                      reg3541 <= $unsigned(wire3507[(3'h5):(3'h4)]);
                    end
                  if ((8'hb7))
                    begin
                      reg3542 <= $unsigned($signed($unsigned($signed(reg3537))));
                      reg3543 <= forvar3547;
                      reg3544 <= reg3528[(4'h8):(1'h1)];
                    end
                  else
                    begin
                      reg3542 <= $signed((($signed(wire3504) && reg3524[(3'h6):(2'h3)]) ?
                          $signed((8'hb5)) : ($unsigned((8'h9e)) ?
                              (reg3518 != reg3526) : forvar3584[(1'h0):(1'h0)])));
                      reg3543 <= $unsigned((8'hac));
                      reg3544 <= forvar3575[(4'h8):(1'h0)];
                    end
                end
              else
                begin
                  if (reg3526[(4'h9):(1'h0)])
                    begin
                      reg3539 <= $unsigned((reg3556 ?
                          (^~(~|reg3589)) : reg3573));
                      reg3540 <= (~^(~|(forvar3579 ?
                          (forvar3512 & reg3518) : $unsigned(reg3529))));
                      reg3541 <= ((~(^(forvar3510 - reg3558))) ?
                          (^~(reg3521 ?
                              $unsigned(reg3551) : (reg3520 ^ reg3533))) : ((&$signed(reg3565)) < $unsigned($signed((8'haa)))));
                      reg3542 <= (+((^~(forvar3554 ?
                          (8'ha8) : reg3543)) >> reg3566));
                    end
                  else
                    begin
                      reg3539 <= $signed(forvar3581[(2'h3):(1'h0)]);
                      reg3540 <= ($signed(reg3566) ?
                          (8'ha5) : $unsigned($signed(reg3557)));
                    end
                  for (forvar3543 = (1'h0); (forvar3543 < (2'h3)); forvar3543 = (forvar3543 + (1'h1)))
                    begin
                      reg3544 <= $signed(forvar3520);
                    end
                  if (reg3580[(3'h5):(3'h5)])
                    begin
                      reg3545 <= (~^$signed({reg3593[(4'ha):(3'h5)]}));
                      reg3546 <= $unsigned((~forvar3547[(2'h2):(2'h2)]));
                      reg3547 <= ($unsigned((forvar3530[(2'h2):(1'h0)] || (forvar3544 ?
                          reg3523 : reg3530))) << {($unsigned(reg3525) >> $unsigned(reg3567))});
                      reg3548 <= $unsigned((forvar3570[(1'h0):(1'h0)] | reg3527[(2'h3):(2'h2)]));
                    end
                  else
                    begin
                      reg3545 <= reg3546[(4'ha):(3'h5)];
                      reg3546 <= $unsigned($unsigned(reg3535[(4'hc):(4'hb)]));
                      reg3547 <= reg3556[(1'h1):(1'h0)];
                      reg3548 <= $signed(({(!reg3591)} ?
                          {(|reg3517)} : forvar3581[(2'h2):(1'h1)]));
                    end
                end
            end
          else
            begin
              for (forvar3539 = (1'h0); (forvar3539 < (1'h0)); forvar3539 = (forvar3539 + (1'h1)))
                begin
                  if ((~&(+(~$signed(forvar3509)))))
                    begin
                      reg3540 <= (&(reg3537 ?
                          $unsigned(forvar3517[(4'ha):(3'h7)]) : ({wire3504} | reg3573)));
                      reg3541 <= (reg3550[(3'h5):(2'h3)] ?
                          reg3574 : $unsigned(((reg3514 ?
                              forvar3524 : reg3580) - ((8'hb8) ?
                              forvar3571 : wire3505))));
                    end
                  else
                    begin
                      reg3540 <= {{forvar3517[(4'hc):(2'h2)]}};
                      reg3541 <= $unsigned({reg3564[(4'hb):(4'h8)]});
                      reg3542 <= ((!(!(^forvar3509))) << $unsigned($unsigned($unsigned(reg3532))));
                    end
                  reg3543 <= {reg3573};
                end
              if ({($unsigned((forvar3519 ? reg3525 : forvar3575)) ?
                      ((forvar3547 ? reg3537 : reg3531) ?
                          $unsigned((8'hb9)) : reg3539[(3'h6):(3'h6)]) : {{reg3573}})})
                begin
                  for (forvar3544 = (1'h0); (forvar3544 < (1'h0)); forvar3544 = (forvar3544 + (1'h1)))
                    begin
                      reg3545 <= ({{reg3545}} ?
                          wire3504[(1'h1):(1'h1)] : {$unsigned($unsigned((8'haa)))});
                    end
                  for (forvar3546 = (1'h0); (forvar3546 < (1'h0)); forvar3546 = (forvar3546 + (1'h1)))
                    begin
                      reg3547 <= $signed(((^$signed(forvar3517)) <<< (forvar3547[(2'h3):(1'h0)] < $unsigned(reg3542))));
                      reg3548 <= ((^((-reg3591) ?
                          {(8'hac)} : (~|forvar3539))) * ($signed($signed(forvar3543)) ^ ((^reg3537) | $signed(reg3558))));
                      reg3549 <= ({(^~(reg3539 ?
                              reg3551 : forvar3532))} || $unsigned(reg3522[(1'h1):(1'h0)]));
                    end
                end
              else
                begin
                  reg3544 <= $unsigned($signed((+reg3569[(1'h0):(1'h0)])));
                  reg3545 <= forvar3546[(2'h3):(1'h0)];
                  for (forvar3546 = (1'h0); (forvar3546 < (1'h0)); forvar3546 = (forvar3546 + (1'h1)))
                    begin
                      reg3547 <= reg3586[(3'h5):(1'h0)];
                      reg3548 <= forvar3532;
                      reg3549 <= reg3571;
                    end
                end
              for (forvar3550 = (1'h0); (forvar3550 < (2'h2)); forvar3550 = (forvar3550 + (1'h1)))
                begin
                  for (forvar3551 = (1'h0); (forvar3551 < (2'h2)); forvar3551 = (forvar3551 + (1'h1)))
                    begin
                      reg3552 <= forvar3514[(3'h7):(1'h1)];
                      reg3553 <= (8'hb8);
                    end
                  reg3554 <= (($unsigned(forvar3543) | reg3569[(3'h5):(1'h0)]) == reg3586);
                  reg3555 <= forvar3543;
                end
              for (forvar3556 = (1'h0); (forvar3556 < (2'h2)); forvar3556 = (forvar3556 + (1'h1)))
                begin
                  for (forvar3557 = (1'h0); (forvar3557 < (1'h1)); forvar3557 = (forvar3557 + (1'h1)))
                    begin
                      reg3558 <= (~reg3514);
                      reg3559 <= (forvar3559 ?
                          (~^({reg3531} >>> (!reg3580))) : ({wire3507} >> wire3503[(3'h5):(1'h1)]));
                      reg3560 <= reg3554;
                    end
                  for (forvar3561 = (1'h0); (forvar3561 < (2'h3)); forvar3561 = (forvar3561 + (1'h1)))
                    begin
                      reg3562 <= forvar3520[(1'h0):(1'h0)];
                    end
                end
            end
          reg3563 <= reg3586[(2'h2):(1'h0)];
        end
      reg3594 <= $unsigned((!$unsigned(((8'hba) ~^ reg3540))));
    end
  assign wire3595 = (($signed({reg3548}) ?
                        ((forvar3539 || forvar3551) >>> (~^forvar3519)) : (reg3532 > reg3528)) > (reg3542[(2'h2):(1'h1)] * $unsigned(forvar3530)));
  assign wire3596 = (8'ha0);
  assign wire3597 = $unsigned(reg3537);
  assign wire3598 = $unsigned($unsigned($signed(forvar3550[(1'h0):(1'h0)])));
  assign wire3599 = $signed(forvar3578);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1764
#( parameter param2748 = ((((^~(8'h9c)) ? ((8'ha8) <<< (8'h9e)) : ((8'hb9) ? (8'ha5) : (8'ha3))) * {{(8'ha6)}}) > (^~(8'hb1))) )
(y, clk, wire1768, wire1767, wire1766, wire1765);
  output wire [(32'h1539):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire1768;
  input wire signed [(4'h9):(1'h0)] wire1767;
  input wire [(5'h10):(1'h0)] wire1766;
  input wire signed [(2'h3):(1'h0)] wire1765;
  wire signed [(3'h7):(1'h0)] wire2747;
  wire signed [(4'hf):(1'h0)] wire2746;
  reg [(4'hf):(1'h0)] reg2745 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2744 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2743 = (1'h0);
  reg [(4'hd):(1'h0)] reg2742 = (1'h0);
  reg [(4'h8):(1'h0)] reg2741 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2740 = (1'h0);
  reg [(4'he):(1'h0)] reg2739 = (1'h0);
  reg [(4'h8):(1'h0)] reg2738 = (1'h0);
  reg [(5'h10):(1'h0)] reg2737 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2736 = (1'h0);
  reg [(4'h9):(1'h0)] reg2735 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2734 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2733 = (1'h0);
  reg [(5'h10):(1'h0)] reg2732 = (1'h0);
  reg [(4'hb):(1'h0)] reg2731 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2730 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2729 = (1'h0);
  reg [(4'hd):(1'h0)] reg2728 = (1'h0);
  reg [(3'h5):(1'h0)] reg2727 = (1'h0);
  reg [(4'hd):(1'h0)] reg2726 = (1'h0);
  reg [(3'h5):(1'h0)] reg2725 = (1'h0);
  reg [(4'hc):(1'h0)] reg2724 = (1'h0);
  reg [(4'hb):(1'h0)] reg2723 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2722 = (1'h0);
  reg [(4'hc):(1'h0)] reg2721 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2720 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2719 = (1'h0);
  reg [(4'ha):(1'h0)] reg2718 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2717 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2716 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2715 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2714 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2713 = (1'h0);
  reg [(2'h3):(1'h0)] reg2712 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2711 = (1'h0);
  reg [(4'h9):(1'h0)] reg2710 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2709 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2708 = (1'h0);
  reg [(4'h9):(1'h0)] reg2707 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2706 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2705 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2680 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2677 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2674 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2672 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2669 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2667 = (1'h0);
  reg [(3'h7):(1'h0)] reg2665 = (1'h0);
  reg [(4'h8):(1'h0)] reg2693 = (1'h0);
  reg [(4'hf):(1'h0)] reg2704 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2703 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2702 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2701 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2700 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2699 = (1'h0);
  reg [(3'h7):(1'h0)] reg2698 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2697 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2696 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2695 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2694 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2693 = (1'h0);
  reg [(3'h6):(1'h0)] reg2676 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2675 = (1'h0);
  reg [(4'hf):(1'h0)] reg2673 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2668 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2666 = (1'h0);
  reg [(4'hf):(1'h0)] reg2692 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2691 = (1'h0);
  reg [(4'hf):(1'h0)] reg2690 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2689 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2688 = (1'h0);
  reg [(5'h10):(1'h0)] reg2687 = (1'h0);
  reg [(3'h6):(1'h0)] reg2686 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2685 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2684 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2683 = (1'h0);
  reg [(4'hb):(1'h0)] reg2682 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2681 = (1'h0);
  reg [(5'h10):(1'h0)] reg2680 = (1'h0);
  reg [(3'h7):(1'h0)] reg2679 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2678 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2677 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2676 = (1'h0);
  reg [(3'h6):(1'h0)] reg2675 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2674 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2673 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2672 = (1'h0);
  reg [(3'h7):(1'h0)] reg2671 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2670 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2669 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2668 = (1'h0);
  reg [(2'h3):(1'h0)] reg2667 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2666 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2665 = (1'h0);
  reg [(4'ha):(1'h0)] reg2664 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2659 = (1'h0);
  reg [(4'hc):(1'h0)] reg2663 = (1'h0);
  reg [(2'h3):(1'h0)] reg2662 = (1'h0);
  reg [(3'h4):(1'h0)] reg2661 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2660 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2659 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2650 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2649 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2658 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2657 = (1'h0);
  reg [(4'hc):(1'h0)] reg2656 = (1'h0);
  reg [(4'he):(1'h0)] forvar2655 = (1'h0);
  reg [(4'hf):(1'h0)] reg2654 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2653 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2652 = (1'h0);
  reg [(3'h5):(1'h0)] reg2651 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2650 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2649 = (1'h0);
  reg [(2'h3):(1'h0)] reg2648 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2647 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2646 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2645 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2644 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2643 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2642 = (1'h0);
  reg [(4'hf):(1'h0)] reg2641 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2640 = (1'h0);
  reg [(5'h10):(1'h0)] reg2639 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2632 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2630 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2638 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2637 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2636 = (1'h0);
  reg [(3'h7):(1'h0)] reg2631 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2629 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2627 = (1'h0);
  reg [(3'h5):(1'h0)] reg2626 = (1'h0);
  reg [(4'hf):(1'h0)] reg2635 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2634 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2633 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2632 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2631 = (1'h0);
  reg [(4'hd):(1'h0)] reg2630 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2629 = (1'h0);
  reg [(4'hb):(1'h0)] reg2628 = (1'h0);
  reg [(2'h3):(1'h0)] reg2627 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2626 = (1'h0);
  reg [(3'h5):(1'h0)] reg2625 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2624 = (1'h0);
  reg [(3'h7):(1'h0)] reg2623 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2622 = (1'h0);
  reg [(3'h7):(1'h0)] reg2621 = (1'h0);
  reg [(4'hd):(1'h0)] reg2620 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2619 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2618 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2617 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2616 = (1'h0);
  reg [(4'hf):(1'h0)] reg2615 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2614 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2613 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2612 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2611 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2610 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2609 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2608 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2607 = (1'h0);
  reg [(4'h8):(1'h0)] reg2606 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2605 = (1'h0);
  reg [(4'ha):(1'h0)] reg2604 = (1'h0);
  reg [(4'ha):(1'h0)] reg2603 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2602 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2601 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2600 = (1'h0);
  reg [(4'hc):(1'h0)] reg2599 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2598 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2597 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2596 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2595 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2594 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2593 = (1'h0);
  reg [(3'h5):(1'h0)] reg2592 = (1'h0);
  reg [(2'h2):(1'h0)] reg2591 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2590 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2588 = (1'h0);
  reg [(3'h5):(1'h0)] reg2590 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2589 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2588 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2587 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2586 = (1'h0);
  wire [(4'ha):(1'h0)] wire2585;
  wire signed [(3'h5):(1'h0)] wire2584;
  wire signed [(3'h5):(1'h0)] wire2582;
  wire signed [(3'h4):(1'h0)] wire2121;
  wire [(4'h9):(1'h0)] wire2120;
  reg [(4'he):(1'h0)] reg2088 = (1'h0);
  reg [(3'h6):(1'h0)] reg2119 = (1'h0);
  reg [(4'h8):(1'h0)] reg2118 = (1'h0);
  reg [(3'h7):(1'h0)] reg2117 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2116 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2115 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2114 = (1'h0);
  reg [(4'hb):(1'h0)] reg2113 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2112 = (1'h0);
  reg [(4'ha):(1'h0)] reg2111 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2110 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2109 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2108 = (1'h0);
  reg [(4'hd):(1'h0)] reg2107 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2106 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2105 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2104 = (1'h0);
  reg [(4'he):(1'h0)] reg2103 = (1'h0);
  reg [(4'ha):(1'h0)] reg2102 = (1'h0);
  reg [(4'hb):(1'h0)] reg2101 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2100 = (1'h0);
  reg [(4'h8):(1'h0)] reg2099 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2098 = (1'h0);
  reg [(4'he):(1'h0)] reg2097 = (1'h0);
  reg [(3'h4):(1'h0)] reg2096 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2095 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2094 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2093 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2092 = (1'h0);
  reg [(4'hf):(1'h0)] reg2091 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2090 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2089 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2088 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2083 = (1'h0);
  reg [(4'he):(1'h0)] reg2078 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2080 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2076 = (1'h0);
  reg [(4'hd):(1'h0)] reg2069 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2087 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2086 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2085 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2084 = (1'h0);
  reg [(2'h2):(1'h0)] reg2083 = (1'h0);
  reg [(3'h5):(1'h0)] reg2082 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2081 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2080 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2079 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2078 = (1'h0);
  reg [(4'h9):(1'h0)] reg2077 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2076 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2075 = (1'h0);
  reg [(3'h4):(1'h0)] reg2074 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2073 = (1'h0);
  reg [(4'ha):(1'h0)] reg2072 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2071 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2070 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2069 = (1'h0);
  reg [(4'ha):(1'h0)] reg2068 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2067 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2065 = (1'h0);
  reg [(4'hc):(1'h0)] reg2066 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2065 = (1'h0);
  reg [(4'h9):(1'h0)] reg2064 = (1'h0);
  reg [(5'h10):(1'h0)] reg2059 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2063 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2062 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2061 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2060 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2059 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2049 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2048 = (1'h0);
  reg [(2'h2):(1'h0)] reg2058 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2057 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2056 = (1'h0);
  reg [(4'h9):(1'h0)] reg2055 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2054 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2053 = (1'h0);
  reg [(4'hb):(1'h0)] reg2052 = (1'h0);
  reg [(5'h10):(1'h0)] reg2051 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2050 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2049 = (1'h0);
  reg [(4'h9):(1'h0)] reg2048 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2047 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2043 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2041 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2047 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2046 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2045 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2044 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2043 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2040 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2042 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2041 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2040 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2039 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2038 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2037 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2036 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2035 = (1'h0);
  reg [(4'he):(1'h0)] forvar2034 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2033 = (1'h0);
  reg [(2'h3):(1'h0)] reg2032 = (1'h0);
  reg [(4'hb):(1'h0)] reg2031 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2030 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2029 = (1'h0);
  reg [(4'h9):(1'h0)] reg2028 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2027 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2026 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2025 = (1'h0);
  reg [(4'he):(1'h0)] forvar2024 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2023 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2022 = (1'h0);
  reg [(3'h4):(1'h0)] reg2021 = (1'h0);
  reg [(3'h5):(1'h0)] reg2020 = (1'h0);
  reg [(4'he):(1'h0)] reg2019 = (1'h0);
  reg [(4'he):(1'h0)] forvar2018 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2017 = (1'h0);
  reg [(2'h2):(1'h0)] reg2011 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2009 = (1'h0);
  reg [(4'he):(1'h0)] forvar2006 = (1'h0);
  reg [(4'he):(1'h0)] reg2016 = (1'h0);
  reg [(2'h3):(1'h0)] reg2015 = (1'h0);
  reg [(4'hd):(1'h0)] reg2014 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2013 = (1'h0);
  reg [(4'h9):(1'h0)] reg2012 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2011 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2010 = (1'h0);
  reg [(4'hb):(1'h0)] reg2009 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2008 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2007 = (1'h0);
  reg [(4'hb):(1'h0)] reg2006 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2005 = (1'h0);
  reg [(4'hb):(1'h0)] reg2004 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2003 = (1'h0);
  reg [(3'h4):(1'h0)] reg2002 = (1'h0);
  reg [(3'h7):(1'h0)] reg2001 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2000 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1999 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1998 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1997 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1996 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1995 = (1'h0);
  reg [(4'hc):(1'h0)] reg1994 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1993 = (1'h0);
  reg [(4'h8):(1'h0)] reg1992 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1991 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1990 = (1'h0);
  reg [(4'hc):(1'h0)] reg1975 = (1'h0);
  reg [(4'hd):(1'h0)] reg1989 = (1'h0);
  reg [(2'h3):(1'h0)] reg1988 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1987 = (1'h0);
  reg [(3'h4):(1'h0)] reg1986 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1985 = (1'h0);
  reg [(4'hb):(1'h0)] reg1984 = (1'h0);
  reg [(4'h8):(1'h0)] reg1983 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1982 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1981 = (1'h0);
  reg [(4'he):(1'h0)] forvar1980 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1979 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1978 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1977 = (1'h0);
  reg [(2'h2):(1'h0)] reg1976 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1975 = (1'h0);
  reg [(3'h7):(1'h0)] reg1974 = (1'h0);
  reg [(4'he):(1'h0)] reg1973 = (1'h0);
  reg [(3'h4):(1'h0)] reg1972 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1971 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1970 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1969 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1968 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1967 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1966 = (1'h0);
  reg [(4'he):(1'h0)] reg1948 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1945 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1965 = (1'h0);
  reg [(3'h6):(1'h0)] reg1964 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1963 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1958 = (1'h0);
  reg [(4'hd):(1'h0)] reg1955 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1962 = (1'h0);
  reg [(3'h7):(1'h0)] reg1961 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1960 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1959 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1958 = (1'h0);
  reg [(4'h9):(1'h0)] reg1957 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1956 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1955 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1954 = (1'h0);
  reg [(2'h2):(1'h0)] reg1953 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1952 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1951 = (1'h0);
  reg [(4'hc):(1'h0)] reg1950 = (1'h0);
  reg [(4'hb):(1'h0)] reg1949 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1948 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1944 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1941 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1940 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1939 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1937 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1947 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1946 = (1'h0);
  reg [(2'h3):(1'h0)] reg1945 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1944 = (1'h0);
  reg [(4'ha):(1'h0)] reg1943 = (1'h0);
  reg [(3'h6):(1'h0)] reg1942 = (1'h0);
  reg [(4'h8):(1'h0)] reg1941 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1940 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1939 = (1'h0);
  reg [(4'h9):(1'h0)] reg1938 = (1'h0);
  reg [(4'he):(1'h0)] reg1937 = (1'h0);
  reg [(5'h10):(1'h0)] reg1936 = (1'h0);
  reg [(2'h3):(1'h0)] reg1935 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1934 = (1'h0);
  reg [(3'h4):(1'h0)] reg1933 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1932 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1927 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1932 = (1'h0);
  reg [(2'h3):(1'h0)] reg1931 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1930 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1929 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1928 = (1'h0);
  reg [(4'ha):(1'h0)] reg1927 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1925 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1924 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1920 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1917 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1913 = (1'h0);
  reg [(2'h3):(1'h0)] reg1926 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1925 = (1'h0);
  reg [(3'h4):(1'h0)] reg1924 = (1'h0);
  reg [(3'h5):(1'h0)] reg1923 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1922 = (1'h0);
  reg [(4'hb):(1'h0)] reg1921 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1920 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1919 = (1'h0);
  reg [(4'he):(1'h0)] reg1918 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1917 = (1'h0);
  reg [(2'h3):(1'h0)] reg1916 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1914 = (1'h0);
  reg [(2'h2):(1'h0)] reg1915 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1914 = (1'h0);
  reg [(4'he):(1'h0)] reg1913 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1912 = (1'h0);
  reg [(4'he):(1'h0)] reg1907 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1906 = (1'h0);
  reg [(4'he):(1'h0)] reg1905 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1904 = (1'h0);
  reg [(4'h8):(1'h0)] reg1911 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1910 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1909 = (1'h0);
  reg [(4'hb):(1'h0)] reg1908 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1907 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1906 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1905 = (1'h0);
  reg [(4'hd):(1'h0)] reg1904 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1901 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1894 = (1'h0);
  reg [(4'ha):(1'h0)] reg1903 = (1'h0);
  reg [(2'h3):(1'h0)] reg1902 = (1'h0);
  reg [(5'h10):(1'h0)] reg1901 = (1'h0);
  reg [(3'h4):(1'h0)] reg1900 = (1'h0);
  reg [(4'hc):(1'h0)] reg1899 = (1'h0);
  reg [(2'h3):(1'h0)] reg1898 = (1'h0);
  reg [(4'ha):(1'h0)] reg1897 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1896 = (1'h0);
  reg [(4'ha):(1'h0)] reg1895 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1894 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1893 = (1'h0);
  reg [(3'h7):(1'h0)] reg1892 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1891 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1890 = (1'h0);
  reg [(3'h5):(1'h0)] reg1889 = (1'h0);
  reg [(3'h4):(1'h0)] reg1888 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1887 = (1'h0);
  reg [(3'h7):(1'h0)] reg1886 = (1'h0);
  reg [(2'h3):(1'h0)] reg1885 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1884 = (1'h0);
  reg [(5'h10):(1'h0)] reg1883 = (1'h0);
  reg [(2'h3):(1'h0)] reg1882 = (1'h0);
  reg [(4'hf):(1'h0)] reg1881 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1880 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1879 = (1'h0);
  reg [(4'hf):(1'h0)] reg1878 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1877 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1876 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1875 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1874 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1873 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1872 = (1'h0);
  reg [(4'hd):(1'h0)] reg1871 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1870 = (1'h0);
  reg [(4'he):(1'h0)] reg1869 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1868 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1867 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1866 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1865 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1864 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1863 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1862 = (1'h0);
  reg [(4'hc):(1'h0)] reg1861 = (1'h0);
  reg [(4'hc):(1'h0)] reg1860 = (1'h0);
  reg [(4'h9):(1'h0)] reg1859 = (1'h0);
  reg [(4'hd):(1'h0)] reg1858 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1857 = (1'h0);
  reg [(4'hb):(1'h0)] reg1856 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1855 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1854 = (1'h0);
  reg [(4'he):(1'h0)] reg1853 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1852 = (1'h0);
  reg [(3'h4):(1'h0)] reg1851 = (1'h0);
  reg [(3'h7):(1'h0)] reg1850 = (1'h0);
  reg [(4'hb):(1'h0)] reg1849 = (1'h0);
  reg [(4'h9):(1'h0)] reg1848 = (1'h0);
  reg [(3'h7):(1'h0)] reg1847 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1846 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1845 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1844 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1843 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1840 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1839 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1838 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1834 = (1'h0);
  reg [(3'h7):(1'h0)] reg1842 = (1'h0);
  reg [(3'h4):(1'h0)] reg1841 = (1'h0);
  reg [(4'h8):(1'h0)] reg1840 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1839 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1838 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1837 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1836 = (1'h0);
  reg [(4'h8):(1'h0)] reg1835 = (1'h0);
  reg [(4'he):(1'h0)] reg1834 = (1'h0);
  reg [(4'hc):(1'h0)] reg1833 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1832 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1831 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1830 = (1'h0);
  reg [(2'h2):(1'h0)] reg1811 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1809 = (1'h0);
  reg [(2'h2):(1'h0)] reg1807 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1806 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1805 = (1'h0);
  reg [(4'he):(1'h0)] forvar1803 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1801 = (1'h0);
  reg [(4'hb):(1'h0)] reg1797 = (1'h0);
  reg [(4'hd):(1'h0)] reg1802 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1799 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1789 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1783 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1775 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1780 = (1'h0);
  reg [(4'h9):(1'h0)] reg1829 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1828 = (1'h0);
  reg [(4'he):(1'h0)] reg1827 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1826 = (1'h0);
  reg [(2'h3):(1'h0)] reg1825 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1824 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1823 = (1'h0);
  reg [(3'h4):(1'h0)] reg1822 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1821 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1820 = (1'h0);
  reg [(4'h9):(1'h0)] reg1819 = (1'h0);
  reg [(2'h3):(1'h0)] reg1818 = (1'h0);
  reg [(4'hd):(1'h0)] reg1817 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1816 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1815 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1814 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1813 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1812 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1811 = (1'h0);
  reg [(4'hd):(1'h0)] reg1810 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1809 = (1'h0);
  reg [(4'hc):(1'h0)] reg1808 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1807 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1806 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1794 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1793 = (1'h0);
  reg [(4'h8):(1'h0)] reg1805 = (1'h0);
  reg [(3'h4):(1'h0)] reg1804 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1803 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1802 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1801 = (1'h0);
  reg [(4'hf):(1'h0)] reg1800 = (1'h0);
  reg [(2'h3):(1'h0)] reg1799 = (1'h0);
  reg [(4'hd):(1'h0)] reg1798 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1797 = (1'h0);
  reg [(4'h9):(1'h0)] reg1796 = (1'h0);
  reg [(3'h4):(1'h0)] reg1795 = (1'h0);
  reg [(5'h10):(1'h0)] reg1794 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1793 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1788 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1787 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1785 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1784 = (1'h0);
  reg [(4'h8):(1'h0)] reg1792 = (1'h0);
  reg [(2'h2):(1'h0)] reg1791 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1790 = (1'h0);
  reg [(5'h10):(1'h0)] reg1789 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1788 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1787 = (1'h0);
  reg [(3'h7):(1'h0)] reg1786 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1785 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1784 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1776 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1783 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1782 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1781 = (1'h0);
  reg [(2'h3):(1'h0)] reg1780 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1779 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1778 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1777 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1776 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1775 = (1'h0);
  wire [(2'h2):(1'h0)] wire1774;
  wire [(3'h7):(1'h0)] wire1773;
  wire [(3'h5):(1'h0)] wire1772;
  wire signed [(4'h8):(1'h0)] wire1771;
  wire [(4'hc):(1'h0)] wire1770;
  wire [(4'ha):(1'h0)] wire1769;
  assign y = {wire2747,
                 wire2746,
                 reg2745,
                 reg2744,
                 reg2743,
                 reg2742,
                 reg2741,
                 reg2740,
                 reg2739,
                 reg2738,
                 reg2737,
                 forvar2736,
                 reg2735,
                 forvar2734,
                 reg2733,
                 reg2732,
                 reg2731,
                 forvar2730,
                 reg2729,
                 reg2728,
                 reg2727,
                 reg2726,
                 reg2725,
                 reg2724,
                 reg2723,
                 reg2722,
                 reg2721,
                 forvar2720,
                 reg2719,
                 reg2718,
                 reg2717,
                 reg2716,
                 forvar2715,
                 reg2714,
                 reg2713,
                 reg2712,
                 reg2711,
                 reg2710,
                 reg2709,
                 forvar2708,
                 reg2707,
                 forvar2706,
                 forvar2705,
                 forvar2680,
                 forvar2677,
                 forvar2674,
                 forvar2672,
                 forvar2669,
                 forvar2667,
                 reg2665,
                 reg2693,
                 reg2704,
                 forvar2703,
                 reg2702,
                 reg2701,
                 reg2700,
                 forvar2699,
                 reg2698,
                 reg2697,
                 reg2696,
                 forvar2695,
                 reg2694,
                 forvar2693,
                 reg2676,
                 forvar2675,
                 reg2673,
                 reg2668,
                 reg2666,
                 reg2692,
                 reg2691,
                 reg2690,
                 reg2689,
                 forvar2688,
                 reg2687,
                 reg2686,
                 reg2685,
                 reg2684,
                 forvar2683,
                 reg2682,
                 reg2681,
                 reg2680,
                 reg2679,
                 reg2678,
                 reg2677,
                 forvar2676,
                 reg2675,
                 reg2674,
                 forvar2673,
                 reg2672,
                 reg2671,
                 reg2670,
                 reg2669,
                 forvar2668,
                 reg2667,
                 forvar2666,
                 forvar2665,
                 reg2664,
                 reg2659,
                 reg2663,
                 reg2662,
                 reg2661,
                 reg2660,
                 forvar2659,
                 reg2650,
                 forvar2649,
                 reg2658,
                 reg2657,
                 reg2656,
                 forvar2655,
                 reg2654,
                 reg2653,
                 reg2652,
                 reg2651,
                 forvar2650,
                 reg2649,
                 reg2648,
                 reg2647,
                 forvar2646,
                 forvar2645,
                 reg2644,
                 reg2643,
                 reg2642,
                 reg2641,
                 forvar2640,
                 reg2639,
                 forvar2632,
                 forvar2630,
                 reg2638,
                 reg2637,
                 reg2636,
                 reg2631,
                 reg2629,
                 forvar2627,
                 reg2626,
                 reg2635,
                 reg2634,
                 reg2633,
                 reg2632,
                 forvar2631,
                 reg2630,
                 forvar2629,
                 reg2628,
                 reg2627,
                 forvar2626,
                 reg2625,
                 forvar2624,
                 reg2623,
                 reg2622,
                 reg2621,
                 reg2620,
                 reg2619,
                 reg2618,
                 reg2617,
                 reg2616,
                 reg2615,
                 forvar2614,
                 reg2613,
                 forvar2612,
                 forvar2611,
                 forvar2610,
                 reg2609,
                 reg2608,
                 reg2607,
                 reg2606,
                 reg2605,
                 reg2604,
                 reg2603,
                 reg2602,
                 reg2601,
                 forvar2600,
                 reg2599,
                 reg2598,
                 reg2597,
                 forvar2596,
                 forvar2595,
                 reg2594,
                 reg2593,
                 reg2592,
                 reg2591,
                 forvar2590,
                 reg2588,
                 reg2590,
                 reg2589,
                 forvar2588,
                 forvar2587,
                 forvar2586,
                 wire2585,
                 wire2584,
                 wire2582,
                 wire2121,
                 wire2120,
                 reg2088,
                 reg2119,
                 reg2118,
                 reg2117,
                 reg2116,
                 reg2115,
                 forvar2114,
                 reg2113,
                 reg2112,
                 reg2111,
                 reg2110,
                 forvar2109,
                 reg2108,
                 reg2107,
                 reg2106,
                 reg2105,
                 forvar2104,
                 reg2103,
                 reg2102,
                 reg2101,
                 forvar2100,
                 reg2099,
                 reg2098,
                 reg2097,
                 reg2096,
                 reg2095,
                 reg2094,
                 reg2093,
                 reg2092,
                 reg2091,
                 reg2090,
                 forvar2089,
                 forvar2088,
                 forvar2083,
                 reg2078,
                 reg2080,
                 forvar2076,
                 reg2069,
                 reg2087,
                 reg2086,
                 reg2085,
                 reg2084,
                 reg2083,
                 reg2082,
                 reg2081,
                 forvar2080,
                 reg2079,
                 forvar2078,
                 reg2077,
                 reg2076,
                 reg2075,
                 reg2074,
                 reg2073,
                 reg2072,
                 reg2071,
                 forvar2070,
                 forvar2069,
                 reg2068,
                 reg2067,
                 forvar2065,
                 reg2066,
                 reg2065,
                 reg2064,
                 reg2059,
                 reg2063,
                 forvar2062,
                 reg2061,
                 reg2060,
                 forvar2059,
                 reg2049,
                 forvar2048,
                 reg2058,
                 forvar2057,
                 reg2056,
                 reg2055,
                 reg2054,
                 reg2053,
                 reg2052,
                 reg2051,
                 reg2050,
                 forvar2049,
                 reg2048,
                 forvar2047,
                 forvar2043,
                 forvar2041,
                 reg2047,
                 reg2046,
                 reg2045,
                 reg2044,
                 reg2043,
                 forvar2040,
                 reg2042,
                 reg2041,
                 reg2040,
                 forvar2039,
                 reg2038,
                 reg2037,
                 reg2036,
                 reg2035,
                 forvar2034,
                 reg2033,
                 reg2032,
                 reg2031,
                 reg2030,
                 forvar2029,
                 reg2028,
                 reg2027,
                 reg2026,
                 reg2025,
                 forvar2024,
                 forvar2023,
                 forvar2022,
                 reg2021,
                 reg2020,
                 reg2019,
                 forvar2018,
                 forvar2017,
                 reg2011,
                 forvar2009,
                 forvar2006,
                 reg2016,
                 reg2015,
                 reg2014,
                 reg2013,
                 reg2012,
                 forvar2011,
                 reg2010,
                 reg2009,
                 reg2008,
                 reg2007,
                 reg2006,
                 reg2005,
                 reg2004,
                 reg2003,
                 reg2002,
                 reg2001,
                 forvar2000,
                 reg1999,
                 forvar1998,
                 forvar1997,
                 forvar1996,
                 reg1995,
                 reg1994,
                 reg1993,
                 reg1992,
                 forvar1991,
                 forvar1990,
                 reg1975,
                 reg1989,
                 reg1988,
                 reg1987,
                 reg1986,
                 reg1985,
                 reg1984,
                 reg1983,
                 reg1982,
                 reg1981,
                 forvar1980,
                 reg1979,
                 reg1978,
                 reg1977,
                 reg1976,
                 forvar1975,
                 reg1974,
                 reg1973,
                 reg1972,
                 reg1971,
                 reg1970,
                 forvar1969,
                 forvar1968,
                 forvar1967,
                 reg1966,
                 reg1948,
                 forvar1945,
                 reg1965,
                 reg1964,
                 forvar1963,
                 forvar1958,
                 reg1955,
                 reg1962,
                 reg1961,
                 reg1960,
                 reg1959,
                 reg1958,
                 reg1957,
                 reg1956,
                 forvar1955,
                 reg1954,
                 reg1953,
                 reg1952,
                 reg1951,
                 reg1950,
                 reg1949,
                 forvar1948,
                 reg1944,
                 forvar1941,
                 reg1940,
                 forvar1939,
                 forvar1937,
                 reg1947,
                 reg1946,
                 reg1945,
                 forvar1944,
                 reg1943,
                 reg1942,
                 reg1941,
                 forvar1940,
                 reg1939,
                 reg1938,
                 reg1937,
                 reg1936,
                 reg1935,
                 reg1934,
                 reg1933,
                 forvar1932,
                 forvar1927,
                 reg1932,
                 reg1931,
                 forvar1930,
                 reg1929,
                 reg1928,
                 reg1927,
                 reg1925,
                 forvar1924,
                 reg1920,
                 forvar1917,
                 forvar1913,
                 reg1926,
                 forvar1925,
                 reg1924,
                 reg1923,
                 forvar1922,
                 reg1921,
                 forvar1920,
                 reg1919,
                 reg1918,
                 reg1917,
                 reg1916,
                 reg1914,
                 reg1915,
                 forvar1914,
                 reg1913,
                 forvar1912,
                 reg1907,
                 forvar1906,
                 reg1905,
                 forvar1904,
                 reg1911,
                 reg1910,
                 reg1909,
                 reg1908,
                 forvar1907,
                 reg1906,
                 forvar1905,
                 reg1904,
                 forvar1901,
                 forvar1894,
                 reg1903,
                 reg1902,
                 reg1901,
                 reg1900,
                 reg1899,
                 reg1898,
                 reg1897,
                 forvar1896,
                 reg1895,
                 reg1894,
                 reg1893,
                 reg1892,
                 reg1891,
                 reg1890,
                 reg1889,
                 reg1888,
                 forvar1887,
                 reg1886,
                 reg1885,
                 forvar1884,
                 reg1883,
                 reg1882,
                 reg1881,
                 reg1880,
                 reg1879,
                 reg1878,
                 reg1877,
                 forvar1876,
                 forvar1875,
                 forvar1874,
                 reg1873,
                 reg1872,
                 reg1871,
                 forvar1870,
                 reg1869,
                 reg1868,
                 forvar1867,
                 forvar1866,
                 reg1865,
                 reg1864,
                 reg1863,
                 reg1862,
                 reg1861,
                 reg1860,
                 reg1859,
                 reg1858,
                 forvar1857,
                 reg1856,
                 reg1855,
                 reg1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 reg1850,
                 reg1849,
                 reg1848,
                 reg1847,
                 reg1846,
                 forvar1845,
                 reg1844,
                 reg1843,
                 forvar1840,
                 forvar1839,
                 reg1838,
                 forvar1834,
                 reg1842,
                 reg1841,
                 reg1840,
                 reg1839,
                 forvar1838,
                 reg1837,
                 reg1836,
                 reg1835,
                 reg1834,
                 reg1833,
                 forvar1832,
                 forvar1831,
                 forvar1830,
                 reg1811,
                 forvar1809,
                 reg1807,
                 reg1806,
                 forvar1805,
                 forvar1803,
                 forvar1801,
                 reg1797,
                 reg1802,
                 forvar1799,
                 forvar1789,
                 forvar1783,
                 reg1775,
                 forvar1780,
                 reg1829,
                 reg1828,
                 reg1827,
                 reg1826,
                 reg1825,
                 forvar1824,
                 reg1823,
                 reg1822,
                 forvar1821,
                 forvar1820,
                 reg1819,
                 reg1818,
                 reg1817,
                 reg1816,
                 reg1815,
                 reg1814,
                 reg1813,
                 reg1812,
                 forvar1811,
                 reg1810,
                 reg1809,
                 reg1808,
                 forvar1807,
                 forvar1806,
                 forvar1794,
                 reg1793,
                 reg1805,
                 reg1804,
                 reg1803,
                 forvar1802,
                 reg1801,
                 reg1800,
                 reg1799,
                 reg1798,
                 forvar1797,
                 reg1796,
                 reg1795,
                 reg1794,
                 forvar1793,
                 forvar1788,
                 reg1787,
                 forvar1785,
                 reg1784,
                 reg1792,
                 reg1791,
                 reg1790,
                 reg1789,
                 reg1788,
                 forvar1787,
                 reg1786,
                 reg1785,
                 forvar1784,
                 reg1776,
                 reg1783,
                 reg1782,
                 reg1781,
                 reg1780,
                 reg1779,
                 reg1778,
                 reg1777,
                 forvar1776,
                 forvar1775,
                 wire1774,
                 wire1773,
                 wire1772,
                 wire1771,
                 wire1770,
                 wire1769,
                 (1'h0)};
  assign wire1769 = (8'h9f);
  assign wire1770 = wire1769;
  assign wire1771 = (wire1769 >>> ($unsigned(wire1767) < wire1768[(3'h6):(3'h5)]));
  assign wire1772 = wire1769[(3'h7):(3'h5)];
  assign wire1773 = $unsigned(wire1768[(4'hb):(1'h0)]);
  assign wire1774 = (({(wire1770 + wire1767)} >>> {(wire1765 ?
                            wire1768 : wire1769)}) ^~ (-((wire1766 * wire1768) && {wire1765})));
  always
    @(posedge clk) begin
      if (((+wire1774[(1'h1):(1'h1)]) || (wire1774 ?
          (wire1774 == (wire1770 ? wire1770 : wire1766)) : $unsigned((wire1773 ?
              (8'ha5) : wire1765)))))
        begin
          for (forvar1775 = (1'h0); (forvar1775 < (1'h0)); forvar1775 = (forvar1775 + (1'h1)))
            begin
              if ((!wire1769[(4'h9):(3'h7)]))
                begin
                  for (forvar1776 = (1'h0); (forvar1776 < (2'h2)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 <= wire1765;
                    end
                  if (($signed(((wire1772 ? wire1772 : wire1772) ?
                          (reg1777 ? reg1777 : wire1772) : (!(8'hb8)))) ?
                      {wire1770} : wire1769[(4'ha):(4'h9)]))
                    begin
                      reg1778 <= ($signed(wire1771[(3'h6):(1'h0)]) - $unsigned($signed(wire1769)));
                      reg1779 <= $signed(wire1771[(1'h1):(1'h1)]);
                      reg1780 <= ({$signed((-wire1774))} >>> $signed(wire1772));
                      reg1781 <= forvar1775;
                    end
                  else
                    begin
                      reg1778 <= (^~wire1774);
                      reg1779 <= {($unsigned(wire1773) + $unsigned({(8'ha7)}))};
                    end
                  if ((wire1771[(2'h2):(1'h0)] ?
                      (^$unsigned(((8'haf) ?
                          wire1774 : wire1770))) : (((|forvar1775) ?
                              (^~wire1766) : wire1769[(1'h0):(1'h0)]) ?
                          wire1774[(1'h1):(1'h0)] : wire1772)))
                    begin
                      reg1782 <= ((8'hb3) ?
                          $signed($signed($unsigned(reg1779))) : wire1773[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1782 <= wire1774[(1'h1):(1'h1)];
                    end
                  reg1783 <= wire1774;
                end
              else
                begin
                  if (wire1770)
                    begin
                      reg1776 <= (reg1781 ?
                          wire1771 : ($unsigned($unsigned(reg1783)) << wire1774[(2'h2):(1'h1)]));
                      reg1777 <= (~{reg1777});
                      reg1778 <= (~&$signed(reg1783));
                      reg1779 <= wire1773;
                    end
                  else
                    begin
                      reg1776 <= {{(8'hae)}};
                      reg1777 <= (|$unsigned($signed((wire1767 ?
                          reg1783 : (8'hb3)))));
                      reg1778 <= $signed((reg1781 ?
                          ($signed(wire1770) ?
                              {wire1771} : (wire1767 ?
                                  reg1781 : wire1765)) : $signed(wire1768[(2'h3):(2'h2)])));
                    end
                  if ($unsigned((+$unsigned((wire1770 & wire1772)))))
                    begin
                      reg1780 <= ((-(wire1770 ?
                          $signed(forvar1775) : ((8'ha5) != wire1774))) <<< (8'hb7));
                      reg1781 <= ($unsigned((~&(forvar1775 >> wire1765))) ?
                          $unsigned((((8'hba) ? wire1767 : reg1781) ?
                              (wire1772 != (8'hb1)) : (reg1776 != reg1776))) : forvar1775[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg1780 <= $unsigned(wire1767[(1'h0):(1'h0)]);
                    end
                end
              if (((reg1776[(3'h5):(3'h5)] ?
                      ((wire1771 & (8'hb4)) ^~ (^~wire1767)) : $signed((wire1768 ?
                          wire1774 : wire1768))) ?
                  $unsigned($unsigned((wire1767 <= wire1770))) : (8'ha0)))
                begin
                  for (forvar1784 = (1'h0); (forvar1784 < (1'h0)); forvar1784 = (forvar1784 + (1'h1)))
                    begin
                      reg1785 <= {$unsigned({(+wire1774)})};
                    end
                  reg1786 <= ((8'had) != (~&$unsigned(wire1771[(1'h1):(1'h1)])));
                  for (forvar1787 = (1'h0); (forvar1787 < (1'h0)); forvar1787 = (forvar1787 + (1'h1)))
                    begin
                      reg1788 <= $unsigned(($unsigned(wire1774[(2'h2):(2'h2)]) ?
                          ($signed(forvar1784) ~^ (forvar1784 ?
                              reg1786 : forvar1775)) : {(wire1767 ?
                                  wire1767 : wire1765)}));
                      reg1789 <= {wire1772};
                    end
                  if (((&wire1767[(2'h2):(1'h0)]) >> ($signed(reg1777[(4'hb):(3'h6)]) ?
                      reg1776 : ((wire1768 ?
                          wire1768 : reg1780) && reg1780[(2'h3):(1'h1)]))))
                    begin
                      reg1790 <= {$unsigned(wire1771[(3'h5):(3'h4)])};
                    end
                  else
                    begin
                      reg1790 <= ($signed($unsigned((forvar1776 || wire1765))) ?
                          $signed($signed(wire1773[(3'h6):(1'h1)])) : $unsigned($unsigned((forvar1776 | reg1780))));
                      reg1791 <= ($signed(((|wire1765) <= wire1767[(2'h2):(1'h1)])) ?
                          $unsigned({(forvar1787 ?
                                  reg1782 : forvar1784)}) : $unsigned($unsigned((8'hb5))));
                      reg1792 <= ($signed($unsigned({reg1783})) ?
                          (!$signed(reg1779[(3'h7):(3'h6)])) : (8'hb8));
                    end
                end
              else
                begin
                  reg1784 <= {{$signed((8'ha6))}};
                  for (forvar1785 = (1'h0); (forvar1785 < (1'h0)); forvar1785 = (forvar1785 + (1'h1)))
                    begin
                      reg1786 <= reg1785[(2'h2):(2'h2)];
                      reg1787 <= reg1788[(1'h1):(1'h1)];
                    end
                  for (forvar1788 = (1'h0); (forvar1788 < (2'h3)); forvar1788 = (forvar1788 + (1'h1)))
                    begin
                      reg1789 <= ((wire1768 ?
                              $signed($unsigned(reg1785)) : $unsigned(wire1765)) ?
                          ({$unsigned(reg1785)} ?
                              $signed((~&wire1769)) : reg1785[(2'h3):(2'h3)]) : $unsigned(wire1773));
                      reg1790 <= wire1773;
                    end
                end
              if ((({(reg1782 * (8'hab))} ?
                  wire1772 : $unsigned((!reg1790))) > $signed((8'hb7))))
                begin
                  for (forvar1793 = (1'h0); (forvar1793 < (2'h3)); forvar1793 = (forvar1793 + (1'h1)))
                    begin
                      reg1794 <= (~|$signed(reg1786));
                      reg1795 <= {(reg1781[(3'h5):(2'h2)] != wire1766)};
                      reg1796 <= $signed({($unsigned(wire1765) ~^ $unsigned(wire1772))});
                    end
                  for (forvar1797 = (1'h0); (forvar1797 < (1'h0)); forvar1797 = (forvar1797 + (1'h1)))
                    begin
                      reg1798 <= (reg1782[(1'h0):(1'h0)] <= ({$signed(wire1771)} >= reg1783));
                      reg1799 <= reg1786;
                      reg1800 <= ({{{forvar1775}}} ?
                          $signed(($signed((8'hb6)) >= $unsigned(reg1799))) : (^~$unsigned($unsigned((8'hae)))));
                      reg1801 <= wire1769[(3'h5):(1'h0)];
                    end
                  for (forvar1802 = (1'h0); (forvar1802 < (1'h1)); forvar1802 = (forvar1802 + (1'h1)))
                    begin
                      reg1803 <= $unsigned(((&(&(8'had))) ?
                          (wire1770[(4'h8):(1'h1)] <<< $signed((8'ha4))) : forvar1787[(2'h2):(1'h0)]));
                      reg1804 <= (^forvar1785[(1'h0):(1'h0)]);
                      reg1805 <= wire1765;
                    end
                end
              else
                begin
                  reg1793 <= (-($signed(((8'ha7) == forvar1785)) - ($unsigned(reg1781) >> (~forvar1793))));
                  for (forvar1794 = (1'h0); (forvar1794 < (2'h3)); forvar1794 = (forvar1794 + (1'h1)))
                    begin
                      reg1795 <= forvar1776;
                    end
                end
              for (forvar1806 = (1'h0); (forvar1806 < (1'h0)); forvar1806 = (forvar1806 + (1'h1)))
                begin
                  for (forvar1807 = (1'h0); (forvar1807 < (1'h0)); forvar1807 = (forvar1807 + (1'h1)))
                    begin
                      reg1808 <= ($signed(reg1804) ?
                          {(|reg1787[(2'h3):(2'h3)])} : ((~^reg1785) * ($signed(reg1777) ?
                              (wire1768 ? (8'ha6) : reg1804) : forvar1797)));
                      reg1809 <= {$signed({$unsigned(reg1800)})};
                    end
                  reg1810 <= $unsigned($unsigned(reg1794[(1'h0):(1'h0)]));
                  for (forvar1811 = (1'h0); (forvar1811 < (1'h1)); forvar1811 = (forvar1811 + (1'h1)))
                    begin
                      reg1812 <= (-$unsigned(reg1778[(2'h3):(2'h3)]));
                      reg1813 <= ({(&reg1799[(2'h3):(2'h2)])} ^ ($signed((8'ha4)) >>> reg1789));
                      reg1814 <= (wire1774[(1'h1):(1'h1)] ?
                          (({reg1799} ?
                                  {(8'h9c)} : (reg1801 ? reg1792 : (8'hb1))) ?
                              {{forvar1793}} : reg1791[(1'h0):(1'h0)]) : (8'ha8));
                      reg1815 <= $signed({{$unsigned(reg1791)}});
                    end
                  if ((reg1796[(1'h0):(1'h0)] ?
                      (+(forvar1785[(2'h2):(1'h1)] && (~&reg1809))) : {wire1767[(4'h9):(1'h1)]}))
                    begin
                      reg1816 <= reg1814;
                    end
                  else
                    begin
                      reg1816 <= wire1766[(1'h1):(1'h1)];
                      reg1817 <= (reg1799[(1'h1):(1'h0)] ?
                          (!reg1776[(4'ha):(2'h2)]) : ($signed((wire1772 ~^ reg1791)) ^ $unsigned(forvar1785[(2'h2):(1'h1)])));
                      reg1818 <= {{(^(^~reg1799))}};
                      reg1819 <= reg1808;
                    end
                end
            end
          for (forvar1820 = (1'h0); (forvar1820 < (1'h0)); forvar1820 = (forvar1820 + (1'h1)))
            begin
              for (forvar1821 = (1'h0); (forvar1821 < (2'h3)); forvar1821 = (forvar1821 + (1'h1)))
                begin
                  if (forvar1793)
                    begin
                      reg1822 <= reg1803[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg1822 <= (~^$unsigned(((reg1787 ? reg1787 : (8'ha6)) ?
                          (reg1800 ?
                              reg1801 : forvar1811) : (reg1822 + (8'hba)))));
                      reg1823 <= reg1800[(4'hf):(3'h5)];
                    end
                  for (forvar1824 = (1'h0); (forvar1824 < (1'h1)); forvar1824 = (forvar1824 + (1'h1)))
                    begin
                      reg1825 <= reg1799;
                      reg1826 <= reg1796;
                    end
                  if ($signed(({(wire1773 ?
                          wire1768 : wire1769)} && $unsigned(reg1790))))
                    begin
                      reg1827 <= {(~$unsigned($unsigned(forvar1821)))};
                      reg1828 <= $signed(reg1799);
                      reg1829 <= ((-reg1813) ?
                          $signed({{reg1795}}) : ({{reg1786}} || $unsigned($signed(reg1800))));
                    end
                  else
                    begin
                      reg1827 <= {{(-{(8'ha1)})}};
                    end
                end
            end
        end
      else
        begin
          if ((wire1770[(3'h5):(3'h5)] ?
              ((reg1816[(4'h9):(3'h6)] != {reg1794}) ?
                  ((wire1774 - forvar1784) ?
                      (wire1768 >>> wire1773) : wire1766[(4'h9):(1'h0)]) : (^~(reg1794 ?
                      forvar1820 : wire1766))) : $signed(forvar1806[(4'hc):(4'hb)])))
            begin
              for (forvar1775 = (1'h0); (forvar1775 < (1'h0)); forvar1775 = (forvar1775 + (1'h1)))
                begin
                  reg1776 <= (~&($unsigned($unsigned(forvar1788)) ?
                      $unsigned(reg1808[(4'ha):(3'h7)]) : (reg1798 == (wire1772 + reg1780))));
                end
              if ((+(-{(|forvar1775)})))
                begin
                  if ((~(reg1788[(3'h7):(3'h4)] * {(!reg1818)})))
                    begin
                      reg1777 <= ({reg1799[(2'h2):(2'h2)]} ^~ $unsigned($unsigned(reg1826)));
                      reg1778 <= reg1787[(3'h5):(1'h1)];
                      reg1779 <= reg1785;
                      reg1780 <= reg1785[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg1777 <= forvar1775;
                      reg1778 <= $signed((~|{{reg1776}}));
                    end
                  if ($unsigned(($unsigned(((8'hb0) ?
                      forvar1807 : (8'h9d))) <<< ((reg1817 ?
                          forvar1794 : (8'hb7)) ?
                      {reg1780} : $unsigned(forvar1802)))))
                    begin
                      reg1781 <= ((reg1823 ? (+{reg1810}) : {(8'hb0)}) ?
                          reg1808[(4'h8):(3'h4)] : $signed(reg1794));
                      reg1782 <= $signed($unsigned(reg1818));
                    end
                  else
                    begin
                      reg1781 <= forvar1776[(3'h6):(3'h6)];
                      reg1782 <= $signed($signed($signed(reg1827[(3'h4):(3'h4)])));
                    end
                  if ($signed(($signed(forvar1793[(3'h4):(1'h1)]) ?
                      ((reg1792 ? forvar1785 : reg1788) ?
                          (reg1816 != reg1800) : (reg1784 < reg1817)) : {(wire1772 | reg1788)})))
                    begin
                      reg1783 <= ($signed($signed(((8'hb6) < reg1819))) ?
                          $unsigned((^(forvar1787 ?
                              (8'had) : reg1794))) : ($signed((~|reg1782)) ?
                              ($unsigned(reg1817) >>> {reg1809}) : $signed((reg1808 ?
                                  reg1813 : forvar1793))));
                    end
                  else
                    begin
                      reg1783 <= (((^$unsigned(wire1771)) ?
                              reg1808 : (^reg1778[(3'h5):(2'h3)])) ?
                          $unsigned((^~(8'hb0))) : reg1808);
                      reg1784 <= forvar1821[(2'h3):(2'h3)];
                      reg1785 <= ($signed($signed((!reg1787))) >> $signed((+$signed(reg1819))));
                      reg1786 <= forvar1784;
                    end
                  for (forvar1787 = (1'h0); (forvar1787 < (1'h1)); forvar1787 = (forvar1787 + (1'h1)))
                    begin
                      reg1788 <= (^~(wire1767 ?
                          reg1814[(1'h0):(1'h0)] : reg1793));
                      reg1789 <= (^reg1784);
                      reg1790 <= (~reg1778[(2'h2):(2'h2)]);
                      reg1791 <= reg1810;
                    end
                end
              else
                begin
                  if (reg1783[(3'h4):(3'h4)])
                    begin
                      reg1777 <= reg1803[(1'h1):(1'h0)];
                      reg1778 <= $unsigned((8'hac));
                      reg1779 <= reg1790[(3'h4):(2'h2)];
                    end
                  else
                    begin
                      reg1777 <= ({reg1795[(2'h3):(1'h1)]} || $unsigned(reg1799));
                      reg1778 <= ((^$unsigned((+forvar1787))) <= $signed(reg1816));
                    end
                  for (forvar1780 = (1'h0); (forvar1780 < (1'h1)); forvar1780 = (forvar1780 + (1'h1)))
                    begin
                      reg1781 <= wire1774[(2'h2):(1'h0)];
                      reg1782 <= $signed({$signed((wire1773 ?
                              wire1767 : (8'haa)))});
                      reg1783 <= $unsigned((|$unsigned(((8'hb4) + forvar1793))));
                    end
                end
            end
          else
            begin
              if ((({(wire1774 & reg1805)} ?
                      reg1776[(2'h3):(1'h1)] : {$unsigned(reg1825)}) ?
                  wire1769[(2'h3):(1'h0)] : reg1819))
                begin
                  if (((forvar1797[(3'h6):(1'h0)] ^ $signed($signed((8'haf)))) ?
                      wire1772[(3'h4):(1'h1)] : (~(!reg1789[(4'he):(2'h3)]))))
                    begin
                      reg1775 <= (^~{(~^$signed(reg1825))});
                      reg1776 <= wire1774[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg1775 <= (reg1788[(1'h0):(1'h0)] ?
                          (8'hae) : (reg1829 ?
                              (^$signed(reg1784)) : forvar1802));
                      reg1776 <= (+$unsigned($signed((reg1817 == reg1782))));
                      reg1777 <= (^($unsigned($unsigned((8'ha1))) ?
                          $unsigned({forvar1775}) : reg1825));
                    end
                end
              else
                begin
                  reg1775 <= $signed((~|((reg1788 ?
                      reg1777 : reg1803) + (forvar1780 < reg1778))));
                  if ($unsigned({((reg1809 <<< reg1816) >= $unsigned(reg1827))}))
                    begin
                      reg1776 <= (reg1812 ?
                          $signed((reg1825 <= $unsigned(reg1779))) : wire1768[(4'hb):(3'h4)]);
                      reg1777 <= forvar1775[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1776 <= forvar1811;
                    end
                  if ((&$signed($signed(wire1773[(2'h2):(1'h0)]))))
                    begin
                      reg1778 <= $unsigned($unsigned((~reg1776)));
                      reg1779 <= $signed($signed(({reg1785} != $signed(reg1786))));
                    end
                  else
                    begin
                      reg1778 <= (($unsigned($signed(forvar1802)) == (forvar1806[(4'hf):(4'ha)] >= $signed(reg1792))) ?
                          reg1823[(2'h2):(2'h2)] : reg1827);
                      reg1779 <= $signed($unsigned((reg1786 ?
                          $unsigned(reg1819) : (reg1799 || reg1819))));
                      reg1780 <= ((reg1812[(2'h2):(1'h1)] ?
                          $unsigned((~&reg1828)) : (~$signed(reg1782))) == forvar1811[(3'h6):(3'h5)]);
                    end
                  reg1781 <= $signed(reg1828);
                end
              if (((8'hb4) < $signed((8'ha6))))
                begin
                  reg1782 <= {{$unsigned((-reg1794))}};
                  for (forvar1783 = (1'h0); (forvar1783 < (2'h3)); forvar1783 = (forvar1783 + (1'h1)))
                    begin
                      reg1784 <= (+reg1775);
                      reg1785 <= $signed({$unsigned((reg1784 ?
                              forvar1793 : forvar1820))});
                    end
                end
              else
                begin
                  if ((8'hb0))
                    begin
                      reg1782 <= ({($signed(reg1793) ?
                                  {reg1826} : $signed(reg1783))} ?
                          $signed(reg1822) : forvar1785);
                    end
                  else
                    begin
                      reg1782 <= ((($signed(reg1819) ?
                              (reg1800 ? (8'hb2) : reg1815) : {forvar1811}) ?
                          wire1773 : ((reg1822 | reg1816) ?
                              $signed(forvar1793) : $signed(reg1794))) | ($unsigned($unsigned(forvar1802)) ?
                          ((forvar1807 ~^ (8'ha9)) ?
                              (|reg1776) : (reg1785 | (8'hae))) : ($unsigned(reg1790) | $signed((8'haa)))));
                      reg1783 <= ((~&(~&((8'hba) >> reg1775))) >>> $signed(({reg1784} ?
                          wire1767[(2'h2):(1'h0)] : $unsigned(reg1799))));
                      reg1784 <= reg1785;
                      reg1785 <= $signed((((forvar1784 ~^ wire1768) + (wire1774 < reg1810)) ?
                          reg1788[(3'h6):(2'h2)] : $signed((|(8'haf)))));
                    end
                  if (reg1786)
                    begin
                      reg1786 <= (~^reg1825);
                      reg1787 <= $unsigned({$unsigned(wire1774)});
                      reg1788 <= ($unsigned((~&reg1777)) ?
                          $signed((^~(reg1793 >= reg1816))) : {wire1766});
                    end
                  else
                    begin
                      reg1786 <= (&reg1826);
                      reg1787 <= reg1809;
                    end
                  for (forvar1789 = (1'h0); (forvar1789 < (2'h3)); forvar1789 = (forvar1789 + (1'h1)))
                    begin
                      reg1790 <= {reg1779};
                      reg1791 <= (!((!reg1795[(1'h0):(1'h0)]) + (8'hba)));
                    end
                  reg1792 <= ($unsigned(reg1829) * $signed((reg1826[(3'h4):(1'h1)] ?
                      reg1790[(2'h3):(2'h3)] : $unsigned(forvar1824))));
                end
            end
          if ((8'hb7))
            begin
              for (forvar1793 = (1'h0); (forvar1793 < (1'h1)); forvar1793 = (forvar1793 + (1'h1)))
                begin
                  for (forvar1794 = (1'h0); (forvar1794 < (2'h3)); forvar1794 = (forvar1794 + (1'h1)))
                    begin
                      reg1795 <= (($unsigned((reg1798 ? reg1823 : reg1813)) ?
                              $signed(forvar1806) : $unsigned(forvar1788)) ?
                          wire1773[(3'h5):(3'h4)] : ($signed((-wire1773)) & (wire1767 ~^ forvar1780)));
                      reg1796 <= (&(reg1785[(3'h5):(2'h2)] ~^ $unsigned(wire1768)));
                    end
                end
              for (forvar1797 = (1'h0); (forvar1797 < (1'h1)); forvar1797 = (forvar1797 + (1'h1)))
                begin
                  reg1798 <= (~|(8'hb8));
                  for (forvar1799 = (1'h0); (forvar1799 < (1'h0)); forvar1799 = (forvar1799 + (1'h1)))
                    begin
                      reg1800 <= forvar1824[(1'h0):(1'h0)];
                      reg1801 <= (reg1794 ?
                          $signed($signed(forvar1793[(2'h3):(2'h2)])) : $unsigned($unsigned(forvar1789[(4'hb):(3'h6)])));
                      reg1802 <= ((~&{(forvar1785 ?
                              (8'ha2) : reg1817)}) >= reg1829);
                      reg1803 <= forvar1784[(4'hf):(2'h2)];
                    end
                end
            end
          else
            begin
              if (reg1775)
                begin
                  if ($signed((~|reg1788)))
                    begin
                      reg1793 <= (~^forvar1811[(1'h0):(1'h0)]);
                      reg1794 <= $unsigned(reg1810);
                    end
                  else
                    begin
                      reg1793 <= forvar1780[(1'h0):(1'h0)];
                    end
                  if (((forvar1785[(2'h2):(1'h0)] ?
                          ($unsigned(reg1781) + (^(8'h9f))) : $unsigned((reg1822 ?
                              reg1785 : (8'hb7)))) ?
                      $signed(((~wire1766) ?
                          {forvar1776} : (wire1774 & (8'hb4)))) : (wire1766 != $unsigned((forvar1789 ?
                          wire1772 : forvar1776)))))
                    begin
                      reg1795 <= ({((reg1819 ? (8'hb4) : reg1778) ?
                                  $signed(forvar1799) : $unsigned(forvar1785))} ?
                          (^~wire1769) : $signed(((wire1769 ?
                                  (8'hac) : forvar1820) ?
                              $signed(reg1809) : {reg1805})));
                      reg1796 <= reg1818;
                    end
                  else
                    begin
                      reg1795 <= reg1789;
                      reg1796 <= ((~&(reg1798 && ((8'ha9) * reg1780))) ?
                          forvar1807[(4'h8):(2'h3)] : reg1818[(1'h1):(1'h1)]);
                      reg1797 <= (~|wire1769);
                    end
                end
              else
                begin
                  for (forvar1793 = (1'h0); (forvar1793 < (2'h3)); forvar1793 = (forvar1793 + (1'h1)))
                    begin
                      reg1794 <= $signed({reg1814});
                      reg1795 <= (~^(-(~^(8'h9e))));
                      reg1796 <= reg1777[(3'h5):(1'h0)];
                    end
                  if ((~&reg1779))
                    begin
                      reg1797 <= ((wire1771[(3'h5):(1'h1)] < $signed(((8'hb6) - reg1810))) ?
                          reg1786[(2'h3):(2'h3)] : (~^{reg1810}));
                      reg1798 <= $unsigned({reg1825});
                      reg1799 <= reg1778[(4'h8):(2'h2)];
                    end
                  else
                    begin
                      reg1797 <= (-(($signed(wire1768) ?
                              ((8'ha1) >= reg1796) : $signed(reg1828)) ?
                          wire1768[(3'h5):(1'h1)] : $signed($signed(forvar1797))));
                      reg1798 <= ((~|reg1780) ?
                          (8'h9e) : (!$signed({(8'ha1)})));
                      reg1799 <= reg1805[(2'h3):(1'h1)];
                      reg1800 <= (reg1825[(2'h2):(1'h0)] ?
                          $signed((~^reg1823[(4'h9):(3'h5)])) : ($unsigned($unsigned((8'h9e))) ?
                              $unsigned((reg1784 << wire1769)) : ((reg1790 ?
                                      forvar1784 : wire1766) ?
                                  (|forvar1780) : (forvar1806 >> reg1783))));
                    end
                  for (forvar1801 = (1'h0); (forvar1801 < (2'h3)); forvar1801 = (forvar1801 + (1'h1)))
                    begin
                      reg1802 <= ($unsigned(forvar1775[(2'h2):(1'h1)]) ?
                          $signed(reg1775[(3'h4):(1'h0)]) : (~^reg1804[(1'h0):(1'h0)]));
                    end
                end
              for (forvar1803 = (1'h0); (forvar1803 < (1'h1)); forvar1803 = (forvar1803 + (1'h1)))
                begin
                  if ((($unsigned($signed(reg1793)) ?
                      forvar1787[(3'h5):(1'h0)] : $signed((wire1767 <<< (8'ha4)))) || $unsigned({wire1771[(1'h1):(1'h0)]})))
                    begin
                      reg1804 <= $unsigned($unsigned(forvar1775[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg1804 <= ($signed(forvar1776[(4'he):(1'h1)]) <<< (reg1826[(3'h4):(1'h1)] & $unsigned($signed(forvar1783))));
                    end
                  for (forvar1805 = (1'h0); (forvar1805 < (1'h1)); forvar1805 = (forvar1805 + (1'h1)))
                    begin
                      reg1806 <= (~|(~{wire1774[(1'h1):(1'h0)]}));
                      reg1807 <= reg1786;
                      reg1808 <= ((~^forvar1776) ~^ $signed((-(reg1822 - reg1793))));
                    end
                  for (forvar1809 = (1'h0); (forvar1809 < (1'h1)); forvar1809 = (forvar1809 + (1'h1)))
                    begin
                      reg1810 <= ((-$unsigned({forvar1776})) ^ (^$unsigned({forvar1805})));
                      reg1811 <= ((($signed((8'ha7)) ?
                              $signed(reg1791) : (reg1796 >> forvar1785)) << reg1798) ?
                          $signed(reg1823[(4'h8):(4'h8)]) : ({((8'ha4) + (8'hb2))} ?
                              reg1806[(3'h5):(1'h1)] : {reg1804[(2'h2):(2'h2)]}));
                    end
                  if ((^~forvar1776[(4'he):(2'h2)]))
                    begin
                      reg1812 <= reg1807;
                    end
                  else
                    begin
                      reg1812 <= $signed(($signed($unsigned(reg1818)) ^~ {reg1829[(3'h5):(3'h4)]}));
                    end
                end
            end
        end
      for (forvar1830 = (1'h0); (forvar1830 < (1'h0)); forvar1830 = (forvar1830 + (1'h1)))
        begin
          if (reg1787)
            begin
              for (forvar1831 = (1'h0); (forvar1831 < (2'h2)); forvar1831 = (forvar1831 + (1'h1)))
                begin
                  for (forvar1832 = (1'h0); (forvar1832 < (2'h3)); forvar1832 = (forvar1832 + (1'h1)))
                    begin
                      reg1833 <= reg1798[(4'h9):(3'h4)];
                      reg1834 <= (reg1827[(4'h8):(3'h6)] | $unsigned($signed(wire1770[(4'hc):(4'h8)])));
                      reg1835 <= {$signed(((forvar1789 ^ (8'ha0)) ^ reg1780[(1'h0):(1'h0)]))};
                      reg1836 <= (~&(($signed(reg1815) ^~ $signed(reg1833)) >= (~|(reg1803 ?
                          wire1774 : reg1815))));
                    end
                  reg1837 <= (((reg1825[(2'h2):(1'h0)] ?
                          (8'had) : (forvar1793 ?
                              (8'hb2) : forvar1820)) != (~forvar1799)) ?
                      {wire1772} : $unsigned($signed(forvar1776)));
                  for (forvar1838 = (1'h0); (forvar1838 < (1'h1)); forvar1838 = (forvar1838 + (1'h1)))
                    begin
                      reg1839 <= $signed((-{forvar1806[(3'h7):(1'h1)]}));
                      reg1840 <= $unsigned((8'hb0));
                      reg1841 <= $unsigned($unsigned($signed(forvar1838)));
                    end
                  reg1842 <= ($signed({(~|(8'ha1))}) | ($signed($signed(reg1779)) ?
                      forvar1832 : ((reg1802 ?
                          reg1806 : forvar1794) || $unsigned(reg1813))));
                end
            end
          else
            begin
              for (forvar1831 = (1'h0); (forvar1831 < (1'h0)); forvar1831 = (forvar1831 + (1'h1)))
                begin
                  for (forvar1832 = (1'h0); (forvar1832 < (1'h1)); forvar1832 = (forvar1832 + (1'h1)))
                    begin
                      reg1833 <= $signed((forvar1802 << forvar1788));
                    end
                  for (forvar1834 = (1'h0); (forvar1834 < (2'h3)); forvar1834 = (forvar1834 + (1'h1)))
                    begin
                      reg1835 <= $unsigned((reg1803[(2'h2):(1'h1)] ?
                          $signed(reg1833[(3'h6):(3'h6)]) : ((reg1795 - forvar1831) + $unsigned(reg1782))));
                      reg1836 <= {$unsigned($signed((|wire1769)))};
                      reg1837 <= forvar1794;
                      reg1838 <= forvar1809;
                    end
                end
              for (forvar1839 = (1'h0); (forvar1839 < (1'h0)); forvar1839 = (forvar1839 + (1'h1)))
                begin
                  for (forvar1840 = (1'h0); (forvar1840 < (2'h3)); forvar1840 = (forvar1840 + (1'h1)))
                    begin
                      reg1841 <= $unsigned((8'h9e));
                      reg1842 <= (!{(^$unsigned(reg1780))});
                      reg1843 <= $signed($unsigned($unsigned(forvar1797[(3'h6):(2'h2)])));
                      reg1844 <= reg1818;
                    end
                  for (forvar1845 = (1'h0); (forvar1845 < (2'h2)); forvar1845 = (forvar1845 + (1'h1)))
                    begin
                      reg1846 <= (forvar1775 ?
                          $signed((reg1805 ?
                              reg1805[(1'h1):(1'h0)] : (wire1769 ?
                                  reg1823 : reg1814))) : (forvar1784[(1'h0):(1'h0)] ?
                              ((reg1816 ?
                                  (8'h9d) : reg1804) && $unsigned(reg1788)) : {(forvar1839 ?
                                      reg1816 : reg1842)}));
                      reg1847 <= reg1801;
                      reg1848 <= forvar1803[(4'he):(3'h4)];
                      reg1849 <= (((~(|(8'hba))) < wire1771[(2'h2):(1'h1)]) ?
                          (reg1802 >>> ({forvar1797} ?
                              reg1840 : reg1814[(1'h0):(1'h0)])) : $signed((forvar1801 ?
                              reg1838 : ((8'ha1) ? reg1825 : (8'ha7)))));
                    end
                  if ($signed(forvar1785[(2'h2):(1'h0)]))
                    begin
                      reg1850 <= $signed((~|$signed(reg1783[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg1850 <= reg1805[(1'h1):(1'h1)];
                      reg1851 <= ((forvar1775[(3'h7):(1'h0)] ?
                          (reg1785 ?
                              (reg1844 ?
                                  reg1787 : reg1839) : forvar1839) : $unsigned(((8'ha9) ~^ wire1774))) & (($signed((8'hb0)) ?
                              $signed(reg1812) : $signed(reg1781)) ?
                          reg1803 : (!$signed(reg1781))));
                      reg1852 <= ((($signed(reg1846) ?
                                  {reg1811} : forvar1787[(3'h5):(1'h0)]) ?
                              $signed({reg1848}) : $signed((reg1793 << reg1781))) ?
                          (!$signed($unsigned(reg1843))) : {(-{wire1771})});
                    end
                  if (reg1798)
                    begin
                      reg1853 <= ($unsigned(reg1838[(2'h2):(1'h1)]) ?
                          forvar1788 : (((~|reg1794) ?
                              $unsigned((8'haf)) : (reg1852 ?
                                  reg1843 : reg1840)) && reg1797[(4'hb):(3'h4)]));
                      reg1854 <= (+reg1788);
                    end
                  else
                    begin
                      reg1853 <= ((~^{forvar1806}) ^~ $signed($signed({reg1853})));
                      reg1854 <= (reg1785 ^~ $signed({reg1782}));
                      reg1855 <= (forvar1839[(2'h2):(1'h0)] > reg1785);
                      reg1856 <= ($unsigned((forvar1831[(3'h6):(1'h0)] <<< $unsigned(reg1848))) + forvar1797);
                    end
                end
              for (forvar1857 = (1'h0); (forvar1857 < (1'h1)); forvar1857 = (forvar1857 + (1'h1)))
                begin
                  reg1858 <= (reg1786[(2'h2):(2'h2)] + $signed((|forvar1783[(3'h6):(3'h6)])));
                  if (wire1771[(3'h6):(3'h4)])
                    begin
                      reg1859 <= (~&{reg1794[(4'he):(3'h5)]});
                      reg1860 <= $signed($signed(forvar1787));
                      reg1861 <= $signed($unsigned($unsigned((&forvar1803))));
                      reg1862 <= $unsigned({$signed((reg1792 ^ reg1778))});
                    end
                  else
                    begin
                      reg1859 <= (reg1811[(2'h2):(1'h0)] >>> reg1816[(4'hd):(4'h9)]);
                      reg1860 <= (((-(forvar1787 || reg1839)) && (reg1814 >>> (reg1812 ?
                              reg1858 : reg1778))) ?
                          $signed($unsigned(forvar1839[(2'h3):(1'h0)])) : ((~|(forvar1824 ?
                                  reg1833 : reg1787)) ?
                              reg1835 : $signed(reg1777)));
                      reg1861 <= (8'hb8);
                      reg1862 <= reg1792[(3'h5):(3'h5)];
                    end
                  if ((!reg1842))
                    begin
                      reg1863 <= $signed($signed(forvar1797[(4'hd):(4'h8)]));
                      reg1864 <= $unsigned((~^($unsigned(reg1825) > (forvar1785 >> reg1786))));
                      reg1865 <= ($unsigned((!reg1825)) ?
                          (8'h9c) : $unsigned(($unsigned(reg1785) < $unsigned(reg1847))));
                    end
                  else
                    begin
                      reg1863 <= (&$unsigned(reg1852[(1'h1):(1'h1)]));
                    end
                end
              for (forvar1866 = (1'h0); (forvar1866 < (2'h2)); forvar1866 = (forvar1866 + (1'h1)))
                begin
                  for (forvar1867 = (1'h0); (forvar1867 < (2'h2)); forvar1867 = (forvar1867 + (1'h1)))
                    begin
                      reg1868 <= (&$signed($unsigned(reg1842[(3'h5):(3'h4)])));
                      reg1869 <= {forvar1793[(1'h1):(1'h0)]};
                    end
                  for (forvar1870 = (1'h0); (forvar1870 < (1'h0)); forvar1870 = (forvar1870 + (1'h1)))
                    begin
                      reg1871 <= ($signed((((8'had) ?
                          reg1810 : reg1787) + (reg1816 <<< forvar1834))) ~^ $unsigned($signed($unsigned(forvar1802))));
                      reg1872 <= reg1863[(3'h4):(2'h3)];
                      reg1873 <= $unsigned($signed((~^$signed(forvar1789))));
                    end
                end
            end
        end
      for (forvar1874 = (1'h0); (forvar1874 < (1'h0)); forvar1874 = (forvar1874 + (1'h1)))
        begin
          for (forvar1875 = (1'h0); (forvar1875 < (1'h0)); forvar1875 = (forvar1875 + (1'h1)))
            begin
              if ((!$signed(wire1765)))
                begin
                  for (forvar1876 = (1'h0); (forvar1876 < (1'h1)); forvar1876 = (forvar1876 + (1'h1)))
                    begin
                      reg1877 <= $signed(reg1792[(3'h6):(2'h2)]);
                      reg1878 <= (reg1785 && reg1853);
                      reg1879 <= (reg1799[(1'h0):(1'h0)] ?
                          (($unsigned(reg1842) & $signed(reg1805)) ?
                              reg1786[(1'h1):(1'h1)] : $signed((reg1804 + forvar1788))) : (^~($signed(reg1840) | ((8'hab) ?
                              reg1826 : (8'hb6)))));
                      reg1880 <= ((^reg1819[(3'h5):(1'h0)]) ?
                          $unsigned(($signed(reg1852) ?
                              (~reg1796) : (~^reg1846))) : $signed(($signed(wire1765) ^ (reg1841 ?
                              reg1854 : reg1782))));
                    end
                  reg1881 <= $signed((&($signed(reg1858) ?
                      $signed(reg1835) : forvar1803)));
                end
              else
                begin
                  for (forvar1876 = (1'h0); (forvar1876 < (1'h1)); forvar1876 = (forvar1876 + (1'h1)))
                    begin
                      reg1877 <= reg1775;
                      reg1878 <= $unsigned(forvar1775);
                      reg1879 <= {reg1850};
                      reg1880 <= {forvar1789[(4'hb):(3'h5)]};
                    end
                  if (((((-forvar1802) ^ $signed(reg1778)) ?
                          ((^reg1846) ?
                              reg1850[(3'h5):(2'h3)] : $unsigned(reg1853)) : reg1817[(4'h8):(3'h7)]) ?
                      (~&$signed((forvar1793 ~^ (8'hae)))) : $signed(reg1796)))
                    begin
                      reg1881 <= $signed((8'ha4));
                      reg1882 <= (reg1814 || reg1788);
                    end
                  else
                    begin
                      reg1881 <= $signed($signed({$unsigned(wire1766)}));
                      reg1882 <= ((!$unsigned({reg1779})) * {reg1823});
                      reg1883 <= $signed({(8'hb6)});
                    end
                  for (forvar1884 = (1'h0); (forvar1884 < (1'h0)); forvar1884 = (forvar1884 + (1'h1)))
                    begin
                      reg1885 <= reg1808[(3'h5):(3'h4)];
                      reg1886 <= {(reg1823[(4'ha):(4'ha)] ?
                              (!$unsigned(reg1849)) : ({forvar1834} ?
                                  (reg1780 ^~ forvar1783) : (forvar1776 & forvar1839)))};
                    end
                end
              for (forvar1887 = (1'h0); (forvar1887 < (1'h1)); forvar1887 = (forvar1887 + (1'h1)))
                begin
                  if (((&(forvar1784 ?
                      reg1865 : (^~forvar1794))) >= (((~|reg1790) ?
                      (~forvar1806) : reg1833) >> $unsigned(((8'hb9) ?
                      forvar1838 : forvar1806)))))
                    begin
                      reg1888 <= (~$unsigned($signed((~^(8'h9e)))));
                      reg1889 <= reg1871;
                      reg1890 <= $unsigned(reg1865[(3'h4):(1'h0)]);
                      reg1891 <= (reg1835[(1'h1):(1'h1)] ?
                          ($unsigned($unsigned((8'ha7))) <<< $unsigned($signed(forvar1807))) : reg1793);
                    end
                  else
                    begin
                      reg1888 <= forvar1787;
                      reg1889 <= reg1840[(1'h0):(1'h0)];
                      reg1890 <= ($unsigned({(reg1888 ?
                                  forvar1867 : reg1790)}) ?
                          {(8'hb0)} : (!$unsigned($unsigned(reg1888))));
                    end
                end
              if (reg1777)
                begin
                  if ($unsigned($signed((&$signed((8'hb9))))))
                    begin
                      reg1892 <= reg1779[(3'h5):(1'h0)];
                      reg1893 <= reg1888;
                      reg1894 <= (reg1889 ? wire1768 : reg1803[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1892 <= ($signed(((!reg1818) ?
                              reg1777 : $signed(reg1789))) ?
                          $signed($signed(forvar1834[(1'h1):(1'h0)])) : (^~($signed(reg1819) && $unsigned(reg1780))));
                      reg1893 <= {((8'ha2) && reg1861[(3'h5):(3'h4)])};
                      reg1894 <= ((&($signed((8'hba)) > (reg1889 <<< reg1795))) != (8'hb4));
                      reg1895 <= (-(((reg1816 & reg1807) ?
                              forvar1776 : $unsigned(reg1792)) ?
                          $unsigned(forvar1794) : reg1864[(1'h0):(1'h0)]));
                    end
                  for (forvar1896 = (1'h0); (forvar1896 < (1'h0)); forvar1896 = (forvar1896 + (1'h1)))
                    begin
                      reg1897 <= reg1789[(4'h9):(4'h9)];
                      reg1898 <= ((((^~reg1850) | $signed(wire1769)) > $unsigned(wire1767)) > $signed((^~$unsigned(reg1801))));
                      reg1899 <= reg1842;
                    end
                  if ((+reg1806[(1'h1):(1'h1)]))
                    begin
                      reg1900 <= {({$unsigned(reg1804)} ?
                              (8'h9e) : (forvar1830[(1'h1):(1'h1)] + reg1890))};
                      reg1901 <= $signed((8'h9d));
                      reg1902 <= reg1833[(4'h8):(3'h6)];
                      reg1903 <= ($unsigned($signed((forvar1801 ?
                          reg1849 : forvar1793))) << ($signed($signed(reg1808)) ?
                          ((reg1837 ~^ reg1852) >= $unsigned(wire1768)) : reg1801));
                    end
                  else
                    begin
                      reg1900 <= $signed($unsigned(reg1890[(2'h2):(1'h0)]));
                      reg1901 <= {(reg1852[(1'h0):(1'h0)] | {{(8'ha5)}})};
                    end
                end
              else
                begin
                  if ($signed(((wire1774 ^~ {reg1792}) ?
                      $signed($unsigned(reg1801)) : reg1838)))
                    begin
                      reg1892 <= (reg1792[(3'h7):(1'h1)] ~^ $unsigned($signed(reg1853)));
                      reg1893 <= reg1775[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1892 <= $signed((((8'h9e) ?
                          ((8'hae) ?
                              reg1828 : forvar1783) : $unsigned(reg1899)) > reg1784[(2'h2):(2'h2)]));
                      reg1893 <= $unsigned($unsigned(forvar1799[(2'h2):(2'h2)]));
                    end
                  for (forvar1894 = (1'h0); (forvar1894 < (1'h0)); forvar1894 = (forvar1894 + (1'h1)))
                    begin
                      reg1895 <= $signed($signed(wire1768));
                    end
                  for (forvar1896 = (1'h0); (forvar1896 < (2'h3)); forvar1896 = (forvar1896 + (1'h1)))
                    begin
                      reg1897 <= {$signed($signed(reg1848[(3'h4):(3'h4)]))};
                      reg1898 <= (~(-($signed(wire1774) ?
                          $signed(reg1898) : reg1809[(4'hb):(2'h3)])));
                      reg1899 <= ($signed(forvar1839[(2'h2):(2'h2)]) << forvar1802);
                      reg1900 <= {reg1890};
                    end
                  for (forvar1901 = (1'h0); (forvar1901 < (2'h2)); forvar1901 = (forvar1901 + (1'h1)))
                    begin
                      reg1902 <= (~|(+{reg1806[(1'h0):(1'h0)]}));
                    end
                end
              if (reg1855)
                begin
                  reg1904 <= $signed({$signed(((8'h9d) ? reg1839 : reg1782))});
                  for (forvar1905 = (1'h0); (forvar1905 < (1'h0)); forvar1905 = (forvar1905 + (1'h1)))
                    begin
                      reg1906 <= $signed(((8'hab) >= reg1840));
                    end
                  for (forvar1907 = (1'h0); (forvar1907 < (1'h1)); forvar1907 = (forvar1907 + (1'h1)))
                    begin
                      reg1908 <= $unsigned(forvar1801);
                      reg1909 <= ((((~^wire1774) == ((8'ha4) ?
                          (8'hb7) : reg1900)) << $signed($signed(reg1889))) ^~ {$signed($signed((8'ha1)))});
                      reg1910 <= forvar1845;
                      reg1911 <= (8'hb9);
                    end
                end
              else
                begin
                  for (forvar1904 = (1'h0); (forvar1904 < (2'h3)); forvar1904 = (forvar1904 + (1'h1)))
                    begin
                      reg1905 <= $unsigned($unsigned(({reg1829} | $unsigned(reg1856))));
                    end
                  for (forvar1906 = (1'h0); (forvar1906 < (2'h3)); forvar1906 = (forvar1906 + (1'h1)))
                    begin
                      reg1907 <= reg1892[(2'h3):(2'h3)];
                      reg1908 <= reg1815;
                      reg1909 <= reg1865;
                      reg1910 <= reg1864;
                    end
                end
            end
        end
      if ({$unsigned(reg1804[(1'h1):(1'h0)])})
        begin
          for (forvar1912 = (1'h0); (forvar1912 < (2'h2)); forvar1912 = (forvar1912 + (1'h1)))
            begin
              if ($signed({{(+forvar1838)}}))
                begin
                  reg1913 <= (~^$unsigned({(reg1847 ? reg1816 : reg1844)}));
                  for (forvar1914 = (1'h0); (forvar1914 < (2'h3)); forvar1914 = (forvar1914 + (1'h1)))
                    begin
                      reg1915 <= (($unsigned((reg1898 < reg1808)) ?
                          {(reg1908 ~^ reg1784)} : (wire1768 ?
                              (wire1771 >>> (8'hba)) : reg1913[(1'h0):(1'h0)])) << forvar1894[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  if (($unsigned($signed($unsigned((8'ha1)))) ?
                      forvar1830 : $unsigned(($signed(reg1839) << {reg1800}))))
                    begin
                      reg1913 <= $unsigned(reg1858[(4'h9):(2'h2)]);
                      reg1914 <= reg1885[(2'h3):(2'h2)];
                      reg1915 <= $unsigned(({reg1850[(3'h6):(3'h4)]} ?
                          $unsigned(reg1809[(4'h9):(3'h7)]) : ($signed(reg1886) ?
                              forvar1904[(1'h0):(1'h0)] : forvar1907)));
                    end
                  else
                    begin
                      reg1913 <= ((8'hb0) & $unsigned($signed((^~(8'hb1)))));
                      reg1914 <= $signed((reg1897 ?
                          $unsigned((|reg1826)) : $signed(reg1841)));
                    end
                  if ((~|reg1903))
                    begin
                      reg1916 <= {reg1852};
                      reg1917 <= (~$signed((forvar1832 > $signed(reg1843))));
                      reg1918 <= (reg1897[(3'h6):(2'h2)] < reg1787);
                      reg1919 <= forvar1907[(3'h7):(1'h0)];
                    end
                  else
                    begin
                      reg1916 <= (^~$signed(((8'hb6) ?
                          forvar1867[(3'h6):(3'h4)] : (wire1770 ?
                              (8'ha4) : reg1807))));
                      reg1917 <= {$signed(((reg1818 ? reg1889 : forvar1780) ?
                              $unsigned(reg1795) : (&reg1782)))};
                      reg1918 <= reg1909[(1'h1):(1'h0)];
                    end
                  for (forvar1920 = (1'h0); (forvar1920 < (2'h2)); forvar1920 = (forvar1920 + (1'h1)))
                    begin
                      reg1921 <= (8'hac);
                    end
                end
              for (forvar1922 = (1'h0); (forvar1922 < (1'h1)); forvar1922 = (forvar1922 + (1'h1)))
                begin
                  reg1923 <= {{$signed((8'ha9))}};
                end
              reg1924 <= reg1800[(4'hf):(4'h8)];
              for (forvar1925 = (1'h0); (forvar1925 < (2'h2)); forvar1925 = (forvar1925 + (1'h1)))
                begin
                  reg1926 <= reg1860;
                end
            end
        end
      else
        begin
          for (forvar1912 = (1'h0); (forvar1912 < (2'h2)); forvar1912 = (forvar1912 + (1'h1)))
            begin
              for (forvar1913 = (1'h0); (forvar1913 < (2'h2)); forvar1913 = (forvar1913 + (1'h1)))
                begin
                  if (({reg1856[(4'h8):(2'h3)]} || (|forvar1824[(1'h1):(1'h1)])))
                    begin
                      reg1914 <= reg1799;
                      reg1915 <= $unsigned((8'haf));
                    end
                  else
                    begin
                      reg1914 <= ((reg1781[(1'h1):(1'h1)] - reg1911) || reg1848);
                      reg1915 <= ({$unsigned(wire1771)} ^ $signed((wire1769[(1'h1):(1'h1)] ~^ $signed(reg1911))));
                      reg1916 <= reg1909;
                    end
                  for (forvar1917 = (1'h0); (forvar1917 < (2'h2)); forvar1917 = (forvar1917 + (1'h1)))
                    begin
                      reg1918 <= $unsigned((reg1815[(4'ha):(3'h7)] | (+$unsigned(reg1778))));
                      reg1919 <= {$signed($unsigned($signed(reg1837)))};
                      reg1920 <= (reg1858[(3'h7):(1'h1)] == reg1818);
                      reg1921 <= (8'ha2);
                    end
                  for (forvar1922 = (1'h0); (forvar1922 < (1'h0)); forvar1922 = (forvar1922 + (1'h1)))
                    begin
                      reg1923 <= (^~(&(forvar1884[(4'ha):(2'h2)] ?
                          (forvar1914 ? (8'h9e) : reg1802) : ((8'hb7) ?
                              reg1805 : reg1793))));
                    end
                  for (forvar1924 = (1'h0); (forvar1924 < (2'h3)); forvar1924 = (forvar1924 + (1'h1)))
                    begin
                      reg1925 <= reg1802;
                      reg1926 <= (forvar1834[(3'h5):(2'h3)] ?
                          ({forvar1805[(4'h8):(3'h5)]} ?
                              $unsigned(((8'hba) ?
                                  (8'ha6) : reg1811)) : $unsigned({reg1905})) : (8'h9c));
                    end
                end
              if ((reg1840[(3'h6):(3'h5)] ? reg1856 : reg1891))
                begin
                  if ((reg1776[(3'h4):(2'h2)] ?
                      $signed(reg1852) : reg1842[(1'h1):(1'h1)]))
                    begin
                      reg1927 <= forvar1811;
                      reg1928 <= (reg1842 && $unsigned((|(reg1883 ~^ reg1869))));
                    end
                  else
                    begin
                      reg1927 <= forvar1821[(3'h4):(1'h1)];
                      reg1928 <= $signed($signed($signed($unsigned(reg1900))));
                      reg1929 <= (reg1789 >> ((^~(~&forvar1924)) <= ((reg1791 ^ reg1925) ?
                          $signed(reg1895) : (forvar1803 ?
                              forvar1801 : wire1766))));
                    end
                  for (forvar1930 = (1'h0); (forvar1930 < (2'h2)); forvar1930 = (forvar1930 + (1'h1)))
                    begin
                      reg1931 <= $signed($signed((+$signed(forvar1794))));
                      reg1932 <= reg1807;
                    end
                end
              else
                begin
                  for (forvar1927 = (1'h0); (forvar1927 < (2'h3)); forvar1927 = (forvar1927 + (1'h1)))
                    begin
                      reg1928 <= $signed($signed(reg1859));
                      reg1929 <= $unsigned(reg1868);
                    end
                  for (forvar1930 = (1'h0); (forvar1930 < (2'h3)); forvar1930 = (forvar1930 + (1'h1)))
                    begin
                      reg1931 <= $unsigned((|(~^$unsigned(forvar1870))));
                    end
                  for (forvar1932 = (1'h0); (forvar1932 < (2'h2)); forvar1932 = (forvar1932 + (1'h1)))
                    begin
                      reg1933 <= forvar1806[(4'h9):(1'h1)];
                      reg1934 <= reg1904;
                      reg1935 <= reg1803[(1'h0):(1'h0)];
                      reg1936 <= $signed(((((8'h9d) != reg1886) ?
                              (~^reg1784) : $signed((8'hb3))) ?
                          $signed(reg1808[(4'hc):(3'h7)]) : (~$signed(reg1787))));
                    end
                end
            end
          if (($unsigned($signed($signed(reg1905))) <<< $unsigned($signed(forvar1866))))
            begin
              if (($unsigned((~&(-reg1931))) >>> reg1804))
                begin
                  if ($unsigned($unsigned((|$unsigned(reg1863)))))
                    begin
                      reg1937 <= {($signed($signed((8'h9e))) ?
                              ((forvar1780 ? forvar1912 : forvar1906) ?
                                  (^~reg1861) : (reg1851 ?
                                      (8'hb6) : (8'hb8))) : reg1916)};
                      reg1938 <= (((8'h9d) ?
                          ($signed(wire1766) ?
                              reg1822 : (reg1849 ^ (8'ha3))) : $unsigned(reg1786)) <<< $signed(((reg1856 & forvar1784) <= (~reg1905))));
                      reg1939 <= forvar1785[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1937 <= $signed(((reg1809[(3'h7):(3'h7)] | reg1781) ?
                          reg1828[(2'h2):(1'h0)] : $unsigned(reg1880[(1'h0):(1'h0)])));
                      reg1938 <= $unsigned((!reg1901));
                      reg1939 <= reg1783[(2'h3):(2'h3)];
                    end
                  for (forvar1940 = (1'h0); (forvar1940 < (1'h0)); forvar1940 = (forvar1940 + (1'h1)))
                    begin
                      reg1941 <= {({$unsigned(wire1769)} ?
                              (reg1906 ^ (reg1923 ?
                                  (8'haf) : reg1799)) : reg1878)};
                      reg1942 <= ({($unsigned(reg1838) ?
                              (forvar1839 ?
                                  reg1905 : reg1828) : (forvar1907 + forvar1787))} < (reg1784 ?
                          ((|reg1897) ?
                              reg1907 : $signed((8'hb5))) : reg1779[(2'h3):(2'h2)]));
                    end
                  reg1943 <= reg1894;
                  for (forvar1944 = (1'h0); (forvar1944 < (2'h2)); forvar1944 = (forvar1944 + (1'h1)))
                    begin
                      reg1945 <= (reg1782[(2'h3):(2'h2)] & $unsigned(($unsigned((8'ha7)) ?
                          forvar1840[(3'h4):(2'h3)] : reg1804[(2'h3):(1'h1)])));
                      reg1946 <= wire1769[(1'h0):(1'h0)];
                      reg1947 <= (reg1853[(2'h3):(1'h1)] ?
                          (8'h9d) : (&{$unsigned(reg1800)}));
                    end
                end
              else
                begin
                  for (forvar1937 = (1'h0); (forvar1937 < (2'h2)); forvar1937 = (forvar1937 + (1'h1)))
                    begin
                      reg1938 <= {(&$signed(reg1947))};
                    end
                  for (forvar1939 = (1'h0); (forvar1939 < (1'h0)); forvar1939 = (forvar1939 + (1'h1)))
                    begin
                      reg1940 <= reg1844;
                    end
                  for (forvar1941 = (1'h0); (forvar1941 < (2'h2)); forvar1941 = (forvar1941 + (1'h1)))
                    begin
                      reg1942 <= {$unsigned((~^(&(8'ha8))))};
                      reg1943 <= (&(~$unsigned(reg1859[(3'h5):(3'h4)])));
                      reg1944 <= (reg1856[(4'h9):(3'h7)] <= ((8'hb5) ?
                          $unsigned(reg1779) : ({reg1858} + forvar1811[(1'h1):(1'h1)])));
                    end
                end
              if (reg1902[(1'h0):(1'h0)])
                begin
                  for (forvar1948 = (1'h0); (forvar1948 < (1'h1)); forvar1948 = (forvar1948 + (1'h1)))
                    begin
                      reg1949 <= $unsigned($signed((~&(-reg1926))));
                      reg1950 <= wire1771[(3'h6):(1'h0)];
                    end
                  reg1951 <= $signed($unsigned({reg1814}));
                end
              else
                begin
                  for (forvar1948 = (1'h0); (forvar1948 < (1'h1)); forvar1948 = (forvar1948 + (1'h1)))
                    begin
                      reg1949 <= $signed($signed(((&(8'hb4)) ?
                          (reg1901 << reg1926) : (reg1938 ?
                              reg1931 : forvar1937))));
                      reg1950 <= ((~(+(-forvar1775))) ?
                          (((^~(8'hb2)) ? $unsigned(forvar1876) : (^reg1901)) ?
                              {(~&forvar1809)} : $signed($signed(forvar1794))) : forvar1793);
                      reg1951 <= forvar1803[(4'hd):(3'h4)];
                      reg1952 <= $signed((($signed(reg1779) ^ reg1877[(4'hb):(1'h0)]) ?
                          ((|reg1883) && $unsigned(reg1871)) : wire1767));
                    end
                  reg1953 <= reg1947;
                  reg1954 <= forvar1930[(3'h4):(2'h2)];
                end
              if ((forvar1905 - (^$unsigned(forvar1830))))
                begin
                  for (forvar1955 = (1'h0); (forvar1955 < (2'h2)); forvar1955 = (forvar1955 + (1'h1)))
                    begin
                      reg1956 <= $unsigned((~reg1794));
                      reg1957 <= ((^~$signed(reg1898)) >> ((~^(-(8'ha5))) ?
                          ($unsigned(forvar1789) != (wire1772 ?
                              (8'hb5) : reg1838)) : $signed(reg1803[(1'h0):(1'h0)])));
                      reg1958 <= (^(({reg1861} ?
                              (^forvar1803) : (forvar1927 ?
                                  forvar1941 : wire1774)) ?
                          reg1913 : {$signed(forvar1824)}));
                    end
                  if (($signed(forvar1807[(3'h6):(1'h1)]) ?
                      $signed(forvar1914[(2'h2):(1'h1)]) : forvar1912))
                    begin
                      reg1959 <= reg1795;
                    end
                  else
                    begin
                      reg1959 <= (({(reg1893 ? reg1865 : wire1770)} & reg1904) ?
                          (((8'hac) ?
                                  reg1893[(2'h2):(2'h2)] : ((8'haf) + (8'had))) ?
                              ((^reg1953) <= $signed(reg1853)) : $unsigned((~&forvar1801))) : {$signed($signed(reg1786))});
                      reg1960 <= ($signed(reg1788[(3'h5):(2'h2)]) < ((8'hac) ?
                          $unsigned($unsigned(wire1767)) : forvar1917));
                      reg1961 <= ((!(reg1883 == (reg1780 + reg1829))) ?
                          {(-reg1878)} : (!((reg1897 <= forvar1811) ?
                              forvar1834[(4'ha):(1'h1)] : $signed(reg1898))));
                      reg1962 <= forvar1789[(5'h10):(5'h10)];
                    end
                end
              else
                begin
                  if ($unsigned(forvar1801[(3'h5):(2'h2)]))
                    begin
                      reg1955 <= $unsigned(((forvar1834 ?
                              $signed(forvar1907) : wire1774[(1'h0):(1'h0)]) ?
                          (|((8'hb5) >>> reg1789)) : ((forvar1820 ?
                                  reg1903 : (8'hb0)) ?
                              (&forvar1776) : $signed(reg1891))));
                      reg1956 <= $unsigned({((^forvar1805) << $unsigned(reg1895))});
                    end
                  else
                    begin
                      reg1955 <= (|((reg1787[(3'h5):(1'h0)] ?
                          {(8'had)} : (reg1935 ?
                              reg1949 : reg1925)) + $signed(((8'h9f) ?
                          reg1810 : (8'ha9)))));
                      reg1956 <= $signed(((!$signed(forvar1920)) ?
                          $unsigned($unsigned((8'ha2))) : reg1781));
                      reg1957 <= {$unsigned($unsigned($unsigned(reg1943)))};
                    end
                  for (forvar1958 = (1'h0); (forvar1958 < (1'h1)); forvar1958 = (forvar1958 + (1'h1)))
                    begin
                      reg1959 <= (reg1897[(3'h7):(3'h7)] ?
                          $unsigned($signed(wire1772)) : {$unsigned((forvar1870 ?
                                  reg1849 : (8'haa)))});
                      reg1960 <= ($unsigned((8'h9e)) && (reg1860[(3'h5):(3'h4)] | $signed((reg1795 ?
                          reg1823 : reg1927))));
                      reg1961 <= $unsigned((8'hac));
                    end
                  reg1962 <= $unsigned(reg1801);
                end
              for (forvar1963 = (1'h0); (forvar1963 < (1'h0)); forvar1963 = (forvar1963 + (1'h1)))
                begin
                  if ((|((forvar1941 || reg1902) ?
                      $signed(reg1905[(4'hd):(4'h8)]) : $unsigned((forvar1784 << forvar1784)))))
                    begin
                      reg1964 <= (^(~{(|reg1782)}));
                      reg1965 <= (^wire1770[(4'hc):(1'h0)]);
                    end
                  else
                    begin
                      reg1964 <= ($signed($signed((reg1799 ?
                          reg1852 : reg1849))) | $unsigned((^~((8'ha1) ?
                          forvar1925 : reg1908))));
                    end
                end
            end
          else
            begin
              if (reg1816[(4'he):(1'h0)])
                begin
                  for (forvar1937 = (1'h0); (forvar1937 < (1'h1)); forvar1937 = (forvar1937 + (1'h1)))
                    begin
                      reg1938 <= reg1790[(3'h6):(2'h3)];
                      reg1939 <= ((({reg1861} ?
                          {reg1803} : forvar1955[(2'h2):(2'h2)]) >= $unsigned((reg1792 << reg1833))) < (^(&{reg1835})));
                      reg1940 <= (~&($signed((^reg1947)) ?
                          ({forvar1887} || (-(8'hb4))) : reg1778));
                      reg1941 <= {(((~|(8'hb0)) && {forvar1887}) ^~ $unsigned((~^(8'ha2))))};
                    end
                  if ($unsigned(reg1782[(3'h5):(2'h3)]))
                    begin
                      reg1942 <= $unsigned((&((reg1854 ?
                          reg1917 : forvar1797) & $unsigned((8'hb6)))));
                      reg1943 <= (|($unsigned($signed(reg1961)) <= $unsigned($signed((8'ha0)))));
                    end
                  else
                    begin
                      reg1942 <= {$unsigned($signed((^~reg1885)))};
                      reg1943 <= ((^~({forvar1912} || (reg1873 + wire1773))) > $signed(forvar1922[(2'h2):(1'h1)]));
                      reg1944 <= (&{forvar1834[(3'h4):(2'h3)]});
                    end
                end
              else
                begin
                  if (reg1949[(1'h0):(1'h0)])
                    begin
                      reg1937 <= reg1895[(2'h3):(1'h0)];
                      reg1938 <= $unsigned(({((8'hb1) >>> reg1804)} << $signed(reg1911[(3'h4):(2'h2)])));
                    end
                  else
                    begin
                      reg1937 <= ((^((reg1910 ~^ reg1893) ?
                          reg1803[(2'h2):(2'h2)] : (+forvar1803))) & $unsigned($unsigned($unsigned(reg1826))));
                      reg1938 <= $unsigned((reg1954 ?
                          $signed($unsigned(reg1942)) : ((8'hb5) ^~ (reg1818 ?
                              reg1787 : reg1933))));
                      reg1939 <= $signed($signed(((reg1949 >= forvar1839) ~^ $unsigned(reg1917))));
                      reg1940 <= (|$unsigned(reg1965));
                    end
                  for (forvar1941 = (1'h0); (forvar1941 < (2'h3)); forvar1941 = (forvar1941 + (1'h1)))
                    begin
                      reg1942 <= (^~(($signed(reg1787) * reg1880[(1'h0):(1'h0)]) ?
                          $signed($unsigned(reg1829)) : $unsigned($unsigned(reg1883))));
                      reg1943 <= (~^reg1941[(3'h5):(1'h1)]);
                      reg1944 <= (((|((8'ha1) - forvar1876)) ?
                          {forvar1867} : {(reg1869 ?
                                  reg1798 : reg1954)}) & (~&$signed(reg1903[(4'h8):(4'h8)])));
                    end
                  for (forvar1945 = (1'h0); (forvar1945 < (1'h0)); forvar1945 = (forvar1945 + (1'h1)))
                    begin
                      reg1946 <= (reg1901[(2'h2):(2'h2)] != {reg1782[(1'h1):(1'h0)]});
                      reg1947 <= reg1886;
                      reg1948 <= $unsigned($unsigned(($unsigned(reg1809) << reg1899)));
                      reg1949 <= {reg1945};
                    end
                end
            end
          reg1966 <= (8'hb9);
          for (forvar1967 = (1'h0); (forvar1967 < (2'h2)); forvar1967 = (forvar1967 + (1'h1)))
            begin
              for (forvar1968 = (1'h0); (forvar1968 < (2'h2)); forvar1968 = (forvar1968 + (1'h1)))
                begin
                  for (forvar1969 = (1'h0); (forvar1969 < (2'h3)); forvar1969 = (forvar1969 + (1'h1)))
                    begin
                      reg1970 <= $unsigned($signed((((8'ha8) ?
                              forvar1839 : reg1851) ?
                          (~&reg1790) : reg1812)));
                      reg1971 <= $unsigned(reg1934[(3'h7):(2'h2)]);
                    end
                  if (forvar1907)
                    begin
                      reg1972 <= $unsigned(reg1872[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1972 <= (8'ha6);
                      reg1973 <= {(^~((8'hab) >= (8'ha0)))};
                      reg1974 <= $unsigned((^~reg1789[(4'hf):(3'h4)]));
                    end
                end
              if ($signed($unsigned($unsigned($signed(reg1801)))))
                begin
                  for (forvar1975 = (1'h0); (forvar1975 < (1'h0)); forvar1975 = (forvar1975 + (1'h1)))
                    begin
                      reg1976 <= reg1931;
                      reg1977 <= $signed(($unsigned($unsigned(reg1799)) ^~ ((reg1855 && reg1886) ~^ (8'hae))));
                      reg1978 <= forvar1793[(2'h3):(2'h3)];
                      reg1979 <= reg1962[(4'hf):(4'he)];
                    end
                  for (forvar1980 = (1'h0); (forvar1980 < (2'h2)); forvar1980 = (forvar1980 + (1'h1)))
                    begin
                      reg1981 <= (~|$signed(reg1813));
                      reg1982 <= reg1879;
                    end
                  if ($signed(reg1840))
                    begin
                      reg1983 <= ({$unsigned(forvar1925[(1'h0):(1'h0)])} ?
                          $signed($signed(reg1955)) : ($signed(reg1941[(3'h4):(1'h1)]) ?
                              reg1835 : reg1899[(3'h5):(1'h0)]));
                      reg1984 <= forvar1783[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg1983 <= ($signed(forvar1805[(3'h5):(2'h2)]) ?
                          ((reg1877[(2'h3):(2'h2)] ?
                                  $unsigned(reg1833) : reg1868[(1'h1):(1'h1)]) ?
                              $unsigned($signed(forvar1788)) : reg1826[(1'h0):(1'h0)]) : $unsigned((!(+reg1787))));
                      reg1984 <= reg1919[(1'h0):(1'h0)];
                      reg1985 <= (((forvar1980[(4'ha):(3'h4)] ?
                              reg1795 : reg1873[(2'h3):(2'h3)]) ~^ (8'hb0)) ?
                          ($unsigned((-(8'hb2))) >>> (!(forvar1904 ?
                              reg1978 : reg1948))) : (~|$signed((reg1947 ?
                              reg1890 : reg1834))));
                    end
                  if (($unsigned(reg1908) || $unsigned(((forvar1809 << (8'ha6)) > $unsigned(reg1802)))))
                    begin
                      reg1986 <= $signed(($signed({(8'ha3)}) ?
                          (forvar1968[(3'h7):(3'h7)] << $unsigned((8'hb2))) : forvar1930));
                      reg1987 <= $signed($signed(reg1917));
                      reg1988 <= (8'hba);
                      reg1989 <= reg1878;
                    end
                  else
                    begin
                      reg1986 <= {((|$unsigned(forvar1802)) ?
                              $signed($unsigned(reg1977)) : (|$signed((8'h9e))))};
                      reg1987 <= forvar1925;
                      reg1988 <= (!$unsigned($unsigned($signed((8'had)))));
                    end
                end
              else
                begin
                  reg1975 <= ((reg1842 > forvar1968[(3'h4):(2'h2)]) ?
                      forvar1958[(2'h2):(1'h0)] : (-(~{(8'hac)})));
                end
              for (forvar1990 = (1'h0); (forvar1990 < (2'h3)); forvar1990 = (forvar1990 + (1'h1)))
                begin
                  for (forvar1991 = (1'h0); (forvar1991 < (2'h2)); forvar1991 = (forvar1991 + (1'h1)))
                    begin
                      reg1992 <= {$signed($signed((forvar1948 >> reg1835)))};
                      reg1993 <= $unsigned(((((8'hae) ^~ reg1961) - $unsigned(reg1849)) ?
                          $unsigned((reg1790 | reg1807)) : $signed((8'hb3))));
                      reg1994 <= $signed(forvar1805);
                      reg1995 <= $signed((reg1853[(4'ha):(4'h9)] >> (reg1863 ?
                          $unsigned(reg1910) : reg1934[(1'h1):(1'h0)])));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1996 = (1'h0); (forvar1996 < (2'h3)); forvar1996 = (forvar1996 + (1'h1)))
        begin
          for (forvar1997 = (1'h0); (forvar1997 < (2'h3)); forvar1997 = (forvar1997 + (1'h1)))
            begin
              if (reg1776)
                begin
                  for (forvar1998 = (1'h0); (forvar1998 < (1'h0)); forvar1998 = (forvar1998 + (1'h1)))
                    begin
                      reg1999 <= (+reg1933[(1'h0):(1'h0)]);
                    end
                  for (forvar2000 = (1'h0); (forvar2000 < (1'h1)); forvar2000 = (forvar2000 + (1'h1)))
                    begin
                      reg2001 <= forvar1783;
                      reg2002 <= (reg1779 ^ reg1825[(2'h3):(2'h2)]);
                      reg2003 <= ($signed((&(reg1794 <= reg1880))) ?
                          (reg1778[(4'h9):(4'h8)] ?
                              {(reg1903 ?
                                      reg1921 : wire1768)} : {$signed(reg1834)}) : reg2001[(3'h7):(3'h7)]);
                      reg2004 <= ((reg1931 ?
                              $unsigned(((8'ha0) || reg1894)) : reg1919) ?
                          ($signed(reg1891) == {forvar1948[(3'h4):(2'h2)]}) : (forvar1789 > $signed({reg1788})));
                    end
                end
              else
                begin
                  for (forvar1998 = (1'h0); (forvar1998 < (1'h0)); forvar1998 = (forvar1998 + (1'h1)))
                    begin
                      reg1999 <= forvar1824;
                    end
                end
              reg2005 <= $unsigned(forvar1912);
              if (reg1970)
                begin
                  if ((($signed((~&reg1982)) ?
                          (~^(&reg1977)) : $signed($unsigned(reg1918))) ?
                      (($unsigned(reg1920) || $signed(forvar1948)) ?
                          ({forvar1932} ?
                              $signed((8'hb6)) : (reg1891 ?
                                  reg1847 : reg1807)) : $unsigned((8'h9f))) : ({(-reg1916)} * $unsigned(reg1925))))
                    begin
                      reg2006 <= (($signed((~|forvar1805)) ?
                              ($signed(reg1841) & (+reg1853)) : {(^(8'ha2))}) ?
                          forvar2000[(3'h4):(3'h4)] : (~^($unsigned(reg1776) ?
                              (reg1908 ~^ reg1989) : ((8'hac) ?
                                  reg1952 : (8'h9d)))));
                    end
                  else
                    begin
                      reg2006 <= {(^~((reg1865 ? (8'hb4) : reg1885) ?
                              (^~reg1790) : (reg1902 ^ reg1994)))};
                      reg2007 <= ($signed($signed((&(8'had)))) ?
                          $signed({(reg1800 ?
                                  reg1959 : reg1983)}) : ({(~^(8'hb0))} && $signed($signed(reg1892))));
                      reg2008 <= ({$signed($signed(reg1903))} ?
                          reg1916[(2'h3):(2'h2)] : ($signed($signed(reg1956)) * reg1802[(3'h5):(2'h2)]));
                      reg2009 <= ($signed((8'ha9)) == forvar1958);
                    end
                  reg2010 <= (^(+$unsigned((~&reg1865))));
                  for (forvar2011 = (1'h0); (forvar2011 < (2'h3)); forvar2011 = (forvar2011 + (1'h1)))
                    begin
                      reg2012 <= forvar1776;
                      reg2013 <= {(~reg1979)};
                      reg2014 <= {forvar1857};
                    end
                  if (reg1903)
                    begin
                      reg2015 <= ({((reg2014 ?
                                  reg1840 : forvar1937) + reg2012[(2'h2):(1'h1)])} ?
                          (~forvar1839) : (+(((8'hb2) ?
                              reg1805 : reg1928) <<< (reg1905 <= forvar1914))));
                    end
                  else
                    begin
                      reg2015 <= $unsigned(reg1862[(2'h3):(1'h0)]);
                      reg2016 <= reg1942[(3'h6):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar2006 = (1'h0); (forvar2006 < (1'h0)); forvar2006 = (forvar2006 + (1'h1)))
                    begin
                      reg2007 <= $signed(($signed(reg1826) ~^ $unsigned((reg1964 ?
                          reg1983 : forvar1896))));
                      reg2008 <= (&((!(!reg1790)) ?
                          $unsigned($unsigned(reg1858)) : (reg1778 ?
                              (8'h9f) : (reg1917 - forvar1820))));
                    end
                  for (forvar2009 = (1'h0); (forvar2009 < (2'h3)); forvar2009 = (forvar2009 + (1'h1)))
                    begin
                      reg2010 <= wire1770[(2'h2):(2'h2)];
                      reg2011 <= forvar1963;
                    end
                  reg2012 <= (~|((reg1999 ?
                      reg1886 : (reg1965 >> reg1940)) ^ $unsigned({forvar1866})));
                end
              for (forvar2017 = (1'h0); (forvar2017 < (1'h1)); forvar2017 = (forvar2017 + (1'h1)))
                begin
                  for (forvar2018 = (1'h0); (forvar2018 < (1'h1)); forvar2018 = (forvar2018 + (1'h1)))
                    begin
                      reg2019 <= reg2010;
                      reg2020 <= (reg1936 ?
                          ((forvar1867 ? ((8'hb8) << reg1907) : reg1812) ?
                              ($unsigned(forvar1937) & $signed((8'ha2))) : (~|(reg2011 <= forvar1805))) : $signed(forvar1830));
                      reg2021 <= (&$signed(reg2007[(1'h1):(1'h1)]));
                    end
                end
            end
          for (forvar2022 = (1'h0); (forvar2022 < (1'h1)); forvar2022 = (forvar2022 + (1'h1)))
            begin
              for (forvar2023 = (1'h0); (forvar2023 < (1'h0)); forvar2023 = (forvar2023 + (1'h1)))
                begin
                  for (forvar2024 = (1'h0); (forvar2024 < (2'h2)); forvar2024 = (forvar2024 + (1'h1)))
                    begin
                      reg2025 <= forvar1793;
                    end
                  if (forvar1876)
                    begin
                      reg2026 <= reg1890[(1'h0):(1'h0)];
                      reg2027 <= $signed((({reg1886} ?
                              forvar2006 : $unsigned(reg1882)) ?
                          (((8'h9d) ? forvar1866 : reg2008) ?
                              reg1803 : forvar1840[(1'h0):(1'h0)]) : reg1818[(1'h0):(1'h0)]));
                      reg2028 <= ($unsigned((+$signed(forvar1914))) ?
                          (reg1903 <= {reg1783[(1'h1):(1'h1)]}) : {(~^{(8'ha7)})});
                    end
                  else
                    begin
                      reg2026 <= (($unsigned((~|forvar1904)) * $signed($unsigned(reg1835))) ?
                          {wire1773} : forvar1788);
                      reg2027 <= $unsigned($unsigned(reg1908[(2'h3):(1'h0)]));
                      reg2028 <= $signed($signed(reg1959[(4'ha):(4'ha)]));
                    end
                  for (forvar2029 = (1'h0); (forvar2029 < (2'h2)); forvar2029 = (forvar2029 + (1'h1)))
                    begin
                      reg2030 <= ((-(^~forvar1834)) ?
                          reg1921[(4'hb):(4'h8)] : $unsigned(($signed(reg1900) >> (forvar1793 >= reg1920))));
                      reg2031 <= reg2011[(2'h2):(1'h0)];
                      reg2032 <= ((((reg1815 * forvar1799) >>> reg1974) & $signed($signed((8'ha7)))) - ($signed(reg1859[(3'h5):(2'h3)]) ?
                          (+(reg1791 ? reg1999 : reg1985)) : reg1950));
                      reg2033 <= (reg1886[(1'h0):(1'h0)] <<< forvar1820);
                    end
                  for (forvar2034 = (1'h0); (forvar2034 < (1'h0)); forvar2034 = (forvar2034 + (1'h1)))
                    begin
                      reg2035 <= (~$signed($unsigned((!(8'hae)))));
                      reg2036 <= (~$signed($unsigned((forvar2022 * (8'hb7)))));
                    end
                end
              reg2037 <= reg1890;
              reg2038 <= (~^({reg1972[(2'h2):(2'h2)]} > reg1810[(4'hc):(2'h2)]));
            end
        end
      for (forvar2039 = (1'h0); (forvar2039 < (1'h0)); forvar2039 = (forvar2039 + (1'h1)))
        begin
          if ((~&(((reg1865 ? reg1782 : reg1862) ?
                  $signed((8'ha0)) : (reg1903 ? forvar1991 : reg1778)) ?
              ($unsigned(forvar1787) >> $unsigned(reg1837)) : $signed(((8'ha3) ?
                  reg2010 : reg1948)))))
            begin
              if (({($unsigned((8'hb9)) <<< forvar1991[(3'h4):(1'h0)])} ?
                  $unsigned($unsigned((forvar1806 ^ forvar1990))) : $signed(reg1782)))
                begin
                  if ($signed($unsigned({{forvar1968}})))
                    begin
                      reg2040 <= (8'hae);
                    end
                  else
                    begin
                      reg2040 <= $unsigned({(^$unsigned((8'hb1)))});
                      reg2041 <= $unsigned((({reg1872} >> reg1815[(4'hf):(3'h4)]) ?
                          ($signed(reg1882) + reg1934) : ((reg1918 ?
                                  forvar1896 : (8'ha3)) ?
                              (reg1892 ?
                                  reg2032 : (8'hb2)) : (reg1818 <= reg1822))));
                    end
                  reg2042 <= (wire1768[(3'h6):(2'h2)] ?
                      $unsigned(reg1946) : $unsigned(($signed((8'h9c)) >>> $signed(reg1958))));
                end
              else
                begin
                  for (forvar2040 = (1'h0); (forvar2040 < (1'h1)); forvar2040 = (forvar2040 + (1'h1)))
                    begin
                      reg2041 <= (~^forvar1832[(1'h1):(1'h0)]);
                      reg2042 <= (~^{((+reg1864) ?
                              (+reg2032) : $signed(forvar1776))});
                      reg2043 <= (~|reg1910);
                    end
                  if ((&$signed((-(reg1971 + reg1854)))))
                    begin
                      reg2044 <= forvar1801[(4'h9):(3'h6)];
                      reg2045 <= {$signed(((~^reg1877) ?
                              reg1872[(1'h1):(1'h1)] : reg1885[(1'h1):(1'h1)]))};
                      reg2046 <= (-$unsigned({$signed(reg1825)}));
                    end
                  else
                    begin
                      reg2044 <= (($signed($signed(forvar1914)) ?
                          (^(reg1987 ?
                              reg2007 : reg1888)) : reg1927) << $signed(({forvar2022} <= (~^forvar1925))));
                    end
                  if (forvar1927[(2'h2):(1'h0)])
                    begin
                      reg2047 <= $signed((({reg1839} ?
                          $unsigned(reg2042) : {forvar2006}) || reg1964[(2'h3):(1'h1)]));
                    end
                  else
                    begin
                      reg2047 <= (^$unsigned((~reg1873[(1'h1):(1'h0)])));
                    end
                end
            end
          else
            begin
              for (forvar2040 = (1'h0); (forvar2040 < (1'h1)); forvar2040 = (forvar2040 + (1'h1)))
                begin
                  for (forvar2041 = (1'h0); (forvar2041 < (2'h3)); forvar2041 = (forvar2041 + (1'h1)))
                    begin
                      reg2042 <= reg1909[(3'h7):(1'h0)];
                    end
                  for (forvar2043 = (1'h0); (forvar2043 < (2'h2)); forvar2043 = (forvar2043 + (1'h1)))
                    begin
                      reg2044 <= (((reg2014 <= (reg1957 || wire1770)) ?
                          $unsigned($signed(reg1881)) : $unsigned((-(8'hb5)))) - $signed($signed({reg1921})));
                      reg2045 <= {(($unsigned(reg1971) ?
                              reg2043[(4'hf):(4'h9)] : {(8'hba)}) ^~ $signed({reg1797}))};
                      reg2046 <= (~(reg1839[(4'ha):(3'h4)] || ($unsigned(reg1901) ?
                          (~forvar1839) : reg2015)));
                    end
                end
              if (forvar2043[(2'h2):(2'h2)])
                begin
                  for (forvar2047 = (1'h0); (forvar2047 < (1'h0)); forvar2047 = (forvar2047 + (1'h1)))
                    begin
                      reg2048 <= (~^($unsigned((^~forvar1904)) & reg1950[(4'h9):(1'h1)]));
                    end
                  for (forvar2049 = (1'h0); (forvar2049 < (1'h0)); forvar2049 = (forvar2049 + (1'h1)))
                    begin
                      reg2050 <= reg1975[(1'h0):(1'h0)];
                      reg2051 <= $unsigned($signed(forvar1884[(2'h3):(1'h0)]));
                      reg2052 <= forvar1896;
                    end
                  if ({(8'hb9)})
                    begin
                      reg2053 <= ((^$signed((-reg1935))) ?
                          ($signed((forvar1930 <<< reg1889)) > ($unsigned(forvar2011) ?
                              (|(8'h9f)) : reg1879)) : {(|reg1928)});
                      reg2054 <= reg2004[(2'h3):(1'h0)];
                      reg2055 <= $signed(forvar1785);
                    end
                  else
                    begin
                      reg2053 <= forvar1783;
                      reg2054 <= $signed(($signed(forvar1912[(2'h2):(1'h1)]) ?
                          reg1934 : (^forvar1789[(4'h9):(4'h9)])));
                      reg2055 <= ($signed(((reg2033 < reg2048) < (~|reg2033))) > $unsigned($signed($signed(reg1977))));
                      reg2056 <= $signed($unsigned((forvar1980 ^~ $signed((8'hb7)))));
                    end
                  for (forvar2057 = (1'h0); (forvar2057 < (1'h1)); forvar2057 = (forvar2057 + (1'h1)))
                    begin
                      reg2058 <= forvar1894;
                    end
                end
              else
                begin
                  reg2047 <= $unsigned((reg2009 << $signed({reg1979})));
                  for (forvar2048 = (1'h0); (forvar2048 < (1'h0)); forvar2048 = (forvar2048 + (1'h1)))
                    begin
                      reg2049 <= reg2011;
                      reg2050 <= (~&((reg2028 * $signed(wire1765)) - ((~^forvar1924) ?
                          {reg1956} : ((8'hb1) ^ reg2042))));
                    end
                end
              if ((({(reg1907 ? reg1851 : reg1784)} ?
                      ({reg1901} << (reg1929 > (8'hb0))) : {(-reg2054)}) ?
                  $unsigned(reg1905[(4'hd):(3'h5)]) : reg1954))
                begin
                  for (forvar2059 = (1'h0); (forvar2059 < (1'h0)); forvar2059 = (forvar2059 + (1'h1)))
                    begin
                      reg2060 <= reg2014[(4'hb):(3'h7)];
                    end
                  reg2061 <= (-(~^{((8'ha9) || reg1801)}));
                  for (forvar2062 = (1'h0); (forvar2062 < (2'h3)); forvar2062 = (forvar2062 + (1'h1)))
                    begin
                      reg2063 <= reg1952;
                    end
                end
              else
                begin
                  if (($signed($signed($unsigned((8'hb0)))) <= (&reg1923)))
                    begin
                      reg2059 <= (reg1981[(3'h7):(3'h7)] + reg2042);
                      reg2060 <= (~&(((~&forvar2062) ?
                          (reg1840 ~^ reg1811) : $unsigned(reg1899)) - $unsigned((reg1804 >>> reg1808))));
                    end
                  else
                    begin
                      reg2059 <= (~&{reg1956});
                    end
                  reg2061 <= reg1838;
                end
            end
          reg2064 <= reg1948;
        end
      if ((reg1932[(3'h7):(2'h3)] ?
          ($unsigned(forvar1955[(2'h2):(1'h1)]) && forvar1963[(1'h0):(1'h0)]) : $signed(reg1925)))
        begin
          reg2065 <= reg1933;
          reg2066 <= ({(8'hae)} ? (8'hb6) : reg2050[(4'hb):(3'h6)]);
        end
      else
        begin
          if ($unsigned(forvar1914))
            begin
              for (forvar2065 = (1'h0); (forvar2065 < (1'h1)); forvar2065 = (forvar2065 + (1'h1)))
                begin
                  reg2066 <= reg1780;
                  if ($unsigned((8'ha1)))
                    begin
                      reg2067 <= (-{reg1817});
                    end
                  else
                    begin
                      reg2067 <= $signed((~|((forvar1784 ? reg1966 : reg1793) ?
                          (forvar1799 ?
                              reg1799 : reg1999) : $unsigned(reg1797))));
                      reg2068 <= reg2004;
                    end
                end
              for (forvar2069 = (1'h0); (forvar2069 < (1'h0)); forvar2069 = (forvar2069 + (1'h1)))
                begin
                  for (forvar2070 = (1'h0); (forvar2070 < (2'h2)); forvar2070 = (forvar2070 + (1'h1)))
                    begin
                      reg2071 <= ($unsigned($signed({forvar1803})) * reg1813);
                      reg2072 <= (~|forvar1787);
                      reg2073 <= ({(-{reg1994})} | (($unsigned(forvar1894) ~^ $signed(reg1783)) + forvar1906[(1'h0):(1'h0)]));
                      reg2074 <= $unsigned(((+$unsigned((8'hb6))) ?
                          (|$unsigned(forvar2011)) : reg2068[(3'h4):(2'h2)]));
                    end
                  if (reg1958)
                    begin
                      reg2075 <= $unsigned($signed((8'ha0)));
                    end
                  else
                    begin
                      reg2075 <= forvar2009[(1'h0):(1'h0)];
                      reg2076 <= ($unsigned(reg2050) > ($signed(reg1911[(2'h2):(2'h2)]) ?
                          $signed($unsigned(forvar1802)) : forvar1917));
                      reg2077 <= $unsigned(reg1935);
                    end
                  for (forvar2078 = (1'h0); (forvar2078 < (1'h0)); forvar2078 = (forvar2078 + (1'h1)))
                    begin
                      reg2079 <= ($signed((&(8'h9f))) << (((reg1786 >= wire1767) ^ reg1960) ?
                          (~(~reg1811)) : $signed($signed(forvar1930))));
                    end
                end
              for (forvar2080 = (1'h0); (forvar2080 < (1'h1)); forvar2080 = (forvar2080 + (1'h1)))
                begin
                  reg2081 <= forvar1789[(3'h5):(3'h5)];
                  reg2082 <= $signed((forvar1794[(4'hd):(3'h5)] >= $unsigned((forvar2047 & reg1926))));
                  if ($unsigned(((reg1785[(3'h7):(2'h2)] ?
                          $unsigned((8'h9c)) : {forvar1811}) ?
                      $unsigned((forvar2048 > reg1956)) : ((reg1795 ?
                          (8'h9d) : reg2019) >>> $unsigned(reg1825)))))
                    begin
                      reg2083 <= {reg2002[(2'h2):(2'h2)]};
                    end
                  else
                    begin
                      reg2083 <= $signed((+($signed((8'hb9)) ?
                          $unsigned(wire1766) : reg1984)));
                    end
                  if (($signed($unsigned($unsigned(forvar1866))) >>> $signed(((reg2036 ?
                      forvar1912 : reg1883) + (+(8'hac))))))
                    begin
                      reg2084 <= $signed(({{reg1945}} == ((wire1771 ?
                          reg1786 : forvar1944) <<< forvar2047[(3'h5):(3'h5)])));
                      reg2085 <= $signed({(~&{reg2051})});
                      reg2086 <= (&(~&$unsigned((^~reg2006))));
                      reg2087 <= {$unsigned(reg2014[(3'h5):(2'h2)])};
                    end
                  else
                    begin
                      reg2084 <= $unsigned(forvar1780[(1'h1):(1'h1)]);
                    end
                end
            end
          else
            begin
              if ((8'ha3))
                begin
                  for (forvar2065 = (1'h0); (forvar2065 < (1'h0)); forvar2065 = (forvar2065 + (1'h1)))
                    begin
                      reg2066 <= (!(($signed(reg1918) > {reg1828}) ^~ (reg1890 <= (forvar1917 ?
                          reg1843 : reg1982))));
                      reg2067 <= (^~reg2003);
                      reg2068 <= reg1791[(1'h1):(1'h1)];
                      reg2069 <= ((|(forvar1811[(3'h7):(2'h3)] && $signed(reg2036))) || reg1891[(1'h0):(1'h0)]);
                    end
                  for (forvar2070 = (1'h0); (forvar2070 < (2'h3)); forvar2070 = (forvar2070 + (1'h1)))
                    begin
                      reg2071 <= forvar2059;
                      reg2072 <= (8'ha1);
                      reg2073 <= (reg2060 ^~ reg1995[(3'h7):(3'h5)]);
                      reg2074 <= $unsigned(((8'hb0) ?
                          ($signed((8'ha7)) > $unsigned(forvar1799)) : reg2028[(2'h2):(2'h2)]));
                    end
                  reg2075 <= ((((reg1815 <<< reg1886) * (reg1981 - reg1858)) >> (reg1945[(1'h0):(1'h0)] != (reg1893 ?
                      reg1960 : forvar2006))) > reg1985);
                end
              else
                begin
                  for (forvar2065 = (1'h0); (forvar2065 < (2'h2)); forvar2065 = (forvar2065 + (1'h1)))
                    begin
                      reg2066 <= ((8'had) ?
                          (((reg1776 ? reg1853 : reg1803) | (reg1970 ?
                                  (8'ha6) : reg2081)) ?
                              (8'hac) : ($unsigned(forvar1821) ^~ (-reg1938))) : reg2010[(2'h2):(1'h1)]);
                      reg2067 <= reg1906[(4'h8):(3'h6)];
                    end
                  reg2068 <= $signed(((^(~&reg2014)) == ((~reg2059) ?
                      {forvar2047} : $unsigned(reg2084))));
                end
              if (({$unsigned((|reg1940))} ?
                  ($unsigned($signed(forvar1980)) & forvar1874[(2'h2):(1'h0)]) : (~|((reg1994 ?
                          wire1773 : forvar1914) ?
                      (reg2001 > reg1878) : (forvar2022 ? reg1834 : (8'ha3))))))
                begin
                  for (forvar2076 = (1'h0); (forvar2076 < (2'h2)); forvar2076 = (forvar2076 + (1'h1)))
                    begin
                      reg2077 <= $unsigned(($unsigned(reg2083[(2'h2):(1'h1)]) ?
                          $unsigned($signed(reg1953)) : ((reg2036 ?
                              forvar1831 : reg2059) >> {reg1977})));
                    end
                  for (forvar2078 = (1'h0); (forvar2078 < (2'h2)); forvar2078 = (forvar2078 + (1'h1)))
                    begin
                      reg2079 <= ($signed($signed(((8'h9c) && forvar1788))) ^~ (((~&(8'h9f)) ?
                          $signed(reg1851) : $signed(reg2031)) > (~|(reg2063 && reg1849))));
                      reg2080 <= (-($signed({reg1964}) ?
                          reg1976[(1'h0):(1'h0)] : reg1836[(4'h9):(1'h0)]));
                    end
                end
              else
                begin
                  if ($signed((!{$signed(reg1906)})))
                    begin
                      reg2076 <= $signed(forvar1838[(2'h3):(2'h2)]);
                      reg2077 <= forvar1937;
                    end
                  else
                    begin
                      reg2076 <= {reg1994};
                      reg2077 <= $unsigned(forvar1838);
                      reg2078 <= $signed((&forvar1832[(1'h1):(1'h0)]));
                      reg2079 <= reg1805;
                    end
                  for (forvar2080 = (1'h0); (forvar2080 < (1'h1)); forvar2080 = (forvar2080 + (1'h1)))
                    begin
                      reg2081 <= (($signed(reg1979) ?
                              reg1966 : $unsigned($signed(reg2075))) ?
                          $signed({(forvar2048 ?
                                  reg1787 : reg1954)}) : ($signed(reg2030[(2'h3):(1'h1)]) ?
                              (~&$unsigned(reg2012)) : ((reg2010 > forvar2048) != forvar2049[(1'h0):(1'h0)])));
                    end
                  reg2082 <= forvar1806[(1'h0):(1'h0)];
                  for (forvar2083 = (1'h0); (forvar2083 < (1'h1)); forvar2083 = (forvar2083 + (1'h1)))
                    begin
                      reg2084 <= {($signed(reg1919) ?
                              reg2010[(2'h2):(1'h0)] : reg1948[(4'hd):(4'hd)])};
                      reg2085 <= (forvar1799[(1'h1):(1'h0)] ?
                          (-$unsigned((reg1803 ?
                              (8'ha9) : (8'ha8)))) : (8'h9d));
                      reg2086 <= (-($unsigned($unsigned(forvar1783)) ?
                          ((forvar1803 ? (8'ha0) : reg1780) ?
                              (reg1914 << forvar1940) : reg2046) : {(^reg2083)}));
                      reg2087 <= reg1878;
                    end
                end
            end
          if ($signed(forvar1905[(4'h9):(1'h0)]))
            begin
              for (forvar2088 = (1'h0); (forvar2088 < (2'h2)); forvar2088 = (forvar2088 + (1'h1)))
                begin
                  for (forvar2089 = (1'h0); (forvar2089 < (2'h2)); forvar2089 = (forvar2089 + (1'h1)))
                    begin
                      reg2090 <= (forvar1784 ?
                          reg1907[(1'h1):(1'h0)] : reg1816);
                      reg2091 <= {{$signed(((8'hb9) ? reg1797 : forvar2041))}};
                      reg2092 <= (!$unsigned(forvar1894));
                      reg2093 <= {((forvar1780[(2'h3):(1'h0)] ?
                              {reg1966} : (8'ha7)) > $unsigned(((8'ha6) ?
                              forvar1912 : reg1803)))};
                    end
                  reg2094 <= (^$unsigned((-reg1840[(4'h8):(3'h5)])));
                  if ((8'hab))
                    begin
                      reg2095 <= (-$unsigned($unsigned($unsigned(reg1989))));
                      reg2096 <= ({{$unsigned(reg1802)}} ?
                          forvar1887[(1'h1):(1'h0)] : reg1907[(2'h2):(2'h2)]);
                      reg2097 <= reg2064[(3'h5):(3'h5)];
                      reg2098 <= reg1939[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg2095 <= ($unsigned($signed((-reg1827))) ^~ {(|(reg1944 ?
                              (8'h9f) : reg2075))});
                      reg2096 <= ($unsigned($unsigned($unsigned(reg1880))) ?
                          {reg1800[(4'he):(4'h8)]} : ((forvar2089[(4'h8):(1'h0)] ?
                                  $unsigned(reg2001) : (forvar1940 ?
                                      reg1917 : reg1787)) ?
                              {$unsigned(wire1773)} : $unsigned($unsigned(reg2001))));
                      reg2097 <= forvar2041;
                    end
                  reg2099 <= ($signed($signed((forvar1801 ?
                      reg1789 : forvar1969))) >>> {$unsigned($signed(reg1933))});
                end
              for (forvar2100 = (1'h0); (forvar2100 < (2'h3)); forvar2100 = (forvar2100 + (1'h1)))
                begin
                  if ($signed((|$unsigned({reg1795}))))
                    begin
                      reg2101 <= (reg2015 < $unsigned({forvar1801}));
                      reg2102 <= ($signed((forvar1907 ?
                              wire1770 : $signed(forvar1958))) ?
                          reg2068[(3'h6):(2'h3)] : (8'hb3));
                    end
                  else
                    begin
                      reg2101 <= $signed(($unsigned(forvar1894) && (reg1868 ?
                          (reg2082 ?
                              reg1986 : reg2021) : reg1813[(5'h10):(3'h5)])));
                    end
                end
              reg2103 <= {($signed({reg1860}) < $signed(reg1878[(4'hc):(3'h7)]))};
              for (forvar2104 = (1'h0); (forvar2104 < (2'h2)); forvar2104 = (forvar2104 + (1'h1)))
                begin
                  if (reg2032)
                    begin
                      reg2105 <= $unsigned($signed({reg2077}));
                      reg2106 <= ({reg1975} + {($signed((8'hae)) | (~^(8'ha3)))});
                      reg2107 <= $unsigned($signed(((~^reg1802) - (~&reg1902))));
                      reg2108 <= reg1795[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2105 <= reg2052;
                      reg2106 <= $signed(forvar1996[(3'h4):(1'h0)]);
                      reg2107 <= ($signed(((+reg2091) ^~ (forvar1967 ?
                          (8'h9f) : (8'h9e)))) | (($signed(reg2063) ^~ $unsigned(reg1989)) ~^ $signed($signed(reg1799))));
                    end
                  for (forvar2109 = (1'h0); (forvar2109 < (2'h3)); forvar2109 = (forvar2109 + (1'h1)))
                    begin
                      reg2110 <= (~&(|(reg2107 ?
                          (forvar1990 >= reg1892) : (&(8'hb8)))));
                      reg2111 <= reg1800[(4'hc):(1'h1)];
                      reg2112 <= ({$signed({reg1939})} && reg2045[(2'h2):(1'h1)]);
                      reg2113 <= $signed((reg1893 ?
                          reg1917 : ($signed(reg1841) >>> $signed(reg1924))));
                    end
                  for (forvar2114 = (1'h0); (forvar2114 < (2'h2)); forvar2114 = (forvar2114 + (1'h1)))
                    begin
                      reg2115 <= (8'hb0);
                      reg2116 <= (((&$signed(forvar1801)) ?
                          reg1862 : reg1783) && $unsigned((~^$unsigned(reg1858))));
                      reg2117 <= ((~$signed(reg2055[(4'h8):(3'h4)])) & forvar1990[(1'h1):(1'h0)]);
                      reg2118 <= (($unsigned($unsigned(reg1816)) & (reg1981[(2'h3):(1'h1)] ?
                          $signed((8'hb8)) : $signed(forvar1785))) << ($signed(forvar1794[(4'he):(3'h7)]) ?
                          reg1905[(4'h9):(3'h5)] : $unsigned(reg2066[(1'h1):(1'h1)])));
                    end
                  reg2119 <= ((($signed(reg2044) ?
                          $unsigned(reg2112) : reg2038[(4'hc):(4'h8)]) ^ {(~|reg2092)}) ?
                      (reg1779[(3'h7):(3'h6)] ^ reg1790) : ({(forvar2024 <= forvar1905)} <<< reg2015));
                end
            end
          else
            begin
              reg2088 <= $signed($unsigned($signed((reg1960 < (8'h9d)))));
            end
        end
    end
  assign wire2120 = (8'hba);
  assign wire2121 = (+$signed((&(^~reg2071))));
  module2122 modinst2583 (wire2582, clk, reg1895, reg2048, reg1927, forvar1867);
  assign wire2584 = ($signed((reg2015 ?
                        (|forvar1775) : (8'haf))) | ($signed({forvar1801}) <<< $unsigned({forvar1783})));
  assign wire2585 = {$signed((!forvar1845))};
  always
    @(posedge clk) begin
      for (forvar2586 = (1'h0); (forvar2586 < (1'h1)); forvar2586 = (forvar2586 + (1'h1)))
        begin
          for (forvar2587 = (1'h0); (forvar2587 < (2'h2)); forvar2587 = (forvar2587 + (1'h1)))
            begin
              if ($unsigned((8'hac)))
                begin
                  for (forvar2588 = (1'h0); (forvar2588 < (1'h0)); forvar2588 = (forvar2588 + (1'h1)))
                    begin
                      reg2589 <= ((^~((forvar1839 ?
                              forvar2049 : reg1892) ^~ reg2098)) ?
                          {$unsigned(forvar1991)} : forvar1794);
                      reg2590 <= $unsigned((~&(reg2058 ? {reg2077} : reg2002)));
                    end
                end
              else
                begin
                  if ((reg1811 ?
                      ($unsigned((reg1823 >= reg1799)) ^~ (~|$unsigned(forvar1917))) : (reg2073 <<< $signed({reg1956}))))
                    begin
                      reg2588 <= (~(($unsigned(forvar2041) * reg2033) ?
                          {(forvar1839 ^~ reg2016)} : ({reg2037} <<< reg1974)));
                      reg2589 <= $signed((8'ha9));
                    end
                  else
                    begin
                      reg2588 <= $unsigned($unsigned(reg1881[(1'h0):(1'h0)]));
                    end
                  for (forvar2590 = (1'h0); (forvar2590 < (2'h2)); forvar2590 = (forvar2590 + (1'h1)))
                    begin
                      reg2591 <= reg2055[(3'h4):(3'h4)];
                      reg2592 <= ($unsigned((wire1765[(2'h3):(2'h2)] ?
                          ((8'h9c) ? reg2026 : reg1914) : (wire2121 ?
                              forvar1834 : reg2015))) ~^ $unsigned(forvar1857[(2'h2):(1'h0)]));
                    end
                  if (reg1977[(2'h2):(1'h0)])
                    begin
                      reg2593 <= {$unsigned(($signed(reg2044) * $signed(reg2105)))};
                      reg2594 <= $signed((8'ha1));
                    end
                  else
                    begin
                      reg2593 <= ((^(reg1888[(1'h0):(1'h0)] ?
                          $signed(forvar2059) : (~|reg1898))) != reg1796[(1'h0):(1'h0)]);
                      reg2594 <= $unsigned({reg1881[(4'hf):(1'h1)]});
                    end
                end
              for (forvar2595 = (1'h0); (forvar2595 < (1'h0)); forvar2595 = (forvar2595 + (1'h1)))
                begin
                  for (forvar2596 = (1'h0); (forvar2596 < (2'h3)); forvar2596 = (forvar2596 + (1'h1)))
                    begin
                      reg2597 <= (reg2073 + (({reg2007} ?
                              reg1952 : forvar2047) ?
                          $unsigned($unsigned(reg1960)) : {$signed(reg1806)}));
                      reg2598 <= (~&(forvar1824 ?
                          (forvar2114 ?
                              {forvar1905} : (8'hb7)) : {(&forvar1945)}));
                      reg2599 <= {reg1841[(3'h4):(1'h1)]};
                    end
                end
              for (forvar2600 = (1'h0); (forvar2600 < (1'h1)); forvar2600 = (forvar2600 + (1'h1)))
                begin
                  if (forvar2022)
                    begin
                      reg2601 <= ($signed($unsigned((reg2108 != forvar1803))) & (reg1934 <= reg1861));
                    end
                  else
                    begin
                      reg2601 <= $signed((reg1966[(1'h1):(1'h0)] ?
                          wire2582 : (forvar1793[(1'h0):(1'h0)] > $unsigned(reg1939))));
                      reg2602 <= {(8'h9e)};
                      reg2603 <= (^~{reg2597[(3'h5):(2'h3)]});
                      reg2604 <= ((reg1784 ?
                          $unsigned($signed(reg1784)) : (~(forvar1784 ?
                              reg2591 : reg2044))) ^ (reg1908 < reg2028[(3'h6):(3'h6)]));
                    end
                  reg2605 <= reg1940[(3'h4):(1'h1)];
                  if ((+((~&(~&(8'hae))) - $signed((reg1941 >>> reg1856)))))
                    begin
                      reg2606 <= reg1854[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg2606 <= (($signed(reg1954) ?
                          reg1890[(1'h0):(1'h0)] : (~(~(8'ha3)))) && ((wire2584 <<< (reg1900 * reg2069)) ?
                          reg1989 : $unsigned((+(8'hb4)))));
                    end
                  if (((($unsigned(reg1836) ?
                              (~^reg1848) : (reg1934 <<< forvar2018)) ?
                          reg2020[(2'h2):(2'h2)] : $unsigned(forvar1925[(3'h5):(2'h2)])) ?
                      $signed(reg1788) : (8'hb7)))
                    begin
                      reg2607 <= $unsigned($signed($unsigned(forvar1967)));
                      reg2608 <= (((reg1860[(4'h9):(3'h5)] ?
                          $unsigned(reg1805) : $unsigned(reg2013)) + (reg1888 * (8'ha3))) ~^ ($signed(forvar1990[(2'h2):(1'h1)]) > ($unsigned(reg1883) >= reg1913)));
                      reg2609 <= ((8'ha6) << {(reg1916 ?
                              reg1844[(3'h6):(1'h0)] : (reg1783 ?
                                  reg1886 : forvar2104))});
                    end
                  else
                    begin
                      reg2607 <= {wire1768};
                      reg2608 <= $unsigned($signed($unsigned((~&wire2585))));
                      reg2609 <= reg1840;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar2610 = (1'h0); (forvar2610 < (2'h2)); forvar2610 = (forvar2610 + (1'h1)))
        begin
          for (forvar2611 = (1'h0); (forvar2611 < (2'h2)); forvar2611 = (forvar2611 + (1'h1)))
            begin
              for (forvar2612 = (1'h0); (forvar2612 < (2'h3)); forvar2612 = (forvar2612 + (1'h1)))
                begin
                  reg2613 <= ($unsigned($signed($unsigned(reg2076))) && (8'hb2));
                  for (forvar2614 = (1'h0); (forvar2614 < (1'h0)); forvar2614 = (forvar2614 + (1'h1)))
                    begin
                      reg2615 <= ((((|forvar1874) << (^~forvar1975)) ?
                          {(&reg2009)} : (reg2014 ?
                              (forvar1776 * reg1840) : forvar1920[(2'h3):(1'h1)])) >= (wire1771[(2'h3):(2'h3)] < ((~|reg2063) ?
                          (reg1865 <= forvar1924) : (reg1946 <= (8'hb0)))));
                      reg2616 <= (8'hb7);
                      reg2617 <= {$signed(reg2117)};
                    end
                  reg2618 <= (-($signed({reg1894}) ?
                      ((-(8'hba)) ?
                          forvar2009[(2'h3):(1'h1)] : reg1865) : ((~^reg2096) ?
                          (8'ha6) : $signed(reg1786))));
                  if ({$unsigned(((-forvar1945) >>> {reg2118}))})
                    begin
                      reg2619 <= ((^$unsigned(forvar2109[(1'h1):(1'h0)])) | ($signed(((8'haa) ?
                              reg1808 : reg1843)) ?
                          $signed(((8'ha1) == reg1901)) : (~|$unsigned(reg2604))));
                    end
                  else
                    begin
                      reg2619 <= reg1995;
                      reg2620 <= (&forvar1840);
                      reg2621 <= (~&$unsigned((((8'hb8) == forvar1780) ?
                          $unsigned((8'ha9)) : (|forvar2009))));
                      reg2622 <= {reg1919[(2'h2):(1'h1)]};
                    end
                end
              reg2623 <= forvar1788;
            end
        end
      for (forvar2624 = (1'h0); (forvar2624 < (1'h1)); forvar2624 = (forvar2624 + (1'h1)))
        begin
          reg2625 <= {reg2603};
          if ((8'hb6))
            begin
              if (($unsigned((|forvar1968[(3'h4):(2'h3)])) ?
                  (!(reg1924 ?
                      reg1812[(3'h4):(2'h3)] : (reg1986 ?
                          (8'hb3) : (8'hb5)))) : (!(~forvar1975))))
                begin
                  for (forvar2626 = (1'h0); (forvar2626 < (2'h2)); forvar2626 = (forvar2626 + (1'h1)))
                    begin
                      reg2627 <= reg1961[(3'h4):(2'h3)];
                    end
                  reg2628 <= $signed(({(&forvar2059)} ?
                      $unsigned($unsigned(reg1986)) : $unsigned((~^reg2006))));
                  for (forvar2629 = (1'h0); (forvar2629 < (2'h2)); forvar2629 = (forvar2629 + (1'h1)))
                    begin
                      reg2630 <= (((+(+(8'hae))) != $unsigned((-(8'hb1)))) ?
                          (($signed(reg1806) ?
                                  (^~wire1769) : $unsigned(reg2028)) ?
                              (wire1769[(2'h2):(1'h1)] <<< (^reg1871)) : ((&(8'ha5)) ?
                                  reg2616[(3'h4):(2'h2)] : ((8'ha8) ?
                                      (8'ha5) : (8'hb7)))) : ((~{reg2040}) ?
                              reg2067[(3'h4):(2'h2)] : ({(8'hb1)} ?
                                  forvar1801[(2'h2):(2'h2)] : (~(8'hab)))));
                    end
                  for (forvar2631 = (1'h0); (forvar2631 < (2'h3)); forvar2631 = (forvar2631 + (1'h1)))
                    begin
                      reg2632 <= reg1871;
                      reg2633 <= ((^~$unsigned((-reg1790))) ^ (!reg2004[(3'h6):(3'h4)]));
                      reg2634 <= ($signed($unsigned((forvar1990 - reg1835))) - (~&reg2083[(1'h0):(1'h0)]));
                      reg2635 <= (reg2621[(3'h7):(1'h0)] ~^ (reg1994 ?
                          ($unsigned(reg2615) ?
                              (reg1797 ?
                                  reg2069 : (8'hae)) : $unsigned(reg2075)) : $signed({reg2072})));
                    end
                end
              else
                begin
                  reg2626 <= $signed(forvar2057[(3'h5):(3'h5)]);
                  for (forvar2627 = (1'h0); (forvar2627 < (1'h1)); forvar2627 = (forvar2627 + (1'h1)))
                    begin
                      reg2628 <= wire2582;
                      reg2629 <= {(^($unsigned((8'h9f)) < ((8'haf) >= reg1940)))};
                      reg2630 <= forvar1998;
                    end
                  reg2631 <= $unsigned($unsigned($signed($unsigned(reg1819))));
                  reg2632 <= forvar1958;
                end
              reg2636 <= $signed(((~^(reg2004 ? forvar1922 : reg1784)) ?
                  $signed($signed((8'hb8))) : ($signed(forvar2039) >>> $unsigned(reg2096))));
              reg2637 <= ($unsigned(reg1959) ?
                  ($signed({reg1827}) ?
                      ($signed(forvar1832) ?
                          reg2007 : (-reg1862)) : (~&reg1889[(3'h4):(1'h0)])) : $signed($unsigned((forvar1969 ?
                      forvar1945 : reg2047))));
              reg2638 <= forvar2011;
            end
          else
            begin
              for (forvar2626 = (1'h0); (forvar2626 < (2'h2)); forvar2626 = (forvar2626 + (1'h1)))
                begin
                  if ($unsigned(({wire2585[(3'h5):(3'h5)]} ?
                      $unsigned((!reg2635)) : (^~reg1979[(4'h8):(3'h6)]))))
                    begin
                      reg2627 <= {forvar2041};
                      reg2628 <= wire2120[(2'h2):(1'h1)];
                      reg2629 <= (~|forvar1925);
                    end
                  else
                    begin
                      reg2627 <= (!($signed((8'hb6)) ?
                          $unsigned((reg1810 && reg2066)) : reg2035));
                      reg2628 <= {(forvar2587[(3'h6):(3'h5)] << $signed((reg2599 ?
                              (8'hb7) : forvar2600)))};
                    end
                  for (forvar2630 = (1'h0); (forvar2630 < (1'h0)); forvar2630 = (forvar2630 + (1'h1)))
                    begin
                      reg2631 <= ((&reg1940[(2'h2):(1'h1)]) < reg2622[(3'h4):(1'h1)]);
                    end
                end
              if ($unsigned($unsigned($unsigned($unsigned(forvar2078)))))
                begin
                  for (forvar2632 = (1'h0); (forvar2632 < (2'h3)); forvar2632 = (forvar2632 + (1'h1)))
                    begin
                      reg2633 <= (reg1934 & reg1942);
                      reg2634 <= reg1954[(2'h2):(1'h1)];
                      reg2635 <= reg2621;
                    end
                  if ($signed(forvar2629[(2'h2):(1'h1)]))
                    begin
                      reg2636 <= ($unsigned(reg2096[(1'h1):(1'h1)]) ?
                          $signed($signed($unsigned(reg2055))) : ({(forvar1887 < reg1823)} ?
                              $unsigned(forvar1980[(4'hd):(4'hb)]) : reg1782[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg2636 <= ($signed(((reg1917 && reg1906) <<< $signed(wire1770))) > {((forvar2600 ?
                                  forvar1785 : reg2064) ?
                              $signed(reg1947) : $unsigned((8'h9d)))});
                      reg2637 <= forvar1937[(1'h0):(1'h0)];
                      reg2638 <= reg1924[(3'h4):(1'h1)];
                    end
                  reg2639 <= reg1783;
                  for (forvar2640 = (1'h0); (forvar2640 < (2'h2)); forvar2640 = (forvar2640 + (1'h1)))
                    begin
                      reg2641 <= (8'h9c);
                      reg2642 <= (!(~&(reg1972[(3'h4):(3'h4)] ?
                          $unsigned(reg1852) : reg1782[(1'h0):(1'h0)])));
                      reg2643 <= ($signed((reg2047 ?
                              reg1882 : $unsigned(forvar2629))) ?
                          (reg1822[(1'h1):(1'h0)] && ((reg2117 ?
                                  (8'ha6) : reg2009) ?
                              forvar1913[(4'h8):(2'h3)] : forvar1787)) : $unsigned($signed($unsigned(reg1945))));
                      reg2644 <= (wire1768 ?
                          reg2601 : $signed((~^(wire1769 ?
                              (8'hb6) : (8'ha1)))));
                    end
                end
              else
                begin
                  reg2632 <= $signed($unsigned(((!(8'hb4)) ^~ (reg1920 ?
                      reg1849 : forvar2024))));
                  reg2633 <= (&reg1823[(3'h5):(1'h0)]);
                  if (((^$unsigned(reg2044[(1'h1):(1'h1)])) <<< $unsigned($unsigned({forvar1907}))))
                    begin
                      reg2634 <= ((&(^~(~|(8'ha3)))) ? forvar1840 : reg1957);
                      reg2635 <= $signed(reg1898);
                      reg2636 <= forvar1845;
                    end
                  else
                    begin
                      reg2634 <= reg2065;
                      reg2635 <= $signed($unsigned(reg1889[(3'h4):(2'h2)]));
                    end
                  if ($signed($signed(reg1879[(2'h2):(1'h1)])))
                    begin
                      reg2637 <= $signed($unsigned((|(reg1822 || (8'hae)))));
                      reg2638 <= ((+((|forvar1887) ?
                          (reg2105 ?
                              reg2036 : forvar1776) : $unsigned(reg2635))) >= reg2101);
                      reg2639 <= reg1905[(4'ha):(2'h2)];
                    end
                  else
                    begin
                      reg2637 <= ({$unsigned((!(8'h9c)))} ?
                          (($unsigned(reg2083) ?
                              (-reg2069) : (forvar1874 ?
                                  reg1899 : forvar2011)) ~^ (forvar2630 ?
                              $unsigned((8'hab)) : $unsigned(reg1893))) : reg2088);
                    end
                end
            end
          for (forvar2645 = (1'h0); (forvar2645 < (1'h0)); forvar2645 = (forvar2645 + (1'h1)))
            begin
              if ((($signed($unsigned(forvar1904)) & (forvar1824[(1'h0):(1'h0)] >= wire1765)) ?
                  (($unsigned(reg2010) != (reg2117 ?
                      reg1929 : reg2613)) == (~$signed((8'hb8)))) : {$signed($signed(reg1964))}))
                begin
                  for (forvar2646 = (1'h0); (forvar2646 < (2'h3)); forvar2646 = (forvar2646 + (1'h1)))
                    begin
                      reg2647 <= forvar2088;
                      reg2648 <= $unsigned($unsigned($unsigned(reg2014[(4'h8):(3'h7)])));
                      reg2649 <= $signed(($signed(reg1928[(1'h1):(1'h0)]) | $unsigned($unsigned(reg1942))));
                    end
                  for (forvar2650 = (1'h0); (forvar2650 < (2'h2)); forvar2650 = (forvar2650 + (1'h1)))
                    begin
                      reg2651 <= $signed($unsigned($unsigned((~^reg1934))));
                      reg2652 <= reg1941;
                      reg2653 <= ($unsigned(forvar2000) != ($unsigned($signed(reg1891)) & $unsigned($signed(forvar2000))));
                      reg2654 <= reg1790;
                    end
                  for (forvar2655 = (1'h0); (forvar2655 < (1'h0)); forvar2655 = (forvar2655 + (1'h1)))
                    begin
                      reg2656 <= ($unsigned((~^(|reg1945))) << ($unsigned($unsigned(reg2037)) ?
                          $signed((reg1792 ?
                              reg1778 : forvar2631)) : $signed(((8'ha4) ?
                              reg2054 : (8'haf)))));
                      reg2657 <= (($signed($unsigned(forvar2630)) * $unsigned((&forvar1803))) * (~^(((8'hb1) & reg1949) < $unsigned(forvar1905))));
                      reg2658 <= (!{reg1840[(2'h2):(1'h1)]});
                    end
                end
              else
                begin
                  for (forvar2646 = (1'h0); (forvar2646 < (2'h2)); forvar2646 = (forvar2646 + (1'h1)))
                    begin
                      reg2647 <= forvar2059;
                      reg2648 <= $signed($signed({$unsigned(reg2007)}));
                    end
                  for (forvar2649 = (1'h0); (forvar2649 < (1'h1)); forvar2649 = (forvar2649 + (1'h1)))
                    begin
                      reg2650 <= $unsigned($unsigned(forvar2009));
                      reg2651 <= reg2030;
                    end
                  if (forvar1876[(1'h0):(1'h0)])
                    begin
                      reg2652 <= $unsigned($unsigned(($unsigned(reg1985) ?
                          reg1921[(3'h7):(1'h1)] : forvar1785)));
                      reg2653 <= (forvar2649 & ($unsigned(reg1863) < {reg2045}));
                      reg2654 <= reg2602[(3'h6):(3'h6)];
                    end
                  else
                    begin
                      reg2652 <= ({$signed({forvar1803})} ?
                          $signed(($unsigned((8'hb3)) ?
                              reg1783 : $signed(reg1851))) : (($unsigned(reg2630) << $unsigned(reg2032)) < forvar1783));
                    end
                end
              if (reg1905)
                begin
                  for (forvar2659 = (1'h0); (forvar2659 < (2'h2)); forvar2659 = (forvar2659 + (1'h1)))
                    begin
                      reg2660 <= reg2076;
                      reg2661 <= (~|((~|reg1904) * reg2012));
                      reg2662 <= ($signed($signed(reg2598)) ?
                          ($signed(forvar1801) >>> (8'hb6)) : reg1950);
                      reg2663 <= (~^reg1914[(2'h2):(1'h1)]);
                    end
                end
              else
                begin
                  reg2659 <= reg1929;
                end
            end
          reg2664 <= $unsigned(reg2639[(4'hd):(4'hc)]);
        end
      if (($unsigned((!$signed((8'hb7)))) - (forvar2076 - ($unsigned(forvar2624) ~^ $signed(forvar1811)))))
        begin
          if (reg1865)
            begin
              for (forvar2665 = (1'h0); (forvar2665 < (1'h1)); forvar2665 = (forvar2665 + (1'h1)))
                begin
                  for (forvar2666 = (1'h0); (forvar2666 < (1'h0)); forvar2666 = (forvar2666 + (1'h1)))
                    begin
                      reg2667 <= (!({(forvar2650 ^ (8'ha8))} | {forvar1783}));
                    end
                  for (forvar2668 = (1'h0); (forvar2668 < (2'h3)); forvar2668 = (forvar2668 + (1'h1)))
                    begin
                      reg2669 <= (!($unsigned(((8'hab) ?
                          reg2091 : reg1975)) ~^ $unsigned((!reg2107))));
                      reg2670 <= reg1902[(1'h0):(1'h0)];
                      reg2671 <= (|$unsigned(((forvar1793 < (8'haa)) ^~ $signed(reg1989))));
                      reg2672 <= (~&(((wire1765 <= (8'h9c)) ?
                          (reg1899 ?
                              forvar2062 : reg2080) : (~^reg2081)) + (^~$unsigned(reg1781))));
                    end
                  for (forvar2673 = (1'h0); (forvar2673 < (2'h2)); forvar2673 = (forvar2673 + (1'h1)))
                    begin
                      reg2674 <= (!reg2592[(1'h1):(1'h1)]);
                      reg2675 <= forvar1780;
                    end
                end
              for (forvar2676 = (1'h0); (forvar2676 < (2'h2)); forvar2676 = (forvar2676 + (1'h1)))
                begin
                  if (reg1806)
                    begin
                      reg2677 <= (~((reg1859 ?
                              (~^reg1860) : $unsigned(forvar2109)) ?
                          {$signed((8'ha8))} : {((8'hb1) ?
                                  reg2598 : reg2099)}));
                    end
                  else
                    begin
                      reg2677 <= $signed($signed((reg1978 >> reg1885)));
                      reg2678 <= reg2113;
                    end
                  if (((forvar1780 ?
                      (reg1843 <= (forvar2057 ?
                          reg2117 : reg1868)) : reg2660) > (($unsigned(reg2013) ?
                      (~^forvar2104) : (+forvar1838)) != ($unsigned(wire1773) ?
                      reg2075 : ((8'hb0) >= forvar2089)))))
                    begin
                      reg2679 <= $unsigned((8'hba));
                    end
                  else
                    begin
                      reg2679 <= $signed($signed((forvar1990 ?
                          (reg2042 ?
                              reg1946 : reg2075) : reg1942[(3'h4):(2'h2)])));
                    end
                  if ({(({forvar2645} & $signed(reg1782)) ?
                          $unsigned({(8'hb2)}) : ($signed(reg1777) << $signed(reg2092)))})
                    begin
                      reg2680 <= $unsigned((forvar2059[(4'h8):(3'h4)] ?
                          {$signed(reg2675)} : ((reg1909 ? (8'hba) : (8'h9f)) ?
                              $unsigned(reg2108) : (reg1913 ?
                                  reg2056 : forvar2057))));
                      reg2681 <= (reg1858 && $unsigned((reg2026[(3'h4):(2'h3)] << {reg1777})));
                    end
                  else
                    begin
                      reg2680 <= {forvar1821};
                      reg2681 <= reg1851;
                      reg2682 <= reg1856;
                    end
                  for (forvar2683 = (1'h0); (forvar2683 < (1'h0)); forvar2683 = (forvar2683 + (1'h1)))
                    begin
                      reg2684 <= $unsigned({((^~reg2006) + $unsigned(reg1937))});
                      reg2685 <= ((|$signed({reg1910})) ^ $signed((^~$signed(wire1766))));
                      reg2686 <= {(forvar2011[(2'h3):(2'h3)] + $unsigned((forvar2006 ^ reg1810)))};
                      reg2687 <= (8'ha8);
                    end
                end
              for (forvar2688 = (1'h0); (forvar2688 < (1'h1)); forvar2688 = (forvar2688 + (1'h1)))
                begin
                  if ($unsigned((forvar2100[(4'hf):(3'h7)] <<< $unsigned((|reg1975)))))
                    begin
                      reg2689 <= $signed((~|$signed(wire1770[(4'h9):(3'h4)])));
                      reg2690 <= $unsigned(($signed((^~(8'hb1))) & reg2001[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg2689 <= $unsigned((reg2021 ?
                          $signed($signed(forvar1787)) : ((forvar2109 ?
                              (8'ha5) : reg1826) | (8'hb8))));
                      reg2690 <= forvar1789;
                      reg2691 <= (^$unsigned($signed((~|reg2661))));
                    end
                end
              reg2692 <= forvar2596[(1'h0):(1'h0)];
            end
          else
            begin
              for (forvar2665 = (1'h0); (forvar2665 < (2'h3)); forvar2665 = (forvar2665 + (1'h1)))
                begin
                  if (reg1895[(2'h2):(2'h2)])
                    begin
                      reg2666 <= reg2682[(4'ha):(4'ha)];
                    end
                  else
                    begin
                      reg2666 <= (&$unsigned($unsigned($unsigned(forvar1876))));
                      reg2667 <= forvar1927;
                    end
                end
              if ({reg2049[(2'h3):(2'h3)]})
                begin
                  reg2668 <= $signed(forvar1884[(1'h1):(1'h0)]);
                end
              else
                begin
                  if (((({reg1957} ^~ ((8'had) ?
                      reg1913 : forvar2668)) ~^ $signed($unsigned(reg1785))) | reg2642))
                    begin
                      reg2668 <= ($signed($unsigned((reg1904 ?
                          reg1935 : forvar1967))) + reg2032);
                      reg2669 <= ((reg1925[(2'h2):(1'h0)] * $unsigned({forvar2673})) ?
                          (^~((~^reg2650) ?
                              (forvar1998 ?
                                  forvar2059 : reg2098) : $signed(reg1859))) : $unsigned($signed((&reg1880))));
                      reg2670 <= (!((^~((8'hb3) ? reg1826 : reg2021)) ?
                          (!(~^reg1809)) : reg2630[(3'h4):(2'h3)]));
                      reg2671 <= ((($unsigned(reg2093) ~^ (forvar1802 ~^ (8'ha5))) ?
                          ({reg2662} ?
                              (-reg2639) : $unsigned(reg1833)) : $unsigned($unsigned(reg2005))) >>> (&(~|(~|(8'ha4)))));
                    end
                  else
                    begin
                      reg2668 <= ($signed({(reg2093 ? forvar1924 : reg2077)}) ?
                          (($signed(reg1891) || (!reg2634)) ?
                              (8'hb3) : ($unsigned(reg1948) != $signed(forvar1991))) : reg2006[(3'h6):(1'h0)]);
                      reg2669 <= (forvar2069[(4'h8):(3'h4)] ?
                          $signed((~reg2633[(1'h0):(1'h0)])) : (~&$signed(((8'h9c) ?
                              reg2074 : reg2689))));
                    end
                  if ((&$signed({{reg1921}})))
                    begin
                      reg2672 <= ((reg2629[(2'h2):(1'h0)] ?
                          ((forvar1998 != reg1897) != ((8'hb6) ?
                              reg1873 : reg1796)) : $signed((forvar2062 == (8'h9d)))) << $signed($unsigned((~^(8'hb6)))));
                      reg2673 <= $signed($unsigned({$signed(reg1861)}));
                      reg2674 <= (({(reg1901 * reg1960)} ?
                          (&(forvar2631 ?
                              (8'hb3) : forvar1920)) : (8'hab)) & reg2690[(3'h7):(1'h1)]);
                    end
                  else
                    begin
                      reg2672 <= ((-((^~forvar1834) > ((8'hac) << (8'haf)))) ?
                          (forvar2076 > (reg2625[(3'h4):(1'h1)] ?
                              {reg1848} : $unsigned(reg1964))) : (~|(wire1769[(3'h7):(1'h0)] ^~ (8'ha5))));
                    end
                  for (forvar2675 = (1'h0); (forvar2675 < (2'h3)); forvar2675 = (forvar2675 + (1'h1)))
                    begin
                      reg2676 <= $signed($signed({reg2021}));
                      reg2677 <= forvar2586[(1'h0):(1'h0)];
                      reg2678 <= (^~forvar1867[(4'hb):(2'h2)]);
                    end
                  if ($signed($unsigned((~^reg1802))))
                    begin
                      reg2679 <= {reg2641};
                      reg2680 <= $signed($unsigned($unsigned(reg1889[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg2679 <= reg2056[(2'h3):(2'h3)];
                      reg2680 <= $unsigned((reg2606 ~^ $signed($unsigned((8'hab)))));
                      reg2681 <= (~&(|({reg1834} <<< $signed(reg2111))));
                    end
                end
            end
          if ((8'hae))
            begin
              for (forvar2693 = (1'h0); (forvar2693 < (2'h3)); forvar2693 = (forvar2693 + (1'h1)))
                begin
                  reg2694 <= {reg2107};
                  for (forvar2695 = (1'h0); (forvar2695 < (2'h3)); forvar2695 = (forvar2695 + (1'h1)))
                    begin
                      reg2696 <= {(reg2691[(1'h0):(1'h0)] ?
                              $unsigned((reg1955 ?
                                  reg2058 : reg2690)) : $signed(reg2098))};
                      reg2697 <= (~|reg1952);
                      reg2698 <= (reg2065 ?
                          $unsigned($unsigned(reg1782[(1'h1):(1'h1)])) : (~|($unsigned(reg1853) < (reg2044 ?
                              reg1962 : forvar2668))));
                    end
                end
              for (forvar2699 = (1'h0); (forvar2699 < (1'h0)); forvar2699 = (forvar2699 + (1'h1)))
                begin
                  reg2700 <= reg1919;
                  reg2701 <= $signed(((!reg1861[(3'h7):(2'h3)]) ?
                      forvar2588 : $unsigned($unsigned(forvar1998))));
                  if (reg2021[(3'h4):(1'h1)])
                    begin
                      reg2702 <= reg1984[(4'ha):(2'h2)];
                    end
                  else
                    begin
                      reg2702 <= reg2081[(3'h6):(1'h0)];
                    end
                  for (forvar2703 = (1'h0); (forvar2703 < (1'h1)); forvar2703 = (forvar2703 + (1'h1)))
                    begin
                      reg2704 <= $unsigned($unsigned((&$unsigned(forvar2632))));
                    end
                end
            end
          else
            begin
              reg2693 <= reg2009[(4'ha):(3'h5)];
            end
        end
      else
        begin
          reg2665 <= ((forvar1776[(4'he):(4'hc)] != reg2630) ~^ $unsigned((reg2106 ?
              (reg2606 != forvar2659) : {reg1833})));
          if ($unsigned(reg2015))
            begin
              for (forvar2666 = (1'h0); (forvar2666 < (2'h2)); forvar2666 = (forvar2666 + (1'h1)))
                begin
                  for (forvar2667 = (1'h0); (forvar2667 < (2'h3)); forvar2667 = (forvar2667 + (1'h1)))
                    begin
                      reg2668 <= reg1871;
                    end
                  for (forvar2669 = (1'h0); (forvar2669 < (2'h3)); forvar2669 = (forvar2669 + (1'h1)))
                    begin
                      reg2670 <= ($unsigned(forvar1807[(3'h5):(2'h2)]) != reg2066[(2'h3):(2'h3)]);
                      reg2671 <= ((!$unsigned({(8'h9d)})) ?
                          (forvar2089[(3'h5):(2'h3)] && (reg1965 || reg1970)) : ($signed((reg1858 ?
                                  reg2588 : reg2088)) ?
                              $signed((-reg1840)) : (forvar2065 ~^ reg1833)));
                    end
                  if ((+($signed((reg1835 ? forvar1914 : forvar1941)) ?
                      {(^(8'ha2))} : wire2582[(2'h3):(2'h3)])))
                    begin
                      reg2672 <= ((|($signed(reg1995) ?
                          (~|reg1886) : reg1816[(4'hc):(4'h9)])) <= (reg1941[(3'h7):(2'h3)] == (^~forvar1997)));
                      reg2673 <= ((($signed(reg1865) <= $signed(reg1869)) ?
                              ({reg2662} ?
                                  {reg2686} : {forvar1799}) : ($signed(reg2684) ?
                                  (~&reg2044) : {reg2071})) ?
                          (&reg1872) : reg1904);
                    end
                  else
                    begin
                      reg2672 <= reg2044[(3'h4):(2'h2)];
                      reg2673 <= $signed({forvar1901});
                    end
                end
            end
          else
            begin
              if (reg2644[(3'h7):(1'h0)])
                begin
                  if ($signed(forvar1969[(2'h3):(1'h1)]))
                    begin
                      reg2666 <= reg2026;
                      reg2667 <= {{$unsigned({reg1789})}};
                      reg2668 <= reg1854;
                    end
                  else
                    begin
                      reg2666 <= (+(8'h9f));
                      reg2667 <= ((^~reg2046) ?
                          {(reg1946[(1'h1):(1'h1)] ?
                                  (reg1833 >> reg2682) : $unsigned(reg2031))} : $signed($unsigned(reg1873)));
                      reg2668 <= ((|((reg1897 ? reg1966 : forvar1896) ?
                              $unsigned(reg2112) : (|reg2667))) ?
                          (reg1932 >>> $signed((reg1891 ?
                              forvar2626 : (8'ha9)))) : {forvar2047});
                    end
                  for (forvar2669 = (1'h0); (forvar2669 < (1'h0)); forvar2669 = (forvar2669 + (1'h1)))
                    begin
                      reg2670 <= $signed($signed($unsigned(forvar2667[(3'h4):(2'h2)])));
                      reg2671 <= ((8'haf) > (((reg1992 >= (8'hb6)) ?
                              $signed(reg2598) : $unsigned(reg1957)) ?
                          ((~&reg2030) > (&reg2111)) : (^reg1872[(1'h0):(1'h0)])));
                      reg2672 <= (~&(^(^{forvar2022})));
                      reg2673 <= (((reg1782 || reg2069[(3'h4):(1'h0)]) ?
                          ((reg1999 + reg1973) ?
                              (forvar2676 != forvar2065) : $signed(forvar1839)) : $signed((reg2093 <<< forvar1809))) < (8'h9f));
                    end
                end
              else
                begin
                  reg2666 <= $unsigned($unsigned((8'ha7)));
                  for (forvar2667 = (1'h0); (forvar2667 < (2'h2)); forvar2667 = (forvar2667 + (1'h1)))
                    begin
                      reg2668 <= {{($unsigned((8'hb5)) & reg1826[(1'h1):(1'h0)])}};
                    end
                  for (forvar2669 = (1'h0); (forvar2669 < (1'h1)); forvar2669 = (forvar2669 + (1'h1)))
                    begin
                      reg2670 <= $signed($signed((reg2058 ?
                          (reg1929 ? reg1962 : reg2682) : wire1772)));
                      reg2671 <= {reg1836};
                    end
                  for (forvar2672 = (1'h0); (forvar2672 < (1'h0)); forvar2672 = (forvar2672 + (1'h1)))
                    begin
                      reg2673 <= ($unsigned(reg2602) - {(((8'ha6) ?
                              forvar1904 : forvar2070) <= (reg1862 ?
                              wire2584 : (8'h9e)))});
                    end
                end
              for (forvar2674 = (1'h0); (forvar2674 < (1'h0)); forvar2674 = (forvar2674 + (1'h1)))
                begin
                  for (forvar2675 = (1'h0); (forvar2675 < (1'h0)); forvar2675 = (forvar2675 + (1'h1)))
                    begin
                      reg2676 <= (forvar1939 ?
                          reg1807[(1'h0):(1'h0)] : ((^(^~forvar1945)) ?
                              forvar2595[(2'h2):(1'h1)] : wire2121[(2'h2):(2'h2)]));
                    end
                  for (forvar2677 = (1'h0); (forvar2677 < (2'h2)); forvar2677 = (forvar2677 + (1'h1)))
                    begin
                      reg2678 <= $signed($signed({(~reg2687)}));
                      reg2679 <= $unsigned((forvar2023[(4'hc):(1'h1)] ^~ ((!reg2010) ?
                          (forvar2703 ? reg1892 : reg2701) : {forvar2626})));
                    end
                  for (forvar2680 = (1'h0); (forvar2680 < (1'h1)); forvar2680 = (forvar2680 + (1'h1)))
                    begin
                      reg2681 <= forvar2688;
                    end
                  reg2682 <= ($signed((~&$signed((8'ha5)))) & reg1995[(3'h7):(2'h2)]);
                end
            end
        end
      for (forvar2705 = (1'h0); (forvar2705 < (1'h0)); forvar2705 = (forvar2705 + (1'h1)))
        begin
          for (forvar2706 = (1'h0); (forvar2706 < (1'h0)); forvar2706 = (forvar2706 + (1'h1)))
            begin
              reg2707 <= ({(((8'hae) >= (8'hb6)) || (reg2642 ?
                          reg1844 : reg2681))} ?
                  forvar1801[(3'h5):(3'h5)] : {(~^(reg2087 && forvar1866))});
              if ((((8'ha2) + (8'haf)) && ($signed(reg2076[(2'h3):(2'h2)]) ?
                  (~&(reg2048 <<< (8'hae))) : forvar2675[(4'h8):(4'h8)])))
                begin
                  for (forvar2708 = (1'h0); (forvar2708 < (1'h1)); forvar2708 = (forvar2708 + (1'h1)))
                    begin
                      reg2709 <= {(&((reg1898 <= wire1772) >>> (~^forvar2022)))};
                    end
                  reg2710 <= reg2067;
                  if ($signed((reg1917 >= ($signed(wire2584) & (reg2644 ?
                      reg2028 : reg1947)))))
                    begin
                      reg2711 <= reg2691;
                      reg2712 <= ((&(reg1900 == (reg2081 ?
                          reg2077 : (8'hba)))) >>> (reg1858[(4'ha):(3'h7)] ^~ forvar1945[(2'h2):(2'h2)]));
                      reg2713 <= reg1949;
                      reg2714 <= (($signed((reg2049 ? reg1956 : reg1899)) ?
                          reg1931[(2'h2):(2'h2)] : wire2585[(3'h5):(2'h2)]) == reg1825[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg2711 <= $signed($signed({(reg1937 ?
                              reg2632 : (8'ha0))}));
                      reg2712 <= ((~|forvar1998) <= $signed((~|(8'ha6))));
                    end
                  for (forvar2715 = (1'h0); (forvar2715 < (1'h0)); forvar2715 = (forvar2715 + (1'h1)))
                    begin
                      reg2716 <= {(&($signed(reg2116) ?
                              reg1933 : (reg2079 ? (8'ha7) : forvar2041)))};
                      reg2717 <= $signed({$signed((reg2073 >> wire1772))});
                      reg2718 <= {$unsigned($unsigned(forvar2673))};
                      reg2719 <= reg1999[(2'h2):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar2708 = (1'h0); (forvar2708 < (1'h1)); forvar2708 = (forvar2708 + (1'h1)))
                    begin
                      reg2709 <= reg2005;
                    end
                end
              for (forvar2720 = (1'h0); (forvar2720 < (2'h2)); forvar2720 = (forvar2720 + (1'h1)))
                begin
                  if ($signed(($signed(forvar1901) != $signed((+reg2719)))))
                    begin
                      reg2721 <= ((8'ha7) ?
                          reg2098[(4'hf):(2'h3)] : ({$unsigned(reg1905)} & $unsigned($unsigned(reg2677))));
                      reg2722 <= (forvar1932[(1'h0):(1'h0)] & ($signed(forvar1980[(4'h9):(4'h8)]) >> $unsigned(reg2659)));
                      reg2723 <= $unsigned(((^~{reg1957}) ~^ reg2059));
                      reg2724 <= (forvar1780[(2'h3):(1'h0)] ?
                          reg2696[(2'h2):(1'h1)] : (8'hb2));
                    end
                  else
                    begin
                      reg2721 <= ((((reg1906 ? reg2115 : reg1946) ?
                                  ((8'hb5) ^ reg1989) : reg2007[(2'h2):(1'h0)]) ?
                              (reg1988[(1'h0):(1'h0)] == (reg1928 | reg2004)) : (forvar1793 < (reg2712 < forvar1940))) ?
                          ((8'h9c) ?
                              $unsigned($signed(reg1854)) : ({forvar1824} ?
                                  {reg2605} : $unsigned(reg1833))) : $unsigned($signed($unsigned(reg2006))));
                    end
                  reg2725 <= ($signed(forvar2034) ?
                      reg1865[(4'h9):(4'h8)] : (reg2031[(3'h4):(2'h2)] | reg2067));
                  if ($signed(forvar2699))
                    begin
                      reg2726 <= $unsigned(reg2684[(3'h6):(3'h4)]);
                      reg2727 <= $unsigned((&((reg1860 ? (8'hb9) : reg2650) ?
                          reg1982[(3'h7):(3'h5)] : {reg2719})));
                      reg2728 <= {$unsigned(forvar1780[(3'h4):(2'h3)])};
                      reg2729 <= ($unsigned(($signed(reg2697) ^ reg1799[(2'h2):(1'h1)])) ?
                          $unsigned(reg2697) : reg2607);
                    end
                  else
                    begin
                      reg2726 <= reg2050;
                    end
                  for (forvar2730 = (1'h0); (forvar2730 < (1'h0)); forvar2730 = (forvar2730 + (1'h1)))
                    begin
                      reg2731 <= (($signed($unsigned(reg1880)) >>> (!(reg2005 ^ forvar2677))) ?
                          $signed(reg2608[(3'h7):(3'h6)]) : (8'ha8));
                      reg2732 <= {$unsigned(reg2663[(2'h3):(1'h0)])};
                      reg2733 <= reg2674[(3'h6):(2'h3)];
                    end
                end
              for (forvar2734 = (1'h0); (forvar2734 < (1'h1)); forvar2734 = (forvar2734 + (1'h1)))
                begin
                  reg2735 <= reg1872;
                  for (forvar2736 = (1'h0); (forvar2736 < (1'h1)); forvar2736 = (forvar2736 + (1'h1)))
                    begin
                      reg2737 <= (((((8'haf) - reg1938) * (!reg2728)) + (reg1865[(2'h3):(2'h3)] ?
                              (~|forvar2673) : ((8'ha7) ? reg2014 : reg2058))) ?
                          $signed(forvar2080[(3'h6):(3'h5)]) : forvar1997);
                      reg2738 <= (~^reg2077);
                      reg2739 <= $signed({reg2006[(4'hb):(3'h7)]});
                      reg2740 <= reg1971[(3'h4):(1'h0)];
                    end
                  if ((~&(~&$unsigned((reg1862 & reg2697)))))
                    begin
                      reg2741 <= $unsigned((reg2071 ~^ (((8'ha1) ?
                              forvar1806 : forvar1939) ?
                          (~&reg2740) : wire1771[(2'h3):(1'h1)])));
                      reg2742 <= {$signed($signed(reg2105))};
                      reg2743 <= $unsigned((reg1913 ?
                          ($unsigned(reg2714) <<< (~(8'ha0))) : ($unsigned(reg1814) ?
                              (forvar1940 <<< reg1979) : $signed((8'ha2)))));
                      reg2744 <= forvar1866;
                    end
                  else
                    begin
                      reg2741 <= $signed($signed($signed((&reg1810))));
                    end
                  reg2745 <= $unsigned($unsigned($signed((reg1790 ?
                      reg2744 : reg1964))));
                end
            end
        end
    end
  assign wire2746 = $signed({forvar2611[(1'h1):(1'h1)]});
  assign wire2747 = $unsigned({$signed($signed((8'h9d)))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module2122  (y, clk, wire2126, wire2125, wire2124, wire2123);
  output wire [(32'h1428):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h9):(1'h0)] wire2126;
  input wire signed [(4'h9):(1'h0)] wire2125;
  input wire signed [(2'h2):(1'h0)] wire2124;
  input wire [(4'he):(1'h0)] wire2123;
  wire [(4'he):(1'h0)] wire2581;
  wire signed [(3'h4):(1'h0)] wire2580;
  wire signed [(4'hf):(1'h0)] wire2579;
  reg [(4'h8):(1'h0)] forvar2550 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2546 = (1'h0);
  reg [(4'he):(1'h0)] reg2544 = (1'h0);
  reg [(4'ha):(1'h0)] reg2542 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2541 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2536 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2531 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2529 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2519 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2520 = (1'h0);
  reg [(3'h5):(1'h0)] reg2578 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2576 = (1'h0);
  reg [(4'hf):(1'h0)] reg2569 = (1'h0);
  reg [(3'h7):(1'h0)] reg2577 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2576 = (1'h0);
  reg [(3'h4):(1'h0)] reg2575 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2574 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2573 = (1'h0);
  reg [(4'he):(1'h0)] reg2572 = (1'h0);
  reg [(4'h9):(1'h0)] reg2571 = (1'h0);
  reg [(4'ha):(1'h0)] reg2570 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2569 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2568 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2567 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2566 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2565 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2564 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2563 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2562 = (1'h0);
  reg [(3'h7):(1'h0)] reg2561 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2560 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2557 = (1'h0);
  reg [(4'hb):(1'h0)] reg2554 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2560 = (1'h0);
  reg [(4'ha):(1'h0)] reg2559 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2558 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2557 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2556 = (1'h0);
  reg [(5'h10):(1'h0)] reg2555 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2554 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2553 = (1'h0);
  reg [(3'h5):(1'h0)] reg2552 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2551 = (1'h0);
  reg [(2'h3):(1'h0)] reg2550 = (1'h0);
  reg [(3'h6):(1'h0)] reg2549 = (1'h0);
  reg [(4'h9):(1'h0)] reg2548 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2547 = (1'h0);
  reg [(3'h6):(1'h0)] reg2546 = (1'h0);
  reg [(3'h6):(1'h0)] reg2545 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2544 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2523 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2521 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2515 = (1'h0);
  reg [(4'h8):(1'h0)] reg2514 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2537 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2535 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2533 = (1'h0);
  reg [(4'ha):(1'h0)] reg2543 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2542 = (1'h0);
  reg [(3'h4):(1'h0)] reg2541 = (1'h0);
  reg [(4'he):(1'h0)] reg2540 = (1'h0);
  reg [(2'h2):(1'h0)] reg2539 = (1'h0);
  reg [(4'h8):(1'h0)] reg2538 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2537 = (1'h0);
  reg [(4'hb):(1'h0)] reg2536 = (1'h0);
  reg [(4'hc):(1'h0)] reg2535 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2534 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2533 = (1'h0);
  reg [(5'h10):(1'h0)] reg2532 = (1'h0);
  reg [(2'h3):(1'h0)] reg2531 = (1'h0);
  reg [(2'h2):(1'h0)] reg2530 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2529 = (1'h0);
  reg [(3'h5):(1'h0)] reg2528 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2527 = (1'h0);
  reg [(4'hd):(1'h0)] reg2526 = (1'h0);
  reg [(4'hb):(1'h0)] reg2525 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2524 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2523 = (1'h0);
  reg [(4'hc):(1'h0)] reg2522 = (1'h0);
  reg [(4'hf):(1'h0)] reg2521 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2520 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2519 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2518 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2517 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2516 = (1'h0);
  reg [(3'h5):(1'h0)] reg2515 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2514 = (1'h0);
  reg [(4'he):(1'h0)] reg2513 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2512 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2502 = (1'h0);
  reg [(4'he):(1'h0)] reg2499 = (1'h0);
  reg [(4'hc):(1'h0)] reg2511 = (1'h0);
  reg [(4'ha):(1'h0)] reg2510 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2509 = (1'h0);
  reg [(4'hb):(1'h0)] reg2508 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2507 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2506 = (1'h0);
  reg [(4'he):(1'h0)] reg2505 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2504 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2503 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2502 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2501 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2500 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2499 = (1'h0);
  reg [(5'h10):(1'h0)] reg2498 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2497 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2496 = (1'h0);
  reg [(4'h9):(1'h0)] reg2495 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2494 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2493 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2492 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2491 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2490 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2489 = (1'h0);
  reg [(3'h6):(1'h0)] reg2488 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2487 = (1'h0);
  reg [(4'ha):(1'h0)] reg2486 = (1'h0);
  reg [(4'hf):(1'h0)] reg2485 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2484 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2483 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2482 = (1'h0);
  reg [(3'h4):(1'h0)] reg2481 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2480 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2479 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2478 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2460 = (1'h0);
  reg [(2'h3):(1'h0)] reg2477 = (1'h0);
  reg [(3'h5):(1'h0)] reg2476 = (1'h0);
  reg [(5'h10):(1'h0)] reg2475 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2474 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2473 = (1'h0);
  reg [(5'h10):(1'h0)] reg2472 = (1'h0);
  reg [(2'h3):(1'h0)] reg2471 = (1'h0);
  reg [(5'h10):(1'h0)] reg2470 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2469 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2468 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2467 = (1'h0);
  reg [(3'h6):(1'h0)] reg2466 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2465 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2456 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2464 = (1'h0);
  reg [(2'h2):(1'h0)] reg2463 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2462 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2461 = (1'h0);
  reg [(3'h5):(1'h0)] reg2460 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2459 = (1'h0);
  reg [(3'h4):(1'h0)] reg2458 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2457 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2456 = (1'h0);
  reg [(3'h6):(1'h0)] reg2455 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2454 = (1'h0);
  reg [(2'h3):(1'h0)] reg2453 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2452 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2451 = (1'h0);
  reg [(4'hc):(1'h0)] reg2446 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2450 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2449 = (1'h0);
  reg [(3'h4):(1'h0)] reg2448 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2447 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2446 = (1'h0);
  reg [(4'hd):(1'h0)] reg2445 = (1'h0);
  reg [(3'h4):(1'h0)] reg2444 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2443 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2442 = (1'h0);
  reg [(4'he):(1'h0)] forvar2441 = (1'h0);
  reg [(4'ha):(1'h0)] reg2440 = (1'h0);
  reg [(4'hf):(1'h0)] reg2439 = (1'h0);
  reg [(3'h4):(1'h0)] reg2438 = (1'h0);
  reg [(3'h6):(1'h0)] reg2437 = (1'h0);
  reg [(3'h6):(1'h0)] reg2436 = (1'h0);
  reg [(5'h10):(1'h0)] reg2435 = (1'h0);
  reg [(4'hc):(1'h0)] reg2434 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2433 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2432 = (1'h0);
  reg [(4'ha):(1'h0)] reg2431 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2430 = (1'h0);
  reg [(3'h6):(1'h0)] forvar2429 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2428 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2427 = (1'h0);
  reg [(4'hc):(1'h0)] reg2426 = (1'h0);
  reg [(4'hf):(1'h0)] forvar2425 = (1'h0);
  reg [(4'h8):(1'h0)] reg2424 = (1'h0);
  reg [(4'ha):(1'h0)] reg2423 = (1'h0);
  reg [(5'h10):(1'h0)] reg2422 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2421 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2420 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2419 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2418 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2417 = (1'h0);
  reg [(2'h3):(1'h0)] reg2416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2415 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2414 = (1'h0);
  reg [(5'h10):(1'h0)] reg2413 = (1'h0);
  reg [(4'hc):(1'h0)] reg2412 = (1'h0);
  reg [(4'h8):(1'h0)] reg2411 = (1'h0);
  reg [(4'hc):(1'h0)] reg2410 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2409 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2408 = (1'h0);
  reg [(2'h3):(1'h0)] reg2407 = (1'h0);
  reg [(4'h9):(1'h0)] reg2406 = (1'h0);
  reg [(4'hd):(1'h0)] reg2405 = (1'h0);
  reg [(4'he):(1'h0)] reg2404 = (1'h0);
  reg [(4'he):(1'h0)] reg2403 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2402 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2401 = (1'h0);
  reg [(3'h5):(1'h0)] reg2400 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2399 = (1'h0);
  reg [(4'h9):(1'h0)] reg2398 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2397 = (1'h0);
  reg [(4'hf):(1'h0)] reg2396 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2395 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2394 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2393 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2392 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2389 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2388 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2386 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2381 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2380 = (1'h0);
  reg [(2'h2):(1'h0)] reg2377 = (1'h0);
  reg [(3'h6):(1'h0)] reg2376 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2375 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2374 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2391 = (1'h0);
  reg [(3'h4):(1'h0)] reg2390 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2389 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2388 = (1'h0);
  reg [(3'h7):(1'h0)] reg2387 = (1'h0);
  reg [(3'h5):(1'h0)] reg2386 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2385 = (1'h0);
  reg [(4'he):(1'h0)] reg2384 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2383 = (1'h0);
  reg [(2'h3):(1'h0)] reg2382 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2381 = (1'h0);
  reg [(4'h8):(1'h0)] reg2380 = (1'h0);
  reg [(3'h5):(1'h0)] reg2379 = (1'h0);
  reg [(3'h4):(1'h0)] reg2378 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2377 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2376 = (1'h0);
  reg [(4'hc):(1'h0)] reg2375 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2374 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2373 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2372 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire2371;
  reg signed [(4'hc):(1'h0)] reg2370 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2356 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2355 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2349 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2358 = (1'h0);
  reg [(2'h3):(1'h0)] reg2369 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2368 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2367 = (1'h0);
  reg [(2'h3):(1'h0)] reg2366 = (1'h0);
  reg [(3'h4):(1'h0)] reg2365 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2364 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2363 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2362 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2361 = (1'h0);
  reg [(4'hf):(1'h0)] reg2360 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2359 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2358 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2353 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2350 = (1'h0);
  reg [(3'h5):(1'h0)] reg2357 = (1'h0);
  reg [(4'h9):(1'h0)] reg2356 = (1'h0);
  reg [(2'h3):(1'h0)] reg2355 = (1'h0);
  reg [(3'h7):(1'h0)] reg2354 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2353 = (1'h0);
  reg [(4'h8):(1'h0)] reg2352 = (1'h0);
  reg [(2'h2):(1'h0)] reg2351 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2350 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2349 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2348 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire2347;
  wire signed [(4'hb):(1'h0)] wire2346;
  reg signed [(2'h2):(1'h0)] reg2335 = (1'h0);
  reg [(4'hf):(1'h0)] reg2332 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2329 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2313 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2300 = (1'h0);
  reg [(2'h3):(1'h0)] reg2305 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2304 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2299 = (1'h0);
  reg [(3'h5):(1'h0)] reg2283 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2297 = (1'h0);
  reg [(3'h7):(1'h0)] reg2294 = (1'h0);
  reg [(4'ha):(1'h0)] reg2291 = (1'h0);
  reg [(3'h4):(1'h0)] reg2286 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2285 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2280 = (1'h0);
  reg [(4'hc):(1'h0)] reg2276 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2345 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2344 = (1'h0);
  reg [(4'he):(1'h0)] reg2343 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2342 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2341 = (1'h0);
  reg [(4'h9):(1'h0)] reg2340 = (1'h0);
  reg [(4'ha):(1'h0)] reg2339 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2338 = (1'h0);
  reg [(2'h2):(1'h0)] reg2337 = (1'h0);
  reg [(3'h5):(1'h0)] reg2336 = (1'h0);
  reg [(4'hb):(1'h0)] forvar2335 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2334 = (1'h0);
  reg [(3'h5):(1'h0)] reg2333 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2332 = (1'h0);
  reg [(2'h3):(1'h0)] reg2331 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2330 = (1'h0);
  reg [(4'hd):(1'h0)] reg2328 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2329 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2328 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2323 = (1'h0);
  reg [(5'h10):(1'h0)] reg2319 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2318 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2316 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2315 = (1'h0);
  reg [(4'h8):(1'h0)] reg2327 = (1'h0);
  reg [(4'h8):(1'h0)] reg2326 = (1'h0);
  reg [(3'h5):(1'h0)] reg2325 = (1'h0);
  reg [(2'h2):(1'h0)] reg2324 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2323 = (1'h0);
  reg [(3'h5):(1'h0)] reg2322 = (1'h0);
  reg [(4'hd):(1'h0)] reg2321 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2320 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2319 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2318 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2317 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2316 = (1'h0);
  reg [(4'he):(1'h0)] reg2315 = (1'h0);
  reg [(2'h2):(1'h0)] forvar2314 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2313 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2312 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2311 = (1'h0);
  reg [(4'hf):(1'h0)] reg2310 = (1'h0);
  reg [(4'hf):(1'h0)] reg2309 = (1'h0);
  reg [(3'h4):(1'h0)] reg2308 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2307 = (1'h0);
  reg [(4'h8):(1'h0)] reg2306 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2305 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2304 = (1'h0);
  reg [(4'hc):(1'h0)] reg2303 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2302 = (1'h0);
  reg [(4'hb):(1'h0)] reg2301 = (1'h0);
  reg [(3'h6):(1'h0)] reg2300 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2299 = (1'h0);
  reg [(4'ha):(1'h0)] reg2298 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2297 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2296 = (1'h0);
  reg [(4'h8):(1'h0)] reg2295 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2294 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2293 = (1'h0);
  reg [(4'h9):(1'h0)] reg2292 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2291 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2290 = (1'h0);
  reg [(4'hd):(1'h0)] reg2289 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2288 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2287 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2286 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2285 = (1'h0);
  reg [(2'h2):(1'h0)] reg2284 = (1'h0);
  reg [(4'he):(1'h0)] forvar2283 = (1'h0);
  reg [(4'hb):(1'h0)] reg2282 = (1'h0);
  reg [(4'hc):(1'h0)] reg2281 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2280 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2277 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2279 = (1'h0);
  reg [(4'ha):(1'h0)] reg2278 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2277 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2276 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2219 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2214 = (1'h0);
  reg [(3'h4):(1'h0)] reg2271 = (1'h0);
  reg [(3'h6):(1'h0)] reg2275 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2274 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2273 = (1'h0);
  reg [(3'h6):(1'h0)] reg2272 = (1'h0);
  reg [(5'h10):(1'h0)] forvar2271 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2270 = (1'h0);
  reg [(4'hc):(1'h0)] reg2269 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2268 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2267 = (1'h0);
  reg [(3'h5):(1'h0)] reg2266 = (1'h0);
  reg [(4'he):(1'h0)] reg2265 = (1'h0);
  reg [(3'h7):(1'h0)] reg2264 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2263 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2262 = (1'h0);
  reg [(3'h7):(1'h0)] reg2261 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2260 = (1'h0);
  reg [(5'h10):(1'h0)] reg2259 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2258 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2257 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2256 = (1'h0);
  reg [(4'h9):(1'h0)] reg2255 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2254 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2253 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2248 = (1'h0);
  reg [(5'h10):(1'h0)] reg2243 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2242 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2252 = (1'h0);
  reg [(5'h10):(1'h0)] reg2251 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2250 = (1'h0);
  reg [(3'h7):(1'h0)] reg2249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2248 = (1'h0);
  reg [(4'h9):(1'h0)] reg2247 = (1'h0);
  reg [(4'h9):(1'h0)] reg2246 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2245 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2244 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar2243 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2242 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2241 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2229 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2224 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2240 = (1'h0);
  reg [(4'hb):(1'h0)] reg2239 = (1'h0);
  reg [(3'h6):(1'h0)] reg2238 = (1'h0);
  reg [(4'h9):(1'h0)] reg2237 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2233 = (1'h0);
  reg [(3'h4):(1'h0)] forvar2232 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2228 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar2227 = (1'h0);
  reg [(3'h4):(1'h0)] reg2236 = (1'h0);
  reg [(4'hc):(1'h0)] reg2235 = (1'h0);
  reg [(3'h4):(1'h0)] reg2234 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2233 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2232 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2231 = (1'h0);
  reg [(4'ha):(1'h0)] reg2230 = (1'h0);
  reg [(5'h10):(1'h0)] reg2229 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2228 = (1'h0);
  reg [(3'h5):(1'h0)] reg2227 = (1'h0);
  reg [(4'hb):(1'h0)] reg2226 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2225 = (1'h0);
  reg [(3'h4):(1'h0)] reg2224 = (1'h0);
  reg [(3'h5):(1'h0)] reg2223 = (1'h0);
  reg [(4'hc):(1'h0)] reg2222 = (1'h0);
  reg [(3'h4):(1'h0)] reg2221 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2220 = (1'h0);
  reg [(3'h7):(1'h0)] reg2219 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2218 = (1'h0);
  reg [(3'h7):(1'h0)] reg2217 = (1'h0);
  reg [(4'h9):(1'h0)] reg2216 = (1'h0);
  reg [(4'he):(1'h0)] reg2215 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2214 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2213 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2212 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2211 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2210 = (1'h0);
  reg [(3'h5):(1'h0)] reg2209 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2208 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2207 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2206 = (1'h0);
  reg [(4'hf):(1'h0)] reg2205 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2204 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2203 = (1'h0);
  reg [(3'h7):(1'h0)] reg2202 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2201 = (1'h0);
  reg [(4'hc):(1'h0)] forvar2200 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg2199 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2198 = (1'h0);
  reg [(4'hc):(1'h0)] reg2197 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2193 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2192 = (1'h0);
  reg [(4'hf):(1'h0)] reg2191 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2187 = (1'h0);
  reg [(4'hb):(1'h0)] reg2195 = (1'h0);
  reg [(4'hf):(1'h0)] reg2196 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2195 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2194 = (1'h0);
  reg [(3'h7):(1'h0)] reg2193 = (1'h0);
  reg [(4'ha):(1'h0)] reg2192 = (1'h0);
  reg [(4'ha):(1'h0)] forvar2191 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2190 = (1'h0);
  reg [(3'h5):(1'h0)] reg2189 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2188 = (1'h0);
  reg [(4'h8):(1'h0)] reg2187 = (1'h0);
  reg [(4'ha):(1'h0)] reg2175 = (1'h0);
  reg [(5'h10):(1'h0)] reg2174 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar2173 = (1'h0);
  reg [(2'h3):(1'h0)] forvar2170 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2165 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2186 = (1'h0);
  reg [(2'h2):(1'h0)] reg2185 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2184 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2183 = (1'h0);
  reg [(3'h5):(1'h0)] reg2182 = (1'h0);
  reg [(4'h8):(1'h0)] reg2181 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2180 = (1'h0);
  reg [(3'h5):(1'h0)] forvar2179 = (1'h0);
  reg [(5'h10):(1'h0)] reg2178 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2177 = (1'h0);
  reg [(5'h10):(1'h0)] reg2176 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar2175 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2174 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg2172 = (1'h0);
  reg [(3'h6):(1'h0)] reg2173 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2172 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2171 = (1'h0);
  reg [(2'h2):(1'h0)] reg2170 = (1'h0);
  reg [(3'h7):(1'h0)] reg2169 = (1'h0);
  reg [(4'h8):(1'h0)] forvar2162 = (1'h0);
  reg [(3'h7):(1'h0)] reg2161 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2159 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2157 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar2137 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2156 = (1'h0);
  reg [(4'hd):(1'h0)] reg2155 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar2152 = (1'h0);
  reg [(4'h9):(1'h0)] reg2150 = (1'h0);
  reg [(3'h7):(1'h0)] reg2148 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar2147 = (1'h0);
  reg [(4'h9):(1'h0)] reg2144 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2141 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar2133 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar2135 = (1'h0);
  reg [(4'h9):(1'h0)] reg2132 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg2168 = (1'h0);
  reg [(3'h7):(1'h0)] reg2167 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2166 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg2163 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2166 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg2165 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg2164 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar2163 = (1'h0);
  reg [(4'hc):(1'h0)] reg2162 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2161 = (1'h0);
  reg [(4'hf):(1'h0)] reg2160 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2159 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg2158 = (1'h0);
  reg [(3'h6):(1'h0)] reg2157 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar2156 = (1'h0);
  reg [(3'h7):(1'h0)] forvar2155 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg2134 = (1'h0);
  reg [(4'hc):(1'h0)] reg2154 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg2153 = (1'h0);
  reg [(3'h5):(1'h0)] reg2152 = (1'h0);
  reg [(2'h2):(1'h0)] reg2151 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar2150 = (1'h0);
  reg [(3'h5):(1'h0)] reg2149 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar2148 = (1'h0);
  reg [(2'h2):(1'h0)] reg2147 = (1'h0);
  reg [(4'he):(1'h0)] reg2146 = (1'h0);
  reg [(4'ha):(1'h0)] reg2145 = (1'h0);
  reg [(4'h9):(1'h0)] forvar2144 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2143 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2142 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg2141 = (1'h0);
  reg signed [(4'he):(1'h0)] reg2140 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar2139 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg2139 = (1'h0);
  reg [(4'hf):(1'h0)] reg2138 = (1'h0);
  reg [(4'h8):(1'h0)] reg2137 = (1'h0);
  reg [(4'hb):(1'h0)] reg2136 = (1'h0);
  reg [(3'h6):(1'h0)] reg2135 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar2134 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg2133 = (1'h0);
  reg [(4'hd):(1'h0)] forvar2132 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg2131 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg2130 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire2129;
  wire signed [(5'h10):(1'h0)] wire2128;
  wire signed [(2'h2):(1'h0)] wire2127;
  assign y = {wire2581,
                 wire2580,
                 wire2579,
                 forvar2550,
                 forvar2546,
                 reg2544,
                 reg2542,
                 forvar2541,
                 forvar2536,
                 forvar2531,
                 forvar2529,
                 forvar2519,
                 reg2520,
                 reg2578,
                 reg2576,
                 reg2569,
                 reg2577,
                 forvar2576,
                 reg2575,
                 reg2574,
                 forvar2573,
                 reg2572,
                 reg2571,
                 reg2570,
                 forvar2569,
                 forvar2568,
                 reg2567,
                 reg2566,
                 reg2565,
                 reg2564,
                 forvar2563,
                 forvar2562,
                 reg2561,
                 forvar2560,
                 forvar2557,
                 reg2554,
                 reg2560,
                 reg2559,
                 reg2558,
                 reg2557,
                 reg2556,
                 reg2555,
                 forvar2554,
                 reg2553,
                 reg2552,
                 forvar2551,
                 reg2550,
                 reg2549,
                 reg2548,
                 reg2547,
                 reg2546,
                 reg2545,
                 forvar2544,
                 reg2523,
                 forvar2521,
                 forvar2515,
                 reg2514,
                 forvar2537,
                 forvar2535,
                 reg2533,
                 reg2543,
                 forvar2542,
                 reg2541,
                 reg2540,
                 reg2539,
                 reg2538,
                 reg2537,
                 reg2536,
                 reg2535,
                 reg2534,
                 forvar2533,
                 reg2532,
                 reg2531,
                 reg2530,
                 reg2529,
                 reg2528,
                 reg2527,
                 reg2526,
                 reg2525,
                 reg2524,
                 forvar2523,
                 reg2522,
                 reg2521,
                 forvar2520,
                 reg2519,
                 reg2518,
                 reg2517,
                 reg2516,
                 reg2515,
                 forvar2514,
                 reg2513,
                 forvar2512,
                 forvar2502,
                 reg2499,
                 reg2511,
                 reg2510,
                 reg2509,
                 reg2508,
                 reg2507,
                 reg2506,
                 reg2505,
                 reg2504,
                 reg2503,
                 reg2502,
                 reg2501,
                 reg2500,
                 forvar2499,
                 reg2498,
                 forvar2497,
                 reg2496,
                 reg2495,
                 reg2494,
                 reg2493,
                 reg2492,
                 reg2491,
                 reg2490,
                 reg2489,
                 reg2488,
                 reg2487,
                 reg2486,
                 reg2485,
                 forvar2484,
                 forvar2483,
                 forvar2482,
                 reg2481,
                 reg2480,
                 forvar2479,
                 reg2478,
                 forvar2460,
                 reg2477,
                 reg2476,
                 reg2475,
                 forvar2474,
                 reg2473,
                 reg2472,
                 reg2471,
                 reg2470,
                 forvar2469,
                 forvar2468,
                 reg2467,
                 reg2466,
                 forvar2465,
                 forvar2456,
                 reg2464,
                 reg2463,
                 reg2462,
                 reg2461,
                 reg2460,
                 reg2459,
                 reg2458,
                 reg2457,
                 reg2456,
                 reg2455,
                 forvar2454,
                 reg2453,
                 forvar2452,
                 forvar2451,
                 reg2446,
                 reg2450,
                 reg2449,
                 reg2448,
                 reg2447,
                 forvar2446,
                 reg2445,
                 reg2444,
                 reg2443,
                 reg2442,
                 forvar2441,
                 reg2440,
                 reg2439,
                 reg2438,
                 reg2437,
                 reg2436,
                 reg2435,
                 reg2434,
                 forvar2433,
                 reg2432,
                 reg2431,
                 reg2430,
                 forvar2429,
                 forvar2428,
                 reg2427,
                 reg2426,
                 forvar2425,
                 reg2424,
                 reg2423,
                 reg2422,
                 forvar2421,
                 forvar2420,
                 forvar2419,
                 reg2418,
                 reg2417,
                 reg2416,
                 reg2415,
                 reg2414,
                 reg2413,
                 reg2412,
                 reg2411,
                 reg2410,
                 reg2409,
                 forvar2408,
                 reg2407,
                 reg2406,
                 reg2405,
                 reg2404,
                 reg2403,
                 reg2402,
                 reg2401,
                 reg2400,
                 forvar2399,
                 reg2398,
                 reg2397,
                 reg2396,
                 forvar2395,
                 reg2394,
                 reg2393,
                 reg2392,
                 forvar2389,
                 reg2388,
                 forvar2386,
                 forvar2381,
                 forvar2380,
                 reg2377,
                 reg2376,
                 forvar2375,
                 reg2374,
                 reg2391,
                 reg2390,
                 reg2389,
                 forvar2388,
                 reg2387,
                 reg2386,
                 reg2385,
                 reg2384,
                 reg2383,
                 reg2382,
                 reg2381,
                 reg2380,
                 reg2379,
                 reg2378,
                 forvar2377,
                 forvar2376,
                 reg2375,
                 forvar2374,
                 forvar2373,
                 forvar2372,
                 wire2371,
                 reg2370,
                 forvar2356,
                 forvar2355,
                 forvar2349,
                 forvar2358,
                 reg2369,
                 reg2368,
                 forvar2367,
                 reg2366,
                 reg2365,
                 reg2364,
                 reg2363,
                 reg2362,
                 reg2361,
                 reg2360,
                 reg2359,
                 reg2358,
                 forvar2353,
                 reg2350,
                 reg2357,
                 reg2356,
                 reg2355,
                 reg2354,
                 reg2353,
                 reg2352,
                 reg2351,
                 forvar2350,
                 reg2349,
                 forvar2348,
                 wire2347,
                 wire2346,
                 reg2335,
                 reg2332,
                 forvar2329,
                 forvar2313,
                 forvar2300,
                 reg2305,
                 forvar2304,
                 forvar2299,
                 reg2283,
                 reg2297,
                 reg2294,
                 reg2291,
                 reg2286,
                 reg2285,
                 forvar2280,
                 reg2276,
                 reg2345,
                 reg2344,
                 reg2343,
                 reg2342,
                 forvar2341,
                 reg2340,
                 reg2339,
                 forvar2338,
                 reg2337,
                 reg2336,
                 forvar2335,
                 reg2334,
                 reg2333,
                 forvar2332,
                 reg2331,
                 reg2330,
                 reg2328,
                 reg2329,
                 forvar2328,
                 reg2323,
                 reg2319,
                 forvar2318,
                 reg2316,
                 forvar2315,
                 reg2327,
                 reg2326,
                 reg2325,
                 reg2324,
                 forvar2323,
                 reg2322,
                 reg2321,
                 reg2320,
                 forvar2319,
                 reg2318,
                 reg2317,
                 forvar2316,
                 reg2315,
                 forvar2314,
                 reg2313,
                 reg2312,
                 reg2311,
                 reg2310,
                 reg2309,
                 reg2308,
                 reg2307,
                 reg2306,
                 forvar2305,
                 reg2304,
                 reg2303,
                 reg2302,
                 reg2301,
                 reg2300,
                 reg2299,
                 reg2298,
                 forvar2297,
                 reg2296,
                 reg2295,
                 forvar2294,
                 forvar2293,
                 reg2292,
                 forvar2291,
                 reg2290,
                 reg2289,
                 reg2288,
                 reg2287,
                 forvar2286,
                 forvar2285,
                 reg2284,
                 forvar2283,
                 reg2282,
                 reg2281,
                 reg2280,
                 forvar2279,
                 reg2277,
                 reg2279,
                 reg2278,
                 forvar2277,
                 forvar2276,
                 forvar2219,
                 forvar2214,
                 reg2271,
                 reg2275,
                 reg2274,
                 reg2273,
                 reg2272,
                 forvar2271,
                 reg2270,
                 reg2269,
                 reg2268,
                 forvar2267,
                 reg2266,
                 reg2265,
                 reg2264,
                 reg2263,
                 reg2262,
                 reg2261,
                 reg2260,
                 reg2259,
                 reg2258,
                 forvar2257,
                 forvar2256,
                 reg2255,
                 reg2254,
                 reg2253,
                 forvar2248,
                 reg2243,
                 forvar2242,
                 reg2252,
                 reg2251,
                 reg2250,
                 reg2249,
                 reg2248,
                 reg2247,
                 reg2246,
                 reg2245,
                 reg2244,
                 forvar2243,
                 reg2242,
                 reg2241,
                 forvar2229,
                 forvar2224,
                 reg2240,
                 reg2239,
                 reg2238,
                 reg2237,
                 reg2233,
                 forvar2232,
                 reg2228,
                 forvar2227,
                 reg2236,
                 reg2235,
                 reg2234,
                 forvar2233,
                 reg2232,
                 reg2231,
                 reg2230,
                 reg2229,
                 forvar2228,
                 reg2227,
                 reg2226,
                 reg2225,
                 reg2224,
                 reg2223,
                 reg2222,
                 reg2221,
                 reg2220,
                 reg2219,
                 reg2218,
                 reg2217,
                 reg2216,
                 reg2215,
                 reg2214,
                 forvar2213,
                 forvar2212,
                 reg2211,
                 reg2210,
                 reg2209,
                 reg2208,
                 reg2207,
                 forvar2206,
                 reg2205,
                 reg2204,
                 reg2203,
                 reg2202,
                 forvar2201,
                 forvar2200,
                 reg2199,
                 forvar2198,
                 reg2197,
                 forvar2193,
                 forvar2192,
                 reg2191,
                 forvar2187,
                 reg2195,
                 reg2196,
                 forvar2195,
                 reg2194,
                 reg2193,
                 reg2192,
                 forvar2191,
                 reg2190,
                 reg2189,
                 reg2188,
                 reg2187,
                 reg2175,
                 reg2174,
                 forvar2173,
                 forvar2170,
                 forvar2165,
                 reg2186,
                 reg2185,
                 reg2184,
                 reg2183,
                 reg2182,
                 reg2181,
                 reg2180,
                 forvar2179,
                 reg2178,
                 reg2177,
                 reg2176,
                 forvar2175,
                 forvar2174,
                 reg2172,
                 reg2173,
                 forvar2172,
                 reg2171,
                 reg2170,
                 reg2169,
                 forvar2162,
                 reg2161,
                 forvar2159,
                 forvar2157,
                 forvar2137,
                 reg2156,
                 reg2155,
                 forvar2152,
                 reg2150,
                 reg2148,
                 forvar2147,
                 reg2144,
                 forvar2141,
                 forvar2133,
                 forvar2135,
                 reg2132,
                 reg2168,
                 reg2167,
                 forvar2166,
                 reg2163,
                 reg2166,
                 reg2165,
                 reg2164,
                 forvar2163,
                 reg2162,
                 forvar2161,
                 reg2160,
                 reg2159,
                 reg2158,
                 reg2157,
                 forvar2156,
                 forvar2155,
                 reg2134,
                 reg2154,
                 reg2153,
                 reg2152,
                 reg2151,
                 forvar2150,
                 reg2149,
                 forvar2148,
                 reg2147,
                 reg2146,
                 reg2145,
                 forvar2144,
                 reg2143,
                 reg2142,
                 reg2141,
                 reg2140,
                 forvar2139,
                 reg2139,
                 reg2138,
                 reg2137,
                 reg2136,
                 reg2135,
                 forvar2134,
                 reg2133,
                 forvar2132,
                 reg2131,
                 reg2130,
                 wire2129,
                 wire2128,
                 wire2127,
                 (1'h0)};
  assign wire2127 = {wire2125};
  assign wire2128 = wire2124[(1'h0):(1'h0)];
  assign wire2129 = wire2126;
  always
    @(posedge clk) begin
      reg2130 <= $signed($signed(wire2129));
      reg2131 <= reg2130[(1'h1):(1'h1)];
      if ($signed((wire2124[(1'h0):(1'h0)] > (-wire2127[(2'h2):(1'h0)]))))
        begin
          if ((((!$unsigned(wire2125)) ?
                  (~|$signed(wire2127)) : wire2123[(4'hc):(3'h4)]) ?
              {wire2129[(2'h2):(2'h2)]} : (8'had)))
            begin
              for (forvar2132 = (1'h0); (forvar2132 < (2'h3)); forvar2132 = (forvar2132 + (1'h1)))
                begin
                  reg2133 <= forvar2132;
                  for (forvar2134 = (1'h0); (forvar2134 < (1'h0)); forvar2134 = (forvar2134 + (1'h1)))
                    begin
                      reg2135 <= ({$unsigned({reg2133})} ?
                          (|forvar2132) : {(~|(forvar2132 ?
                                  wire2124 : forvar2132))});
                      reg2136 <= ($signed($unsigned(wire2127[(1'h1):(1'h1)])) ?
                          ((8'hb0) ?
                              $signed(((8'hb1) >> wire2127)) : wire2125[(2'h3):(2'h2)]) : ($signed(forvar2134[(3'h5):(3'h5)]) * {wire2124}));
                    end
                  reg2137 <= (^~{((^wire2129) ?
                          $signed(forvar2134) : (~&(8'ha7)))});
                  reg2138 <= $signed({(wire2129[(1'h1):(1'h1)] ^ $unsigned(wire2128))});
                end
              if ({($signed(wire2124[(1'h1):(1'h1)]) ?
                      wire2123[(3'h4):(2'h2)] : wire2129)})
                begin
                  reg2139 <= wire2127[(2'h2):(2'h2)];
                end
              else
                begin
                  for (forvar2139 = (1'h0); (forvar2139 < (2'h2)); forvar2139 = (forvar2139 + (1'h1)))
                    begin
                      reg2140 <= wire2123[(4'hd):(3'h6)];
                      reg2141 <= (|(((reg2139 + (8'ha4)) ?
                          wire2126[(3'h5):(3'h5)] : wire2127[(2'h2):(1'h1)]) >>> $unsigned(wire2125)));
                      reg2142 <= $signed(reg2135);
                      reg2143 <= ($signed({{reg2139}}) >>> $signed((forvar2132[(4'ha):(3'h5)] ?
                          (+(8'h9d)) : $signed((8'hb8)))));
                    end
                end
              for (forvar2144 = (1'h0); (forvar2144 < (1'h1)); forvar2144 = (forvar2144 + (1'h1)))
                begin
                  if ($unsigned($unsigned(((reg2130 || wire2126) ?
                      (reg2130 ? reg2137 : wire2125) : reg2131))))
                    begin
                      reg2145 <= (8'ha8);
                      reg2146 <= $signed(((&reg2133[(1'h0):(1'h0)]) ?
                          $unsigned(reg2131) : $unsigned({(8'h9f)})));
                      reg2147 <= $unsigned(($unsigned((reg2130 ?
                          reg2145 : forvar2139)) * wire2125[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg2145 <= $unsigned($signed(($unsigned(reg2146) ?
                          $signed(reg2145) : forvar2132[(4'h8):(4'h8)])));
                      reg2146 <= $unsigned((+forvar2132[(3'h6):(2'h2)]));
                    end
                end
              for (forvar2148 = (1'h0); (forvar2148 < (1'h0)); forvar2148 = (forvar2148 + (1'h1)))
                begin
                  reg2149 <= $signed(wire2124[(2'h2):(2'h2)]);
                  for (forvar2150 = (1'h0); (forvar2150 < (1'h1)); forvar2150 = (forvar2150 + (1'h1)))
                    begin
                      reg2151 <= wire2127[(1'h1):(1'h0)];
                    end
                  if ((&((^$signed(reg2149)) ?
                      (|((8'hb8) == reg2139)) : $unsigned((reg2143 ?
                          forvar2148 : forvar2150)))))
                    begin
                      reg2152 <= (((^~((8'haf) * reg2137)) > (wire2128 != (!(8'haa)))) - wire2123[(3'h4):(3'h4)]);
                      reg2153 <= $unsigned((((reg2139 || reg2136) + (~^reg2141)) ~^ $signed(((8'ha7) ?
                          reg2139 : wire2127))));
                    end
                  else
                    begin
                      reg2152 <= $unsigned(reg2130);
                      reg2153 <= ((~|reg2152[(2'h3):(2'h3)]) ~^ $unsigned(($unsigned(forvar2144) ^~ (reg2139 == reg2149))));
                      reg2154 <= (!reg2138);
                    end
                end
            end
          else
            begin
              for (forvar2132 = (1'h0); (forvar2132 < (2'h2)); forvar2132 = (forvar2132 + (1'h1)))
                begin
                  if (reg2140)
                    begin
                      reg2133 <= reg2145;
                      reg2134 <= (!{($unsigned((8'hb7)) << $unsigned(wire2124))});
                      reg2135 <= {$unsigned($signed((~forvar2132)))};
                      reg2136 <= $signed((reg2145 <<< wire2127));
                    end
                  else
                    begin
                      reg2133 <= {(^((reg2130 ?
                              wire2125 : reg2137) != (8'hb9)))};
                      reg2134 <= {$unsigned($unsigned($signed(wire2129)))};
                      reg2135 <= ({{$unsigned((8'hb7))}} ?
                          wire2126 : reg2131[(3'h6):(3'h6)]);
                      reg2136 <= reg2141;
                    end
                  reg2137 <= {((reg2138 ?
                          $signed(reg2153) : $unsigned(reg2139)) ^ ((reg2153 ?
                              reg2154 : reg2136) ?
                          (forvar2148 <<< (8'ha0)) : reg2145))};
                  if ($unsigned($unsigned(wire2123[(3'h4):(2'h2)])))
                    begin
                      reg2138 <= (!$signed((^(~(8'hb9)))));
                    end
                  else
                    begin
                      reg2138 <= {forvar2148};
                      reg2139 <= $signed(((((8'haf) ?
                              wire2125 : reg2151) <<< forvar2134[(2'h2):(1'h1)]) ?
                          $unsigned($signed(reg2139)) : $unsigned((+reg2143))));
                    end
                end
              reg2140 <= reg2134[(1'h1):(1'h1)];
            end
          for (forvar2155 = (1'h0); (forvar2155 < (1'h1)); forvar2155 = (forvar2155 + (1'h1)))
            begin
              for (forvar2156 = (1'h0); (forvar2156 < (1'h1)); forvar2156 = (forvar2156 + (1'h1)))
                begin
                  if ({(8'hb7)})
                    begin
                      reg2157 <= reg2130[(2'h3):(1'h1)];
                      reg2158 <= (^~$unsigned($signed((wire2126 ?
                          reg2136 : forvar2156))));
                    end
                  else
                    begin
                      reg2157 <= (~|(&wire2126));
                      reg2158 <= reg2141;
                      reg2159 <= ((8'hb1) & reg2157);
                      reg2160 <= (!($signed($signed(reg2141)) ?
                          reg2143[(3'h5):(2'h3)] : (~|(reg2135 ?
                              wire2127 : reg2142))));
                    end
                end
              if (forvar2155[(3'h6):(2'h3)])
                begin
                  for (forvar2161 = (1'h0); (forvar2161 < (2'h3)); forvar2161 = (forvar2161 + (1'h1)))
                    begin
                      reg2162 <= $signed($unsigned({reg2146[(4'hd):(4'h9)]}));
                    end
                  for (forvar2163 = (1'h0); (forvar2163 < (2'h2)); forvar2163 = (forvar2163 + (1'h1)))
                    begin
                      reg2164 <= {({$signed(reg2142)} - (+$signed((8'ha9))))};
                      reg2165 <= ({((^reg2145) & $unsigned(reg2159))} == (reg2130 ?
                          forvar2132 : {(^~reg2135)}));
                      reg2166 <= (+$unsigned({wire2126}));
                    end
                end
              else
                begin
                  for (forvar2161 = (1'h0); (forvar2161 < (2'h3)); forvar2161 = (forvar2161 + (1'h1)))
                    begin
                      reg2162 <= (~^((!(reg2134 ?
                          reg2159 : reg2138)) >= (^~reg2142[(4'hb):(2'h3)])));
                      reg2163 <= (((reg2143 && (^reg2137)) >= ((!forvar2134) <<< $unsigned(forvar2144))) ?
                          $unsigned(({reg2141} ?
                              reg2142 : reg2135)) : forvar2144);
                    end
                  if ($signed(wire2128))
                    begin
                      reg2164 <= ((($signed(reg2163) ~^ (reg2131 ?
                              reg2142 : forvar2144)) | (^(wire2124 ?
                              forvar2148 : reg2152))) ?
                          $signed({(reg2165 ?
                                  reg2142 : reg2164)}) : (((~(8'h9f)) ?
                                  reg2164 : (reg2154 ? reg2140 : reg2153)) ?
                              {{(8'hb1)}} : ((reg2163 ? wire2126 : reg2130) ?
                                  {(8'hb6)} : wire2123[(4'h8):(3'h5)])));
                    end
                  else
                    begin
                      reg2164 <= {(wire2129 ?
                              (-forvar2144) : $unsigned((+wire2126)))};
                    end
                  reg2165 <= forvar2132[(2'h2):(2'h2)];
                  for (forvar2166 = (1'h0); (forvar2166 < (2'h2)); forvar2166 = (forvar2166 + (1'h1)))
                    begin
                      reg2167 <= $signed($signed(reg2140));
                    end
                end
            end
          reg2168 <= (forvar2134 && ((+(forvar2161 ? reg2142 : (8'ha6))) ?
              (reg2140 < $signed(reg2159)) : $signed($unsigned(reg2162))));
        end
      else
        begin
          if (((^~$unsigned((reg2145 & reg2166))) ?
              reg2149[(1'h0):(1'h0)] : forvar2132[(3'h6):(3'h5)]))
            begin
              if ($signed({($signed((8'ha9)) ? reg2158 : {reg2136})}))
                begin
                  if ($unsigned($unsigned(reg2131[(3'h5):(1'h1)])))
                    begin
                      reg2132 <= reg2137[(3'h5):(2'h2)];
                      reg2133 <= $signed($signed(wire2127[(1'h1):(1'h1)]));
                      reg2134 <= ((!($signed((8'hb0)) ?
                          (reg2146 || wire2127) : reg2133)) >= ({(wire2129 ^ (8'hb0))} >> ((reg2152 & reg2158) ?
                          (wire2123 ^~ reg2152) : $signed(reg2137))));
                    end
                  else
                    begin
                      reg2132 <= ($signed($unsigned((wire2124 ?
                          reg2162 : (8'haa)))) * ($signed({reg2154}) >> (!(reg2162 < reg2140))));
                      reg2133 <= reg2165[(1'h1):(1'h1)];
                      reg2134 <= (^~(-{{forvar2134}}));
                    end
                  for (forvar2135 = (1'h0); (forvar2135 < (2'h2)); forvar2135 = (forvar2135 + (1'h1)))
                    begin
                      reg2136 <= (((+(reg2139 ? forvar2139 : (8'ha6))) ?
                              ((reg2132 & reg2151) & {reg2142}) : ($signed(forvar2150) ^ $unsigned(reg2143))) ?
                          (wire2123[(1'h1):(1'h0)] ?
                              reg2141[(3'h4):(2'h3)] : reg2166) : $unsigned(forvar2150));
                      reg2137 <= ((~$signed(((8'hb7) - (8'hba)))) ?
                          (~^(|(reg2139 | reg2140))) : $unsigned($signed((forvar2163 * (8'hb0)))));
                      reg2138 <= $signed($unsigned(forvar2139));
                    end
                end
              else
                begin
                  reg2132 <= ($unsigned(({reg2165} ?
                          $unsigned(forvar2166) : (|reg2137))) ?
                      $unsigned($signed($unsigned(reg2137))) : reg2142);
                  for (forvar2133 = (1'h0); (forvar2133 < (1'h0)); forvar2133 = (forvar2133 + (1'h1)))
                    begin
                      reg2134 <= (~|reg2143);
                      reg2135 <= ((((reg2168 <<< reg2152) * (reg2142 * wire2129)) ?
                              wire2127 : reg2157) ?
                          $unsigned((~&reg2140[(4'hb):(3'h5)])) : wire2127);
                      reg2136 <= {{(8'hb4)}};
                    end
                  if ($signed((((8'h9f) * $unsigned(reg2140)) | reg2130[(1'h0):(1'h0)])))
                    begin
                      reg2137 <= ($unsigned($signed((8'hb7))) <<< ($unsigned($unsigned(reg2160)) && $signed($signed((8'hb7)))));
                      reg2138 <= ($signed(((wire2129 | reg2141) << (forvar2161 ?
                          reg2136 : forvar2135))) != reg2135[(2'h3):(2'h2)]);
                      reg2139 <= $signed($unsigned($unsigned((reg2165 < (8'hb0)))));
                      reg2140 <= $signed((reg2131[(1'h1):(1'h1)] ?
                          reg2168[(1'h1):(1'h1)] : {(forvar2166 <<< wire2127)}));
                    end
                  else
                    begin
                      reg2137 <= $unsigned((|$signed(wire2125)));
                      reg2138 <= $signed($unsigned({(reg2166 ?
                              reg2140 : wire2124)}));
                      reg2139 <= ((($unsigned(forvar2150) + (forvar2148 >> reg2154)) ?
                              (reg2141[(1'h0):(1'h0)] == {(8'hb1)}) : ((~&(8'had)) ?
                                  (+(8'hb2)) : (~|reg2153))) ?
                          forvar2133 : $signed($signed((forvar2144 ?
                              wire2123 : forvar2133))));
                    end
                end
              for (forvar2141 = (1'h0); (forvar2141 < (2'h3)); forvar2141 = (forvar2141 + (1'h1)))
                begin
                  if ($unsigned({reg2163}))
                    begin
                      reg2142 <= $unsigned(forvar2161);
                      reg2143 <= {({$unsigned(wire2124)} * (&reg2149[(1'h0):(1'h0)]))};
                      reg2144 <= (reg2153 ?
                          forvar2134 : $unsigned(forvar2134[(3'h5):(3'h5)]));
                      reg2145 <= $unsigned({(~(reg2141 ?
                              forvar2156 : forvar2156))});
                    end
                  else
                    begin
                      reg2142 <= ((8'ha5) >> (~|($signed((8'hb6)) >= reg2164)));
                      reg2143 <= {$unsigned(reg2162)};
                      reg2144 <= ($signed((~(forvar2148 ? reg2157 : reg2145))) ?
                          ((reg2151 ^ (reg2151 ? reg2153 : reg2149)) ?
                              ((^reg2136) & ((8'ha7) ?
                                  forvar2150 : reg2134)) : {(reg2146 * reg2130)}) : ({(wire2127 ?
                                      wire2125 : wire2124)} ?
                              reg2146 : $unsigned({(8'hb5)})));
                    end
                  reg2146 <= $signed(($signed((reg2166 ^ (8'ha3))) << wire2127));
                  for (forvar2147 = (1'h0); (forvar2147 < (2'h3)); forvar2147 = (forvar2147 + (1'h1)))
                    begin
                      reg2148 <= reg2149[(2'h2):(1'h0)];
                      reg2149 <= $unsigned((-$unsigned($signed(forvar2144))));
                      reg2150 <= reg2159[(3'h4):(3'h4)];
                      reg2151 <= ((^(reg2136[(3'h6):(3'h4)] ?
                          (reg2146 >= wire2127) : forvar2139)) * reg2137);
                    end
                  for (forvar2152 = (1'h0); (forvar2152 < (1'h0)); forvar2152 = (forvar2152 + (1'h1)))
                    begin
                      reg2153 <= forvar2152;
                      reg2154 <= (~|(reg2147 ?
                          ($unsigned(wire2129) * $signed(reg2135)) : (forvar2147 * reg2163)));
                      reg2155 <= $signed($signed(forvar2144));
                      reg2156 <= forvar2144[(3'h6):(1'h1)];
                    end
                end
            end
          else
            begin
              if ((8'ha7))
                begin
                  reg2132 <= reg2156[(4'hd):(4'h9)];
                  reg2133 <= $unsigned(reg2142);
                  reg2134 <= reg2132[(1'h1):(1'h1)];
                end
              else
                begin
                  reg2132 <= reg2135;
                  for (forvar2133 = (1'h0); (forvar2133 < (2'h2)); forvar2133 = (forvar2133 + (1'h1)))
                    begin
                      reg2134 <= ((-((forvar2155 ~^ forvar2155) && (~|reg2166))) ?
                          {($signed((8'hb2)) ?
                                  $unsigned(reg2136) : (reg2139 ?
                                      reg2137 : reg2137))} : ((~&(reg2167 <= reg2144)) ?
                              reg2150[(1'h0):(1'h0)] : {reg2156[(4'he):(3'h6)]}));
                      reg2135 <= ((({forvar2148} << (reg2138 ?
                              forvar2144 : reg2144)) * {(forvar2161 && (8'hb4))}) ?
                          reg2133 : (reg2167[(2'h2):(2'h2)] ?
                              $unsigned(((8'h9f) ?
                                  reg2140 : reg2131)) : $signed((forvar2141 ?
                                  reg2141 : reg2132))));
                      reg2136 <= (forvar2135 ? (8'hab) : forvar2133);
                    end
                end
              for (forvar2137 = (1'h0); (forvar2137 < (2'h3)); forvar2137 = (forvar2137 + (1'h1)))
                begin
                  reg2138 <= $signed(({(reg2152 ?
                          reg2133 : wire2127)} ^ reg2153[(3'h4):(1'h0)]));
                end
              reg2139 <= forvar2161;
              reg2140 <= {(forvar2141[(3'h4):(1'h0)] >= forvar2141[(4'hb):(3'h4)])};
            end
          for (forvar2157 = (1'h0); (forvar2157 < (1'h1)); forvar2157 = (forvar2157 + (1'h1)))
            begin
              reg2158 <= (reg2156[(1'h0):(1'h0)] ?
                  $signed(forvar2155[(3'h7):(3'h6)]) : (!reg2145));
              for (forvar2159 = (1'h0); (forvar2159 < (2'h3)); forvar2159 = (forvar2159 + (1'h1)))
                begin
                  reg2160 <= {reg2151};
                  reg2161 <= ($signed((+(-forvar2155))) ?
                      $unsigned(reg2165[(4'h9):(3'h5)]) : reg2163);
                  for (forvar2162 = (1'h0); (forvar2162 < (2'h2)); forvar2162 = (forvar2162 + (1'h1)))
                    begin
                      reg2163 <= $signed($unsigned($unsigned((reg2138 ?
                          (8'haf) : reg2166))));
                      reg2164 <= reg2166[(4'hc):(3'h4)];
                    end
                end
            end
          if ((8'ha9))
            begin
              if (($signed($signed($signed(reg2164))) ?
                  reg2167[(3'h5):(2'h2)] : (~|reg2168)))
                begin
                  if (wire2128[(3'h4):(2'h2)])
                    begin
                      reg2165 <= reg2154[(2'h3):(2'h3)];
                      reg2166 <= (|(~^$unsigned(((8'ha6) >> (8'ha8)))));
                      reg2167 <= (~wire2126[(2'h3):(1'h1)]);
                      reg2168 <= $unsigned($signed($signed((forvar2135 == forvar2148))));
                    end
                  else
                    begin
                      reg2165 <= reg2166[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  if ($signed(reg2160))
                    begin
                      reg2165 <= {$signed($signed((forvar2132 ?
                              (8'hb6) : reg2144)))};
                      reg2166 <= forvar2148;
                    end
                  else
                    begin
                      reg2165 <= ((8'hb4) ?
                          $signed($signed($unsigned(reg2139))) : forvar2132[(4'h9):(1'h0)]);
                      reg2166 <= {$signed(reg2153[(2'h3):(2'h3)])};
                      reg2167 <= ($unsigned(forvar2152) ?
                          $unsigned((8'hba)) : ($unsigned(reg2149[(1'h0):(1'h0)]) ?
                              ({reg2151} && $signed(forvar2144)) : $unsigned((~|reg2166))));
                      reg2168 <= ({$unsigned((~|reg2131))} >>> (~^(!(8'hb7))));
                    end
                  if ($signed($unsigned($unsigned($unsigned(reg2130)))))
                    begin
                      reg2169 <= (~^((~reg2134) && $signed((reg2145 ?
                          forvar2144 : reg2162))));
                      reg2170 <= ((~|forvar2135) >>> forvar2163);
                    end
                  else
                    begin
                      reg2169 <= ((((reg2141 >= forvar2155) ~^ $unsigned(reg2133)) == ((8'hb7) == $signed(wire2123))) ?
                          (({reg2132} >> $signed(wire2124)) ?
                              wire2125[(3'h4):(1'h0)] : reg2147) : (~|$unsigned(reg2140[(1'h1):(1'h0)])));
                      reg2170 <= reg2166;
                      reg2171 <= ((8'hb0) >= $signed($unsigned({forvar2150})));
                    end
                end
              if (((8'hb6) & (^reg2132[(3'h6):(2'h3)])))
                begin
                  for (forvar2172 = (1'h0); (forvar2172 < (1'h0)); forvar2172 = (forvar2172 + (1'h1)))
                    begin
                      reg2173 <= reg2152[(3'h5):(1'h0)];
                    end
                end
              else
                begin
                  reg2172 <= wire2124;
                end
              for (forvar2174 = (1'h0); (forvar2174 < (2'h3)); forvar2174 = (forvar2174 + (1'h1)))
                begin
                  for (forvar2175 = (1'h0); (forvar2175 < (2'h2)); forvar2175 = (forvar2175 + (1'h1)))
                    begin
                      reg2176 <= $signed(reg2166[(3'h7):(2'h3)]);
                      reg2177 <= $unsigned((8'hb3));
                      reg2178 <= $unsigned((((-wire2125) <= {reg2151}) ?
                          reg2152 : reg2161[(3'h4):(1'h1)]));
                    end
                  for (forvar2179 = (1'h0); (forvar2179 < (2'h3)); forvar2179 = (forvar2179 + (1'h1)))
                    begin
                      reg2180 <= $unsigned($signed((~^forvar2141)));
                      reg2181 <= (~|(reg2131[(3'h7):(2'h2)] - $signed($unsigned(reg2159))));
                      reg2182 <= {reg2164};
                    end
                  if ((^~forvar2179))
                    begin
                      reg2183 <= ((~|(forvar2135 ?
                              (reg2144 || reg2172) : (reg2173 >> reg2152))) ?
                          ($unsigned($signed(wire2125)) == reg2182) : ($signed((forvar2134 ?
                                  reg2143 : reg2169)) ?
                              ((-reg2178) ^ (reg2173 ^ (8'hba))) : $unsigned($unsigned((8'hab)))));
                      reg2184 <= ($unsigned(($signed(wire2129) ?
                              $unsigned(reg2160) : reg2156[(1'h0):(1'h0)])) ?
                          $unsigned($signed((-forvar2141))) : (|reg2161[(1'h1):(1'h1)]));
                      reg2185 <= $unsigned($signed(((reg2182 ?
                              forvar2175 : reg2149) ?
                          $signed(forvar2139) : {reg2130})));
                      reg2186 <= {(&((8'ha6) ?
                              reg2140[(2'h3):(2'h2)] : reg2149))};
                    end
                  else
                    begin
                      reg2183 <= ((^reg2150) ?
                          reg2165[(1'h0):(1'h0)] : ((!((8'had) ?
                              (8'hb3) : (8'hb7))) >> $unsigned((reg2148 ^~ reg2168))));
                      reg2184 <= $signed($unsigned(({(8'had)} ?
                          (reg2139 ? reg2158 : reg2145) : $signed((8'h9e)))));
                      reg2185 <= wire2125[(2'h2):(2'h2)];
                    end
                end
            end
          else
            begin
              for (forvar2165 = (1'h0); (forvar2165 < (2'h3)); forvar2165 = (forvar2165 + (1'h1)))
                begin
                  for (forvar2166 = (1'h0); (forvar2166 < (2'h2)); forvar2166 = (forvar2166 + (1'h1)))
                    begin
                      reg2167 <= $unsigned($unsigned({reg2160[(4'he):(1'h1)]}));
                      reg2168 <= (((~^(^~reg2148)) ? (-(~reg2141)) : (8'had)) ?
                          $unsigned(forvar2175[(1'h0):(1'h0)]) : ($unsigned(reg2151[(1'h1):(1'h0)]) != $signed(forvar2134[(1'h1):(1'h0)])));
                      reg2169 <= reg2182;
                    end
                end
              if (forvar2134)
                begin
                  for (forvar2170 = (1'h0); (forvar2170 < (2'h3)); forvar2170 = (forvar2170 + (1'h1)))
                    begin
                      reg2171 <= (-forvar2159[(3'h7):(3'h5)]);
                      reg2172 <= (((reg2159[(2'h3):(1'h0)] << $signed(reg2141)) ?
                          {{reg2181}} : (^(reg2185 ?
                              reg2141 : reg2133))) >> (($signed(forvar2152) ?
                          (wire2124 ^ reg2165) : {reg2160}) * reg2162[(4'hb):(4'hb)]));
                    end
                  for (forvar2173 = (1'h0); (forvar2173 < (2'h2)); forvar2173 = (forvar2173 + (1'h1)))
                    begin
                      reg2174 <= $unsigned(($unsigned($unsigned(reg2142)) == $signed((reg2151 ?
                          (8'hb6) : wire2124))));
                      reg2175 <= $signed(reg2132);
                      reg2176 <= ((reg2175 ?
                              ((~^reg2133) <= $signed((8'haf))) : $signed({reg2165})) ?
                          (~|$unsigned((~&reg2169))) : $unsigned((~&$unsigned(reg2165))));
                      reg2177 <= $signed($unsigned(reg2173[(1'h1):(1'h1)]));
                    end
                  reg2178 <= (!forvar2172);
                  for (forvar2179 = (1'h0); (forvar2179 < (2'h2)); forvar2179 = (forvar2179 + (1'h1)))
                    begin
                      reg2180 <= (|$signed(reg2139));
                      reg2181 <= $signed($signed((!(reg2143 == (8'hb6)))));
                    end
                end
              else
                begin
                  if (((forvar2155[(3'h7):(3'h6)] ?
                      {(forvar2179 && forvar2163)} : $signed($signed(reg2180))) ^~ (($signed((8'hae)) ~^ (reg2182 ^ reg2168)) ?
                      forvar2174 : wire2129[(4'h8):(3'h7)])))
                    begin
                      reg2170 <= ({(-((8'hb3) ?
                              reg2177 : reg2156))} << (|$unsigned(forvar2155)));
                      reg2171 <= (reg2153[(2'h3):(2'h2)] <<< (((wire2126 ?
                          reg2183 : reg2147) - (~^reg2166)) != {(^reg2149)}));
                      reg2172 <= ($signed($unsigned((wire2127 + reg2149))) ^ $unsigned((forvar2179 ?
                          (!(8'hb5)) : (reg2182 <<< reg2156))));
                      reg2173 <= (reg2138 ?
                          ($unsigned((+reg2139)) ?
                              reg2162[(3'h5):(1'h0)] : reg2171[(1'h0):(1'h0)]) : $unsigned($unsigned($signed(forvar2135))));
                    end
                  else
                    begin
                      reg2170 <= (wire2124 ?
                          forvar2133[(1'h1):(1'h1)] : $signed(reg2132[(2'h2):(1'h1)]));
                    end
                  if ($unsigned($unsigned(forvar2166)))
                    begin
                      reg2174 <= ($signed(($signed(reg2185) << reg2145)) ?
                          $unsigned(forvar2165) : ((~(forvar2166 ?
                                  reg2174 : reg2165)) ?
                              (^~$signed(reg2172)) : ({reg2152} == (~reg2169))));
                      reg2175 <= {{((forvar2144 ?
                                  (8'h9c) : reg2141) & $signed((8'hb6)))}};
                    end
                  else
                    begin
                      reg2174 <= $signed(reg2139[(4'hb):(3'h5)]);
                      reg2175 <= ($unsigned($signed($signed(reg2156))) * $signed($signed((reg2136 < forvar2166))));
                    end
                  if ($signed(forvar2134))
                    begin
                      reg2176 <= (^{({reg2133} ?
                              wire2128[(4'hf):(2'h3)] : (reg2178 ?
                                  (8'haa) : reg2142))});
                      reg2177 <= $signed(forvar2163[(4'h8):(2'h3)]);
                    end
                  else
                    begin
                      reg2176 <= {(~$unsigned((~^reg2155)))};
                      reg2177 <= (~^$signed(forvar2137));
                      reg2178 <= ($signed($signed($unsigned(reg2175))) ?
                          forvar2135[(1'h1):(1'h1)] : forvar2161[(3'h4):(1'h0)]);
                    end
                end
              reg2182 <= ($signed((~|reg2170[(1'h0):(1'h0)])) * (wire2125[(1'h1):(1'h0)] <= $unsigned($signed(reg2174))));
            end
          if (reg2152[(3'h4):(2'h2)])
            begin
              if ({(($signed(reg2134) + (reg2178 || reg2164)) + $signed(reg2153))})
                begin
                  if ($signed((~|$unsigned((reg2156 ? reg2183 : reg2152)))))
                    begin
                      reg2187 <= $signed(forvar2159);
                      reg2188 <= reg2175[(4'h9):(3'h5)];
                      reg2189 <= $signed((forvar2165 ?
                          $signed(reg2144[(1'h1):(1'h1)]) : reg2161[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg2187 <= ((8'h9d) <<< (((wire2128 ?
                              reg2175 : reg2185) >> $unsigned((8'h9f))) ?
                          reg2177 : (~^$signed(reg2160))));
                      reg2188 <= (8'ha7);
                      reg2189 <= $signed($unsigned((8'h9f)));
                      reg2190 <= {(reg2134 ?
                              ((reg2180 > reg2186) ?
                                  forvar2162[(2'h2):(1'h1)] : (wire2126 ?
                                      reg2169 : wire2125)) : $signed((~reg2177)))};
                    end
                end
              else
                begin
                  if (((~reg2180[(4'h9):(3'h6)]) > (8'ha7)))
                    begin
                      reg2187 <= forvar2157[(4'hb):(2'h3)];
                      reg2188 <= $signed($signed($signed((!reg2157))));
                    end
                  else
                    begin
                      reg2187 <= (reg2184[(2'h3):(2'h2)] ?
                          $unsigned({(8'h9d)}) : $signed(((~&(8'hb6)) ?
                              ((8'haf) + reg2166) : $unsigned(wire2126))));
                      reg2188 <= $signed(($unsigned((reg2159 | reg2141)) ?
                          (reg2186[(1'h0):(1'h0)] << $signed(forvar2132)) : reg2151));
                      reg2189 <= $signed(forvar2152);
                    end
                end
              if (reg2138[(3'h4):(1'h0)])
                begin
                  for (forvar2191 = (1'h0); (forvar2191 < (1'h1)); forvar2191 = (forvar2191 + (1'h1)))
                    begin
                      reg2192 <= $unsigned(reg2158);
                      reg2193 <= (~(reg2167[(3'h6):(3'h5)] | (((8'haf) >= reg2192) ?
                          forvar2173 : (^reg2177))));
                    end
                  reg2194 <= $unsigned(((((8'hb6) ? forvar2148 : reg2160) ?
                          $unsigned(forvar2132) : $unsigned(reg2184)) ?
                      $signed((^~wire2129)) : $signed(wire2124[(1'h0):(1'h0)])));
                  for (forvar2195 = (1'h0); (forvar2195 < (2'h3)); forvar2195 = (forvar2195 + (1'h1)))
                    begin
                      reg2196 <= $signed((((forvar2155 & reg2148) || $unsigned(forvar2159)) ?
                          {forvar2174[(3'h6):(3'h6)]} : reg2140));
                    end
                end
              else
                begin
                  for (forvar2191 = (1'h0); (forvar2191 < (1'h1)); forvar2191 = (forvar2191 + (1'h1)))
                    begin
                      reg2192 <= (!forvar2170[(1'h1):(1'h1)]);
                      reg2193 <= reg2154;
                      reg2194 <= reg2154;
                      reg2195 <= (!reg2190[(4'hd):(4'hd)]);
                    end
                  reg2196 <= ($unsigned(((~^wire2127) >>> $signed(reg2173))) ?
                      $unsigned((-{forvar2150})) : reg2147);
                end
            end
          else
            begin
              for (forvar2187 = (1'h0); (forvar2187 < (2'h3)); forvar2187 = (forvar2187 + (1'h1)))
                begin
                  if ((($signed({forvar2156}) * (-(reg2168 >>> forvar2150))) * ({{forvar2155}} ?
                      forvar2166 : reg2162[(3'h7):(2'h2)])))
                    begin
                      reg2188 <= (^~(((reg2150 ?
                          reg2134 : reg2192) || {reg2133}) * (~^reg2157[(1'h0):(1'h0)])));
                      reg2189 <= (~|$unsigned($unsigned($unsigned(reg2175))));
                      reg2190 <= $unsigned(forvar2135[(1'h1):(1'h0)]);
                      reg2191 <= (reg2141 >> $signed(forvar2144));
                    end
                  else
                    begin
                      reg2188 <= ((~^(~forvar2175)) >>> {forvar2172});
                      reg2189 <= $signed((~^($unsigned(forvar2141) ?
                          wire2126 : ((8'hb1) << forvar2147))));
                    end
                end
              if ($unsigned({reg2135}))
                begin
                  for (forvar2192 = (1'h0); (forvar2192 < (2'h3)); forvar2192 = (forvar2192 + (1'h1)))
                    begin
                      reg2193 <= ((^~(^{(8'h9f)})) << $unsigned(((forvar2139 ?
                          forvar2148 : reg2190) ^~ $unsigned(wire2125))));
                      reg2194 <= reg2131;
                      reg2195 <= $unsigned($unsigned(reg2176[(3'h5):(1'h0)]));
                    end
                end
              else
                begin
                  reg2192 <= reg2193;
                  for (forvar2193 = (1'h0); (forvar2193 < (2'h2)); forvar2193 = (forvar2193 + (1'h1)))
                    begin
                      reg2194 <= (8'had);
                      reg2195 <= $unsigned(($unsigned(forvar2141[(4'h9):(4'h8)]) & reg2159[(2'h3):(1'h0)]));
                      reg2196 <= $unsigned((reg2130 && $unsigned((forvar2133 >>> reg2147))));
                      reg2197 <= $signed(wire2128);
                    end
                  for (forvar2198 = (1'h0); (forvar2198 < (2'h3)); forvar2198 = (forvar2198 + (1'h1)))
                    begin
                      reg2199 <= (-forvar2139[(3'h7):(3'h6)]);
                    end
                end
              for (forvar2200 = (1'h0); (forvar2200 < (2'h2)); forvar2200 = (forvar2200 + (1'h1)))
                begin
                  for (forvar2201 = (1'h0); (forvar2201 < (1'h1)); forvar2201 = (forvar2201 + (1'h1)))
                    begin
                      reg2202 <= (~reg2190[(4'hd):(3'h6)]);
                      reg2203 <= $signed(($unsigned({forvar2179}) & forvar2161));
                      reg2204 <= $unsigned((|$signed((forvar2162 ?
                          reg2142 : reg2168))));
                      reg2205 <= (-$signed(forvar2166[(2'h3):(2'h3)]));
                    end
                  for (forvar2206 = (1'h0); (forvar2206 < (2'h3)); forvar2206 = (forvar2206 + (1'h1)))
                    begin
                      reg2207 <= reg2196;
                      reg2208 <= forvar2161[(3'h5):(1'h0)];
                      reg2209 <= reg2182;
                      reg2210 <= (({(reg2199 ?
                              (8'hb8) : reg2151)} <= {$unsigned((8'hb6))}) >> ((forvar2152 ?
                          (~forvar2195) : reg2203) < forvar2152));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if (forvar2141)
        begin
          reg2211 <= (^~({reg2194[(3'h7):(3'h6)]} + $unsigned(((8'ha6) ^ reg2147))));
          for (forvar2212 = (1'h0); (forvar2212 < (2'h3)); forvar2212 = (forvar2212 + (1'h1)))
            begin
              for (forvar2213 = (1'h0); (forvar2213 < (1'h1)); forvar2213 = (forvar2213 + (1'h1)))
                begin
                  if ($signed((forvar2150 ?
                      (wire2125 ?
                          $signed((8'hba)) : (forvar2159 ?
                              reg2192 : forvar2166)) : forvar2162)))
                    begin
                      reg2214 <= ((reg2147 ?
                          $unsigned($signed(reg2145)) : forvar2135[(1'h1):(1'h0)]) || $unsigned(reg2188[(1'h0):(1'h0)]));
                      reg2215 <= (~|(((reg2196 ?
                              reg2190 : reg2184) << ((8'ha7) > reg2193)) ?
                          $unsigned($signed(reg2192)) : (8'hb0)));
                    end
                  else
                    begin
                      reg2214 <= $unsigned(($unsigned($signed((8'hab))) > $signed({reg2140})));
                      reg2215 <= forvar2198[(4'h8):(3'h6)];
                      reg2216 <= ((~^$unsigned((reg2189 != forvar2200))) && ((~$signed(reg2172)) >> reg2171));
                      reg2217 <= reg2163[(3'h5):(2'h3)];
                    end
                  if ($unsigned($signed((wire2125[(3'h4):(2'h2)] ?
                      {reg2189} : ((8'hb3) < forvar2165)))))
                    begin
                      reg2218 <= (8'ha9);
                      reg2219 <= $signed(forvar2159);
                      reg2220 <= $unsigned(forvar2159);
                      reg2221 <= (forvar2213[(1'h1):(1'h1)] ?
                          $unsigned($signed({reg2130})) : $signed(forvar2144[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg2218 <= (~|reg2205[(3'h7):(1'h1)]);
                      reg2219 <= $signed(forvar2174);
                    end
                end
              reg2222 <= {$signed($signed($unsigned(reg2194)))};
            end
          if ((!((~|(forvar2175 ?
              reg2161 : (8'ha5))) ~^ $unsigned((^~reg2190)))))
            begin
              if ({(($signed(reg2159) ? $unsigned(reg2154) : reg2165) ?
                      (~&reg2203) : ($unsigned(reg2154) ?
                          {(8'h9e)} : (forvar2132 >>> reg2142)))})
                begin
                  reg2223 <= reg2215;
                  if ((!$unsigned(reg2141[(3'h7):(3'h5)])))
                    begin
                      reg2224 <= $unsigned(($unsigned(((8'ha8) * forvar2135)) ^~ $unsigned((reg2182 >> (8'hb0)))));
                    end
                  else
                    begin
                      reg2224 <= (+$unsigned($signed(((8'ha4) != reg2195))));
                      reg2225 <= (^~reg2149);
                    end
                end
              else
                begin
                  if ((8'hab))
                    begin
                      reg2223 <= (reg2220 ?
                          reg2142 : $unsigned(forvar2156[(3'h5):(2'h2)]));
                      reg2224 <= (forvar2134 <<< $signed($unsigned(reg2222)));
                      reg2225 <= $unsigned($signed($unsigned({reg2196})));
                      reg2226 <= (reg2162[(2'h3):(1'h1)] ?
                          $signed((reg2202 ^ (&forvar2155))) : forvar2161[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg2223 <= {reg2161};
                      reg2224 <= ((reg2161 >>> reg2181[(3'h6):(1'h0)]) - ($unsigned(reg2166) || ((reg2154 ^ reg2141) || reg2134)));
                      reg2225 <= (|{((reg2226 < reg2216) ?
                              $unsigned((8'hab)) : $signed(forvar2165))});
                    end
                end
              if ($unsigned((reg2211 ~^ $signed(reg2174[(3'h4):(2'h2)]))))
                begin
                  reg2227 <= ({(reg2157[(3'h5):(1'h1)] == forvar2135[(1'h0):(1'h0)])} ?
                      (forvar2159[(3'h4):(2'h3)] ?
                          $unsigned(reg2207[(2'h2):(2'h2)]) : ($unsigned((8'hb0)) ?
                              forvar2200 : $signed(reg2214))) : (|wire2125));
                  for (forvar2228 = (1'h0); (forvar2228 < (2'h2)); forvar2228 = (forvar2228 + (1'h1)))
                    begin
                      reg2229 <= reg2134;
                      reg2230 <= (~|reg2139);
                      reg2231 <= forvar2175[(2'h2):(2'h2)];
                      reg2232 <= (&$signed(($unsigned(forvar2135) ~^ (!forvar2150))));
                    end
                  for (forvar2233 = (1'h0); (forvar2233 < (1'h0)); forvar2233 = (forvar2233 + (1'h1)))
                    begin
                      reg2234 <= {reg2195[(3'h6):(2'h3)]};
                      reg2235 <= $signed($signed(({reg2232} ?
                          (reg2193 == reg2173) : (~(8'hae)))));
                      reg2236 <= reg2195[(4'ha):(3'h6)];
                    end
                end
              else
                begin
                  for (forvar2227 = (1'h0); (forvar2227 < (2'h3)); forvar2227 = (forvar2227 + (1'h1)))
                    begin
                      reg2228 <= ((forvar2150[(3'h5):(2'h2)] ?
                          ({reg2196} ?
                              (^~reg2149) : (~^reg2191)) : {{reg2142}}) < (^~(-(reg2224 ?
                          (8'haf) : forvar2166))));
                      reg2229 <= wire2125;
                    end
                  reg2230 <= $signed((((forvar2201 ? reg2210 : (8'hb6)) ?
                      (forvar2161 ?
                          forvar2155 : reg2195) : (~^reg2229)) >>> (~&reg2142)));
                  reg2231 <= $unsigned((reg2163[(3'h6):(1'h1)] ?
                      (reg2202[(2'h3):(1'h0)] ?
                          reg2214[(4'he):(4'ha)] : $signed(reg2210)) : $unsigned(((8'hac) ?
                          (8'hb2) : (8'ha2)))));
                  for (forvar2232 = (1'h0); (forvar2232 < (2'h3)); forvar2232 = (forvar2232 + (1'h1)))
                    begin
                      reg2233 <= wire2128[(4'hf):(3'h6)];
                      reg2234 <= (((reg2199[(3'h4):(3'h4)] ?
                          (reg2151 ?
                              reg2180 : reg2192) : (&reg2177)) < {$unsigned(reg2139)}) & (reg2190 & forvar2206));
                    end
                end
              if ($unsigned($unsigned(forvar2228[(3'h5):(3'h4)])))
                begin
                  if ($signed(forvar2134[(2'h3):(2'h3)]))
                    begin
                      reg2237 <= (8'ha7);
                    end
                  else
                    begin
                      reg2237 <= {reg2209};
                      reg2238 <= (~^$signed(reg2151[(2'h2):(1'h0)]));
                      reg2239 <= $unsigned((|$signed((forvar2170 ?
                          forvar2201 : forvar2141))));
                      reg2240 <= reg2184;
                    end
                end
              else
                begin
                  if (($unsigned($signed($signed(reg2228))) || $signed($signed((forvar2195 ?
                      forvar2165 : reg2133)))))
                    begin
                      reg2237 <= forvar2206[(1'h1):(1'h0)];
                      reg2238 <= (&(((~|forvar2195) - forvar2175) << $unsigned($unsigned(reg2190))));
                      reg2239 <= reg2155[(4'ha):(2'h2)];
                      reg2240 <= $signed($signed({$signed(reg2190)}));
                    end
                  else
                    begin
                      reg2237 <= (~$unsigned($unsigned((reg2218 ?
                          forvar2161 : reg2234))));
                      reg2238 <= reg2236[(1'h0):(1'h0)];
                    end
                end
            end
          else
            begin
              reg2223 <= (|reg2232);
              if ((($unsigned(reg2219) * (^reg2139[(4'h9):(1'h0)])) ?
                  (~|(+(^~reg2167))) : reg2234))
                begin
                  for (forvar2224 = (1'h0); (forvar2224 < (2'h2)); forvar2224 = (forvar2224 + (1'h1)))
                    begin
                      reg2225 <= $unsigned((reg2131[(1'h0):(1'h0)] ^~ $unsigned($unsigned(forvar2193))));
                    end
                  reg2226 <= {(~^$signed((reg2192 ? forvar2147 : reg2219)))};
                  for (forvar2227 = (1'h0); (forvar2227 < (2'h2)); forvar2227 = (forvar2227 + (1'h1)))
                    begin
                      reg2228 <= forvar2224[(3'h7):(3'h5)];
                    end
                end
              else
                begin
                  for (forvar2224 = (1'h0); (forvar2224 < (2'h2)); forvar2224 = (forvar2224 + (1'h1)))
                    begin
                      reg2225 <= $unsigned((~^$unsigned($signed(reg2230))));
                      reg2226 <= (reg2196[(4'he):(1'h1)] ?
                          ($signed((~forvar2133)) ?
                              (^~$unsigned(forvar2232)) : forvar2232[(2'h3):(1'h1)]) : $unsigned(($unsigned(reg2159) ?
                              (reg2236 ?
                                  forvar2141 : forvar2159) : $signed(wire2125))));
                    end
                end
              if ((~|((-reg2207) << (reg2218 ?
                  wire2123[(2'h3):(2'h2)] : (reg2236 ? forvar2144 : reg2240)))))
                begin
                  for (forvar2229 = (1'h0); (forvar2229 < (2'h3)); forvar2229 = (forvar2229 + (1'h1)))
                    begin
                      reg2230 <= $unsigned(forvar2150);
                      reg2231 <= {{reg2230}};
                      reg2232 <= forvar2228[(2'h3):(1'h0)];
                      reg2233 <= forvar2161[(1'h1):(1'h0)];
                    end
                  if ($signed({(|$signed(forvar2148))}))
                    begin
                      reg2234 <= (-$signed(forvar2155));
                    end
                  else
                    begin
                      reg2234 <= (reg2157[(3'h5):(2'h2)] ?
                          $unsigned($unsigned($unsigned(reg2167))) : reg2155);
                      reg2235 <= {$unsigned($unsigned($unsigned(reg2193)))};
                      reg2236 <= ($signed(((forvar2173 >>> reg2145) ^~ (forvar2132 ?
                              reg2231 : reg2134))) ?
                          (((reg2236 ? forvar2147 : reg2234) ?
                              reg2163[(3'h5):(3'h5)] : (reg2220 != wire2123)) >> $signed($signed(forvar2213))) : forvar2173);
                    end
                  if (reg2175)
                    begin
                      reg2237 <= {(+$signed((+reg2191)))};
                    end
                  else
                    begin
                      reg2237 <= $unsigned($signed(forvar2165));
                    end
                end
              else
                begin
                  if ($signed((forvar2224[(2'h2):(1'h0)] & $unsigned($signed((8'hb8))))))
                    begin
                      reg2229 <= (({(forvar2175 ? reg2172 : reg2227)} ?
                              $unsigned((reg2183 ?
                                  reg2187 : reg2178)) : $signed({reg2166})) ?
                          $signed(forvar2198) : {{(reg2211 * wire2123)}});
                      reg2230 <= {($signed($unsigned(forvar2172)) ?
                              $signed(forvar2224[(3'h7):(3'h5)]) : (^(reg2183 <= reg2143)))};
                      reg2231 <= $unsigned(reg2151[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg2229 <= ((($signed((8'ha9)) || reg2220[(3'h5):(2'h3)]) || forvar2201[(4'ha):(3'h6)]) > $signed(((reg2171 ?
                              reg2229 : (8'ha2)) ?
                          forvar2134 : reg2142[(4'he):(4'h8)])));
                    end
                  if ((|(-$unsigned(forvar2134))))
                    begin
                      reg2232 <= reg2170;
                      reg2233 <= $signed($signed(forvar2172[(3'h4):(1'h1)]));
                      reg2234 <= forvar2174[(4'hd):(3'h5)];
                    end
                  else
                    begin
                      reg2232 <= $signed((^$signed(reg2153)));
                      reg2233 <= reg2160;
                    end
                end
            end
          if ((forvar2172[(2'h2):(2'h2)] ^ $signed(($unsigned(reg2228) <= $signed(reg2154)))))
            begin
              reg2241 <= (reg2159 != ({(8'ha6)} <= reg2234[(2'h2):(2'h2)]));
            end
          else
            begin
              reg2241 <= (reg2167 ?
                  (forvar2139 ?
                      $unsigned(((8'hb3) - (8'hb3))) : $unsigned((reg2228 <<< reg2199))) : (|$signed(reg2216)));
              if ((^~$signed((8'hb6))))
                begin
                  reg2242 <= ($unsigned($signed($signed(reg2226))) >>> reg2209[(3'h4):(3'h4)]);
                  for (forvar2243 = (1'h0); (forvar2243 < (1'h0)); forvar2243 = (forvar2243 + (1'h1)))
                    begin
                      reg2244 <= (reg2189 & $signed(reg2152[(1'h0):(1'h0)]));
                      reg2245 <= $signed({(|$signed((8'hba)))});
                      reg2246 <= $unsigned((~(^~$unsigned((8'h9e)))));
                      reg2247 <= {$signed($unsigned((reg2181 ?
                              reg2226 : (8'ha9))))};
                    end
                  if (({reg2221} >= (~reg2190[(3'h5):(2'h3)])))
                    begin
                      reg2248 <= (reg2219[(1'h0):(1'h0)] == $unsigned($unsigned((reg2230 ?
                          reg2226 : reg2193))));
                      reg2249 <= reg2191;
                    end
                  else
                    begin
                      reg2248 <= $signed($unsigned({$unsigned(reg2171)}));
                      reg2249 <= $unsigned((|(8'haf)));
                    end
                  if (forvar2172[(2'h3):(2'h3)])
                    begin
                      reg2250 <= (|$unsigned($signed($unsigned(reg2233))));
                      reg2251 <= forvar2233;
                    end
                  else
                    begin
                      reg2250 <= reg2250[(2'h2):(2'h2)];
                      reg2251 <= reg2181;
                      reg2252 <= ((reg2176[(5'h10):(4'hf)] | (&$unsigned(reg2219))) ?
                          $signed(((reg2188 ?
                              (8'hae) : reg2169) ~^ forvar2206[(1'h1):(1'h1)])) : $signed(($unsigned((8'haa)) ?
                              (reg2188 << forvar2187) : reg2202[(2'h3):(2'h3)])));
                    end
                end
              else
                begin
                  for (forvar2242 = (1'h0); (forvar2242 < (2'h3)); forvar2242 = (forvar2242 + (1'h1)))
                    begin
                      reg2243 <= (+$unsigned(reg2218));
                      reg2244 <= $signed(((8'hb5) - reg2224));
                      reg2245 <= forvar2228[(3'h4):(1'h0)];
                      reg2246 <= $signed({(^~{reg2161})});
                    end
                  reg2247 <= $signed(wire2123[(2'h3):(1'h1)]);
                  for (forvar2248 = (1'h0); (forvar2248 < (1'h1)); forvar2248 = (forvar2248 + (1'h1)))
                    begin
                      reg2249 <= (((~(!reg2150)) ?
                              reg2228 : (reg2158[(4'he):(4'h9)] ^ {reg2183})) ?
                          reg2204 : (~&{$signed(reg2171)}));
                      reg2250 <= forvar2206[(4'hd):(1'h1)];
                      reg2251 <= reg2174;
                    end
                  if ((reg2248[(3'h4):(2'h3)] ~^ {forvar2233[(3'h4):(2'h3)]}))
                    begin
                      reg2252 <= (8'ha3);
                    end
                  else
                    begin
                      reg2252 <= $signed(forvar2155);
                      reg2253 <= reg2226;
                      reg2254 <= ((((forvar2163 <<< reg2176) >>> (-forvar2163)) + reg2196[(4'hb):(3'h5)]) <<< $signed($unsigned(reg2241)));
                      reg2255 <= $signed((reg2132 ?
                          $unsigned($unsigned(forvar2150)) : wire2126[(1'h1):(1'h0)]));
                    end
                end
              for (forvar2256 = (1'h0); (forvar2256 < (2'h2)); forvar2256 = (forvar2256 + (1'h1)))
                begin
                  for (forvar2257 = (1'h0); (forvar2257 < (1'h1)); forvar2257 = (forvar2257 + (1'h1)))
                    begin
                      reg2258 <= ((^reg2208[(3'h4):(2'h3)]) >> reg2234);
                      reg2259 <= reg2195[(4'hb):(4'hb)];
                      reg2260 <= (8'ha3);
                    end
                  reg2261 <= ({(8'ha6)} && reg2134);
                end
              if (reg2137)
                begin
                  if ($signed($unsigned(reg2214)))
                    begin
                      reg2262 <= ($signed({(wire2126 ^~ forvar2156)}) ?
                          reg2154[(4'h9):(3'h6)] : (~^forvar2229[(3'h7):(1'h0)]));
                      reg2263 <= {(reg2233[(2'h3):(1'h1)] ?
                              $signed((reg2235 ?
                                  forvar2148 : (8'hb1))) : ($unsigned((8'had)) ?
                                  forvar2192[(4'hc):(4'ha)] : reg2131))};
                      reg2264 <= reg2246;
                      reg2265 <= (forvar2173[(1'h1):(1'h1)] || $signed($signed((reg2263 ?
                          reg2196 : forvar2200))));
                    end
                  else
                    begin
                      reg2262 <= {($signed(reg2224) ?
                              reg2177[(3'h6):(1'h0)] : {$signed((8'hb6))})};
                      reg2263 <= (~|(reg2165 - forvar2161));
                      reg2264 <= reg2139;
                    end
                  reg2266 <= (~&{reg2164[(1'h0):(1'h0)]});
                  for (forvar2267 = (1'h0); (forvar2267 < (2'h3)); forvar2267 = (forvar2267 + (1'h1)))
                    begin
                      reg2268 <= (~^{(+(~|(8'hae)))});
                      reg2269 <= reg2193[(1'h1):(1'h0)];
                      reg2270 <= ((reg2136[(4'h9):(3'h7)] ?
                              forvar2150 : (~forvar2191)) ?
                          $unsigned((8'h9e)) : {{$unsigned(forvar2166)}});
                    end
                  for (forvar2271 = (1'h0); (forvar2271 < (2'h3)); forvar2271 = (forvar2271 + (1'h1)))
                    begin
                      reg2272 <= $signed(forvar2228);
                      reg2273 <= reg2199[(2'h3):(2'h3)];
                      reg2274 <= reg2236;
                      reg2275 <= $signed(($signed($signed(forvar2147)) << $unsigned($unsigned(reg2237))));
                    end
                end
              else
                begin
                  if (reg2218[(2'h2):(1'h1)])
                    begin
                      reg2262 <= reg2148;
                      reg2263 <= $unsigned($unsigned(reg2211));
                    end
                  else
                    begin
                      reg2262 <= (-(|reg2197[(1'h1):(1'h0)]));
                      reg2263 <= {forvar2206};
                    end
                  if ($unsigned(({reg2149[(3'h5):(3'h5)]} - $unsigned($signed(reg2152)))))
                    begin
                      reg2264 <= reg2246[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg2264 <= (^~$signed(reg2134));
                      reg2265 <= forvar2191;
                    end
                  reg2266 <= $signed(forvar2195[(2'h2):(1'h1)]);
                  for (forvar2267 = (1'h0); (forvar2267 < (2'h2)); forvar2267 = (forvar2267 + (1'h1)))
                    begin
                      reg2268 <= $signed(reg2174[(3'h6):(3'h4)]);
                      reg2269 <= reg2149[(1'h1):(1'h0)];
                      reg2270 <= (^(((forvar2163 ?
                          forvar2147 : reg2220) <<< (-reg2140)) >>> (&reg2258)));
                      reg2271 <= (($signed(reg2139[(4'hd):(2'h3)]) << wire2123[(4'hb):(3'h5)]) ?
                          ((8'ha9) <= ((reg2228 | reg2153) == (wire2126 * reg2219))) : {(((8'ha8) > forvar2193) + $unsigned(forvar2144))});
                    end
                end
            end
        end
      else
        begin
          reg2211 <= $unsigned((~&(reg2139[(3'h4):(2'h3)] + reg2228[(5'h10):(2'h2)])));
          for (forvar2212 = (1'h0); (forvar2212 < (1'h0)); forvar2212 = (forvar2212 + (1'h1)))
            begin
              for (forvar2213 = (1'h0); (forvar2213 < (1'h0)); forvar2213 = (forvar2213 + (1'h1)))
                begin
                  for (forvar2214 = (1'h0); (forvar2214 < (1'h0)); forvar2214 = (forvar2214 + (1'h1)))
                    begin
                      reg2215 <= ($signed($signed($signed(reg2216))) ?
                          reg2163[(3'h5):(3'h4)] : {$signed({reg2272})});
                      reg2216 <= reg2207[(1'h0):(1'h0)];
                      reg2217 <= $unsigned((reg2210[(3'h5):(3'h4)] == (((8'hb6) <<< reg2215) ?
                          (|reg2249) : (!reg2174))));
                      reg2218 <= wire2126[(4'h8):(3'h7)];
                    end
                  for (forvar2219 = (1'h0); (forvar2219 < (2'h3)); forvar2219 = (forvar2219 + (1'h1)))
                    begin
                      reg2220 <= reg2208[(3'h5):(1'h1)];
                    end
                  if ($signed(reg2222))
                    begin
                      reg2221 <= {(($unsigned(reg2150) >>> $unsigned((8'h9f))) ?
                              (8'ha8) : reg2237)};
                    end
                  else
                    begin
                      reg2221 <= (({$signed(reg2136)} >= forvar2224[(1'h0):(1'h0)]) ?
                          $unsigned(($signed(reg2268) & (reg2150 ?
                              forvar2212 : reg2239))) : forvar2248);
                      reg2222 <= $unsigned(($signed((reg2165 ?
                          forvar2191 : forvar2166)) >>> ($unsigned((8'hb5)) - (&reg2239))));
                    end
                  reg2223 <= {forvar2170};
                end
              if (reg2156[(4'hb):(4'hb)])
                begin
                  for (forvar2224 = (1'h0); (forvar2224 < (1'h1)); forvar2224 = (forvar2224 + (1'h1)))
                    begin
                      reg2225 <= (forvar2248[(2'h2):(2'h2)] ^ reg2211[(4'hb):(4'ha)]);
                      reg2226 <= reg2221;
                      reg2227 <= (+((^~$unsigned(reg2145)) ?
                          ($unsigned(forvar2135) ?
                              (reg2217 ?
                                  reg2220 : reg2186) : $signed(reg2251)) : reg2173[(3'h6):(1'h0)]));
                      reg2228 <= (~({$unsigned((8'hab))} * (~|forvar2172[(4'hc):(1'h0)])));
                    end
                  for (forvar2229 = (1'h0); (forvar2229 < (1'h1)); forvar2229 = (forvar2229 + (1'h1)))
                    begin
                      reg2230 <= $signed((8'ha6));
                    end
                end
              else
                begin
                  for (forvar2224 = (1'h0); (forvar2224 < (1'h0)); forvar2224 = (forvar2224 + (1'h1)))
                    begin
                      reg2225 <= ({((+reg2268) == $signed(reg2205))} ?
                          forvar2200 : (!reg2147[(1'h0):(1'h0)]));
                      reg2226 <= (~|(+reg2274[(3'h6):(2'h3)]));
                      reg2227 <= (8'ha0);
                    end
                end
            end
        end
      if ($unsigned((($unsigned(reg2244) <= $unsigned(reg2142)) ?
          ({forvar2228} >>> $unsigned((8'ha6))) : ((forvar2165 ?
                  reg2246 : forvar2161) ?
              forvar2179[(3'h4):(1'h1)] : (reg2209 ? reg2187 : reg2245)))))
        begin
          for (forvar2276 = (1'h0); (forvar2276 < (2'h3)); forvar2276 = (forvar2276 + (1'h1)))
            begin
              if ((reg2231 ?
                  $unsigned((reg2227[(2'h2):(1'h0)] ?
                      (^~reg2248) : (reg2193 >>> reg2133))) : $unsigned($unsigned((reg2152 ^ (8'hba))))))
                begin
                  for (forvar2277 = (1'h0); (forvar2277 < (2'h2)); forvar2277 = (forvar2277 + (1'h1)))
                    begin
                      reg2278 <= $unsigned((&{reg2247[(4'h9):(3'h6)]}));
                      reg2279 <= $unsigned(($unsigned((reg2173 | forvar2192)) && reg2214));
                    end
                end
              else
                begin
                  reg2277 <= (((~|(8'ha1)) == reg2172[(3'h6):(2'h2)]) >> reg2165);
                  reg2278 <= $signed(reg2140[(3'h7):(3'h5)]);
                  for (forvar2279 = (1'h0); (forvar2279 < (1'h0)); forvar2279 = (forvar2279 + (1'h1)))
                    begin
                      reg2280 <= (^~(({forvar2133} ^~ reg2211) ?
                          ((reg2242 && reg2165) ?
                              $unsigned(forvar2224) : reg2260) : forvar2134));
                      reg2281 <= {$unsigned($signed((forvar2213 == reg2199)))};
                      reg2282 <= ($unsigned(($unsigned(reg2269) ?
                              ((8'ha5) ?
                                  (8'hae) : (8'ha1)) : $signed(forvar2200))) ?
                          $unsigned(($signed(reg2135) && {(8'haf)})) : ((|{wire2127}) | $signed((forvar2191 > reg2204))));
                    end
                  for (forvar2283 = (1'h0); (forvar2283 < (2'h2)); forvar2283 = (forvar2283 + (1'h1)))
                    begin
                      reg2284 <= ($signed((((8'had) ? forvar2147 : reg2227) ?
                          reg2261[(2'h2):(1'h1)] : $signed((8'hb6)))) ~^ (|$signed((reg2218 && (8'ha7)))));
                    end
                end
              for (forvar2285 = (1'h0); (forvar2285 < (1'h1)); forvar2285 = (forvar2285 + (1'h1)))
                begin
                  for (forvar2286 = (1'h0); (forvar2286 < (2'h2)); forvar2286 = (forvar2286 + (1'h1)))
                    begin
                      reg2287 <= (reg2157 ?
                          ($unsigned((&reg2263)) ?
                              {(reg2181 ?
                                      reg2157 : reg2242)} : forvar2161) : $signed(reg2139[(3'h4):(2'h2)]));
                    end
                  if ((^(($unsigned(reg2264) && {forvar2156}) ?
                      ($unsigned((8'ha0)) ?
                          $unsigned(forvar2279) : {forvar2214}) : reg2176[(5'h10):(3'h6)])))
                    begin
                      reg2288 <= ((^$signed($unsigned(forvar2174))) ?
                          $unsigned($signed(reg2185)) : $signed($unsigned($unsigned((8'hb5)))));
                    end
                  else
                    begin
                      reg2288 <= $unsigned(($signed((reg2202 - (8'hac))) <= reg2150));
                      reg2289 <= $signed(((&$signed((8'ha7))) << ((reg2176 ?
                              reg2167 : forvar2277) ?
                          reg2269[(2'h3):(1'h1)] : forvar2156[(4'hc):(4'hc)])));
                      reg2290 <= $unsigned(((~|(&forvar2286)) ?
                          (+(reg2241 - reg2169)) : (-(~^(8'hb2)))));
                    end
                end
            end
          for (forvar2291 = (1'h0); (forvar2291 < (1'h0)); forvar2291 = (forvar2291 + (1'h1)))
            begin
              reg2292 <= {(~|($signed(wire2129) ^~ reg2226[(4'h9):(1'h1)]))};
              for (forvar2293 = (1'h0); (forvar2293 < (1'h1)); forvar2293 = (forvar2293 + (1'h1)))
                begin
                  for (forvar2294 = (1'h0); (forvar2294 < (2'h3)); forvar2294 = (forvar2294 + (1'h1)))
                    begin
                      reg2295 <= reg2269[(2'h3):(2'h2)];
                      reg2296 <= forvar2200[(3'h6):(3'h4)];
                    end
                  for (forvar2297 = (1'h0); (forvar2297 < (1'h1)); forvar2297 = (forvar2297 + (1'h1)))
                    begin
                      reg2298 <= ({((~|(8'ha7)) ?
                                  forvar2228 : $unsigned((8'hb5)))} ?
                          (&$unsigned($signed(forvar2170))) : reg2164);
                      reg2299 <= $unsigned((+$signed((reg2187 <<< forvar2172))));
                      reg2300 <= ((^reg2132[(3'h4):(2'h3)]) ?
                          (reg2166 ?
                              (-(~|reg2188)) : (reg2251[(2'h3):(1'h0)] ?
                                  reg2155[(4'h9):(3'h7)] : (reg2139 <<< (8'ha6)))) : reg2203[(3'h7):(1'h0)]);
                    end
                  if ($signed(({reg2152[(1'h1):(1'h1)]} ?
                      $signed({reg2133}) : ((reg2248 <= reg2223) ?
                          reg2236[(2'h3):(1'h0)] : (~|reg2251)))))
                    begin
                      reg2301 <= $signed(reg2230);
                      reg2302 <= forvar2174[(2'h3):(2'h3)];
                      reg2303 <= (reg2247[(3'h7):(1'h1)] >= (^~$signed(reg2205)));
                      reg2304 <= (forvar2165 | forvar2283);
                    end
                  else
                    begin
                      reg2301 <= reg2247[(1'h0):(1'h0)];
                    end
                end
              for (forvar2305 = (1'h0); (forvar2305 < (1'h0)); forvar2305 = (forvar2305 + (1'h1)))
                begin
                  if (reg2208[(3'h6):(1'h1)])
                    begin
                      reg2306 <= (|$signed((~&forvar2213)));
                      reg2307 <= $unsigned((8'hab));
                    end
                  else
                    begin
                      reg2306 <= reg2217[(3'h7):(1'h0)];
                      reg2307 <= forvar2305;
                      reg2308 <= $signed((((reg2225 ? forvar2228 : forvar2242) ?
                              $signed(reg2235) : (8'hac)) ?
                          ($unsigned(reg2172) ?
                              reg2138[(4'hb):(3'h4)] : (reg2269 << forvar2198)) : $unsigned(forvar2159[(4'h8):(2'h3)])));
                      reg2309 <= ((((reg2245 ? forvar2294 : reg2242) ?
                                  forvar2150[(4'h8):(2'h2)] : {reg2241}) ?
                              (^~(~^reg2194)) : (~^(8'hb1))) ?
                          {{$unsigned(forvar2172)}} : (+((reg2141 ?
                                  (8'hb4) : reg2162) ?
                              (forvar2206 - reg2308) : (forvar2192 > (8'hb6)))));
                    end
                  if (forvar2191)
                    begin
                      reg2310 <= reg2235;
                      reg2311 <= reg2148;
                    end
                  else
                    begin
                      reg2310 <= reg2225[(2'h2):(1'h1)];
                      reg2311 <= $unsigned((!$signed($unsigned(forvar2293))));
                      reg2312 <= $unsigned($signed($unsigned($signed(reg2214))));
                      reg2313 <= $unsigned(reg2133);
                    end
                end
            end
          for (forvar2314 = (1'h0); (forvar2314 < (2'h2)); forvar2314 = (forvar2314 + (1'h1)))
            begin
              if ($signed((((reg2192 ? reg2155 : reg2224) - $signed(reg2310)) ?
                  (reg2178 & wire2128) : {reg2152})))
                begin
                  reg2315 <= (forvar2228[(4'h8):(2'h2)] || ($unsigned((reg2244 ?
                      reg2277 : (8'ha5))) || (reg2196[(4'ha):(2'h3)] - $signed(forvar2206))));
                  for (forvar2316 = (1'h0); (forvar2316 < (1'h0)); forvar2316 = (forvar2316 + (1'h1)))
                    begin
                      reg2317 <= (~&(8'haa));
                      reg2318 <= $signed(($unsigned((reg2192 ^~ reg2209)) <<< reg2205));
                    end
                  for (forvar2319 = (1'h0); (forvar2319 < (2'h2)); forvar2319 = (forvar2319 + (1'h1)))
                    begin
                      reg2320 <= (8'h9d);
                      reg2321 <= reg2312[(2'h3):(1'h1)];
                      reg2322 <= ((+(&(reg2214 ?
                          reg2152 : reg2309))) <<< (reg2262 >> reg2224));
                    end
                  for (forvar2323 = (1'h0); (forvar2323 < (2'h2)); forvar2323 = (forvar2323 + (1'h1)))
                    begin
                      reg2324 <= ($unsigned((reg2250 ?
                              reg2140 : (reg2151 <= (8'had)))) ?
                          forvar2229 : $unsigned(((reg2174 ?
                                  (8'hb6) : forvar2267) ?
                              {(8'hba)} : (reg2130 ? reg2202 : forvar2212))));
                      reg2325 <= (|(reg2139[(1'h1):(1'h0)] ?
                          ((~&forvar2133) ?
                              forvar2271 : $unsigned(reg2321)) : (~((8'ha3) ?
                              forvar2141 : reg2258))));
                      reg2326 <= (reg2219[(3'h7):(2'h2)] << $unsigned((reg2288[(3'h5):(1'h1)] ?
                          (-forvar2170) : $signed(reg2222))));
                      reg2327 <= (8'hb3);
                    end
                end
              else
                begin
                  for (forvar2315 = (1'h0); (forvar2315 < (1'h1)); forvar2315 = (forvar2315 + (1'h1)))
                    begin
                      reg2316 <= reg2181;
                      reg2317 <= $unsigned(reg2155);
                    end
                  for (forvar2318 = (1'h0); (forvar2318 < (2'h3)); forvar2318 = (forvar2318 + (1'h1)))
                    begin
                      reg2319 <= $unsigned({(^((8'hb0) ?
                              forvar2162 : forvar2187))});
                      reg2320 <= {((8'haa) ~^ reg2251)};
                      reg2321 <= reg2263[(3'h4):(1'h1)];
                      reg2322 <= $signed((($signed((8'hb7)) < reg2208[(2'h2):(1'h1)]) ?
                          reg2205[(1'h0):(1'h0)] : $unsigned((~^(8'hb9)))));
                    end
                  if ({($unsigned({reg2310}) ?
                          $unsigned(reg2216) : (+(reg2136 > reg2225)))})
                    begin
                      reg2323 <= (reg2281[(2'h3):(2'h3)] | (($signed(reg2134) & $signed(reg2219)) <= (-forvar2166[(1'h0):(1'h0)])));
                      reg2324 <= (~&(forvar2286 ?
                          $unsigned((reg2157 ?
                              reg2157 : reg2227)) : forvar2224[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg2323 <= $signed(reg2264[(3'h7):(3'h6)]);
                      reg2324 <= reg2236;
                      reg2325 <= $signed(reg2279);
                    end
                end
              if (($signed($unsigned((forvar2150 ^ forvar2233))) == (reg2167[(1'h0):(1'h0)] > $signed($signed(forvar2156)))))
                begin
                  for (forvar2328 = (1'h0); (forvar2328 < (1'h1)); forvar2328 = (forvar2328 + (1'h1)))
                    begin
                      reg2329 <= reg2141[(4'ha):(2'h3)];
                    end
                end
              else
                begin
                  reg2328 <= reg2245;
                  if ((&reg2307[(4'hc):(4'hb)]))
                    begin
                      reg2329 <= reg2190[(3'h6):(1'h1)];
                      reg2330 <= ($unsigned(reg2136) ?
                          $unsigned(reg2180) : forvar2318[(3'h5):(1'h0)]);
                      reg2331 <= ({wire2125} ?
                          $signed((forvar2141[(4'ha):(3'h7)] >>> $unsigned(reg2249))) : (reg2134 << {{reg2281}}));
                    end
                  else
                    begin
                      reg2329 <= ($unsigned(forvar2165[(1'h1):(1'h1)]) >>> (~&$signed(((8'ha4) ?
                          (8'hb3) : (8'hae)))));
                      reg2330 <= ($unsigned((forvar2277[(4'hc):(3'h7)] ?
                          ((8'ha0) ?
                              reg2180 : reg2331) : $signed(reg2231))) == {$unsigned(reg2260)});
                      reg2331 <= reg2205[(3'h4):(1'h1)];
                    end
                  for (forvar2332 = (1'h0); (forvar2332 < (2'h2)); forvar2332 = (forvar2332 + (1'h1)))
                    begin
                      reg2333 <= (~&forvar2191[(3'h4):(3'h4)]);
                    end
                  reg2334 <= (reg2253 ?
                      {(^$signed(forvar2137))} : reg2331[(1'h1):(1'h1)]);
                end
              if ($unsigned((^~{(8'hb4)})))
                begin
                  for (forvar2335 = (1'h0); (forvar2335 < (1'h0)); forvar2335 = (forvar2335 + (1'h1)))
                    begin
                      reg2336 <= (forvar2228 ^ $signed($unsigned((^~reg2135))));
                    end
                end
              else
                begin
                  for (forvar2335 = (1'h0); (forvar2335 < (1'h1)); forvar2335 = (forvar2335 + (1'h1)))
                    begin
                      reg2336 <= forvar2294;
                      reg2337 <= reg2153[(2'h3):(2'h2)];
                    end
                  for (forvar2338 = (1'h0); (forvar2338 < (1'h1)); forvar2338 = (forvar2338 + (1'h1)))
                    begin
                      reg2339 <= (reg2177[(3'h6):(3'h6)] != $unsigned((8'ha2)));
                      reg2340 <= {(8'ha4)};
                    end
                  for (forvar2341 = (1'h0); (forvar2341 < (1'h1)); forvar2341 = (forvar2341 + (1'h1)))
                    begin
                      reg2342 <= $signed(reg2304);
                      reg2343 <= (~&{forvar2293[(3'h5):(2'h3)]});
                      reg2344 <= $signed({forvar2286[(4'hc):(2'h3)]});
                    end
                  reg2345 <= ((|(forvar2148[(2'h2):(1'h1)] >= (forvar2283 ?
                      forvar2297 : reg2171))) || (($signed(reg2269) ?
                          reg2316[(2'h3):(2'h2)] : reg2224[(1'h1):(1'h1)]) ?
                      (-forvar2294) : (reg2169[(1'h0):(1'h0)] ?
                          reg2308 : $signed(forvar2187))));
                end
            end
        end
      else
        begin
          if ((&$unsigned(((reg2258 && reg2251) >= {forvar2277}))))
            begin
              reg2276 <= (^reg2147);
              for (forvar2277 = (1'h0); (forvar2277 < (1'h1)); forvar2277 = (forvar2277 + (1'h1)))
                begin
                  if (reg2196)
                    begin
                      reg2278 <= $unsigned(reg2161);
                      reg2279 <= (((~$signed(reg2233)) * ((reg2140 || reg2191) ^ $unsigned(reg2265))) ?
                          $signed(((reg2236 ? forvar2213 : reg2176) ?
                              reg2188[(1'h1):(1'h0)] : (reg2203 ?
                                  reg2136 : reg2261))) : reg2135[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg2278 <= (~^(($unsigned(reg2241) ?
                              {reg2327} : (reg2159 < reg2168)) ?
                          reg2301[(3'h5):(2'h3)] : (~&$unsigned(forvar2286))));
                      reg2279 <= (reg2340[(1'h0):(1'h0)] ?
                          ((^forvar2150[(3'h6):(3'h4)]) && reg2251[(4'h9):(1'h1)]) : reg2233[(4'hd):(3'h5)]);
                    end
                  for (forvar2280 = (1'h0); (forvar2280 < (1'h1)); forvar2280 = (forvar2280 + (1'h1)))
                    begin
                      reg2281 <= forvar2172[(4'hd):(3'h7)];
                      reg2282 <= reg2168;
                    end
                end
              if ((((reg2253[(3'h6):(2'h3)] ?
                  (-(8'ha0)) : {reg2175}) >> forvar2279) >= reg2340[(3'h4):(2'h2)]))
                begin
                  for (forvar2283 = (1'h0); (forvar2283 < (2'h3)); forvar2283 = (forvar2283 + (1'h1)))
                    begin
                      reg2284 <= ($signed((-(forvar2286 | forvar2280))) ?
                          ($signed(reg2224[(1'h1):(1'h0)]) ?
                              $signed(wire2124) : (reg2278[(3'h4):(3'h4)] + (-reg2220))) : ($unsigned(forvar2133) ^~ reg2219[(3'h7):(3'h6)]));
                      reg2285 <= reg2312[(1'h0):(1'h0)];
                    end
                  if ((8'ha9))
                    begin
                      reg2286 <= $unsigned({(reg2258[(2'h2):(2'h2)] == $signed(forvar2341))});
                      reg2287 <= (forvar2161[(1'h0):(1'h0)] | ({(reg2334 ?
                              forvar2193 : reg2344)} == (~|reg2192)));
                    end
                  else
                    begin
                      reg2286 <= {{($signed((8'ha6)) ?
                                  $signed((8'hb0)) : (forvar2157 ?
                                      reg2171 : reg2304))}};
                    end
                  if ($unsigned($signed({{reg2307}})))
                    begin
                      reg2288 <= ((^$signed(reg2152)) < (+reg2281[(3'h7):(2'h3)]));
                    end
                  else
                    begin
                      reg2288 <= {(+(((8'h9d) && reg2261) ?
                              (forvar2141 ^~ reg2313) : $unsigned(reg2161)))};
                    end
                  if (forvar2319)
                    begin
                      reg2289 <= {(8'hb4)};
                      reg2290 <= reg2218;
                      reg2291 <= ($unsigned($unsigned((reg2318 ?
                              reg2149 : forvar2201))) ?
                          reg2189 : (((&forvar2335) ?
                              {wire2125} : reg2202) >= ((forvar2328 ^~ reg2263) ?
                              forvar2213 : (~forvar2162))));
                    end
                  else
                    begin
                      reg2289 <= (+$unsigned($unsigned(forvar2135)));
                    end
                end
              else
                begin
                  for (forvar2283 = (1'h0); (forvar2283 < (2'h2)); forvar2283 = (forvar2283 + (1'h1)))
                    begin
                      reg2284 <= (8'ha9);
                    end
                  for (forvar2285 = (1'h0); (forvar2285 < (1'h1)); forvar2285 = (forvar2285 + (1'h1)))
                    begin
                      reg2286 <= (reg2302 == ({(forvar2132 ~^ reg2219)} ?
                          $unsigned(forvar2141) : (reg2220[(3'h5):(3'h4)] >>> (8'hb9))));
                      reg2287 <= (((~&reg2269) ?
                          (^(reg2323 ?
                              reg2193 : reg2248)) : reg2233[(3'h6):(2'h3)]) + $signed(((reg2266 ?
                          reg2141 : (8'haf)) + $signed((8'hb8)))));
                    end
                  if (reg2276)
                    begin
                      reg2288 <= ($unsigned($signed($unsigned(reg2173))) | (((~&forvar2165) ?
                          forvar2328[(1'h0):(1'h0)] : reg2264[(3'h5):(1'h1)]) & $signed((reg2159 * reg2317))));
                      reg2289 <= ((!{forvar2166}) ?
                          reg2178 : reg2323[(2'h2):(2'h2)]);
                      reg2290 <= forvar2159[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg2288 <= $unsigned((($unsigned(reg2321) & (reg2149 || reg2173)) & (~$signed(reg2261))));
                      reg2289 <= reg2239[(3'h6):(3'h6)];
                      reg2290 <= $signed(reg2331);
                      reg2291 <= (&(~|$signed(forvar2291)));
                    end
                  reg2292 <= ((8'ha9) ?
                      ((forvar2139 ?
                          reg2227[(2'h3):(1'h1)] : $signed(forvar2256)) > ((reg2236 || (8'hb6)) ?
                          $signed(forvar2232) : {reg2164})) : (~&(reg2280 < reg2306[(2'h2):(1'h0)])));
                end
              for (forvar2293 = (1'h0); (forvar2293 < (1'h0)); forvar2293 = (forvar2293 + (1'h1)))
                begin
                  if (forvar2318[(1'h1):(1'h1)])
                    begin
                      reg2294 <= {$unsigned($unsigned(reg2303))};
                    end
                  else
                    begin
                      reg2294 <= (reg2184 <<< $signed({(reg2260 & (8'hb5))}));
                      reg2295 <= reg2180;
                    end
                  if (((8'ha5) - forvar2175))
                    begin
                      reg2296 <= $unsigned((~^$unsigned($unsigned(reg2282))));
                    end
                  else
                    begin
                      reg2296 <= $unsigned((((+reg2254) ?
                          forvar2283 : forvar2156) <<< reg2167[(2'h2):(1'h1)]));
                      reg2297 <= (8'ha7);
                      reg2298 <= $unsigned(reg2272);
                    end
                end
            end
          else
            begin
              if ((reg2317[(2'h2):(1'h1)] <= $unsigned((8'ha7))))
                begin
                  if ($signed(forvar2294))
                    begin
                      reg2276 <= $unsigned(reg2237[(3'h7):(3'h5)]);
                      reg2277 <= reg2164[(1'h0):(1'h0)];
                      reg2278 <= (($signed(reg2154[(3'h4):(1'h0)]) && reg2302) + $signed(reg2195));
                    end
                  else
                    begin
                      reg2276 <= (reg2232[(1'h1):(1'h0)] - (+(~|(8'ha5))));
                      reg2277 <= $unsigned((!{$unsigned(forvar2224)}));
                      reg2278 <= (!reg2272);
                      reg2279 <= reg2306;
                    end
                  for (forvar2280 = (1'h0); (forvar2280 < (2'h3)); forvar2280 = (forvar2280 + (1'h1)))
                    begin
                      reg2281 <= (forvar2335[(4'hb):(4'ha)] + (^reg2209));
                    end
                end
              else
                begin
                  for (forvar2276 = (1'h0); (forvar2276 < (2'h3)); forvar2276 = (forvar2276 + (1'h1)))
                    begin
                      reg2277 <= reg2238[(3'h4):(1'h0)];
                    end
                  if (reg2248)
                    begin
                      reg2278 <= {reg2345};
                    end
                  else
                    begin
                      reg2278 <= ({{$signed(forvar2283)}} ?
                          $unsigned(((reg2142 ~^ (8'ha8)) < (reg2130 ?
                              reg2138 : forvar2155))) : ($unsigned(reg2140[(4'he):(1'h0)]) ?
                              (8'haa) : $unsigned({reg2342})));
                      reg2279 <= (8'h9e);
                      reg2280 <= $unsigned($signed(((reg2214 ^~ (8'hac)) ?
                          reg2248 : (forvar2135 ? (8'hba) : reg2193))));
                    end
                  if ({(8'ha1)})
                    begin
                      reg2281 <= (^~(!({reg2307} ?
                          reg2170[(1'h1):(1'h0)] : forvar2161[(2'h2):(1'h0)])));
                      reg2282 <= $signed({$unsigned(reg2285)});
                      reg2283 <= (&$signed(((reg2196 && forvar2257) * reg2255[(3'h6):(3'h6)])));
                      reg2284 <= ((&($signed(forvar2332) & (+reg2342))) ^~ $signed($signed((reg2273 >> reg2156))));
                    end
                  else
                    begin
                      reg2281 <= reg2287[(2'h3):(1'h1)];
                      reg2282 <= (((((8'had) * reg2244) < {reg2180}) ?
                              ((^~reg2299) ?
                                  reg2151 : (reg2302 >= (8'ha7))) : $unsigned((reg2189 ?
                                  reg2218 : reg2202))) ?
                          $unsigned($signed(reg2191)) : reg2216[(2'h3):(1'h1)]);
                      reg2283 <= $signed(((((8'hb9) <<< reg2218) ^ $signed(reg2203)) >>> (^~forvar2213[(2'h3):(2'h2)])));
                      reg2284 <= ((reg2255 ?
                              ($signed(forvar2294) ?
                                  (reg2260 ^~ reg2151) : reg2167[(3'h4):(1'h0)]) : $signed(forvar2141[(4'ha):(3'h6)])) ?
                          reg2306 : ($signed(reg2230) ?
                              $unsigned(reg2197[(4'hc):(2'h3)]) : reg2310));
                    end
                end
            end
          for (forvar2299 = (1'h0); (forvar2299 < (1'h0)); forvar2299 = (forvar2299 + (1'h1)))
            begin
              if (forvar2141)
                begin
                  if ({$signed(((reg2191 ?
                          reg2290 : reg2171) + $unsigned(reg2286)))})
                    begin
                      reg2300 <= (($unsigned(reg2302) ?
                              ((&forvar2172) ?
                                  reg2242[(1'h0):(1'h0)] : $unsigned(forvar2227)) : $signed($unsigned(reg2281))) ?
                          ($signed($signed(reg2237)) ?
                              forvar2279[(2'h3):(2'h2)] : (!$unsigned(forvar2155))) : $unsigned(reg2161));
                      reg2301 <= ($signed(reg2311) <= (-reg2234));
                      reg2302 <= (({(reg2274 ?
                                  reg2171 : reg2163)} - $unsigned(reg2268)) ?
                          reg2164 : reg2284[(2'h2):(1'h0)]);
                      reg2303 <= forvar2279;
                    end
                  else
                    begin
                      reg2300 <= $unsigned($signed($signed(reg2137)));
                      reg2301 <= {(reg2163[(4'ha):(4'h9)] ?
                              $unsigned(forvar2243[(2'h2):(1'h0)]) : $signed((!reg2140)))};
                    end
                  for (forvar2304 = (1'h0); (forvar2304 < (2'h3)); forvar2304 = (forvar2304 + (1'h1)))
                    begin
                      reg2305 <= (^reg2202);
                      reg2306 <= $signed(forvar2335);
                      reg2307 <= ($signed((8'ha0)) * $signed(reg2238[(3'h6):(2'h2)]));
                    end
                  reg2308 <= {reg2325};
                  if ((~&(((reg2193 | forvar2162) ?
                      reg2298[(4'h8):(4'h8)] : (reg2251 ^ reg2223)) ^~ reg2248[(1'h0):(1'h0)])))
                    begin
                      reg2309 <= reg2304;
                      reg2310 <= reg2266[(1'h0):(1'h0)];
                      reg2311 <= reg2207;
                      reg2312 <= $signed($signed(($signed((8'h9c)) ?
                          $signed((8'ha9)) : $signed(forvar2318))));
                    end
                  else
                    begin
                      reg2309 <= ($unsigned($signed($signed(forvar2135))) ?
                          (($unsigned(forvar2277) ?
                                  (forvar2213 - reg2316) : $unsigned(reg2295)) ?
                              reg2210[(2'h3):(2'h2)] : forvar2155) : $unsigned((forvar2229 ?
                              (reg2282 ?
                                  reg2169 : forvar2175) : (+forvar2161))));
                      reg2310 <= reg2262;
                    end
                end
              else
                begin
                  for (forvar2300 = (1'h0); (forvar2300 < (1'h1)); forvar2300 = (forvar2300 + (1'h1)))
                    begin
                      reg2301 <= $unsigned(forvar2191);
                      reg2302 <= ((forvar2193 ?
                          reg2292[(2'h2):(2'h2)] : reg2250) ^ forvar2316);
                      reg2303 <= $unsigned($unsigned($signed({(8'hb3)})));
                      reg2304 <= {(reg2169 >> forvar2291)};
                    end
                  reg2305 <= reg2225;
                  if (((~^$unsigned((reg2175 ? reg2232 : reg2163))) ?
                      (((forvar2157 ? reg2260 : (8'ha3)) && reg2279) ?
                          (forvar2229 ?
                              $signed(reg2313) : forvar2243) : forvar2304[(2'h3):(2'h3)]) : reg2327[(3'h4):(2'h3)]))
                    begin
                      reg2306 <= $unsigned((forvar2150 < forvar2157));
                      reg2307 <= (($unsigned($signed(reg2155)) - (~(^~reg2322))) ?
                          reg2238 : forvar2341);
                    end
                  else
                    begin
                      reg2306 <= (reg2158 + (-forvar2267[(4'hd):(4'ha)]));
                      reg2307 <= forvar2200;
                      reg2308 <= ((reg2247[(1'h0):(1'h0)] + reg2161) ?
                          (8'hb6) : reg2236);
                      reg2309 <= $signed((&(reg2282[(4'h8):(4'h8)] | $signed(reg2282))));
                    end
                end
              for (forvar2313 = (1'h0); (forvar2313 < (1'h1)); forvar2313 = (forvar2313 + (1'h1)))
                begin
                  for (forvar2314 = (1'h0); (forvar2314 < (1'h1)); forvar2314 = (forvar2314 + (1'h1)))
                    begin
                      reg2315 <= (({reg2316} ?
                          (^(forvar2214 ? reg2296 : (8'ha2))) : ((~reg2180) ?
                              $unsigned(reg2207) : reg2188)) ^~ reg2334);
                      reg2316 <= forvar2243[(3'h4):(1'h1)];
                      reg2317 <= reg2136[(4'ha):(3'h5)];
                    end
                  if (($unsigned({reg2166[(1'h1):(1'h0)]}) ?
                      (^$signed(forvar2299[(3'h4):(2'h3)])) : $unsigned(reg2131)))
                    begin
                      reg2318 <= $unsigned((~^(8'hb0)));
                      reg2319 <= (+{(reg2339[(1'h1):(1'h0)] ?
                              forvar2212 : (-reg2145))});
                    end
                  else
                    begin
                      reg2318 <= reg2278[(2'h3):(2'h3)];
                    end
                  if ((8'haa))
                    begin
                      reg2320 <= (reg2162 > (((~|reg2325) && $unsigned(reg2225)) ?
                          (~|(reg2249 <= reg2211)) : (~&reg2334[(2'h2):(1'h1)])));
                      reg2321 <= reg2296[(4'h8):(1'h0)];
                      reg2322 <= $signed($unsigned((8'h9e)));
                    end
                  else
                    begin
                      reg2320 <= $signed(reg2218);
                      reg2321 <= ($unsigned((~^(wire2124 >>> reg2273))) ?
                          reg2139 : $signed($unsigned({reg2226})));
                      reg2322 <= {(~^(reg2145 == $signed(reg2217)))};
                    end
                end
              for (forvar2323 = (1'h0); (forvar2323 < (2'h3)); forvar2323 = (forvar2323 + (1'h1)))
                begin
                  if (($signed($signed(reg2230)) * (^~$unsigned((reg2185 << reg2274)))))
                    begin
                      reg2324 <= (+((&$signed(reg2144)) && {(reg2155 ^~ reg2327)}));
                      reg2325 <= (({(|(8'h9f))} >= ($signed(forvar2335) >>> reg2334[(4'ha):(4'ha)])) ?
                          reg2204[(2'h3):(1'h0)] : (^((reg2161 ^~ reg2182) | {reg2247})));
                      reg2326 <= {reg2284};
                      reg2327 <= $unsigned($signed((^~(!reg2318))));
                    end
                  else
                    begin
                      reg2324 <= forvar2271[(3'h4):(3'h4)];
                    end
                end
            end
          for (forvar2328 = (1'h0); (forvar2328 < (2'h3)); forvar2328 = (forvar2328 + (1'h1)))
            begin
              for (forvar2329 = (1'h0); (forvar2329 < (2'h3)); forvar2329 = (forvar2329 + (1'h1)))
                begin
                  if ($signed((reg2291[(3'h6):(1'h1)] ?
                      reg2142[(2'h2):(2'h2)] : ((reg2210 ?
                          forvar2193 : (8'had)) * reg2182[(3'h4):(1'h0)]))))
                    begin
                      reg2330 <= (((reg2159 ?
                                  $unsigned(forvar2201) : (reg2282 | reg2271)) ?
                              (forvar2314 * forvar2213) : reg2229[(2'h2):(2'h2)]) ?
                          ($unsigned({reg2274}) ?
                              {((8'haa) * reg2210)} : reg2297[(4'hc):(3'h5)]) : (reg2162 <<< reg2172));
                      reg2331 <= (~|forvar2323[(3'h6):(1'h1)]);
                      reg2332 <= {{$signed((reg2146 | reg2248))}};
                      reg2333 <= $signed(reg2250[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg2330 <= reg2147;
                    end
                  reg2334 <= reg2249;
                  reg2335 <= (!{{(reg2184 > (8'hb7))}});
                  reg2336 <= $signed((^$signed($signed(reg2248))));
                end
            end
        end
    end
  assign wire2346 = $signed(((8'hae) < (~(8'ha3))));
  assign wire2347 = forvar2198;
  always
    @(posedge clk) begin
      for (forvar2348 = (1'h0); (forvar2348 < (2'h2)); forvar2348 = (forvar2348 + (1'h1)))
        begin
          if ({reg2228})
            begin
              reg2349 <= (($signed($signed(forvar2206)) ~^ {reg2345[(3'h5):(1'h0)]}) < reg2147);
              if (forvar2191)
                begin
                  for (forvar2350 = (1'h0); (forvar2350 < (1'h0)); forvar2350 = (forvar2350 + (1'h1)))
                    begin
                      reg2351 <= reg2283;
                      reg2352 <= reg2276[(3'h7):(3'h7)];
                      reg2353 <= forvar2319;
                    end
                  reg2354 <= ((reg2310 >>> reg2326) ~^ (reg2178[(4'hf):(4'h8)] & ((forvar2144 < reg2339) <<< forvar2285)));
                  if (reg2345)
                    begin
                      reg2355 <= (8'ha4);
                      reg2356 <= ((forvar2323 ?
                              ((~^forvar2206) <<< (reg2263 ?
                                  reg2272 : wire2123)) : forvar2213[(2'h2):(2'h2)]) ?
                          $signed({forvar2280}) : {$unsigned(forvar2329[(1'h0):(1'h0)])});
                      reg2357 <= (reg2171 ?
                          ($unsigned(forvar2227[(3'h4):(2'h2)]) & ($unsigned(forvar2293) && (forvar2170 >= forvar2305))) : ($signed($signed(forvar2150)) ?
                              (+reg2237) : (8'hac)));
                    end
                  else
                    begin
                      reg2355 <= forvar2224;
                      reg2356 <= (reg2130[(3'h7):(2'h3)] ?
                          {$unsigned((-(8'hac)))} : $unsigned($unsigned((8'h9d))));
                      reg2357 <= $unsigned(reg2182[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  reg2350 <= ($signed($signed((reg2131 ?
                      reg2220 : reg2304))) ~^ $signed({$signed(reg2274)}));
                  reg2351 <= ((forvar2285[(1'h0):(1'h0)] <<< ({reg2215} ?
                      (-reg2336) : forvar2187)) > forvar2173[(3'h5):(2'h3)]);
                  reg2352 <= ($signed((reg2144 || forvar2315)) <<< ($unsigned(reg2303[(4'ha):(4'h8)]) * ((reg2269 ?
                          reg2301 : forvar2299) ?
                      forvar2299 : {reg2197})));
                  for (forvar2353 = (1'h0); (forvar2353 < (2'h3)); forvar2353 = (forvar2353 + (1'h1)))
                    begin
                      reg2354 <= $signed(reg2210);
                      reg2355 <= ((((!reg2323) ?
                              reg2159 : {reg2182}) ^~ (~^$signed(reg2262))) ?
                          (~((~&forvar2173) ?
                              $unsigned(forvar2232) : (!reg2236))) : $unsigned($signed(reg2237)));
                    end
                end
              if ((^~(^~(reg2263[(3'h6):(2'h2)] ? forvar2323 : {reg2303}))))
                begin
                  if ((((~(reg2335 - (8'ha3))) > (((8'ha0) && forvar2200) ?
                          (~|reg2274) : (reg2255 >>> reg2299))) ?
                      (-(+(^forvar2243))) : (forvar2291[(2'h2):(1'h0)] ?
                          $signed(reg2189) : reg2161[(1'h1):(1'h1)])))
                    begin
                      reg2358 <= reg2211[(4'ha):(1'h0)];
                      reg2359 <= ((~&{(!forvar2155)}) + {(8'h9c)});
                      reg2360 <= forvar2341[(3'h7):(3'h7)];
                      reg2361 <= reg2325[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg2358 <= $unsigned({($unsigned(reg2215) ?
                              $signed(forvar2242) : reg2154[(3'h4):(2'h2)])});
                      reg2359 <= reg2196;
                      reg2360 <= $signed(reg2226);
                      reg2361 <= reg2169[(1'h1):(1'h1)];
                    end
                  if (($unsigned($signed((reg2316 ? forvar2156 : forvar2214))) ?
                      $unsigned(({reg2340} > (!reg2325))) : reg2254))
                    begin
                      reg2362 <= ({($unsigned((8'ha5)) & ((8'haa) >>> reg2216))} || forvar2304);
                      reg2363 <= reg2233;
                    end
                  else
                    begin
                      reg2362 <= reg2162;
                      reg2363 <= ((+(8'hb8)) || forvar2141);
                      reg2364 <= $unsigned(reg2310[(2'h3):(2'h3)]);
                      reg2365 <= ((~(reg2265 == (reg2330 ?
                          (8'hb6) : reg2248))) | reg2186);
                    end
                  reg2366 <= (reg2243 <= $signed($signed($unsigned((8'hab)))));
                  for (forvar2367 = (1'h0); (forvar2367 < (1'h1)); forvar2367 = (forvar2367 + (1'h1)))
                    begin
                      reg2368 <= $signed((($unsigned(reg2151) ?
                          reg2197 : ((8'ha3) ?
                              reg2180 : reg2205)) && (+{reg2344})));
                      reg2369 <= ($unsigned(reg2294) << {$unsigned($unsigned(reg2194))});
                    end
                end
              else
                begin
                  for (forvar2358 = (1'h0); (forvar2358 < (2'h3)); forvar2358 = (forvar2358 + (1'h1)))
                    begin
                      reg2359 <= ($unsigned($unsigned($unsigned(reg2268))) ?
                          $signed(((reg2333 ?
                              reg2249 : reg2231) > (|reg2361))) : (~(reg2302[(3'h6):(1'h1)] & $unsigned(reg2187))));
                      reg2360 <= reg2155;
                      reg2361 <= $unsigned((~wire2128[(4'h8):(2'h2)]));
                      reg2362 <= $signed($signed(reg2276[(3'h6):(2'h3)]));
                    end
                end
            end
          else
            begin
              for (forvar2349 = (1'h0); (forvar2349 < (2'h3)); forvar2349 = (forvar2349 + (1'h1)))
                begin
                  reg2350 <= (&((forvar2338 & reg2345) ^ ((reg2336 ?
                          reg2209 : wire2347) ?
                      forvar2198 : $signed(wire2125))));
                  if ($unsigned({(8'h9f)}))
                    begin
                      reg2351 <= wire2123[(1'h0):(1'h0)];
                      reg2352 <= {(reg2182 ?
                              reg2207[(2'h3):(2'h3)] : $signed(reg2211[(4'h8):(3'h6)]))};
                      reg2353 <= $signed((reg2194[(4'hc):(1'h0)] && reg2209));
                      reg2354 <= $signed(reg2320);
                    end
                  else
                    begin
                      reg2351 <= ({((!reg2300) * (reg2266 ?
                              (8'haa) : reg2300))} <<< {reg2277});
                      reg2352 <= $signed({$signed($signed((8'hba)))});
                    end
                end
              for (forvar2355 = (1'h0); (forvar2355 < (2'h2)); forvar2355 = (forvar2355 + (1'h1)))
                begin
                  for (forvar2356 = (1'h0); (forvar2356 < (1'h0)); forvar2356 = (forvar2356 + (1'h1)))
                    begin
                      reg2357 <= $signed(forvar2243);
                    end
                end
            end
        end
      reg2370 <= (!forvar2166);
    end
  assign wire2371 = $signed({forvar2271});
  always
    @(posedge clk) begin
      for (forvar2372 = (1'h0); (forvar2372 < (2'h2)); forvar2372 = (forvar2372 + (1'h1)))
        begin
          if ($unsigned($signed(reg2354[(3'h7):(2'h3)])))
            begin
              for (forvar2373 = (1'h0); (forvar2373 < (2'h2)); forvar2373 = (forvar2373 + (1'h1)))
                begin
                  for (forvar2374 = (1'h0); (forvar2374 < (2'h2)); forvar2374 = (forvar2374 + (1'h1)))
                    begin
                      reg2375 <= $signed((~$signed((reg2147 ?
                          reg2184 : reg2134))));
                    end
                end
              for (forvar2376 = (1'h0); (forvar2376 < (1'h0)); forvar2376 = (forvar2376 + (1'h1)))
                begin
                  for (forvar2377 = (1'h0); (forvar2377 < (2'h3)); forvar2377 = (forvar2377 + (1'h1)))
                    begin
                      reg2378 <= $unsigned($unsigned(((reg2303 ^ reg2322) ?
                          forvar2374 : {reg2187})));
                      reg2379 <= forvar2192;
                      reg2380 <= $signed(reg2229);
                    end
                  if (reg2356)
                    begin
                      reg2381 <= $signed($signed(((reg2252 ?
                          reg2180 : reg2245) ^~ reg2262[(1'h1):(1'h0)])));
                      reg2382 <= {(~{((8'ha4) <= reg2203)})};
                      reg2383 <= {(!(+$signed(forvar2156)))};
                    end
                  else
                    begin
                      reg2381 <= ($unsigned(($unsigned(reg2259) << (forvar2141 <<< forvar2219))) >>> (~^$unsigned((forvar2137 ?
                          forvar2256 : reg2163))));
                      reg2382 <= reg2164;
                    end
                  if (forvar2227)
                    begin
                      reg2384 <= reg2143[(3'h6):(2'h2)];
                      reg2385 <= ((((wire2346 <= (8'h9f)) ?
                              reg2137[(4'h8):(3'h6)] : {reg2180}) ?
                          (reg2148 ?
                              {reg2180} : reg2266[(1'h0):(1'h0)]) : wire2347) >>> $signed($unsigned({reg2148})));
                    end
                  else
                    begin
                      reg2384 <= (^forvar2155[(2'h3):(2'h3)]);
                      reg2385 <= (forvar2286 ? $unsigned(reg2281) : reg2142);
                      reg2386 <= reg2152[(1'h0):(1'h0)];
                    end
                end
              if ((reg2326[(4'h8):(2'h3)] <= (~^(~(reg2230 ?
                  forvar2165 : reg2150)))))
                begin
                  reg2387 <= (^(8'hab));
                  for (forvar2388 = (1'h0); (forvar2388 < (2'h2)); forvar2388 = (forvar2388 + (1'h1)))
                    begin
                      reg2389 <= $signed((((reg2236 ^ forvar2315) ?
                          {forvar2271} : (^reg2161)) - $unsigned($unsigned((8'ha3)))));
                    end
                  reg2390 <= (8'hb9);
                end
              else
                begin
                  reg2387 <= $unsigned($signed((-{forvar2191})));
                  for (forvar2388 = (1'h0); (forvar2388 < (2'h2)); forvar2388 = (forvar2388 + (1'h1)))
                    begin
                      reg2389 <= (^forvar2179[(1'h1):(1'h1)]);
                    end
                end
              reg2391 <= reg2146;
            end
          else
            begin
              for (forvar2373 = (1'h0); (forvar2373 < (1'h1)); forvar2373 = (forvar2373 + (1'h1)))
                begin
                  reg2374 <= (reg2233[(4'he):(4'h8)] != ((~&reg2133) >> $unsigned($unsigned(reg2234))));
                  for (forvar2375 = (1'h0); (forvar2375 < (1'h1)); forvar2375 = (forvar2375 + (1'h1)))
                    begin
                      reg2376 <= reg2246;
                      reg2377 <= reg2223;
                      reg2378 <= reg2243;
                      reg2379 <= (+reg2349);
                    end
                end
              for (forvar2380 = (1'h0); (forvar2380 < (2'h3)); forvar2380 = (forvar2380 + (1'h1)))
                begin
                  for (forvar2381 = (1'h0); (forvar2381 < (2'h3)); forvar2381 = (forvar2381 + (1'h1)))
                    begin
                      reg2382 <= $signed((&{$unsigned(reg2166)}));
                      reg2383 <= ((|$unsigned(reg2180)) > (~^(|reg2232)));
                      reg2384 <= ($signed(($unsigned((8'h9e)) > $unsigned(reg2357))) * forvar2243);
                      reg2385 <= ((reg2167 ?
                          $unsigned((forvar2276 >>> forvar2323)) : $unsigned(forvar2201[(2'h2):(2'h2)])) + reg2250[(4'ha):(3'h6)]);
                    end
                  for (forvar2386 = (1'h0); (forvar2386 < (2'h2)); forvar2386 = (forvar2386 + (1'h1)))
                    begin
                      reg2387 <= reg2315;
                      reg2388 <= (reg2320 ?
                          forvar2161[(1'h1):(1'h0)] : (($unsigned(reg2327) ^ reg2337[(1'h0):(1'h0)]) >>> $signed(reg2298)));
                    end
                  for (forvar2389 = (1'h0); (forvar2389 < (1'h0)); forvar2389 = (forvar2389 + (1'h1)))
                    begin
                      reg2390 <= reg2237[(3'h5):(2'h3)];
                      reg2391 <= $unsigned($signed({reg2187[(2'h2):(1'h0)]}));
                      reg2392 <= $signed(($unsigned($unsigned(wire2346)) > reg2272));
                    end
                  if ((^~$unsigned($signed(reg2278))))
                    begin
                      reg2393 <= (&({$unsigned(reg2230)} || reg2248[(2'h3):(2'h3)]));
                      reg2394 <= ((reg2269[(3'h5):(2'h2)] ^~ {(forvar2367 ?
                              forvar2280 : reg2217)}) && ((forvar2285[(1'h1):(1'h0)] & (forvar2376 || reg2330)) >> reg2150[(4'h8):(2'h3)]));
                    end
                  else
                    begin
                      reg2393 <= {$unsigned((reg2229[(4'he):(4'ha)] + (8'ha4)))};
                    end
                end
              for (forvar2395 = (1'h0); (forvar2395 < (1'h0)); forvar2395 = (forvar2395 + (1'h1)))
                begin
                  if ($unsigned((forvar2174[(4'hd):(3'h7)] ?
                      reg2130 : $signed({(8'h9f)}))))
                    begin
                      reg2396 <= reg2307;
                      reg2397 <= {$signed((-(reg2207 ? reg2165 : reg2326)))};
                      reg2398 <= (~&($unsigned(reg2144) ^ $unsigned(reg2339[(3'h5):(3'h5)])));
                    end
                  else
                    begin
                      reg2396 <= (({$unsigned(forvar2173)} ?
                              ($signed(reg2291) ?
                                  (wire2127 ^ forvar2377) : wire2125[(3'h4):(2'h3)]) : ((reg2380 ~^ reg2207) * (forvar2201 ?
                                  reg2299 : reg2397))) ?
                          reg2355[(1'h0):(1'h0)] : $unsigned(reg2301[(2'h3):(2'h2)]));
                    end
                  for (forvar2399 = (1'h0); (forvar2399 < (1'h0)); forvar2399 = (forvar2399 + (1'h1)))
                    begin
                      reg2400 <= $unsigned($unsigned(({(8'hba)} ?
                          (^(8'hba)) : $unsigned(reg2290))));
                      reg2401 <= (8'hb2);
                      reg2402 <= (+reg2370);
                      reg2403 <= $unsigned(reg2171);
                    end
                  if ($unsigned((+$unsigned((forvar2380 ? (8'hb1) : reg2192)))))
                    begin
                      reg2404 <= forvar2372;
                      reg2405 <= reg2239[(4'hb):(4'ha)];
                      reg2406 <= (~^($unsigned($unsigned(reg2244)) & (&reg2174[(4'hf):(4'hd)])));
                    end
                  else
                    begin
                      reg2404 <= (+reg2216);
                      reg2405 <= $signed(reg2204);
                      reg2406 <= $signed((forvar2228[(3'h7):(1'h1)] != $signed($unsigned(forvar2313))));
                      reg2407 <= ((|((&reg2224) ?
                              (wire2124 ?
                                  forvar2381 : forvar2191) : (forvar2155 ?
                                  forvar2233 : forvar2341))) ?
                          $signed(reg2369) : $unsigned(({forvar2314} >> $signed((8'h9e)))));
                    end
                end
              for (forvar2408 = (1'h0); (forvar2408 < (1'h0)); forvar2408 = (forvar2408 + (1'h1)))
                begin
                  if ((~|$unsigned((~^reg2211[(1'h1):(1'h0)]))))
                    begin
                      reg2409 <= $unsigned((forvar2380 >= ($signed(reg2291) || reg2269[(3'h5):(2'h2)])));
                      reg2410 <= (reg2214 ?
                          reg2388 : ((~(reg2243 ?
                              wire2129 : reg2142)) && (forvar2286[(4'hc):(4'ha)] ?
                              {reg2332} : reg2315)));
                      reg2411 <= reg2393;
                      reg2412 <= $unsigned(($unsigned((reg2196 <<< reg2254)) ?
                          ((~^(8'hac)) ?
                              (!reg2156) : {reg2239}) : $unsigned(forvar2212)));
                    end
                  else
                    begin
                      reg2409 <= reg2284[(1'h1):(1'h0)];
                    end
                  reg2413 <= reg2149;
                  if ({{(~forvar2200[(1'h0):(1'h0)])}})
                    begin
                      reg2414 <= reg2236;
                      reg2415 <= $signed(({forvar2305} ?
                          (reg2316 || $unsigned((8'hb0))) : {$unsigned(reg2141)}));
                      reg2416 <= {reg2226[(3'h5):(2'h2)]};
                      reg2417 <= ($unsigned(((forvar2172 * reg2192) ?
                          (reg2154 ? reg2248 : reg2265) : (reg2415 ?
                              forvar2353 : reg2315))) >>> wire2371[(4'h9):(3'h7)]);
                    end
                  else
                    begin
                      reg2414 <= {reg2331[(1'h1):(1'h1)]};
                    end
                  reg2418 <= ($signed((!(forvar2150 << reg2252))) | reg2402);
                end
            end
          for (forvar2419 = (1'h0); (forvar2419 < (1'h1)); forvar2419 = (forvar2419 + (1'h1)))
            begin
              for (forvar2420 = (1'h0); (forvar2420 < (1'h1)); forvar2420 = (forvar2420 + (1'h1)))
                begin
                  for (forvar2421 = (1'h0); (forvar2421 < (1'h0)); forvar2421 = (forvar2421 + (1'h1)))
                    begin
                      reg2422 <= $signed(((^(!forvar2376)) * {$unsigned((8'hb8))}));
                      reg2423 <= {(^~forvar2201)};
                      reg2424 <= $signed(reg2400[(3'h4):(3'h4)]);
                    end
                  for (forvar2425 = (1'h0); (forvar2425 < (1'h0)); forvar2425 = (forvar2425 + (1'h1)))
                    begin
                      reg2426 <= reg2354[(3'h4):(2'h2)];
                      reg2427 <= (~forvar2332);
                    end
                end
              for (forvar2428 = (1'h0); (forvar2428 < (1'h0)); forvar2428 = (forvar2428 + (1'h1)))
                begin
                  for (forvar2429 = (1'h0); (forvar2429 < (1'h0)); forvar2429 = (forvar2429 + (1'h1)))
                    begin
                      reg2430 <= $signed($unsigned((forvar2165 > $unsigned(reg2306))));
                      reg2431 <= forvar2159[(3'h6):(1'h0)];
                      reg2432 <= ({$signed(reg2180)} >>> $unsigned(($signed(reg2426) >> reg2202[(3'h6):(2'h3)])));
                    end
                  for (forvar2433 = (1'h0); (forvar2433 < (1'h0)); forvar2433 = (forvar2433 + (1'h1)))
                    begin
                      reg2434 <= {(forvar2433[(2'h2):(1'h0)] << $signed($signed(reg2163)))};
                      reg2435 <= (($signed((reg2196 != reg2174)) ?
                          (forvar2349[(2'h2):(1'h1)] ?
                              ((8'ha4) ?
                                  forvar2156 : (8'h9e)) : (reg2140 == forvar2219)) : reg2323) < $unsigned((|$signed((8'hb8)))));
                      reg2436 <= forvar2358[(2'h3):(2'h3)];
                      reg2437 <= reg2147[(1'h0):(1'h0)];
                    end
                  if ((reg2436[(2'h3):(2'h2)] == ($unsigned(reg2390[(3'h4):(1'h0)]) + reg2330[(1'h0):(1'h0)])))
                    begin
                      reg2438 <= reg2223[(3'h4):(2'h2)];
                      reg2439 <= ($signed($signed(reg2315)) <= ({reg2306[(3'h6):(2'h3)]} ~^ $signed((|reg2242))));
                      reg2440 <= $signed(($unsigned(((8'h9f) ?
                              (8'ha1) : forvar2297)) ?
                          reg2135 : (reg2310[(2'h3):(1'h0)] ?
                              (!(8'hb4)) : (forvar2408 ? (8'h9f) : reg2379))));
                    end
                  else
                    begin
                      reg2438 <= (-reg2223);
                      reg2439 <= $signed(reg2276);
                      reg2440 <= ((({reg2424} ?
                          (-reg2409) : (~|reg2407)) != reg2276[(2'h3):(1'h1)]) << ($unsigned((~&reg2194)) & (reg2438 || reg2432[(1'h1):(1'h1)])));
                    end
                end
              if ({$unsigned(reg2368[(4'hd):(3'h6)])})
                begin
                  for (forvar2441 = (1'h0); (forvar2441 < (1'h0)); forvar2441 = (forvar2441 + (1'h1)))
                    begin
                      reg2442 <= (&({forvar2380[(3'h5):(2'h3)]} | {(reg2265 <<< reg2339)}));
                      reg2443 <= {(!((reg2312 ?
                              reg2321 : reg2158) == (forvar2212 != forvar2139)))};
                      reg2444 <= (^((8'hb9) << $unsigned($unsigned(reg2131))));
                      reg2445 <= reg2180;
                    end
                  for (forvar2446 = (1'h0); (forvar2446 < (2'h2)); forvar2446 = (forvar2446 + (1'h1)))
                    begin
                      reg2447 <= ((!forvar2229) ?
                          ((^~(^~reg2133)) ?
                              ((-reg2217) - $signed(forvar2332)) : $unsigned(forvar2201[(2'h2):(1'h1)])) : $signed((reg2443[(1'h1):(1'h1)] ?
                              (reg2317 ? reg2276 : reg2396) : reg2170)));
                      reg2448 <= (~$unsigned(($unsigned(forvar2446) ~^ (8'ha1))));
                      reg2449 <= (8'ha7);
                      reg2450 <= forvar2219[(3'h4):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar2441 = (1'h0); (forvar2441 < (2'h2)); forvar2441 = (forvar2441 + (1'h1)))
                    begin
                      reg2442 <= reg2317;
                      reg2443 <= forvar2421[(5'h10):(4'hf)];
                      reg2444 <= ((8'hb5) ?
                          forvar2313 : (reg2199[(3'h7):(3'h6)] ^~ {$unsigned(reg2369)}));
                      reg2445 <= ((~$signed((^~forvar2429))) ?
                          {(reg2155 >= $signed(reg2157))} : {{$signed(wire2347)}});
                    end
                  reg2446 <= (8'hb3);
                end
            end
        end
      for (forvar2451 = (1'h0); (forvar2451 < (1'h1)); forvar2451 = (forvar2451 + (1'h1)))
        begin
          if ((({(^reg2403)} ?
                  (^reg2281[(2'h2):(1'h1)]) : forvar2179[(3'h5):(1'h1)]) ?
              (~forvar2377) : reg2237))
            begin
              for (forvar2452 = (1'h0); (forvar2452 < (1'h1)); forvar2452 = (forvar2452 + (1'h1)))
                begin
                  reg2453 <= ($unsigned($unsigned(reg2342[(1'h1):(1'h1)])) <= (+$signed((~^reg2304))));
                  for (forvar2454 = (1'h0); (forvar2454 < (2'h3)); forvar2454 = (forvar2454 + (1'h1)))
                    begin
                      reg2455 <= $signed($signed($unsigned((reg2311 << reg2190))));
                    end
                end
              if (({(~&reg2436)} - reg2333[(1'h0):(1'h0)]))
                begin
                  if ({$signed(((forvar2399 != reg2449) ?
                          reg2196[(4'hd):(4'h8)] : $signed(reg2252)))})
                    begin
                      reg2456 <= reg2449;
                      reg2457 <= ($signed(reg2382) != forvar2372);
                      reg2458 <= (~$signed(reg2191));
                      reg2459 <= (($unsigned(reg2167) ?
                          $signed($signed(reg2311)) : reg2324[(1'h1):(1'h0)]) >> (((reg2247 ?
                              reg2356 : (8'hb0)) <<< $unsigned(forvar2228)) ?
                          reg2357 : $unsigned((&reg2226))));
                    end
                  else
                    begin
                      reg2456 <= reg2176;
                      reg2457 <= $unsigned({{$unsigned(reg2434)}});
                    end
                  reg2460 <= $signed((~|((-reg2263) ?
                      (~|(8'ha9)) : $unsigned(forvar2300))));
                  if ($unsigned((reg2443[(4'he):(1'h0)] || (^reg2144))))
                    begin
                      reg2461 <= (reg2141[(4'h9):(1'h0)] * (($signed((8'hb5)) < {reg2272}) ?
                          $unsigned($unsigned(reg2306)) : forvar2315));
                      reg2462 <= (reg2276[(1'h1):(1'h0)] >>> reg2328);
                      reg2463 <= {(~|reg2368)};
                      reg2464 <= ((reg2354[(3'h4):(1'h1)] ?
                              $signed((+reg2280)) : reg2434[(3'h4):(2'h2)]) ?
                          (reg2169 >>> $signed((-forvar2294))) : (&(8'ha8)));
                    end
                  else
                    begin
                      reg2461 <= $signed($signed(reg2360));
                      reg2462 <= forvar2161[(2'h3):(1'h0)];
                      reg2463 <= ($unsigned((reg2264 + (reg2442 ?
                              forvar2144 : (8'h9c)))) ?
                          wire2126[(2'h2):(1'h0)] : (^~$signed((reg2405 ?
                              forvar2381 : reg2405))));
                      reg2464 <= (reg2242[(1'h0):(1'h0)] ?
                          (reg2374 != reg2319[(5'h10):(3'h4)]) : reg2443);
                    end
                end
              else
                begin
                  for (forvar2456 = (1'h0); (forvar2456 < (1'h0)); forvar2456 = (forvar2456 + (1'h1)))
                    begin
                      reg2457 <= forvar2170[(1'h0):(1'h0)];
                      reg2458 <= ($signed($signed({forvar2323})) + $unsigned(reg2261));
                      reg2459 <= forvar2135[(1'h1):(1'h1)];
                    end
                end
              for (forvar2465 = (1'h0); (forvar2465 < (2'h3)); forvar2465 = (forvar2465 + (1'h1)))
                begin
                  if ((!reg2186))
                    begin
                      reg2466 <= (~|((forvar2451 ?
                          $unsigned((8'ha5)) : (8'had)) ~^ ($signed(forvar2191) <= (wire2347 ?
                          forvar2367 : reg2324))));
                      reg2467 <= reg2204;
                    end
                  else
                    begin
                      reg2466 <= $unsigned((reg2216[(3'h6):(3'h4)] ?
                          $signed(reg2461) : $unsigned(reg2245)));
                    end
                end
              for (forvar2468 = (1'h0); (forvar2468 < (1'h0)); forvar2468 = (forvar2468 + (1'h1)))
                begin
                  for (forvar2469 = (1'h0); (forvar2469 < (2'h2)); forvar2469 = (forvar2469 + (1'h1)))
                    begin
                      reg2470 <= ((!$signed($signed(wire2123))) ?
                          $signed(((+(8'h9f)) != $signed(reg2303))) : {((|reg2172) == forvar2381)});
                      reg2471 <= (^{(^~$signed((8'h9f)))});
                      reg2472 <= ((((forvar2214 - reg2383) > $signed(reg2449)) << (-reg2157[(2'h3):(2'h3)])) ?
                          reg2385 : forvar2162);
                      reg2473 <= $signed({{reg2248[(1'h0):(1'h0)]}});
                    end
                  for (forvar2474 = (1'h0); (forvar2474 < (2'h3)); forvar2474 = (forvar2474 + (1'h1)))
                    begin
                      reg2475 <= $signed(forvar2191[(3'h5):(2'h3)]);
                    end
                  reg2476 <= $signed({$unsigned((~|forvar2314))});
                  reg2477 <= ((reg2301 ?
                          {(reg2339 <= reg2172)} : $signed($unsigned(forvar2399))) ?
                      $signed(((forvar2137 >> forvar2293) ?
                          (reg2449 <= reg2431) : $unsigned((8'hb1)))) : ($signed((reg2390 <<< reg2140)) ?
                          (^~((8'hba) ? (8'had) : reg2168)) : {(~^wire2124)}));
                end
            end
          else
            begin
              for (forvar2452 = (1'h0); (forvar2452 < (1'h1)); forvar2452 = (forvar2452 + (1'h1)))
                begin
                  reg2453 <= $signed(($signed((forvar2243 ?
                      reg2193 : (8'ha8))) || ($signed((8'hba)) ?
                      (^reg2157) : reg2255[(1'h0):(1'h0)])));
                end
              for (forvar2454 = (1'h0); (forvar2454 < (1'h0)); forvar2454 = (forvar2454 + (1'h1)))
                begin
                  if (((((reg2288 ? forvar2408 : reg2202) ?
                              (reg2144 ? reg2384 : (8'hae)) : (-reg2185)) ?
                          $signed(reg2238[(2'h2):(2'h2)]) : (reg2270 << (reg2379 > forvar2134))) ?
                      reg2471[(1'h1):(1'h0)] : forvar2192[(2'h2):(2'h2)]))
                    begin
                      reg2455 <= $unsigned(((^~$signed(reg2181)) ?
                          forvar2323 : $unsigned($unsigned(reg2280))));
                      reg2456 <= ((8'hb3) >> $signed(reg2277));
                      reg2457 <= $signed(({(reg2161 ? reg2151 : reg2193)} ?
                          (~^$signed(forvar2314)) : $signed((reg2411 - (8'hb3)))));
                    end
                  else
                    begin
                      reg2455 <= ((forvar2446[(3'h5):(2'h3)] ?
                              reg2246 : forvar2314[(1'h0):(1'h0)]) ?
                          forvar2374 : forvar2212);
                      reg2456 <= (~^$signed(reg2156));
                      reg2457 <= forvar2389;
                    end
                  if (reg2238[(2'h2):(1'h1)])
                    begin
                      reg2458 <= reg2136;
                      reg2459 <= (((reg2182 <<< (reg2329 ~^ (8'ha0))) ?
                              {reg2336} : ((^~reg2230) | $signed(forvar2386))) ?
                          (^~((!reg2424) ^ (reg2333 << reg2274))) : reg2357);
                    end
                  else
                    begin
                      reg2458 <= ({$signed($signed(reg2362))} ?
                          forvar2135[(2'h2):(1'h0)] : reg2431[(4'ha):(4'h9)]);
                      reg2459 <= $signed($signed($unsigned(forvar2341[(4'h8):(1'h0)])));
                    end
                  for (forvar2460 = (1'h0); (forvar2460 < (1'h0)); forvar2460 = (forvar2460 + (1'h1)))
                    begin
                      reg2461 <= {(((forvar2315 & reg2386) > reg2397) ?
                              (+forvar2356) : (+(reg2351 > reg2151)))};
                      reg2462 <= reg2249[(1'h0):(1'h0)];
                      reg2463 <= (^$unsigned(((forvar2465 ? reg2383 : (8'hb4)) ?
                          (8'hb5) : reg2229[(2'h2):(1'h1)])));
                      reg2464 <= (reg2284 ?
                          (((reg2398 ? reg2389 : reg2158) ?
                              reg2189 : reg2444[(2'h2):(1'h0)]) && reg2228[(3'h4):(1'h0)]) : $signed(reg2296));
                    end
                end
            end
          reg2478 <= $unsigned((reg2135[(3'h4):(3'h4)] ^~ (!(forvar2297 ?
              reg2175 : reg2177))));
          for (forvar2479 = (1'h0); (forvar2479 < (2'h2)); forvar2479 = (forvar2479 + (1'h1)))
            begin
              if ({reg2291})
                begin
                  reg2480 <= wire2124[(1'h0):(1'h0)];
                  reg2481 <= (reg2168 ?
                      $signed(($signed(forvar2429) >> (~^reg2170))) : (($unsigned(reg2253) ?
                              (reg2297 ^ (8'hb6)) : (~^(8'hb9))) ?
                          reg2251 : $signed($unsigned(reg2218))));
                end
              else
                begin
                  if ((((((8'had) || reg2153) ?
                      $unsigned((8'haa)) : (reg2430 | (8'h9f))) || (reg2275 ?
                      $unsigned(reg2251) : $unsigned(reg2236))) >= $unsigned($signed(((8'h9f) ?
                      reg2263 : reg2438)))))
                    begin
                      reg2480 <= reg2386[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg2480 <= $unsigned($signed(((~^reg2143) - $signed(reg2417))));
                      reg2481 <= (({(reg2260 ? reg2358 : reg2318)} ?
                          $signed($unsigned(reg2378)) : {reg2310}) - {$signed((&(8'hb3)))});
                    end
                end
            end
          for (forvar2482 = (1'h0); (forvar2482 < (2'h3)); forvar2482 = (forvar2482 + (1'h1)))
            begin
              for (forvar2483 = (1'h0); (forvar2483 < (2'h2)); forvar2483 = (forvar2483 + (1'h1)))
                begin
                  for (forvar2484 = (1'h0); (forvar2484 < (1'h1)); forvar2484 = (forvar2484 + (1'h1)))
                    begin
                      reg2485 <= ({($unsigned(reg2459) ?
                                  reg2202[(3'h4):(3'h4)] : (-reg2148))} ?
                          $signed($signed($unsigned((8'hb3)))) : reg2432);
                      reg2486 <= ($unsigned($unsigned(forvar2195)) ?
                          reg2246 : ((|$signed(reg2208)) ?
                              forvar2132 : $unsigned(reg2427)));
                      reg2487 <= ($signed(forvar2313[(1'h1):(1'h1)]) ?
                          forvar2429[(1'h0):(1'h0)] : {($signed((8'h9c)) | $signed((8'ha5)))});
                      reg2488 <= $signed($unsigned($signed({forvar2376})));
                    end
                  if ((reg2400[(3'h4):(1'h1)] ?
                      reg2444[(1'h0):(1'h0)] : $unsigned(((reg2487 ?
                              reg2216 : forvar2191) ?
                          (|(8'h9d)) : {(8'hb4)}))))
                    begin
                      reg2489 <= $unsigned(($unsigned($signed(reg2309)) < reg2177));
                      reg2490 <= reg2466;
                      reg2491 <= reg2336[(3'h4):(3'h4)];
                      reg2492 <= ((((&forvar2267) ?
                              $unsigned(reg2136) : reg2411[(1'h1):(1'h1)]) & $signed($unsigned((8'hb9)))) ?
                          $signed(reg2388[(4'h8):(3'h5)]) : reg2325[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg2489 <= $signed((-$unsigned(reg2218)));
                      reg2490 <= (reg2311[(4'hf):(1'h1)] ?
                          forvar2349 : $signed($signed({reg2278})));
                      reg2491 <= ($unsigned(reg2158) > ((~^(reg2301 - (8'hb3))) <= (reg2424 << $signed((8'hb0)))));
                    end
                  if ({{reg2426[(3'h5):(3'h5)]}})
                    begin
                      reg2493 <= $signed(forvar2373[(4'h8):(2'h3)]);
                      reg2494 <= (^~(reg2289 ?
                          (-$unsigned(reg2273)) : reg2326));
                      reg2495 <= forvar2319;
                      reg2496 <= (reg2402[(1'h0):(1'h0)] | {reg2374[(3'h7):(3'h4)]});
                    end
                  else
                    begin
                      reg2493 <= $unsigned((8'ha6));
                    end
                end
              if (reg2188)
                begin
                  for (forvar2497 = (1'h0); (forvar2497 < (2'h3)); forvar2497 = (forvar2497 + (1'h1)))
                    begin
                      reg2498 <= {reg2331[(1'h1):(1'h0)]};
                    end
                  for (forvar2499 = (1'h0); (forvar2499 < (1'h0)); forvar2499 = (forvar2499 + (1'h1)))
                    begin
                      reg2500 <= $signed(reg2207);
                      reg2501 <= reg2361;
                      reg2502 <= (~|(reg2170 >>> reg2391));
                      reg2503 <= {(+(+(forvar2134 ? reg2427 : reg2228)))};
                    end
                  if ($signed(forvar2316[(1'h0):(1'h0)]))
                    begin
                      reg2504 <= $signed($signed((-(reg2357 ?
                          forvar2451 : reg2376))));
                      reg2505 <= reg2491[(4'h9):(1'h1)];
                      reg2506 <= {(reg2199 == $unsigned($signed(reg2376)))};
                      reg2507 <= reg2165[(4'ha):(4'h9)];
                    end
                  else
                    begin
                      reg2504 <= ({((forvar2305 != reg2383) ?
                              (~|reg2184) : (~|forvar2150))} ~^ ((-$signed(forvar2152)) ?
                          ((reg2146 ? forvar2155 : (8'haa)) ?
                              forvar2267[(3'h5):(2'h2)] : {reg2263}) : $unsigned($signed(forvar2283))));
                      reg2505 <= (reg2277[(4'hd):(3'h7)] ?
                          $unsigned($signed({reg2463})) : (reg2306[(1'h1):(1'h1)] != ((-(8'hb0)) ?
                              (reg2403 <= (8'ha8)) : (~^forvar2139))));
                    end
                  if ((reg2449 << $signed($signed($unsigned((8'ha0))))))
                    begin
                      reg2508 <= forvar2335[(3'h4):(1'h1)];
                      reg2509 <= forvar2242;
                      reg2510 <= (~^(~&(+$unsigned(reg2506))));
                      reg2511 <= reg2164[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg2508 <= (~|(($signed(reg2142) ^ reg2245[(3'h4):(2'h3)]) ?
                          $signed(reg2471) : (&reg2404)));
                      reg2509 <= (((&$signed((8'hb8))) * (reg2296 <<< $unsigned(reg2291))) ?
                          $signed($signed($signed(reg2337))) : reg2323[(1'h1):(1'h1)]);
                      reg2510 <= (^({(reg2135 << forvar2452)} ?
                          reg2377 : $signed($signed(reg2320))));
                    end
                end
              else
                begin
                  for (forvar2497 = (1'h0); (forvar2497 < (1'h1)); forvar2497 = (forvar2497 + (1'h1)))
                    begin
                      reg2498 <= reg2321;
                      reg2499 <= $signed(reg2340[(3'h7):(3'h7)]);
                      reg2500 <= forvar2376;
                      reg2501 <= (^~(((^(8'ha1)) && (reg2149 >= forvar2232)) && ((reg2357 | (8'had)) ?
                          reg2189 : (~^reg2283))));
                    end
                  for (forvar2502 = (1'h0); (forvar2502 < (1'h0)); forvar2502 = (forvar2502 + (1'h1)))
                    begin
                      reg2503 <= (~&reg2505);
                      reg2504 <= $unsigned((reg2222[(1'h0):(1'h0)] ?
                          $unsigned($unsigned(reg2445)) : reg2283));
                      reg2505 <= reg2417;
                    end
                end
              for (forvar2512 = (1'h0); (forvar2512 < (2'h2)); forvar2512 = (forvar2512 + (1'h1)))
                begin
                  reg2513 <= ($unsigned({$unsigned(reg2434)}) ?
                      forvar2271[(4'ha):(1'h0)] : reg2461[(1'h0):(1'h0)]);
                end
            end
        end
      if (((((reg2436 ? reg2232 : reg2171) ?
              (reg2431 ? reg2503 : (8'h9c)) : (~|reg2253)) != ((reg2297 ?
              reg2331 : (8'h9c)) ^ (reg2377 || (8'hac)))) ?
          reg2237 : ((+(reg2197 << forvar2315)) != ($signed((8'haa)) ?
              ((8'ha1) ? (8'hb7) : forvar2155) : forvar2214[(4'hb):(4'h8)]))))
        begin
          if ($signed((((wire2125 >= reg2366) ?
              (^~reg2364) : (reg2171 ? reg2478 : forvar2198)) <<< (reg2356 ?
              $unsigned(forvar2267) : (forvar2256 ? reg2467 : reg2276)))))
            begin
              for (forvar2514 = (1'h0); (forvar2514 < (1'h1)); forvar2514 = (forvar2514 + (1'h1)))
                begin
                  if ($signed(reg2189))
                    begin
                      reg2515 <= ($unsigned($unsigned((reg2492 ?
                          reg2197 : forvar2152))) < $unsigned(((reg2139 == forvar2243) >>> (reg2281 > forvar2229))));
                      reg2516 <= $signed($unsigned((~|reg2376)));
                    end
                  else
                    begin
                      reg2515 <= (^reg2248[(3'h4):(2'h3)]);
                      reg2516 <= forvar2514;
                      reg2517 <= forvar2267[(4'h8):(1'h1)];
                      reg2518 <= (^$unsigned(($signed(reg2481) ?
                          reg2169[(1'h0):(1'h0)] : $unsigned(reg2473))));
                    end
                  reg2519 <= (reg2503 && (reg2392 >> ((forvar2395 * reg2400) ?
                      (forvar2305 | reg2220) : reg2167)));
                  for (forvar2520 = (1'h0); (forvar2520 < (1'h0)); forvar2520 = (forvar2520 + (1'h1)))
                    begin
                      reg2521 <= $signed(reg2223);
                      reg2522 <= $unsigned((reg2271 ?
                          $signed((!reg2490)) : $signed($signed(reg2411))));
                    end
                  for (forvar2523 = (1'h0); (forvar2523 < (2'h2)); forvar2523 = (forvar2523 + (1'h1)))
                    begin
                      reg2524 <= $signed((^reg2164));
                    end
                end
              if (forvar2408[(2'h2):(1'h1)])
                begin
                  if ((reg2403[(4'he):(1'h1)] - $signed(($unsigned((8'haa)) | reg2268[(1'h0):(1'h0)]))))
                    begin
                      reg2525 <= forvar2232[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg2525 <= ($signed($unsigned((reg2415 >>> reg2335))) * reg2349);
                      reg2526 <= $signed($unsigned((forvar2315[(3'h4):(2'h3)] & reg2351[(1'h1):(1'h1)])));
                    end
                  reg2527 <= $unsigned(reg2491[(4'h8):(2'h3)]);
                  reg2528 <= $signed($unsigned((~^(8'hb5))));
                end
              else
                begin
                  if ({(8'h9f)})
                    begin
                      reg2525 <= reg2496;
                      reg2526 <= (reg2157 ^~ forvar2174[(4'h8):(3'h6)]);
                      reg2527 <= $signed(((~^forvar2367[(2'h3):(1'h1)]) || $signed((reg2313 >= reg2177))));
                    end
                  else
                    begin
                      reg2525 <= ((($signed(reg2335) ?
                              (~reg2170) : (reg2130 ?
                                  reg2406 : (8'h9e))) <= reg2328) ?
                          (8'h9c) : (^reg2525));
                      reg2526 <= forvar2456[(2'h2):(1'h1)];
                      reg2527 <= (($unsigned((reg2377 ? reg2189 : (8'hab))) ?
                          {$signed(reg2390)} : reg2440) >= (~|reg2516));
                      reg2528 <= reg2417;
                    end
                  reg2529 <= ((^~$signed((~&reg2323))) != (^~(reg2315 > {reg2279})));
                  if (reg2252[(3'h4):(2'h3)])
                    begin
                      reg2530 <= $unsigned($unsigned($signed(reg2447[(4'h8):(3'h7)])));
                    end
                  else
                    begin
                      reg2530 <= forvar2294;
                    end
                end
              if (forvar2497)
                begin
                  if ($signed((^((reg2159 | reg2316) ?
                      $signed((8'hb8)) : {reg2137}))))
                    begin
                      reg2531 <= $unsigned((|(~|(forvar2213 ?
                          reg2295 : reg2287))));
                    end
                  else
                    begin
                      reg2531 <= ((!$unsigned($unsigned((8'hb5)))) != reg2369);
                      reg2532 <= (^$signed($signed((~|forvar2148))));
                    end
                  for (forvar2533 = (1'h0); (forvar2533 < (2'h3)); forvar2533 = (forvar2533 + (1'h1)))
                    begin
                      reg2534 <= (8'hb5);
                      reg2535 <= ({(-forvar2152[(1'h1):(1'h0)])} == (($unsigned(reg2459) * (^~(8'hb3))) ?
                          forvar2150 : {reg2218[(2'h2):(1'h1)]}));
                      reg2536 <= {{$unsigned(forvar2329[(3'h6):(3'h5)])}};
                      reg2537 <= (reg2261[(2'h3):(1'h1)] ?
                          (($unsigned(forvar2133) ?
                              (reg2358 ? (8'ha1) : (8'ha3)) : ((8'hba) ?
                                  reg2322 : reg2184)) ^ ((reg2345 <<< forvar2133) ?
                              $signed((8'hb1)) : $signed(reg2444))) : $unsigned($unsigned((^reg2345))));
                    end
                  if (((reg2276 ?
                      forvar2338[(1'h1):(1'h1)] : (8'ha7)) > forvar2191))
                    begin
                      reg2538 <= (($unsigned((reg2184 ?
                              reg2487 : reg2494)) != $unsigned($unsigned(wire2347))) ?
                          reg2473[(3'h5):(1'h1)] : $signed((forvar2433 >>> {reg2331})));
                      reg2539 <= $signed(forvar2141[(4'hd):(4'h8)]);
                      reg2540 <= forvar2358[(3'h5):(1'h1)];
                      reg2541 <= ((reg2492 ~^ $unsigned((|reg2498))) & ($signed($signed(reg2297)) < ({reg2345} || (reg2255 ?
                          (8'h9e) : reg2315))));
                    end
                  else
                    begin
                      reg2538 <= ((~&($signed((8'h9e)) ?
                              (+reg2511) : forvar2267[(4'hc):(3'h4)])) ?
                          $signed((^~(!(8'hba)))) : (|(reg2319[(4'ha):(3'h7)] ?
                              reg2311[(3'h6):(2'h2)] : $signed(reg2340))));
                    end
                  for (forvar2542 = (1'h0); (forvar2542 < (2'h3)); forvar2542 = (forvar2542 + (1'h1)))
                    begin
                      reg2543 <= ((!(reg2302 ?
                              $signed(forvar2499) : $unsigned(reg2351))) ?
                          reg2504 : (8'hb2));
                    end
                end
              else
                begin
                  if (reg2270)
                    begin
                      reg2531 <= $unsigned($signed($unsigned((-reg2186))));
                      reg2532 <= ({forvar2452[(3'h6):(2'h3)]} & (+(forvar2214[(4'h8):(2'h3)] ?
                          (reg2518 >>> reg2378) : reg2133)));
                    end
                  else
                    begin
                      reg2531 <= (($signed((reg2534 ^ reg2453)) ?
                          reg2152[(1'h1):(1'h0)] : (&((8'ha3) ?
                              reg2413 : reg2447))) ^~ {reg2509[(4'ha):(1'h1)]});
                      reg2532 <= $signed({(+$signed(forvar2465))});
                      reg2533 <= {{$unsigned((reg2204 ?
                                  forvar2256 : reg2538))}};
                      reg2534 <= ($signed($signed((reg2197 < reg2543))) - reg2131[(2'h2):(1'h1)]);
                    end
                  for (forvar2535 = (1'h0); (forvar2535 < (1'h0)); forvar2535 = (forvar2535 + (1'h1)))
                    begin
                      reg2536 <= (~(forvar2428[(1'h1):(1'h1)] > $signed($signed(reg2220))));
                    end
                  for (forvar2537 = (1'h0); (forvar2537 < (1'h0)); forvar2537 = (forvar2537 + (1'h1)))
                    begin
                      reg2538 <= ({{forvar2214[(3'h4):(3'h4)]}} || reg2243[(5'h10):(2'h2)]);
                      reg2539 <= $signed($unsigned($unsigned({reg2423})));
                      reg2540 <= forvar2482;
                    end
                end
            end
          else
            begin
              if ($signed((forvar2175 ?
                  (reg2219 * (forvar2367 << (8'ha0))) : ($unsigned(reg2286) ?
                      (&reg2356) : (reg2432 ? (8'hb3) : reg2513)))))
                begin
                  if (forvar2191)
                    begin
                      reg2514 <= $unsigned(reg2353);
                    end
                  else
                    begin
                      reg2514 <= $unsigned($signed(reg2263));
                    end
                  for (forvar2515 = (1'h0); (forvar2515 < (1'h0)); forvar2515 = (forvar2515 + (1'h1)))
                    begin
                      reg2516 <= forvar2421[(1'h1):(1'h1)];
                      reg2517 <= reg2466;
                      reg2518 <= (^~(~&reg2155[(4'hb):(3'h6)]));
                    end
                end
              else
                begin
                  if ((&$signed(((~|forvar2380) ?
                      (reg2143 ?
                          reg2226 : forvar2441) : (forvar2285 <= forvar2280)))))
                    begin
                      reg2514 <= {(+(reg2235[(4'ha):(4'ha)] ?
                              reg2402[(3'h4):(3'h4)] : $signed(reg2325)))};
                    end
                  else
                    begin
                      reg2514 <= (~($unsigned(reg2353[(1'h1):(1'h1)]) ^ (forvar2537[(1'h0):(1'h0)] ?
                          (!reg2130) : (reg2131 ? forvar2389 : (8'ha8)))));
                      reg2515 <= ($unsigned(reg2321[(4'hd):(3'h7)]) | reg2230);
                    end
                end
              reg2519 <= (($signed({(8'hac)}) || $unsigned(((8'hb4) ?
                  reg2476 : reg2416))) != (((reg2503 ?
                  forvar2315 : forvar2315) <<< reg2513[(2'h2):(2'h2)]) >> {$unsigned(forvar2232)}));
              for (forvar2520 = (1'h0); (forvar2520 < (1'h1)); forvar2520 = (forvar2520 + (1'h1)))
                begin
                  for (forvar2521 = (1'h0); (forvar2521 < (1'h0)); forvar2521 = (forvar2521 + (1'h1)))
                    begin
                      reg2522 <= (forvar2428 ?
                          $unsigned(reg2336[(2'h2):(1'h1)]) : reg2217);
                      reg2523 <= $unsigned(forvar2429);
                      reg2524 <= ({(8'hba)} ?
                          ($unsigned($signed(forvar2338)) ?
                              reg2209[(1'h0):(1'h0)] : $signed(reg2410)) : $unsigned($signed($signed(wire2126))));
                    end
                  if ($unsigned({$signed((^~(8'hb1)))}))
                    begin
                      reg2525 <= ($signed($unsigned($unsigned(reg2415))) ?
                          $signed(($signed(forvar2367) >> reg2324)) : (reg2170 * ((~&forvar2419) | reg2315[(3'h6):(3'h4)])));
                      reg2526 <= {(reg2358[(3'h5):(3'h5)] ?
                              $signed($unsigned(reg2344)) : forvar2468[(3'h4):(1'h1)])};
                    end
                  else
                    begin
                      reg2525 <= forvar2175;
                      reg2526 <= reg2489;
                    end
                  if (({reg2277} ?
                      $signed($unsigned((+forvar2195))) : $unsigned((8'hae))))
                    begin
                      reg2527 <= $unsigned((forvar2381[(2'h3):(2'h3)] ?
                          reg2538[(1'h1):(1'h0)] : (&(forvar2483 || (8'ha7)))));
                    end
                  else
                    begin
                      reg2527 <= reg2294[(3'h7):(3'h5)];
                      reg2528 <= {(&(((8'ha6) > reg2540) ?
                              ((8'ha8) ?
                                  reg2318 : (8'ha6)) : reg2297[(4'he):(4'he)]))};
                      reg2529 <= $signed({reg2405});
                      reg2530 <= ((~&$signed(forvar2305)) || reg2235);
                    end
                  if ((reg2254[(4'h9):(3'h4)] < reg2192[(3'h7):(2'h3)]))
                    begin
                      reg2531 <= (forvar2474 ?
                          (((8'hab) ? $signed(reg2275) : (&forvar2300)) ?
                              reg2168[(1'h0):(1'h0)] : ($unsigned(forvar2191) >= $signed(forvar2294))) : reg2342[(4'hb):(2'h2)]);
                      reg2532 <= ((~$signed((forvar2479 ?
                          reg2526 : reg2317))) || (^~$unsigned((forvar2161 < (8'ha1)))));
                      reg2533 <= $signed(($unsigned(reg2426) >>> reg2326));
                    end
                  else
                    begin
                      reg2531 <= (reg2466[(3'h5):(3'h4)] ?
                          reg2525 : (+reg2358[(1'h0):(1'h0)]));
                      reg2532 <= $unsigned(reg2533[(4'h9):(3'h5)]);
                      reg2533 <= ($unsigned($unsigned(forvar2367[(2'h3):(2'h3)])) || $signed($signed($unsigned(reg2268))));
                      reg2534 <= $unsigned(($unsigned((|forvar2421)) | (reg2337[(1'h1):(1'h1)] ?
                          (forvar2133 - reg2171) : $signed((8'ha8)))));
                    end
                end
            end
          for (forvar2544 = (1'h0); (forvar2544 < (1'h1)); forvar2544 = (forvar2544 + (1'h1)))
            begin
              reg2545 <= reg2393[(4'hb):(4'hb)];
              if ((~($unsigned(wire2347) <= (~reg2228[(1'h1):(1'h0)]))))
                begin
                  if ($unsigned(wire2123))
                    begin
                      reg2546 <= (&($signed((forvar2338 == reg2195)) != forvar2148));
                      reg2547 <= (($signed(reg2313) & forvar2468[(4'h9):(2'h3)]) >>> ($unsigned(reg2130[(3'h6):(2'h2)]) > $signed($unsigned(reg2493))));
                      reg2548 <= $unsigned(((^~$signed(reg2184)) ?
                          ((forvar2399 ? reg2164 : reg2302) ?
                              (~|(8'hb7)) : (!(8'hae))) : (((8'ha1) ?
                              forvar2381 : forvar2206) - (reg2427 & reg2141))));
                      reg2549 <= $unsigned($unsigned((((8'hb8) ?
                              reg2134 : reg2282) ?
                          (reg2255 && reg2140) : reg2243[(4'hb):(4'h8)])));
                    end
                  else
                    begin
                      reg2546 <= (((forvar2353 ?
                          $signed(forvar2271) : (+(8'hba))) >> reg2318[(1'h0):(1'h0)]) - (&((!forvar2286) & $signed((8'hb7)))));
                      reg2547 <= (($signed($signed(reg2253)) <<< $signed({reg2387})) ?
                          $unsigned($unsigned(reg2166)) : $unsigned(forvar2381[(3'h5):(2'h2)]));
                      reg2548 <= (8'ha8);
                    end
                  if ({$signed({((8'hb5) ? (8'h9e) : reg2308)})})
                    begin
                      reg2550 <= $unsigned((-(|reg2502)));
                    end
                  else
                    begin
                      reg2550 <= (reg2313 ?
                          reg2261 : ((|(!reg2154)) << ((reg2383 ?
                              reg2541 : reg2434) <<< wire2129)));
                    end
                end
              else
                begin
                  reg2546 <= ($signed(reg2333[(1'h0):(1'h0)]) <= $signed(((reg2310 | reg2171) ?
                      {reg2301} : (reg2526 <= (8'hba)))));
                end
              if ((+{(reg2230[(1'h1):(1'h0)] <<< reg2193[(3'h5):(2'h3)])}))
                begin
                  for (forvar2551 = (1'h0); (forvar2551 < (2'h2)); forvar2551 = (forvar2551 + (1'h1)))
                    begin
                      reg2552 <= (($unsigned(reg2279) ?
                              {$signed(reg2211)} : $signed((forvar2299 >= forvar2451))) ?
                          ($signed($unsigned(forvar2162)) ?
                              ($signed((8'hae)) ?
                                  {forvar2372} : {forvar2395}) : reg2402) : (((reg2320 ?
                                  (8'hb2) : reg2159) ?
                              (reg2349 ?
                                  (8'haa) : (8'ha0)) : (-reg2525)) * reg2239[(3'h4):(1'h0)]));
                      reg2553 <= $signed({((reg2324 & reg2379) ^~ (reg2225 << forvar2156))});
                    end
                  for (forvar2554 = (1'h0); (forvar2554 < (2'h2)); forvar2554 = (forvar2554 + (1'h1)))
                    begin
                      reg2555 <= reg2384;
                      reg2556 <= {(~&reg2185)};
                      reg2557 <= $unsigned((reg2368[(1'h1):(1'h0)] ?
                          reg2345 : $unsigned((^reg2203))));
                      reg2558 <= (8'hb0);
                    end
                  if (reg2132[(2'h3):(2'h2)])
                    begin
                      reg2559 <= reg2275[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg2559 <= $unsigned((reg2552 ?
                          forvar2133[(2'h3):(2'h3)] : $signed(((8'haf) != reg2383))));
                      reg2560 <= $signed(reg2329[(3'h6):(3'h5)]);
                    end
                end
              else
                begin
                  for (forvar2551 = (1'h0); (forvar2551 < (2'h3)); forvar2551 = (forvar2551 + (1'h1)))
                    begin
                      reg2552 <= (8'hae);
                      reg2553 <= ($unsigned({reg2303}) << reg2300);
                      reg2554 <= (~^reg2161[(2'h3):(1'h1)]);
                      reg2555 <= ((-reg2537) ?
                          $signed($signed($unsigned(reg2450))) : (reg2462 ?
                              $signed($signed(forvar2134)) : {$signed(forvar2256)}));
                    end
                  if ($unsigned((8'hb7)))
                    begin
                      reg2556 <= ($signed(forvar2551) ?
                          reg2344 : $unsigned((&(~&forvar2314))));
                    end
                  else
                    begin
                      reg2556 <= reg2411;
                    end
                  for (forvar2557 = (1'h0); (forvar2557 < (2'h3)); forvar2557 = (forvar2557 + (1'h1)))
                    begin
                      reg2558 <= $unsigned(reg2486);
                      reg2559 <= $signed($unsigned((~|forvar2256[(1'h0):(1'h0)])));
                    end
                  for (forvar2560 = (1'h0); (forvar2560 < (2'h2)); forvar2560 = (forvar2560 + (1'h1)))
                    begin
                      reg2561 <= (($signed(((8'hae) && reg2349)) ?
                              $unsigned(reg2296) : forvar2174[(1'h0):(1'h0)]) ?
                          {{forvar2367[(1'h1):(1'h1)]}} : ({(reg2207 * reg2283)} << (((8'hae) ?
                                  forvar2452 : forvar2544) ?
                              $unsigned((8'hb3)) : reg2250)));
                    end
                end
              for (forvar2562 = (1'h0); (forvar2562 < (2'h2)); forvar2562 = (forvar2562 + (1'h1)))
                begin
                  for (forvar2563 = (1'h0); (forvar2563 < (1'h0)); forvar2563 = (forvar2563 + (1'h1)))
                    begin
                      reg2564 <= (((~^(reg2470 ?
                              forvar2286 : forvar2377)) == {reg2165[(1'h0):(1'h0)]}) ?
                          (8'h9c) : $signed(forvar2213[(2'h3):(1'h0)]));
                    end
                  if (($signed(((^~reg2131) ?
                      forvar2201 : $unsigned(reg2487))) >>> (^($unsigned(forvar2152) >= $unsigned(reg2344)))))
                    begin
                      reg2565 <= $signed({reg2455[(2'h2):(1'h1)]});
                      reg2566 <= reg2369;
                      reg2567 <= (reg2560 * {(((8'hab) < reg2140) ?
                              $signed(reg2243) : (reg2251 ~^ (8'hb3)))});
                    end
                  else
                    begin
                      reg2565 <= reg2488[(3'h5):(2'h3)];
                      reg2566 <= reg2392;
                      reg2567 <= {reg2137[(2'h3):(1'h0)]};
                    end
                end
            end
          for (forvar2568 = (1'h0); (forvar2568 < (1'h0)); forvar2568 = (forvar2568 + (1'h1)))
            begin
              if (reg2131[(4'h9):(2'h2)])
                begin
                  for (forvar2569 = (1'h0); (forvar2569 < (2'h2)); forvar2569 = (forvar2569 + (1'h1)))
                    begin
                      reg2570 <= reg2558[(2'h3):(2'h3)];
                      reg2571 <= reg2413;
                      reg2572 <= (((((8'h9f) ? forvar2441 : (8'had)) ?
                              {reg2157} : reg2436) <<< (forvar2297[(1'h1):(1'h0)] ~^ $signed(reg2431))) ?
                          ($unsigned($unsigned(reg2307)) + ($signed((8'hae)) | $signed(reg2350))) : ((forvar2232[(3'h4):(2'h3)] ?
                              (8'hb4) : $signed(reg2161)) >>> reg2255));
                    end
                  for (forvar2573 = (1'h0); (forvar2573 < (1'h0)); forvar2573 = (forvar2573 + (1'h1)))
                    begin
                      reg2574 <= $signed((^~(reg2207[(2'h2):(1'h0)] + $signed(reg2250))));
                      reg2575 <= $signed($unsigned(((^~reg2271) ^~ $unsigned((8'h9c)))));
                    end
                  for (forvar2576 = (1'h0); (forvar2576 < (2'h3)); forvar2576 = (forvar2576 + (1'h1)))
                    begin
                      reg2577 <= reg2536[(4'h8):(3'h4)];
                    end
                end
              else
                begin
                  if ($signed(reg2279[(1'h0):(1'h0)]))
                    begin
                      reg2569 <= reg2487[(1'h1):(1'h1)];
                      reg2570 <= reg2444[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2569 <= (-($unsigned(reg2554[(1'h1):(1'h1)]) ?
                          ((reg2486 ?
                              forvar2173 : reg2330) & $signed((8'ha1))) : ($signed(reg2288) ?
                              (forvar2515 != (8'haf)) : $unsigned((8'ha3)))));
                      reg2570 <= $signed($unsigned(reg2473));
                      reg2571 <= (reg2500[(2'h2):(1'h0)] | forvar2166[(1'h0):(1'h0)]);
                      reg2572 <= $unsigned((+((8'hb0) >> (~&reg2223))));
                    end
                  for (forvar2573 = (1'h0); (forvar2573 < (1'h0)); forvar2573 = (forvar2573 + (1'h1)))
                    begin
                      reg2574 <= (forvar2465[(3'h5):(2'h2)] ?
                          reg2300 : (reg2180 ?
                              $unsigned((reg2339 ?
                                  forvar2499 : reg2382)) : {{forvar2433}}));
                      reg2575 <= ($signed(forvar2163[(3'h4):(2'h2)]) ?
                          (($unsigned(reg2499) > forvar2165) ^ {$signed(reg2291)}) : $signed((^(reg2358 ?
                              reg2470 : reg2250))));
                    end
                  reg2576 <= $unsigned(reg2167[(3'h4):(1'h1)]);
                end
            end
          reg2578 <= reg2168[(1'h0):(1'h0)];
        end
      else
        begin
          for (forvar2514 = (1'h0); (forvar2514 < (2'h2)); forvar2514 = (forvar2514 + (1'h1)))
            begin
              reg2515 <= $unsigned((-{(forvar2376 ? reg2131 : reg2260)}));
              if ((reg2574[(3'h5):(3'h4)] ?
                  reg2467 : forvar2377[(3'h5):(3'h5)]))
                begin
                  if (reg2578)
                    begin
                      reg2516 <= forvar2499[(1'h1):(1'h0)];
                      reg2517 <= {reg2189[(2'h2):(2'h2)]};
                      reg2518 <= $unsigned((reg2203[(1'h1):(1'h0)] ~^ $signed((&(8'hb7)))));
                      reg2519 <= reg2406[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg2516 <= (+{(((8'haf) ?
                              reg2218 : reg2369) * forvar2353)});
                      reg2517 <= (reg2574 ?
                          ((((8'ha2) ?
                              reg2332 : wire2129) != (~reg2571)) < (-reg2400)) : (-$signed(reg2280[(1'h1):(1'h1)])));
                    end
                  reg2520 <= reg2272[(3'h4):(1'h0)];
                  if ((8'ha2))
                    begin
                      reg2521 <= (({reg2496} ?
                              (!{(8'ha7)}) : $signed((-reg2530))) ?
                          (~(&{(8'ha5)})) : ($unsigned(forvar2468) ?
                              ((reg2310 ~^ reg2318) ?
                                  ((8'had) ?
                                      forvar2386 : reg2546) : {reg2308}) : $signed((-reg2331))));
                    end
                  else
                    begin
                      reg2521 <= reg2254;
                      reg2522 <= $unsigned(forvar2367[(2'h3):(2'h3)]);
                    end
                end
              else
                begin
                  if ((-forvar2191))
                    begin
                      reg2516 <= {$signed((!((8'hb1) ? reg2277 : reg2254)))};
                      reg2517 <= $unsigned(reg2263[(3'h4):(3'h4)]);
                    end
                  else
                    begin
                      reg2516 <= $signed(reg2456);
                      reg2517 <= (&forvar2137[(4'hb):(4'h8)]);
                      reg2518 <= {(|(~(reg2222 ? (8'hb9) : reg2387)))};
                    end
                  for (forvar2519 = (1'h0); (forvar2519 < (2'h3)); forvar2519 = (forvar2519 + (1'h1)))
                    begin
                      reg2520 <= reg2537;
                      reg2521 <= $unsigned((reg2446[(4'hc):(4'hb)] != {{reg2467}}));
                      reg2522 <= (($unsigned(((8'ha0) ? (8'ha9) : reg2561)) ?
                              (forvar2386[(2'h3):(1'h1)] ?
                                  (8'hb5) : $unsigned(reg2366)) : (&(~&reg2402))) ?
                          reg2506 : reg2553);
                    end
                  for (forvar2523 = (1'h0); (forvar2523 < (1'h1)); forvar2523 = (forvar2523 + (1'h1)))
                    begin
                      reg2524 <= forvar2304[(3'h4):(1'h1)];
                      reg2525 <= ($signed((|(reg2511 ? reg2181 : (8'ha0)))) ?
                          (reg2354[(1'h0):(1'h0)] | reg2499) : $signed(forvar2243[(3'h4):(2'h2)]));
                      reg2526 <= {reg2494[(1'h1):(1'h0)]};
                      reg2527 <= reg2356[(3'h4):(1'h1)];
                    end
                end
              reg2528 <= $signed($unsigned(reg2208));
            end
          for (forvar2529 = (1'h0); (forvar2529 < (1'h0)); forvar2529 = (forvar2529 + (1'h1)))
            begin
              reg2530 <= (((~|reg2259[(4'h8):(2'h3)]) | (reg2334[(4'h9):(3'h7)] == {reg2531})) >> reg2517);
              if ((^forvar2134[(3'h7):(3'h7)]))
                begin
                  for (forvar2531 = (1'h0); (forvar2531 < (1'h1)); forvar2531 = (forvar2531 + (1'h1)))
                    begin
                      reg2532 <= $signed($unsigned(forvar2358[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  if ({($signed($signed(reg2459)) ?
                          reg2310 : $unsigned(reg2548[(1'h1):(1'h1)]))})
                    begin
                      reg2531 <= (+(&reg2396[(4'he):(2'h2)]));
                    end
                  else
                    begin
                      reg2531 <= $unsigned(forvar2560);
                      reg2532 <= $signed(((8'haa) >>> $signed((reg2447 > reg2359))));
                    end
                end
            end
          for (forvar2533 = (1'h0); (forvar2533 < (2'h2)); forvar2533 = (forvar2533 + (1'h1)))
            begin
              reg2534 <= (8'ha2);
            end
          for (forvar2535 = (1'h0); (forvar2535 < (1'h1)); forvar2535 = (forvar2535 + (1'h1)))
            begin
              for (forvar2536 = (1'h0); (forvar2536 < (1'h1)); forvar2536 = (forvar2536 + (1'h1)))
                begin
                  for (forvar2537 = (1'h0); (forvar2537 < (1'h0)); forvar2537 = (forvar2537 + (1'h1)))
                    begin
                      reg2538 <= $signed((^reg2218[(2'h2):(1'h0)]));
                    end
                  if (forvar2329[(4'h8):(1'h0)])
                    begin
                      reg2539 <= forvar2469;
                    end
                  else
                    begin
                      reg2539 <= $unsigned(((^~(reg2299 ?
                          reg2575 : (8'h9c))) & $unsigned((reg2278 ?
                          reg2144 : forvar2134))));
                      reg2540 <= $unsigned((|((reg2216 ? reg2535 : reg2170) ?
                          reg2136[(3'h7):(3'h4)] : $unsigned(forvar2134))));
                    end
                  for (forvar2541 = (1'h0); (forvar2541 < (2'h3)); forvar2541 = (forvar2541 + (1'h1)))
                    begin
                      reg2542 <= reg2514[(3'h4):(2'h3)];
                      reg2543 <= ((reg2146 && {(8'hb8)}) ?
                          reg2197 : (|reg2461));
                      reg2544 <= $unsigned((&((&forvar2148) ?
                          {reg2184} : forvar2356[(3'h7):(3'h5)])));
                      reg2545 <= wire2347;
                    end
                  for (forvar2546 = (1'h0); (forvar2546 < (1'h0)); forvar2546 = (forvar2546 + (1'h1)))
                    begin
                      reg2547 <= forvar2419;
                      reg2548 <= {reg2158};
                      reg2549 <= (|{$unsigned(forvar2465)});
                    end
                end
              for (forvar2550 = (1'h0); (forvar2550 < (2'h2)); forvar2550 = (forvar2550 + (1'h1)))
                begin
                  for (forvar2551 = (1'h0); (forvar2551 < (2'h3)); forvar2551 = (forvar2551 + (1'h1)))
                    begin
                      reg2552 <= $unsigned(((8'ha9) ?
                          ($unsigned((8'hae)) ?
                              (~^reg2538) : reg2475[(3'h6):(2'h2)]) : ((forvar2465 ?
                                  forvar2388 : forvar2318) ?
                              (reg2172 << reg2361) : $signed((8'had)))));
                    end
                end
              reg2553 <= reg2142;
            end
        end
    end
  assign wire2579 = ((!(^~(forvar2482 - reg2368))) >>> (~&(forvar2456 ?
                        (^reg2247) : (&reg2480))));
  assign wire2580 = $signed($unsigned((8'h9e)));
  assign wire2581 = {{($unsigned((8'ha8)) ?
                                {forvar2219} : (reg2300 != reg2370))}};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4572
#( parameter param7005 = {({(8'hb9)} ? ((~(8'hac)) == ((8'ha3) ? (8'hb0) : (8'ha5))) : {((8'hb2) ^~ (8'hb5))})} )
(y, clk, wire4573, wire4574, wire4575, wire4576);
  output wire [(32'h2cc2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire4573;
  input wire [(4'hc):(1'h0)] wire4574;
  input wire [(2'h3):(1'h0)] wire4575;
  input wire signed [(3'h4):(1'h0)] wire4576;
  reg [(3'h5):(1'h0)] reg7004 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg7003 = (1'h0);
  reg [(4'hd):(1'h0)] reg7002 = (1'h0);
  reg [(4'hc):(1'h0)] reg7001 = (1'h0);
  reg [(4'hf):(1'h0)] reg7000 = (1'h0);
  reg [(4'hc):(1'h0)] reg6999 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6998 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6997 = (1'h0);
  reg [(4'h8):(1'h0)] reg6996 = (1'h0);
  reg [(4'h8):(1'h0)] reg6995 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6994 = (1'h0);
  reg [(2'h2):(1'h0)] reg6993 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6992 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6991 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6990 = (1'h0);
  reg [(5'h10):(1'h0)] reg6989 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6988 = (1'h0);
  reg [(3'h7):(1'h0)] reg6987 = (1'h0);
  reg [(4'hb):(1'h0)] reg6986 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6985 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6984 = (1'h0);
  reg [(3'h6):(1'h0)] reg6983 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6982 = (1'h0);
  reg [(3'h7):(1'h0)] reg6981 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6980 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6979 = (1'h0);
  reg [(4'hc):(1'h0)] reg6978 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6977 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6976 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6975 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6974 = (1'h0);
  reg [(4'hf):(1'h0)] reg6973 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6972 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6971 = (1'h0);
  reg [(3'h6):(1'h0)] reg6970 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6969 = (1'h0);
  reg [(4'ha):(1'h0)] reg6968 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6967 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6966 = (1'h0);
  reg [(5'h10):(1'h0)] reg6965 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6964 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6963 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6962 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6961 = (1'h0);
  reg [(4'h9):(1'h0)] reg6960 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6959 = (1'h0);
  reg [(2'h2):(1'h0)] forvar6958 = (1'h0);
  reg [(3'h4):(1'h0)] reg6957 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6956 = (1'h0);
  reg [(4'hb):(1'h0)] reg6955 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6954 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6953 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6952 = (1'h0);
  reg [(2'h2):(1'h0)] reg6951 = (1'h0);
  reg [(2'h2):(1'h0)] reg6944 = (1'h0);
  reg [(4'he):(1'h0)] reg6950 = (1'h0);
  reg [(4'hb):(1'h0)] reg6949 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6948 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6947 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6946 = (1'h0);
  reg [(4'hb):(1'h0)] reg6945 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6944 = (1'h0);
  reg [(5'h10):(1'h0)] reg6943 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6942 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6941 = (1'h0);
  reg [(3'h7):(1'h0)] reg6938 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6936 = (1'h0);
  reg [(2'h3):(1'h0)] reg6940 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6939 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6938 = (1'h0);
  reg [(3'h6):(1'h0)] reg6937 = (1'h0);
  reg [(3'h5):(1'h0)] reg6936 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6935 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6934 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6933 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6932 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6931 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6930 = (1'h0);
  reg [(5'h10):(1'h0)] reg6929 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6928 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6927 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6926 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6925 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6924 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6923 = (1'h0);
  reg [(2'h3):(1'h0)] reg6922 = (1'h0);
  reg [(2'h2):(1'h0)] reg6921 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6920 = (1'h0);
  reg [(2'h2):(1'h0)] forvar6919 = (1'h0);
  reg [(5'h10):(1'h0)] reg6918 = (1'h0);
  reg [(4'hc):(1'h0)] reg6917 = (1'h0);
  reg [(4'hf):(1'h0)] reg6916 = (1'h0);
  reg [(3'h7):(1'h0)] reg6915 = (1'h0);
  reg [(4'hb):(1'h0)] reg6914 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6913 = (1'h0);
  reg [(5'h10):(1'h0)] reg6912 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6911 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6910 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6909 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6908 = (1'h0);
  reg [(3'h7):(1'h0)] reg6907 = (1'h0);
  reg [(4'h9):(1'h0)] reg6906 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6905 = (1'h0);
  reg [(4'hc):(1'h0)] reg6904 = (1'h0);
  reg [(3'h7):(1'h0)] reg6903 = (1'h0);
  reg [(4'hc):(1'h0)] reg6902 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6901 = (1'h0);
  reg [(5'h10):(1'h0)] reg6900 = (1'h0);
  reg [(4'he):(1'h0)] forvar6899 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6898 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6898 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6897 = (1'h0);
  reg [(3'h5):(1'h0)] reg6896 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6877 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6874 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6871 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6895 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6890 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6886 = (1'h0);
  reg [(3'h4):(1'h0)] reg6885 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6894 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6893 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6892 = (1'h0);
  reg [(2'h2):(1'h0)] reg6891 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6890 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6889 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6888 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6887 = (1'h0);
  reg [(4'h9):(1'h0)] reg6886 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6885 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6882 = (1'h0);
  reg [(3'h7):(1'h0)] reg6880 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6884 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6883 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6882 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6881 = (1'h0);
  reg [(4'hb):(1'h0)] forvar6880 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6879 = (1'h0);
  reg [(4'h9):(1'h0)] reg6878 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6877 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6876 = (1'h0);
  reg [(5'h10):(1'h0)] reg6875 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6874 = (1'h0);
  reg [(3'h4):(1'h0)] reg6873 = (1'h0);
  reg [(4'hd):(1'h0)] reg6872 = (1'h0);
  reg [(4'hc):(1'h0)] reg6871 = (1'h0);
  reg [(2'h3):(1'h0)] reg6870 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6869 = (1'h0);
  reg [(5'h10):(1'h0)] reg6868 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6867 = (1'h0);
  wire signed [(3'h4):(1'h0)] wire6866;
  wire [(3'h4):(1'h0)] wire6865;
  wire signed [(4'h9):(1'h0)] wire6864;
  reg [(4'h8):(1'h0)] reg4577 = (1'h0);
  reg [(3'h7):(1'h0)] reg4578 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4579 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4580 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4581 = (1'h0);
  reg [(2'h2):(1'h0)] reg4582 = (1'h0);
  reg [(5'h10):(1'h0)] reg4583 = (1'h0);
  reg [(4'he):(1'h0)] reg4584 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4585 = (1'h0);
  reg [(4'ha):(1'h0)] reg4586 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4587 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4588 = (1'h0);
  reg [(3'h7):(1'h0)] reg4589 = (1'h0);
  reg [(4'h9):(1'h0)] reg4590 = (1'h0);
  reg [(3'h5):(1'h0)] reg4591 = (1'h0);
  reg [(4'ha):(1'h0)] reg4592 = (1'h0);
  reg [(4'hf):(1'h0)] reg4579 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4580 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4581 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4593 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4594 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4595 = (1'h0);
  reg [(3'h7):(1'h0)] reg4596 = (1'h0);
  reg [(4'hb):(1'h0)] reg4597 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4598 = (1'h0);
  reg [(4'hd):(1'h0)] reg4599 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4600 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4601 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4602 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4603 = (1'h0);
  reg [(3'h6):(1'h0)] reg4604 = (1'h0);
  reg [(5'h10):(1'h0)] reg4605 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4594 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4602 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4603 = (1'h0);
  reg [(3'h7):(1'h0)] reg4606 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4607 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4608 = (1'h0);
  reg [(4'ha):(1'h0)] reg4609 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4577 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4578 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4584 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4591 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4592 = (1'h0);
  reg [(3'h4):(1'h0)] reg4593 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4598 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4604 = (1'h0);
  reg [(4'ha):(1'h0)] reg4607 = (1'h0);
  reg [(4'he):(1'h0)] reg4608 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4610 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4611 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4612 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4613 = (1'h0);
  reg [(3'h4):(1'h0)] reg4614 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4610 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4611 = (1'h0);
  reg [(4'he):(1'h0)] forvar4613 = (1'h0);
  reg [(3'h5):(1'h0)] reg4615 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4609 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4616 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4617 = (1'h0);
  reg [(3'h5):(1'h0)] reg4618 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4619 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4620 = (1'h0);
  reg [(2'h3):(1'h0)] reg4621 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4622 = (1'h0);
  reg [(4'hd):(1'h0)] reg4623 = (1'h0);
  reg [(3'h6):(1'h0)] reg4624 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4625 = (1'h0);
  reg [(2'h2):(1'h0)] reg4626 = (1'h0);
  reg [(4'hb):(1'h0)] reg4627 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4628 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4624 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4629 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4630 = (1'h0);
  reg [(4'h9):(1'h0)] reg4631 = (1'h0);
  reg [(2'h3):(1'h0)] reg4632 = (1'h0);
  reg [(3'h4):(1'h0)] reg4633 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4634 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4635 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4636 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4637 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4638 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4636 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4639 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4640 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4641 = (1'h0);
  reg [(4'ha):(1'h0)] reg4642 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4643 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4644 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4645 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4646 = (1'h0);
  reg [(3'h6):(1'h0)] reg4647 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4648 = (1'h0);
  reg [(3'h7):(1'h0)] reg4649 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4650 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4651 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4642 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4643 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4645 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4652 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4653 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4654 = (1'h0);
  reg [(4'h8):(1'h0)] reg4655 = (1'h0);
  reg [(3'h5):(1'h0)] reg4656 = (1'h0);
  reg [(4'hf):(1'h0)] reg4657 = (1'h0);
  reg [(4'hc):(1'h0)] reg4658 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4654 = (1'h0);
  reg [(4'he):(1'h0)] forvar4656 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4659 = (1'h0);
  reg [(4'h9):(1'h0)] reg4660 = (1'h0);
  reg [(5'h10):(1'h0)] reg4661 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4662 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4663 = (1'h0);
  reg [(4'hf):(1'h0)] reg4664 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4665 = (1'h0);
  reg [(4'hb):(1'h0)] reg4666 = (1'h0);
  reg [(4'hd):(1'h0)] reg4667 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4668 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4669 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4670 = (1'h0);
  reg [(3'h4):(1'h0)] reg4671 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4672 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4673 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4674 = (1'h0);
  reg [(4'h9):(1'h0)] reg4675 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4676 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4677 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4678 = (1'h0);
  reg [(5'h10):(1'h0)] reg4679 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4680 = (1'h0);
  reg [(3'h4):(1'h0)] reg4676 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4681 = (1'h0);
  reg [(3'h5):(1'h0)] reg4682 = (1'h0);
  reg [(2'h3):(1'h0)] reg4683 = (1'h0);
  reg [(4'he):(1'h0)] reg4684 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4685 = (1'h0);
  reg [(4'h9):(1'h0)] reg4686 = (1'h0);
  reg [(4'hd):(1'h0)] reg4687 = (1'h0);
  reg [(4'hd):(1'h0)] reg4688 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4689 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4688 = (1'h0);
  reg [(4'hc):(1'h0)] reg4690 = (1'h0);
  reg [(4'ha):(1'h0)] reg4691 = (1'h0);
  reg [(4'ha):(1'h0)] reg4692 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4689 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4693 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4694 = (1'h0);
  reg [(4'ha):(1'h0)] reg4695 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4696 = (1'h0);
  reg [(3'h6):(1'h0)] reg4697 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4698 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4699 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4700 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4701 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4702 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4703 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4704 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4705 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4706 = (1'h0);
  reg [(4'hd):(1'h0)] reg4707 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4708 = (1'h0);
  reg [(5'h10):(1'h0)] reg4709 = (1'h0);
  reg [(3'h4):(1'h0)] reg4710 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4711 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4712 = (1'h0);
  reg [(4'h9):(1'h0)] reg4713 = (1'h0);
  reg [(4'h9):(1'h0)] reg4714 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4715 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4716 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4717 = (1'h0);
  reg [(4'h9):(1'h0)] reg4718 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4719 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4720 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4721 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4722 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4723 = (1'h0);
  reg [(4'hc):(1'h0)] reg4724 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4715 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4725 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4726 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4727 = (1'h0);
  reg [(4'ha):(1'h0)] reg4728 = (1'h0);
  reg [(3'h7):(1'h0)] reg4729 = (1'h0);
  reg [(4'hc):(1'h0)] reg4730 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4731 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4732 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4733 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4734 = (1'h0);
  reg [(4'h9):(1'h0)] reg4735 = (1'h0);
  reg [(2'h3):(1'h0)] reg4736 = (1'h0);
  reg [(2'h3):(1'h0)] reg4725 = (1'h0);
  reg [(3'h4):(1'h0)] reg4727 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4731 = (1'h0);
  reg [(4'hd):(1'h0)] reg4733 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4737 = (1'h0);
  reg [(2'h2):(1'h0)] reg4738 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4739 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4740 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4738 = (1'h0);
  reg [(3'h6):(1'h0)] reg4741 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4742 = (1'h0);
  reg [(4'h8):(1'h0)] reg4743 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4744 = (1'h0);
  reg [(3'h7):(1'h0)] forvar4745 = (1'h0);
  reg [(3'h6):(1'h0)] reg4746 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4747 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4748 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4749 = (1'h0);
  reg [(3'h7):(1'h0)] reg4750 = (1'h0);
  reg [(3'h4):(1'h0)] reg4751 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4752 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4753 = (1'h0);
  reg [(4'ha):(1'h0)] reg4754 = (1'h0);
  reg [(2'h2):(1'h0)] reg4755 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4756 = (1'h0);
  reg [(4'hb):(1'h0)] reg4757 = (1'h0);
  reg [(3'h6):(1'h0)] reg4758 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4759 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4760 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4761 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4762 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4763 = (1'h0);
  reg [(4'hc):(1'h0)] reg4764 = (1'h0);
  reg [(3'h6):(1'h0)] reg4765 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4766 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4758 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4759 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4763 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4767 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4768 = (1'h0);
  reg [(3'h6):(1'h0)] reg4769 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4770 = (1'h0);
  reg [(4'hd):(1'h0)] reg4771 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4772 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4773 = (1'h0);
  reg [(4'ha):(1'h0)] reg4774 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4775 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4776 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4777 = (1'h0);
  reg [(3'h5):(1'h0)] reg4778 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4745 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4746 = (1'h0);
  reg [(5'h10):(1'h0)] reg4749 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4753 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4755 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4779 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4780 = (1'h0);
  reg [(3'h6):(1'h0)] reg4781 = (1'h0);
  reg [(2'h3):(1'h0)] reg4782 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4783 = (1'h0);
  reg [(5'h10):(1'h0)] reg4784 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4785 = (1'h0);
  reg [(4'he):(1'h0)] forvar4786 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4787 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4788 = (1'h0);
  reg [(3'h7):(1'h0)] reg4789 = (1'h0);
  reg [(4'hf):(1'h0)] reg4790 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4786 = (1'h0);
  reg [(4'hd):(1'h0)] reg4791 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4792 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4793 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4794 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4795 = (1'h0);
  reg [(3'h6):(1'h0)] reg4796 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4797 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4741 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4744 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4748 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4750 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4760 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4770 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4775 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4777 = (1'h0);
  reg [(2'h2):(1'h0)] reg4779 = (1'h0);
  reg [(3'h5):(1'h0)] reg4780 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4766 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4768 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4781 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4789 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar4771 = (1'h0);
  reg [(5'h10):(1'h0)] reg4773 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire4798;
  wire signed [(2'h3):(1'h0)] wire4799;
  reg [(4'h9):(1'h0)] reg4800 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4801 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4802 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4803 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4804 = (1'h0);
  reg [(3'h6):(1'h0)] reg4805 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4806 = (1'h0);
  reg [(4'h9):(1'h0)] reg4807 = (1'h0);
  reg [(2'h3):(1'h0)] reg4808 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4809 = (1'h0);
  reg [(3'h7):(1'h0)] reg4810 = (1'h0);
  reg [(4'ha):(1'h0)] reg4811 = (1'h0);
  reg [(4'h9):(1'h0)] reg4812 = (1'h0);
  reg [(4'he):(1'h0)] forvar4813 = (1'h0);
  reg [(4'h8):(1'h0)] forvar4814 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4815 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4816 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4817 = (1'h0);
  reg [(3'h5):(1'h0)] reg4818 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4819 = (1'h0);
  reg [(4'h9):(1'h0)] reg4820 = (1'h0);
  reg [(4'hb):(1'h0)] reg4821 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4822 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4823 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4824 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4825 = (1'h0);
  reg [(2'h3):(1'h0)] forvar4826 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4827 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4828 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4829 = (1'h0);
  reg [(4'ha):(1'h0)] reg4830 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4831 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4832 = (1'h0);
  reg [(4'he):(1'h0)] reg4833 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4834 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4835 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4836 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4837 = (1'h0);
  reg [(3'h7):(1'h0)] reg4838 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4839 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4840 = (1'h0);
  reg [(5'h10):(1'h0)] reg4841 = (1'h0);
  reg [(5'h10):(1'h0)] reg4842 = (1'h0);
  reg [(4'he):(1'h0)] forvar4843 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4844 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4845 = (1'h0);
  reg [(4'hf):(1'h0)] reg4846 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4847 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4848 = (1'h0);
  reg [(3'h4):(1'h0)] reg4849 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4850 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4851 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4852 = (1'h0);
  reg [(3'h7):(1'h0)] reg4853 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4837 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4839 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4840 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4843 = (1'h0);
  reg [(4'hf):(1'h0)] reg4848 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4849 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4850 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4851 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4854 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4855 = (1'h0);
  reg [(4'hb):(1'h0)] reg4856 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4857 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4858 = (1'h0);
  reg [(4'hd):(1'h0)] reg4859 = (1'h0);
  reg [(4'hb):(1'h0)] reg4860 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4861 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg4862 = (1'h0);
  reg [(5'h10):(1'h0)] reg4863 = (1'h0);
  reg [(4'hf):(1'h0)] reg4864 = (1'h0);
  reg [(3'h4):(1'h0)] reg4865 = (1'h0);
  reg [(3'h6):(1'h0)] reg4866 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4867 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar4864 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4868 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4869 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4870 = (1'h0);
  reg [(4'h9):(1'h0)] reg4871 = (1'h0);
  reg [(2'h3):(1'h0)] reg4872 = (1'h0);
  reg [(4'hb):(1'h0)] reg4873 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4869 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar4874 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg4875 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4876 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4877 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4878 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4879 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg4880 = (1'h0);
  reg [(4'hf):(1'h0)] reg4881 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4882 = (1'h0);
  reg [(2'h3):(1'h0)] reg4883 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar4884 = (1'h0);
  reg [(2'h2):(1'h0)] reg4885 = (1'h0);
  reg [(4'hc):(1'h0)] reg4886 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4887 = (1'h0);
  reg [(2'h3):(1'h0)] reg4888 = (1'h0);
  reg [(4'hc):(1'h0)] reg4889 = (1'h0);
  reg [(4'hf):(1'h0)] reg4879 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4890 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4891 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4892 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4893 = (1'h0);
  reg [(4'hb):(1'h0)] reg4894 = (1'h0);
  reg [(2'h3):(1'h0)] reg4895 = (1'h0);
  reg [(4'h9):(1'h0)] reg4896 = (1'h0);
  reg [(4'ha):(1'h0)] reg4897 = (1'h0);
  reg [(2'h3):(1'h0)] reg4898 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4899 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4900 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4901 = (1'h0);
  reg [(5'h10):(1'h0)] reg4902 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4903 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4904 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4905 = (1'h0);
  reg [(3'h6):(1'h0)] reg4906 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4907 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4908 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4909 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4910 = (1'h0);
  reg [(3'h7):(1'h0)] reg4911 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4912 = (1'h0);
  reg [(4'hb):(1'h0)] forvar4913 = (1'h0);
  reg [(3'h6):(1'h0)] reg4914 = (1'h0);
  reg [(4'he):(1'h0)] reg4915 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4916 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4917 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4918 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4919 = (1'h0);
  reg [(4'hd):(1'h0)] reg4920 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4921 = (1'h0);
  reg [(4'hb):(1'h0)] reg4922 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar4923 = (1'h0);
  reg [(4'hc):(1'h0)] reg4924 = (1'h0);
  reg [(4'hf):(1'h0)] reg4925 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4926 = (1'h0);
  reg [(4'hc):(1'h0)] reg4927 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg4928 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4929 = (1'h0);
  reg [(4'hc):(1'h0)] reg4930 = (1'h0);
  reg [(4'h8):(1'h0)] reg4931 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4932 = (1'h0);
  reg [(4'he):(1'h0)] reg4933 = (1'h0);
  reg [(5'h10):(1'h0)] forvar4929 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4908 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4911 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4912 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar4914 = (1'h0);
  reg [(3'h7):(1'h0)] reg4918 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4920 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4931 = (1'h0);
  reg [(3'h5):(1'h0)] forvar4933 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4934 = (1'h0);
  reg [(4'he):(1'h0)] reg4935 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4936 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4937 = (1'h0);
  reg [(4'he):(1'h0)] reg4938 = (1'h0);
  reg [(4'hc):(1'h0)] reg4939 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4909 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4913 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4910 = (1'h0);
  reg [(4'ha):(1'h0)] forvar4915 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire4940;
  reg signed [(4'hd):(1'h0)] reg4941 = (1'h0);
  reg [(3'h7):(1'h0)] reg4942 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg4943 = (1'h0);
  reg [(4'hc):(1'h0)] forvar4944 = (1'h0);
  reg [(2'h2):(1'h0)] reg4945 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar4946 = (1'h0);
  reg [(4'hb):(1'h0)] reg4947 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4948 = (1'h0);
  reg [(3'h7):(1'h0)] reg4949 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4950 = (1'h0);
  reg [(4'hc):(1'h0)] reg4951 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4952 = (1'h0);
  reg [(4'ha):(1'h0)] reg4953 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4954 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4955 = (1'h0);
  reg [(3'h6):(1'h0)] reg4956 = (1'h0);
  reg [(3'h4):(1'h0)] forvar4957 = (1'h0);
  reg [(2'h2):(1'h0)] forvar4958 = (1'h0);
  reg [(4'h9):(1'h0)] reg4959 = (1'h0);
  reg [(3'h6):(1'h0)] reg4960 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4961 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4941 = (1'h0);
  reg [(4'hc):(1'h0)] reg4944 = (1'h0);
  reg [(4'hd):(1'h0)] reg4946 = (1'h0);
  reg [(4'ha):(1'h0)] reg4952 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4962 = (1'h0);
  reg [(4'h8):(1'h0)] reg4963 = (1'h0);
  reg [(4'h8):(1'h0)] reg4964 = (1'h0);
  reg [(4'ha):(1'h0)] reg4962 = (1'h0);
  reg [(4'hf):(1'h0)] forvar4965 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4966 = (1'h0);
  reg [(4'hd):(1'h0)] reg4967 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4968 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4969 = (1'h0);
  reg [(3'h6):(1'h0)] reg4970 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4971 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4972 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4973 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4974 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4975 = (1'h0);
  reg signed [(4'he):(1'h0)] reg4976 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4977 = (1'h0);
  reg [(4'h9):(1'h0)] reg4978 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4979 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar4980 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg4981 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4982 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4983 = (1'h0);
  reg [(3'h4):(1'h0)] reg4984 = (1'h0);
  reg [(3'h4):(1'h0)] reg4985 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4965 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg4966 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar4969 = (1'h0);
  reg [(4'hb):(1'h0)] reg4972 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4973 = (1'h0);
  reg [(4'he):(1'h0)] forvar4975 = (1'h0);
  reg [(3'h5):(1'h0)] reg4977 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg4980 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar4986 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4987 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4988 = (1'h0);
  reg [(4'h9):(1'h0)] reg4989 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg4990 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg4991 = (1'h0);
  reg [(2'h2):(1'h0)] reg4992 = (1'h0);
  reg [(4'hd):(1'h0)] reg4993 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg4994 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4991 = (1'h0);
  reg [(4'h9):(1'h0)] reg4995 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg4996 = (1'h0);
  reg [(3'h6):(1'h0)] reg4997 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar4998 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar4999 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5000 = (1'h0);
  reg [(5'h10):(1'h0)] reg5001 = (1'h0);
  reg [(2'h2):(1'h0)] reg5002 = (1'h0);
  reg [(2'h2):(1'h0)] reg5003 = (1'h0);
  reg [(2'h2):(1'h0)] reg5004 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5005 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar4995 = (1'h0);
  reg [(4'hd):(1'h0)] forvar4996 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg4998 = (1'h0);
  reg [(3'h4):(1'h0)] reg4999 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5001 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5006 = (1'h0);
  reg [(2'h3):(1'h0)] reg5007 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5008 = (1'h0);
  reg [(2'h3):(1'h0)] reg5009 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5010 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5009 = (1'h0);
  reg [(4'hf):(1'h0)] reg5011 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5012 = (1'h0);
  reg [(3'h5):(1'h0)] reg5013 = (1'h0);
  reg [(4'h8):(1'h0)] reg5014 = (1'h0);
  reg [(5'h10):(1'h0)] reg5015 = (1'h0);
  reg [(5'h10):(1'h0)] reg5016 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5017 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5018 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5019 = (1'h0);
  reg [(3'h6):(1'h0)] reg5020 = (1'h0);
  reg [(2'h2):(1'h0)] reg5021 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5022 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5023 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5024 = (1'h0);
  reg [(4'hc):(1'h0)] reg5025 = (1'h0);
  reg [(4'hc):(1'h0)] reg5026 = (1'h0);
  reg [(4'h8):(1'h0)] reg5027 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5028 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5029 = (1'h0);
  reg [(4'hb):(1'h0)] reg5030 = (1'h0);
  reg [(3'h6):(1'h0)] reg5031 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5032 = (1'h0);
  reg [(2'h2):(1'h0)] reg5033 = (1'h0);
  reg [(2'h3):(1'h0)] reg5034 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5029 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4970 = (1'h0);
  reg [(3'h6):(1'h0)] forvar4974 = (1'h0);
  reg [(3'h6):(1'h0)] reg4986 = (1'h0);
  reg [(4'h9):(1'h0)] forvar4967 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg4988 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar4989 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5003 = (1'h0);
  reg [(3'h6):(1'h0)] reg5006 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5002 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5005 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5008 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5011 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5015 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5019 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5020 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5035 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5036 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5037 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5038 = (1'h0);
  reg [(4'h8):(1'h0)] reg5039 = (1'h0);
  reg [(2'h2):(1'h0)] reg5040 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5035 = (1'h0);
  reg [(3'h7):(1'h0)] reg5036 = (1'h0);
  reg [(4'hc):(1'h0)] reg5041 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5042 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5043 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5044 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5045 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5046 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5047 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5048 = (1'h0);
  reg [(3'h5):(1'h0)] reg5049 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5050 = (1'h0);
  reg [(4'hc):(1'h0)] reg5051 = (1'h0);
  reg [(4'hc):(1'h0)] reg5052 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5053 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5054 = (1'h0);
  reg [(4'hf):(1'h0)] reg5055 = (1'h0);
  reg [(3'h7):(1'h0)] reg5056 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5057 = (1'h0);
  reg [(4'ha):(1'h0)] reg5058 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5059 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5060 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5061 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5062 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5063 = (1'h0);
  reg [(4'he):(1'h0)] forvar5064 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5065 = (1'h0);
  reg [(4'hc):(1'h0)] reg5066 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5067 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5068 = (1'h0);
  reg [(4'hc):(1'h0)] reg5069 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5070 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5071 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5072 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5073 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5074 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5075 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5076 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5077 = (1'h0);
  reg [(3'h4):(1'h0)] reg5078 = (1'h0);
  reg [(4'hc):(1'h0)] reg5079 = (1'h0);
  reg [(4'he):(1'h0)] reg5080 = (1'h0);
  reg [(3'h7):(1'h0)] reg5081 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5039 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5043 = (1'h0);
  reg [(3'h4):(1'h0)] reg5048 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5049 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5054 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5059 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5051 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5053 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5082 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5083 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5084 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5085 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5086 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5087 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5088 = (1'h0);
  reg [(3'h5):(1'h0)] reg5089 = (1'h0);
  reg [(4'h9):(1'h0)] reg5090 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5091 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5092 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5089 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5093 = (1'h0);
  reg [(5'h10):(1'h0)] reg5094 = (1'h0);
  reg [(4'h8):(1'h0)] reg5095 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5096 = (1'h0);
  reg [(4'hf):(1'h0)] reg5097 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5098 = (1'h0);
  reg [(3'h5):(1'h0)] reg5099 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5100 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5101 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5102 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5103 = (1'h0);
  reg [(4'h8):(1'h0)] reg5104 = (1'h0);
  reg [(3'h7):(1'h0)] reg5105 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5082 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5083 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5084 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5088 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5090 = (1'h0);
  reg [(4'hf):(1'h0)] reg5093 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5106 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5107 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5108 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5109 = (1'h0);
  reg [(4'h9):(1'h0)] reg5110 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5111 = (1'h0);
  reg [(5'h10):(1'h0)] reg5112 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5085 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5091 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5104 = (1'h0);
  reg [(3'h7):(1'h0)] reg5106 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5108 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5113 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5114 = (1'h0);
  reg [(4'he):(1'h0)] reg5115 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5116 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5117 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5117 = (1'h0);
  reg [(2'h3):(1'h0)] reg5118 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5119 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5120 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5111 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5121 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5122 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5123 = (1'h0);
  reg [(3'h5):(1'h0)] reg5124 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5125 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5126 = (1'h0);
  reg [(3'h7):(1'h0)] reg5127 = (1'h0);
  reg [(2'h3):(1'h0)] reg5128 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5129 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5130 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5130 = (1'h0);
  reg [(4'he):(1'h0)] reg5131 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5132 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5133 = (1'h0);
  reg [(4'hf):(1'h0)] reg5134 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5135 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5136 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5137 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5138 = (1'h0);
  reg [(4'hb):(1'h0)] reg5139 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5140 = (1'h0);
  reg [(4'hc):(1'h0)] reg5141 = (1'h0);
  reg [(4'h8):(1'h0)] reg5142 = (1'h0);
  reg [(4'ha):(1'h0)] reg5143 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5144 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5145 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5138 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5143 = (1'h0);
  reg [(3'h4):(1'h0)] reg5146 = (1'h0);
  reg [(4'h8):(1'h0)] reg5147 = (1'h0);
  reg [(4'he):(1'h0)] reg5148 = (1'h0);
  reg [(3'h7):(1'h0)] reg5149 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5150 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5151 = (1'h0);
  reg [(5'h10):(1'h0)] reg5152 = (1'h0);
  reg [(3'h4):(1'h0)] reg5153 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5149 = (1'h0);
  reg [(5'h10):(1'h0)] reg5150 = (1'h0);
  reg [(2'h3):(1'h0)] reg5154 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5155 = (1'h0);
  reg [(5'h10):(1'h0)] reg5156 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5157 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5158 = (1'h0);
  reg [(3'h7):(1'h0)] reg5159 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5160 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5161 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5162 = (1'h0);
  reg [(4'hb):(1'h0)] reg5163 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5164 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5165 = (1'h0);
  reg [(4'he):(1'h0)] forvar5166 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5167 = (1'h0);
  reg [(4'hd):(1'h0)] reg5168 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5169 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5170 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5171 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5172 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5173 = (1'h0);
  reg [(5'h10):(1'h0)] reg5174 = (1'h0);
  reg [(4'he):(1'h0)] forvar5175 = (1'h0);
  reg [(2'h3):(1'h0)] reg5176 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5178 = (1'h0);
  reg [(4'h8):(1'h0)] reg5179 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5180 = (1'h0);
  reg [(3'h4):(1'h0)] reg5181 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5182 = (1'h0);
  reg [(4'he):(1'h0)] reg5183 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5184 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5185 = (1'h0);
  reg [(4'hd):(1'h0)] reg5186 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5187 = (1'h0);
  reg [(4'hc):(1'h0)] reg5188 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5189 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5190 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5191 = (1'h0);
  reg [(2'h2):(1'h0)] reg5192 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5185 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5186 = (1'h0);
  reg [(5'h10):(1'h0)] reg5187 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5189 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5193 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5194 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5148 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire5195;
  wire [(3'h7):(1'h0)] wire5196;
  wire signed [(5'h10):(1'h0)] wire5197;
  reg [(4'ha):(1'h0)] forvar5198 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5199 = (1'h0);
  reg [(4'hb):(1'h0)] reg5200 = (1'h0);
  reg [(4'hc):(1'h0)] reg5201 = (1'h0);
  reg [(4'hc):(1'h0)] reg5202 = (1'h0);
  reg [(4'hf):(1'h0)] reg5199 = (1'h0);
  reg [(3'h6):(1'h0)] reg5203 = (1'h0);
  reg [(3'h4):(1'h0)] reg5204 = (1'h0);
  reg [(4'h9):(1'h0)] reg5205 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5206 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5207 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5208 = (1'h0);
  reg [(4'h9):(1'h0)] reg5209 = (1'h0);
  reg [(3'h4):(1'h0)] reg5210 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5211 = (1'h0);
  reg [(4'hd):(1'h0)] reg5206 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5208 = (1'h0);
  reg [(4'hf):(1'h0)] reg5212 = (1'h0);
  reg [(4'hb):(1'h0)] reg5213 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5214 = (1'h0);
  reg [(4'h8):(1'h0)] reg5215 = (1'h0);
  reg [(4'hf):(1'h0)] reg5216 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5217 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5218 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5219 = (1'h0);
  reg [(3'h7):(1'h0)] reg5220 = (1'h0);
  reg [(4'h9):(1'h0)] reg5221 = (1'h0);
  reg [(4'hb):(1'h0)] reg5222 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5223 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5224 = (1'h0);
  reg [(5'h10):(1'h0)] reg5225 = (1'h0);
  reg [(5'h10):(1'h0)] reg5226 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5200 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5227 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5228 = (1'h0);
  reg [(4'hc):(1'h0)] reg5229 = (1'h0);
  reg [(3'h7):(1'h0)] reg5230 = (1'h0);
  reg [(4'hb):(1'h0)] reg5231 = (1'h0);
  reg [(3'h6):(1'h0)] reg5232 = (1'h0);
  reg [(4'he):(1'h0)] reg5233 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5234 = (1'h0);
  reg [(3'h7):(1'h0)] reg5235 = (1'h0);
  reg [(3'h4):(1'h0)] reg5236 = (1'h0);
  reg [(4'hd):(1'h0)] reg5237 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5238 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5239 = (1'h0);
  reg [(5'h10):(1'h0)] reg5240 = (1'h0);
  reg [(5'h10):(1'h0)] reg5241 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5242 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5234 = (1'h0);
  reg [(5'h10):(1'h0)] reg5228 = (1'h0);
  reg [(3'h6):(1'h0)] reg5243 = (1'h0);
  reg [(3'h5):(1'h0)] reg5244 = (1'h0);
  reg [(4'h9):(1'h0)] reg5245 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5245 = (1'h0);
  reg [(3'h5):(1'h0)] reg5246 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5247 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5248 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5249 = (1'h0);
  reg [(4'ha):(1'h0)] reg5250 = (1'h0);
  reg [(4'ha):(1'h0)] reg5251 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5252 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5253 = (1'h0);
  reg [(4'ha):(1'h0)] reg5254 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5243 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5247 = (1'h0);
  reg [(4'he):(1'h0)] reg5248 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5252 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5255 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5256 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5257 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5258 = (1'h0);
  reg [(4'hd):(1'h0)] reg5259 = (1'h0);
  reg [(4'h9):(1'h0)] reg5260 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5261 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5262 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5263 = (1'h0);
  reg [(3'h4):(1'h0)] reg5264 = (1'h0);
  reg [(4'hb):(1'h0)] reg5265 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5266 = (1'h0);
  reg [(4'he):(1'h0)] reg5267 = (1'h0);
  reg [(3'h4):(1'h0)] reg5268 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5269 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5229 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5231 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5238 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5270 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5271 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5272 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5273 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5274 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5275 = (1'h0);
  reg [(4'hd):(1'h0)] reg5276 = (1'h0);
  reg [(4'he):(1'h0)] reg5277 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5278 = (1'h0);
  reg [(4'h9):(1'h0)] reg5279 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5280 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5281 = (1'h0);
  reg [(3'h7):(1'h0)] reg5282 = (1'h0);
  reg [(4'he):(1'h0)] reg5283 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5284 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5285 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5286 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5287 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5288 = (1'h0);
  reg [(2'h2):(1'h0)] reg5289 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5290 = (1'h0);
  reg [(4'h8):(1'h0)] reg5291 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5292 = (1'h0);
  reg [(4'he):(1'h0)] reg5293 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5294 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5295 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5296 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5297 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5298 = (1'h0);
  reg [(3'h6):(1'h0)] reg5299 = (1'h0);
  reg [(2'h3):(1'h0)] reg5300 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5292 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5297 = (1'h0);
  reg [(4'h8):(1'h0)] reg5298 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5301 = (1'h0);
  reg [(2'h3):(1'h0)] reg5302 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5272 = (1'h0);
  reg [(4'he):(1'h0)] reg5274 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5277 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5280 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5281 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5284 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5285 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5301 = (1'h0);
  reg [(3'h4):(1'h0)] reg5303 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5304 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5305 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5302 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5306 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5307 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5308 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5309 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5310 = (1'h0);
  reg [(4'h8):(1'h0)] reg5311 = (1'h0);
  reg [(4'ha):(1'h0)] reg5312 = (1'h0);
  reg [(4'hb):(1'h0)] reg5313 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5314 = (1'h0);
  reg [(4'hd):(1'h0)] reg5315 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5316 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5317 = (1'h0);
  reg [(4'he):(1'h0)] reg5318 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5319 = (1'h0);
  reg [(3'h7):(1'h0)] reg5320 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5321 = (1'h0);
  reg [(4'h9):(1'h0)] reg5322 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5314 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5323 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5324 = (1'h0);
  reg [(4'h9):(1'h0)] reg5325 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5326 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5327 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5328 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5329 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5331 = (1'h0);
  reg [(4'h9):(1'h0)] reg5332 = (1'h0);
  reg [(2'h2):(1'h0)] reg5333 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5334 = (1'h0);
  reg [(2'h3):(1'h0)] reg5335 = (1'h0);
  reg [(4'hf):(1'h0)] reg5336 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5337 = (1'h0);
  reg [(2'h3):(1'h0)] reg5338 = (1'h0);
  reg [(2'h2):(1'h0)] reg5339 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5340 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5341 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5342 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5343 = (1'h0);
  reg [(4'h9):(1'h0)] reg5344 = (1'h0);
  reg [(4'hc):(1'h0)] reg5345 = (1'h0);
  reg [(2'h2):(1'h0)] reg5346 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5347 = (1'h0);
  reg [(4'hb):(1'h0)] reg5348 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5349 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5350 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5351 = (1'h0);
  reg [(4'hf):(1'h0)] reg5352 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5353 = (1'h0);
  reg [(4'hc):(1'h0)] reg5354 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5355 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5356 = (1'h0);
  reg [(4'hb):(1'h0)] reg5357 = (1'h0);
  reg [(4'he):(1'h0)] reg5358 = (1'h0);
  reg [(5'h10):(1'h0)] reg5359 = (1'h0);
  reg [(4'hd):(1'h0)] reg5360 = (1'h0);
  reg [(5'h10):(1'h0)] reg5361 = (1'h0);
  reg [(3'h4):(1'h0)] reg5362 = (1'h0);
  reg [(4'he):(1'h0)] reg5355 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5363 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5364 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5365 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5366 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5367 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5368 = (1'h0);
  reg [(3'h4):(1'h0)] reg5369 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5370 = (1'h0);
  reg [(4'hf):(1'h0)] reg5371 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5372 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5373 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5374 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5375 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5376 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5377 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5378 = (1'h0);
  reg [(3'h5):(1'h0)] reg5379 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5380 = (1'h0);
  reg [(5'h10):(1'h0)] reg5381 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5382 = (1'h0);
  reg [(4'hd):(1'h0)] reg5383 = (1'h0);
  reg [(4'he):(1'h0)] reg5384 = (1'h0);
  reg [(5'h10):(1'h0)] reg5385 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5376 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5377 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5380 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5386 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5382 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5387 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar5388 = (1'h0);
  reg [(4'h9):(1'h0)] reg5389 = (1'h0);
  reg [(2'h2):(1'h0)] reg5390 = (1'h0);
  reg [(3'h4):(1'h0)] reg5391 = (1'h0);
  reg [(3'h4):(1'h0)] reg5392 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5393 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5394 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5395 = (1'h0);
  reg [(4'he):(1'h0)] reg5396 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5397 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5398 = (1'h0);
  reg [(3'h5):(1'h0)] reg5399 = (1'h0);
  reg [(4'hb):(1'h0)] reg5400 = (1'h0);
  reg [(4'hb):(1'h0)] reg5401 = (1'h0);
  reg [(4'h9):(1'h0)] reg5402 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5403 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5404 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5405 = (1'h0);
  reg [(2'h2):(1'h0)] reg5406 = (1'h0);
  reg [(4'hd):(1'h0)] reg5407 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5408 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5409 = (1'h0);
  reg [(4'hb):(1'h0)] reg5410 = (1'h0);
  reg [(4'he):(1'h0)] reg5411 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5412 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5413 = (1'h0);
  reg [(4'ha):(1'h0)] reg5414 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5415 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5416 = (1'h0);
  reg [(3'h7):(1'h0)] reg5417 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5418 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5419 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5420 = (1'h0);
  reg [(4'h8):(1'h0)] reg5421 = (1'h0);
  reg [(4'he):(1'h0)] reg5422 = (1'h0);
  reg [(2'h3):(1'h0)] reg5423 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5424 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5425 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5426 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5427 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5423 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5427 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5428 = (1'h0);
  reg [(4'hd):(1'h0)] reg5429 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5430 = (1'h0);
  reg [(2'h3):(1'h0)] reg5431 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5432 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5433 = (1'h0);
  reg [(3'h7):(1'h0)] reg5434 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5435 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5436 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5437 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5438 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5439 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5440 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5441 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5442 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5443 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5444 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5445 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5446 = (1'h0);
  reg [(2'h3):(1'h0)] reg5447 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5448 = (1'h0);
  reg [(4'hd):(1'h0)] reg5449 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5450 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5451 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5452 = (1'h0);
  reg [(4'ha):(1'h0)] reg5350 = (1'h0);
  reg [(4'hf):(1'h0)] reg5349 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5353 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5360 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5362 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5363 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5364 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5366 = (1'h0);
  reg [(4'h9):(1'h0)] reg5368 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5370 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5372 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5369 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5375 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5378 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5379 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5383 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5388 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5391 = (1'h0);
  reg [(4'hc):(1'h0)] reg5393 = (1'h0);
  reg [(2'h2):(1'h0)] reg5395 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5373 = (1'h0);
  reg [(4'he):(1'h0)] forvar5396 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5398 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5453 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5454 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5455 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5456 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5457 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5458 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5459 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5460 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5461 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5462 = (1'h0);
  reg [(4'hc):(1'h0)] reg5463 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5464 = (1'h0);
  reg [(4'h9):(1'h0)] reg5465 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5466 = (1'h0);
  reg [(4'h8):(1'h0)] reg5467 = (1'h0);
  reg [(2'h3):(1'h0)] reg5468 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5466 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5467 = (1'h0);
  reg [(2'h2):(1'h0)] reg5469 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5470 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5471 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5472 = (1'h0);
  reg [(4'hb):(1'h0)] reg5473 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5474 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5475 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5476 = (1'h0);
  reg [(2'h3):(1'h0)] reg5477 = (1'h0);
  reg [(4'h8):(1'h0)] reg5478 = (1'h0);
  reg [(4'hc):(1'h0)] reg5479 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5480 = (1'h0);
  reg [(2'h3):(1'h0)] reg5481 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5482 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5483 = (1'h0);
  reg [(4'hb):(1'h0)] reg5484 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5485 = (1'h0);
  reg [(4'h8):(1'h0)] reg5486 = (1'h0);
  reg [(4'h8):(1'h0)] reg5487 = (1'h0);
  reg [(2'h3):(1'h0)] reg5488 = (1'h0);
  reg [(2'h3):(1'h0)] reg5489 = (1'h0);
  reg [(4'h8):(1'h0)] reg5490 = (1'h0);
  reg [(3'h7):(1'h0)] reg5491 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5492 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5480 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5484 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5493 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5494 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5495 = (1'h0);
  reg [(3'h6):(1'h0)] reg5496 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5497 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5498 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5499 = (1'h0);
  reg [(3'h4):(1'h0)] reg5500 = (1'h0);
  reg [(4'he):(1'h0)] reg5501 = (1'h0);
  reg [(3'h4):(1'h0)] reg5502 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5503 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5504 = (1'h0);
  wire [(4'h9):(1'h0)] wire6862;
  assign y = {reg7004,
                 reg7003,
                 reg7002,
                 reg7001,
                 reg7000,
                 reg6999,
                 reg6998,
                 forvar6997,
                 reg6996,
                 reg6995,
                 reg6994,
                 reg6993,
                 reg6992,
                 reg6991,
                 reg6990,
                 reg6989,
                 reg6988,
                 reg6987,
                 reg6986,
                 forvar6985,
                 reg6984,
                 reg6983,
                 reg6982,
                 reg6981,
                 reg6980,
                 reg6979,
                 reg6978,
                 forvar6977,
                 reg6976,
                 reg6975,
                 reg6974,
                 reg6973,
                 forvar6972,
                 forvar6971,
                 reg6970,
                 reg6969,
                 reg6968,
                 reg6967,
                 forvar6966,
                 reg6965,
                 forvar6964,
                 reg6963,
                 reg6962,
                 reg6961,
                 reg6960,
                 reg6959,
                 forvar6958,
                 reg6957,
                 reg6956,
                 reg6955,
                 forvar6954,
                 forvar6953,
                 forvar6952,
                 reg6951,
                 reg6944,
                 reg6950,
                 reg6949,
                 reg6948,
                 reg6947,
                 reg6946,
                 reg6945,
                 forvar6944,
                 reg6943,
                 reg6942,
                 reg6941,
                 reg6938,
                 forvar6936,
                 reg6940,
                 reg6939,
                 forvar6938,
                 reg6937,
                 reg6936,
                 reg6935,
                 forvar6934,
                 reg6933,
                 forvar6932,
                 reg6931,
                 reg6930,
                 reg6929,
                 forvar6928,
                 reg6927,
                 reg6926,
                 forvar6925,
                 reg6924,
                 reg6923,
                 reg6922,
                 reg6921,
                 forvar6920,
                 forvar6919,
                 reg6918,
                 reg6917,
                 reg6916,
                 reg6915,
                 reg6914,
                 forvar6913,
                 reg6912,
                 reg6911,
                 forvar6910,
                 forvar6909,
                 reg6908,
                 reg6907,
                 reg6906,
                 forvar6905,
                 reg6904,
                 reg6903,
                 reg6902,
                 reg6901,
                 reg6900,
                 forvar6899,
                 forvar6898,
                 reg6898,
                 forvar6897,
                 reg6896,
                 forvar6877,
                 reg6874,
                 forvar6871,
                 reg6895,
                 forvar6890,
                 forvar6886,
                 reg6885,
                 reg6894,
                 reg6893,
                 forvar6892,
                 reg6891,
                 reg6890,
                 reg6889,
                 reg6888,
                 reg6887,
                 reg6886,
                 forvar6885,
                 reg6882,
                 reg6880,
                 reg6884,
                 reg6883,
                 forvar6882,
                 reg6881,
                 forvar6880,
                 reg6879,
                 reg6878,
                 reg6877,
                 reg6876,
                 reg6875,
                 forvar6874,
                 reg6873,
                 reg6872,
                 reg6871,
                 reg6870,
                 forvar6869,
                 reg6868,
                 forvar6867,
                 wire6866,
                 wire6865,
                 wire6864,
                 reg4577,
                 reg4578,
                 forvar4579,
                 reg4580,
                 reg4581,
                 reg4582,
                 reg4583,
                 reg4584,
                 reg4585,
                 reg4586,
                 reg4587,
                 forvar4588,
                 reg4589,
                 reg4590,
                 reg4591,
                 reg4592,
                 reg4579,
                 forvar4580,
                 forvar4581,
                 forvar4593,
                 forvar4594,
                 reg4595,
                 reg4596,
                 reg4597,
                 reg4598,
                 reg4599,
                 reg4600,
                 reg4601,
                 forvar4602,
                 reg4603,
                 reg4604,
                 reg4605,
                 reg4594,
                 reg4602,
                 forvar4603,
                 reg4606,
                 forvar4607,
                 forvar4608,
                 reg4609,
                 forvar4577,
                 forvar4578,
                 forvar4584,
                 forvar4591,
                 forvar4592,
                 reg4593,
                 forvar4598,
                 forvar4604,
                 reg4607,
                 reg4608,
                 reg4610,
                 forvar4611,
                 reg4612,
                 reg4613,
                 reg4614,
                 forvar4610,
                 reg4611,
                 forvar4613,
                 reg4615,
                 forvar4609,
                 forvar4616,
                 forvar4617,
                 reg4618,
                 reg4619,
                 reg4620,
                 reg4621,
                 reg4622,
                 reg4623,
                 reg4624,
                 reg4625,
                 reg4626,
                 reg4627,
                 reg4628,
                 forvar4624,
                 reg4629,
                 reg4630,
                 reg4631,
                 reg4632,
                 reg4633,
                 reg4634,
                 reg4635,
                 reg4636,
                 reg4637,
                 reg4638,
                 forvar4636,
                 reg4639,
                 forvar4640,
                 reg4641,
                 reg4642,
                 forvar4643,
                 reg4644,
                 reg4645,
                 reg4646,
                 reg4647,
                 forvar4648,
                 reg4649,
                 forvar4650,
                 reg4651,
                 forvar4642,
                 reg4643,
                 forvar4645,
                 forvar4652,
                 forvar4653,
                 reg4654,
                 reg4655,
                 reg4656,
                 reg4657,
                 reg4658,
                 forvar4654,
                 forvar4656,
                 forvar4659,
                 reg4660,
                 reg4661,
                 reg4662,
                 forvar4663,
                 reg4664,
                 reg4665,
                 reg4666,
                 reg4667,
                 reg4668,
                 reg4669,
                 reg4670,
                 reg4671,
                 forvar4672,
                 forvar4673,
                 forvar4674,
                 reg4675,
                 forvar4676,
                 reg4677,
                 reg4678,
                 reg4679,
                 reg4680,
                 reg4676,
                 forvar4681,
                 reg4682,
                 reg4683,
                 reg4684,
                 reg4685,
                 reg4686,
                 reg4687,
                 reg4688,
                 reg4689,
                 forvar4688,
                 reg4690,
                 reg4691,
                 reg4692,
                 forvar4689,
                 reg4693,
                 forvar4694,
                 reg4695,
                 forvar4696,
                 reg4697,
                 forvar4698,
                 reg4699,
                 reg4700,
                 reg4701,
                 reg4702,
                 reg4703,
                 reg4704,
                 forvar4705,
                 reg4706,
                 reg4707,
                 reg4708,
                 reg4709,
                 reg4710,
                 reg4711,
                 forvar4712,
                 reg4713,
                 reg4714,
                 forvar4715,
                 reg4716,
                 forvar4717,
                 reg4718,
                 reg4719,
                 reg4720,
                 reg4721,
                 reg4722,
                 reg4723,
                 reg4724,
                 reg4715,
                 forvar4725,
                 reg4726,
                 forvar4727,
                 reg4728,
                 reg4729,
                 reg4730,
                 reg4731,
                 reg4732,
                 forvar4733,
                 reg4734,
                 reg4735,
                 reg4736,
                 reg4725,
                 reg4727,
                 forvar4731,
                 reg4733,
                 forvar4737,
                 reg4738,
                 reg4739,
                 reg4740,
                 forvar4738,
                 reg4741,
                 reg4742,
                 reg4743,
                 reg4744,
                 forvar4745,
                 reg4746,
                 reg4747,
                 reg4748,
                 forvar4749,
                 reg4750,
                 reg4751,
                 reg4752,
                 reg4753,
                 reg4754,
                 reg4755,
                 reg4756,
                 reg4757,
                 reg4758,
                 forvar4759,
                 reg4760,
                 reg4761,
                 reg4762,
                 forvar4763,
                 reg4764,
                 reg4765,
                 reg4766,
                 forvar4758,
                 reg4759,
                 reg4763,
                 reg4767,
                 reg4768,
                 reg4769,
                 forvar4770,
                 reg4771,
                 reg4772,
                 forvar4773,
                 reg4774,
                 forvar4775,
                 reg4776,
                 reg4777,
                 reg4778,
                 reg4745,
                 forvar4746,
                 reg4749,
                 forvar4753,
                 forvar4755,
                 forvar4779,
                 forvar4780,
                 reg4781,
                 reg4782,
                 reg4783,
                 reg4784,
                 forvar4785,
                 forvar4786,
                 reg4787,
                 reg4788,
                 reg4789,
                 reg4790,
                 reg4786,
                 reg4791,
                 reg4792,
                 reg4793,
                 reg4794,
                 forvar4795,
                 reg4796,
                 reg4797,
                 forvar4741,
                 forvar4744,
                 forvar4748,
                 forvar4750,
                 forvar4760,
                 reg4770,
                 reg4775,
                 forvar4777,
                 reg4779,
                 reg4780,
                 forvar4766,
                 forvar4768,
                 forvar4781,
                 forvar4789,
                 forvar4771,
                 reg4773,
                 wire4798,
                 wire4799,
                 reg4800,
                 forvar4801,
                 forvar4802,
                 reg4803,
                 reg4804,
                 reg4805,
                 forvar4806,
                 reg4807,
                 reg4808,
                 forvar4809,
                 reg4810,
                 reg4811,
                 reg4812,
                 forvar4813,
                 forvar4814,
                 forvar4815,
                 reg4816,
                 forvar4817,
                 reg4818,
                 forvar4819,
                 reg4820,
                 reg4821,
                 reg4822,
                 reg4823,
                 forvar4824,
                 reg4825,
                 forvar4826,
                 forvar4827,
                 reg4828,
                 forvar4829,
                 reg4830,
                 reg4831,
                 reg4832,
                 reg4833,
                 reg4834,
                 reg4835,
                 reg4836,
                 reg4837,
                 reg4838,
                 forvar4839,
                 reg4840,
                 reg4841,
                 reg4842,
                 forvar4843,
                 reg4844,
                 reg4845,
                 reg4846,
                 reg4847,
                 forvar4848,
                 reg4849,
                 forvar4850,
                 forvar4851,
                 reg4852,
                 reg4853,
                 forvar4837,
                 reg4839,
                 forvar4840,
                 reg4843,
                 reg4848,
                 forvar4849,
                 reg4850,
                 reg4851,
                 reg4854,
                 reg4855,
                 reg4856,
                 reg4857,
                 forvar4858,
                 reg4859,
                 reg4860,
                 reg4861,
                 reg4862,
                 reg4863,
                 reg4864,
                 reg4865,
                 reg4866,
                 reg4867,
                 forvar4864,
                 reg4868,
                 forvar4869,
                 reg4870,
                 reg4871,
                 reg4872,
                 reg4873,
                 reg4869,
                 forvar4874,
                 reg4875,
                 forvar4876,
                 forvar4877,
                 reg4878,
                 forvar4879,
                 reg4880,
                 reg4881,
                 reg4882,
                 reg4883,
                 forvar4884,
                 reg4885,
                 reg4886,
                 reg4887,
                 reg4888,
                 reg4889,
                 reg4879,
                 forvar4890,
                 reg4891,
                 reg4892,
                 reg4893,
                 reg4894,
                 reg4895,
                 reg4896,
                 reg4897,
                 reg4898,
                 forvar4899,
                 reg4900,
                 reg4901,
                 reg4902,
                 reg4903,
                 reg4904,
                 reg4905,
                 reg4906,
                 reg4907,
                 forvar4908,
                 forvar4909,
                 reg4910,
                 reg4911,
                 forvar4912,
                 forvar4913,
                 reg4914,
                 reg4915,
                 reg4916,
                 reg4917,
                 forvar4918,
                 reg4919,
                 reg4920,
                 reg4921,
                 reg4922,
                 forvar4923,
                 reg4924,
                 reg4925,
                 reg4926,
                 reg4927,
                 reg4928,
                 reg4929,
                 reg4930,
                 reg4931,
                 reg4932,
                 reg4933,
                 forvar4929,
                 reg4908,
                 forvar4911,
                 reg4912,
                 forvar4914,
                 reg4918,
                 forvar4920,
                 forvar4931,
                 forvar4933,
                 reg4934,
                 reg4935,
                 reg4936,
                 reg4937,
                 reg4938,
                 reg4939,
                 reg4909,
                 reg4913,
                 forvar4910,
                 forvar4915,
                 wire4940,
                 reg4941,
                 reg4942,
                 reg4943,
                 forvar4944,
                 reg4945,
                 forvar4946,
                 reg4947,
                 reg4948,
                 reg4949,
                 reg4950,
                 reg4951,
                 forvar4952,
                 reg4953,
                 reg4954,
                 reg4955,
                 reg4956,
                 forvar4957,
                 forvar4958,
                 reg4959,
                 reg4960,
                 reg4961,
                 forvar4941,
                 reg4944,
                 reg4946,
                 reg4952,
                 forvar4962,
                 reg4963,
                 reg4964,
                 reg4962,
                 forvar4965,
                 forvar4966,
                 reg4967,
                 reg4968,
                 reg4969,
                 reg4970,
                 reg4971,
                 forvar4972,
                 reg4973,
                 reg4974,
                 reg4975,
                 reg4976,
                 forvar4977,
                 reg4978,
                 reg4979,
                 forvar4980,
                 reg4981,
                 reg4982,
                 reg4983,
                 reg4984,
                 reg4985,
                 reg4965,
                 reg4966,
                 forvar4969,
                 reg4972,
                 forvar4973,
                 forvar4975,
                 reg4977,
                 reg4980,
                 forvar4986,
                 reg4987,
                 forvar4988,
                 reg4989,
                 reg4990,
                 reg4991,
                 reg4992,
                 reg4993,
                 reg4994,
                 forvar4991,
                 reg4995,
                 reg4996,
                 reg4997,
                 forvar4998,
                 forvar4999,
                 reg5000,
                 reg5001,
                 reg5002,
                 reg5003,
                 reg5004,
                 reg5005,
                 forvar4995,
                 forvar4996,
                 reg4998,
                 reg4999,
                 forvar5001,
                 forvar5006,
                 reg5007,
                 reg5008,
                 reg5009,
                 reg5010,
                 forvar5009,
                 reg5011,
                 reg5012,
                 reg5013,
                 reg5014,
                 reg5015,
                 reg5016,
                 reg5017,
                 reg5018,
                 forvar5019,
                 reg5020,
                 reg5021,
                 reg5022,
                 reg5023,
                 reg5024,
                 reg5025,
                 reg5026,
                 reg5027,
                 reg5028,
                 forvar5029,
                 reg5030,
                 reg5031,
                 reg5032,
                 reg5033,
                 reg5034,
                 reg5029,
                 forvar4970,
                 forvar4974,
                 reg4986,
                 forvar4967,
                 reg4988,
                 forvar4989,
                 forvar5003,
                 reg5006,
                 forvar5002,
                 forvar5005,
                 forvar5008,
                 forvar5011,
                 forvar5015,
                 reg5019,
                 forvar5020,
                 reg5035,
                 forvar5036,
                 reg5037,
                 reg5038,
                 reg5039,
                 reg5040,
                 forvar5035,
                 reg5036,
                 reg5041,
                 reg5042,
                 reg5043,
                 reg5044,
                 reg5045,
                 reg5046,
                 reg5047,
                 forvar5048,
                 reg5049,
                 reg5050,
                 reg5051,
                 reg5052,
                 forvar5053,
                 forvar5054,
                 reg5055,
                 reg5056,
                 reg5057,
                 reg5058,
                 forvar5059,
                 reg5060,
                 reg5061,
                 forvar5062,
                 forvar5063,
                 forvar5064,
                 reg5065,
                 reg5066,
                 reg5067,
                 forvar5068,
                 reg5069,
                 reg5070,
                 reg5071,
                 reg5072,
                 reg5073,
                 reg5074,
                 forvar5075,
                 forvar5076,
                 reg5077,
                 reg5078,
                 reg5079,
                 reg5080,
                 reg5081,
                 forvar5039,
                 forvar5043,
                 reg5048,
                 forvar5049,
                 reg5054,
                 reg5059,
                 forvar5051,
                 reg5053,
                 forvar5082,
                 reg5083,
                 forvar5084,
                 reg5085,
                 reg5086,
                 reg5087,
                 reg5088,
                 reg5089,
                 reg5090,
                 reg5091,
                 reg5092,
                 forvar5089,
                 forvar5093,
                 reg5094,
                 reg5095,
                 reg5096,
                 reg5097,
                 forvar5098,
                 reg5099,
                 reg5100,
                 reg5101,
                 forvar5102,
                 reg5103,
                 reg5104,
                 reg5105,
                 reg5082,
                 forvar5083,
                 reg5084,
                 forvar5088,
                 forvar5090,
                 reg5093,
                 forvar5106,
                 reg5107,
                 forvar5108,
                 forvar5109,
                 reg5110,
                 reg5111,
                 reg5112,
                 forvar5085,
                 forvar5091,
                 forvar5104,
                 reg5106,
                 reg5108,
                 reg5113,
                 forvar5114,
                 reg5115,
                 reg5116,
                 reg5117,
                 forvar5117,
                 reg5118,
                 reg5119,
                 reg5120,
                 forvar5111,
                 reg5114,
                 reg5121,
                 reg5122,
                 reg5123,
                 reg5124,
                 reg5125,
                 forvar5126,
                 reg5127,
                 reg5128,
                 reg5129,
                 reg5130,
                 forvar5130,
                 reg5131,
                 reg5132,
                 reg5133,
                 reg5134,
                 forvar5135,
                 reg5136,
                 reg5137,
                 forvar5138,
                 reg5139,
                 reg5140,
                 reg5141,
                 reg5142,
                 reg5143,
                 reg5144,
                 reg5145,
                 reg5138,
                 forvar5143,
                 reg5146,
                 reg5147,
                 reg5148,
                 reg5149,
                 forvar5150,
                 reg5151,
                 reg5152,
                 reg5153,
                 forvar5149,
                 reg5150,
                 reg5154,
                 reg5155,
                 reg5156,
                 forvar5157,
                 reg5158,
                 reg5159,
                 reg5160,
                 reg5161,
                 forvar5162,
                 reg5163,
                 reg5164,
                 forvar5165,
                 forvar5166,
                 reg5167,
                 reg5168,
                 reg5169,
                 forvar5170,
                 forvar5171,
                 reg5172,
                 reg5173,
                 reg5174,
                 forvar5175,
                 reg5176,
                 forvar5177,
                 reg5178,
                 reg5179,
                 reg5180,
                 reg5181,
                 reg5182,
                 reg5183,
                 reg5184,
                 forvar5185,
                 reg5186,
                 forvar5187,
                 reg5188,
                 forvar5189,
                 reg5190,
                 reg5191,
                 reg5192,
                 reg5185,
                 forvar5186,
                 reg5187,
                 reg5189,
                 reg5193,
                 reg5194,
                 forvar5148,
                 wire5195,
                 wire5196,
                 wire5197,
                 forvar5198,
                 forvar5199,
                 reg5200,
                 reg5201,
                 reg5202,
                 reg5199,
                 reg5203,
                 reg5204,
                 reg5205,
                 forvar5206,
                 reg5207,
                 forvar5208,
                 reg5209,
                 reg5210,
                 reg5211,
                 reg5206,
                 reg5208,
                 reg5212,
                 reg5213,
                 reg5214,
                 reg5215,
                 reg5216,
                 forvar5217,
                 forvar5218,
                 reg5219,
                 reg5220,
                 reg5221,
                 reg5222,
                 reg5223,
                 forvar5224,
                 reg5225,
                 reg5226,
                 forvar5200,
                 reg5227,
                 forvar5228,
                 reg5229,
                 reg5230,
                 reg5231,
                 reg5232,
                 reg5233,
                 forvar5234,
                 reg5235,
                 reg5236,
                 reg5237,
                 forvar5238,
                 reg5239,
                 reg5240,
                 reg5241,
                 reg5242,
                 reg5234,
                 reg5228,
                 reg5243,
                 reg5244,
                 reg5245,
                 forvar5245,
                 reg5246,
                 reg5247,
                 forvar5248,
                 reg5249,
                 reg5250,
                 reg5251,
                 reg5252,
                 reg5253,
                 reg5254,
                 forvar5243,
                 forvar5247,
                 reg5248,
                 forvar5252,
                 reg5255,
                 reg5256,
                 forvar5257,
                 reg5258,
                 reg5259,
                 reg5260,
                 forvar5261,
                 reg5262,
                 reg5263,
                 reg5264,
                 reg5265,
                 forvar5266,
                 reg5267,
                 reg5268,
                 reg5269,
                 forvar5229,
                 forvar5231,
                 reg5238,
                 forvar5270,
                 reg5271,
                 forvar5272,
                 reg5273,
                 forvar5274,
                 reg5275,
                 reg5276,
                 reg5277,
                 reg5278,
                 reg5279,
                 forvar5280,
                 forvar5281,
                 reg5282,
                 reg5283,
                 reg5284,
                 forvar5285,
                 reg5286,
                 reg5287,
                 reg5288,
                 reg5289,
                 reg5290,
                 reg5291,
                 reg5292,
                 reg5293,
                 reg5294,
                 reg5295,
                 reg5296,
                 reg5297,
                 forvar5298,
                 reg5299,
                 reg5300,
                 forvar5292,
                 forvar5297,
                 reg5298,
                 reg5301,
                 reg5302,
                 reg5272,
                 reg5274,
                 forvar5277,
                 reg5280,
                 reg5281,
                 forvar5284,
                 reg5285,
                 forvar5301,
                 reg5303,
                 reg5304,
                 reg5305,
                 forvar5302,
                 forvar5306,
                 forvar5307,
                 reg5308,
                 reg5309,
                 reg5310,
                 reg5311,
                 reg5312,
                 reg5313,
                 forvar5314,
                 reg5315,
                 reg5316,
                 reg5317,
                 reg5318,
                 reg5319,
                 reg5320,
                 reg5321,
                 reg5322,
                 reg5314,
                 forvar5323,
                 reg5324,
                 reg5325,
                 forvar5326,
                 reg5327,
                 forvar5328,
                 reg5329,
                 reg5330,
                 reg5331,
                 reg5332,
                 reg5333,
                 reg5334,
                 reg5335,
                 reg5336,
                 reg5337,
                 reg5338,
                 reg5339,
                 forvar5340,
                 forvar5341,
                 reg5342,
                 reg5343,
                 reg5344,
                 reg5345,
                 reg5346,
                 reg5347,
                 reg5348,
                 forvar5349,
                 forvar5350,
                 reg5351,
                 reg5352,
                 reg5353,
                 reg5354,
                 forvar5355,
                 reg5356,
                 reg5357,
                 reg5358,
                 reg5359,
                 reg5360,
                 reg5361,
                 reg5362,
                 reg5355,
                 forvar5363,
                 reg5364,
                 reg5365,
                 reg5366,
                 reg5367,
                 forvar5368,
                 reg5369,
                 forvar5370,
                 reg5371,
                 forvar5372,
                 reg5373,
                 reg5374,
                 forvar5375,
                 reg5376,
                 forvar5377,
                 reg5378,
                 reg5379,
                 forvar5380,
                 reg5381,
                 reg5382,
                 reg5383,
                 reg5384,
                 reg5385,
                 forvar5376,
                 reg5377,
                 reg5380,
                 reg5386,
                 forvar5382,
                 forvar5387,
                 forvar5388,
                 reg5389,
                 reg5390,
                 reg5391,
                 reg5392,
                 forvar5393,
                 reg5394,
                 forvar5395,
                 reg5396,
                 reg5397,
                 reg5398,
                 reg5399,
                 reg5400,
                 reg5401,
                 reg5402,
                 forvar5403,
                 forvar5404,
                 forvar5405,
                 reg5406,
                 reg5407,
                 reg5408,
                 forvar5409,
                 reg5410,
                 reg5411,
                 reg5412,
                 reg5413,
                 reg5414,
                 reg5415,
                 forvar5416,
                 reg5417,
                 reg5418,
                 reg5419,
                 forvar5420,
                 reg5421,
                 reg5422,
                 reg5423,
                 forvar5424,
                 reg5425,
                 reg5426,
                 reg5427,
                 forvar5423,
                 forvar5427,
                 reg5428,
                 reg5429,
                 reg5430,
                 reg5431,
                 reg5432,
                 reg5433,
                 reg5434,
                 forvar5435,
                 forvar5436,
                 reg5437,
                 forvar5438,
                 reg5439,
                 forvar5440,
                 reg5441,
                 forvar5442,
                 reg5443,
                 reg5444,
                 reg5445,
                 reg5446,
                 reg5447,
                 reg5448,
                 reg5449,
                 forvar5450,
                 reg5451,
                 reg5452,
                 reg5350,
                 reg5349,
                 forvar5353,
                 forvar5360,
                 forvar5362,
                 reg5363,
                 forvar5364,
                 forvar5366,
                 reg5368,
                 reg5370,
                 reg5372,
                 forvar5369,
                 reg5375,
                 forvar5378,
                 forvar5379,
                 forvar5383,
                 reg5388,
                 forvar5391,
                 reg5393,
                 reg5395,
                 forvar5373,
                 forvar5396,
                 forvar5398,
                 forvar5453,
                 forvar5454,
                 forvar5455,
                 reg5456,
                 reg5457,
                 forvar5458,
                 reg5459,
                 forvar5460,
                 reg5461,
                 reg5462,
                 reg5463,
                 reg5464,
                 reg5465,
                 forvar5466,
                 reg5467,
                 reg5468,
                 reg5466,
                 forvar5467,
                 reg5469,
                 reg5470,
                 reg5471,
                 forvar5472,
                 reg5473,
                 forvar5474,
                 reg5475,
                 forvar5476,
                 reg5477,
                 reg5478,
                 reg5479,
                 forvar5480,
                 reg5481,
                 reg5482,
                 reg5483,
                 reg5484,
                 reg5485,
                 reg5486,
                 reg5487,
                 reg5488,
                 reg5489,
                 reg5490,
                 reg5491,
                 reg5492,
                 reg5480,
                 forvar5484,
                 forvar5493,
                 reg5494,
                 reg5495,
                 reg5496,
                 forvar5497,
                 reg5498,
                 reg5499,
                 reg5500,
                 reg5501,
                 reg5502,
                 forvar5503,
                 reg5504,
                 wire6862,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (((wire4574 << wire4576[(2'h2):(2'h2)]) ^~ {(8'hb6)}))
        begin
          reg4577 <= wire4576[(3'h4):(1'h0)];
          reg4578 <= $signed($signed(($signed(wire4576) ?
              $unsigned(wire4574) : $unsigned(wire4574))));
          if (wire4575[(1'h1):(1'h1)])
            begin
              for (forvar4579 = (1'h0); (forvar4579 < (1'h0)); forvar4579 = (forvar4579 + (1'h1)))
                begin
                  reg4580 <= wire4576[(3'h4):(2'h2)];
                  if ((wire4573[(1'h1):(1'h0)] <<< ($unsigned(wire4573[(2'h3):(2'h3)]) ?
                      wire4574 : $signed(((8'hb3) <<< forvar4579)))))
                    begin
                      reg4581 <= wire4576;
                      reg4582 <= wire4576;
                      reg4583 <= {((8'ha3) + (^~wire4574[(3'h7):(2'h3)]))};
                      reg4584 <= wire4574[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg4581 <= {(&(8'ha1))};
                    end
                  if (forvar4579[(1'h0):(1'h0)])
                    begin
                      reg4585 <= ((reg4580[(3'h7):(1'h1)] <= $signed((~^reg4578))) ?
                          $signed(((forvar4579 ?
                              wire4574 : reg4580) >>> $unsigned(reg4583))) : reg4584[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg4585 <= ((+reg4578[(1'h1):(1'h1)]) ?
                          {($signed((8'ha3)) ?
                                  $unsigned(reg4585) : (8'hb6))} : {(reg4582[(2'h2):(2'h2)] ?
                                  (~^reg4581) : wire4576[(1'h0):(1'h0)])});
                      reg4586 <= {(({wire4573} || $unsigned(reg4577)) ?
                              wire4575 : ((reg4584 ? reg4584 : (8'ha7)) ?
                                  $unsigned(reg4577) : (^reg4577)))};
                      reg4587 <= (($unsigned($signed(reg4583)) < $unsigned((8'hb8))) ^~ ((&{reg4586}) ?
                          (+reg4582) : ($unsigned(wire4574) ?
                              wire4576 : (wire4573 ? wire4574 : (8'hb3)))));
                    end
                  for (forvar4588 = (1'h0); (forvar4588 < (2'h3)); forvar4588 = (forvar4588 + (1'h1)))
                    begin
                      reg4589 <= reg4578;
                      reg4590 <= $unsigned((($unsigned(reg4587) ~^ $unsigned(reg4586)) ?
                          $signed(reg4585[(3'h4):(1'h1)]) : (-$unsigned(reg4585))));
                      reg4591 <= $signed($signed((^$signed(wire4576))));
                    end
                end
              reg4592 <= wire4573;
            end
          else
            begin
              reg4579 <= (($signed({reg4577}) ^ (reg4581[(3'h7):(1'h0)] >> reg4582)) || (-$unsigned($unsigned(reg4581))));
              for (forvar4580 = (1'h0); (forvar4580 < (2'h3)); forvar4580 = (forvar4580 + (1'h1)))
                begin
                  for (forvar4581 = (1'h0); (forvar4581 < (2'h2)); forvar4581 = (forvar4581 + (1'h1)))
                    begin
                      reg4582 <= reg4591;
                      reg4583 <= $signed($signed($signed((~reg4584))));
                      reg4584 <= $unsigned(forvar4581);
                    end
                  reg4585 <= ((8'hb4) ?
                      {reg4581[(4'hd):(2'h3)]} : {reg4586[(1'h0):(1'h0)]});
                  reg4586 <= $unsigned({((^~reg4581) ? reg4587 : reg4590)});
                end
            end
          if ($unsigned(forvar4579[(2'h2):(2'h2)]))
            begin
              for (forvar4593 = (1'h0); (forvar4593 < (1'h1)); forvar4593 = (forvar4593 + (1'h1)))
                begin
                  for (forvar4594 = (1'h0); (forvar4594 < (2'h3)); forvar4594 = (forvar4594 + (1'h1)))
                    begin
                      reg4595 <= ((~forvar4580[(1'h1):(1'h1)]) - (^(+reg4592[(3'h4):(2'h3)])));
                    end
                  if ((($signed(forvar4588) ?
                          $signed($unsigned(forvar4593)) : wire4575) ?
                      $unsigned($unsigned($unsigned(wire4575))) : (&($signed((8'hab)) ?
                          (8'hb5) : ((8'hb3) >>> reg4589)))))
                    begin
                      reg4596 <= (~|(~&$signed(reg4585[(3'h7):(3'h5)])));
                      reg4597 <= {($unsigned((forvar4593 <<< reg4596)) ?
                              $signed((reg4591 ?
                                  reg4584 : reg4585)) : {(reg4592 > reg4580)})};
                    end
                  else
                    begin
                      reg4596 <= $unsigned($signed(reg4590[(1'h1):(1'h1)]));
                      reg4597 <= $signed((~&reg4579[(4'he):(3'h5)]));
                    end
                  if (reg4590[(2'h3):(2'h3)])
                    begin
                      reg4598 <= (reg4591 ?
                          forvar4580[(3'h7):(3'h5)] : ($signed({reg4597}) ?
                              (|forvar4593) : forvar4593));
                      reg4599 <= $signed($unsigned($signed(reg4596)));
                      reg4600 <= $signed(($unsigned((8'ha7)) ?
                          $signed($unsigned((8'ha4))) : $unsigned((8'hb0))));
                      reg4601 <= (8'h9f);
                    end
                  else
                    begin
                      reg4598 <= reg4596[(2'h2):(1'h0)];
                      reg4599 <= (($unsigned((&reg4580)) ?
                          $signed(reg4589[(3'h5):(2'h2)]) : $unsigned($unsigned(reg4601))) && (~&(~&{reg4584})));
                      reg4600 <= (+reg4580[(4'ha):(4'h9)]);
                    end
                  for (forvar4602 = (1'h0); (forvar4602 < (2'h2)); forvar4602 = (forvar4602 + (1'h1)))
                    begin
                      reg4603 <= reg4585[(3'h6):(1'h1)];
                      reg4604 <= $signed(reg4599[(4'ha):(3'h5)]);
                    end
                end
              reg4605 <= $signed(reg4595[(1'h1):(1'h1)]);
            end
          else
            begin
              if ((((~|reg4604) << (~&(forvar4602 ?
                  reg4589 : reg4599))) | wire4575))
                begin
                  for (forvar4593 = (1'h0); (forvar4593 < (1'h1)); forvar4593 = (forvar4593 + (1'h1)))
                    begin
                      reg4594 <= $unsigned((^~reg4604[(3'h5):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar4593 = (1'h0); (forvar4593 < (1'h0)); forvar4593 = (forvar4593 + (1'h1)))
                    begin
                      reg4594 <= reg4590[(3'h4):(3'h4)];
                      reg4595 <= $signed((((8'ha1) < reg4600) >= {$unsigned((8'hb9))}));
                      reg4596 <= (8'hab);
                      reg4597 <= $signed({(reg4594 ^~ (&reg4585))});
                    end
                  reg4598 <= $signed((|($signed(forvar4580) + wire4574)));
                  if ($unsigned((reg4578[(1'h0):(1'h0)] ?
                      (!reg4591[(1'h0):(1'h0)]) : forvar4580[(1'h1):(1'h1)])))
                    begin
                      reg4599 <= ((forvar4580[(3'h4):(1'h0)] <= wire4576) <= ($signed(((8'hb2) << reg4581)) >>> (|(~|reg4589))));
                      reg4600 <= $signed((forvar4588[(4'h9):(4'h9)] ?
                          reg4598[(3'h6):(3'h5)] : $signed(reg4585)));
                      reg4601 <= (|((((8'h9d) ^ wire4573) != {(8'h9d)}) == $unsigned({reg4586})));
                      reg4602 <= (!forvar4588);
                    end
                  else
                    begin
                      reg4599 <= ($unsigned(($signed(reg4583) + (forvar4588 - reg4587))) > wire4575[(2'h2):(1'h0)]);
                    end
                  for (forvar4603 = (1'h0); (forvar4603 < (2'h2)); forvar4603 = (forvar4603 + (1'h1)))
                    begin
                      reg4604 <= $signed($signed((8'h9e)));
                    end
                end
              reg4605 <= forvar4594[(4'h8):(3'h7)];
              reg4606 <= $signed((wire4576[(1'h0):(1'h0)] + reg4601));
              for (forvar4607 = (1'h0); (forvar4607 < (2'h2)); forvar4607 = (forvar4607 + (1'h1)))
                begin
                  for (forvar4608 = (1'h0); (forvar4608 < (1'h0)); forvar4608 = (forvar4608 + (1'h1)))
                    begin
                      reg4609 <= reg4584;
                    end
                end
            end
        end
      else
        begin
          for (forvar4577 = (1'h0); (forvar4577 < (2'h2)); forvar4577 = (forvar4577 + (1'h1)))
            begin
              for (forvar4578 = (1'h0); (forvar4578 < (1'h0)); forvar4578 = (forvar4578 + (1'h1)))
                begin
                  reg4579 <= $signed(($unsigned($unsigned(reg4600)) ?
                      {$unsigned(reg4577)} : $signed($unsigned(reg4602))));
                  reg4580 <= $unsigned((((reg4609 || reg4604) ?
                      (!forvar4593) : reg4597[(1'h0):(1'h0)]) && reg4599[(3'h4):(2'h2)]));
                  if ($unsigned((~^wire4575)))
                    begin
                      reg4581 <= $unsigned($unsigned((^~{forvar4578})));
                      reg4582 <= ((8'hba) ?
                          (8'hb9) : $signed((reg4583 ?
                              (-forvar4578) : $unsigned(wire4576))));
                      reg4583 <= $signed($signed(((reg4586 ?
                              wire4576 : reg4606) ?
                          forvar4607 : (reg4583 <= forvar4593))));
                    end
                  else
                    begin
                      reg4581 <= reg4581;
                      reg4582 <= {($unsigned(reg4595) != wire4575)};
                    end
                  for (forvar4584 = (1'h0); (forvar4584 < (1'h1)); forvar4584 = (forvar4584 + (1'h1)))
                    begin
                      reg4585 <= $signed($unsigned($signed($signed(reg4577))));
                      reg4586 <= ((-forvar4603[(2'h3):(2'h2)]) <<< (^~$unsigned($signed(reg4589))));
                      reg4587 <= $unsigned($unsigned($signed((reg4603 ?
                          reg4582 : reg4609))));
                    end
                end
              for (forvar4588 = (1'h0); (forvar4588 < (2'h3)); forvar4588 = (forvar4588 + (1'h1)))
                begin
                  if ($signed(((forvar4584 ?
                          reg4578[(2'h3):(1'h0)] : $unsigned(forvar4580)) ?
                      forvar4608 : (&(8'haa)))))
                    begin
                      reg4589 <= $unsigned(reg4578[(3'h7):(2'h3)]);
                    end
                  else
                    begin
                      reg4589 <= (~^$unsigned($unsigned(forvar4577[(3'h6):(1'h0)])));
                      reg4590 <= (8'hb4);
                    end
                end
              for (forvar4591 = (1'h0); (forvar4591 < (1'h1)); forvar4591 = (forvar4591 + (1'h1)))
                begin
                  for (forvar4592 = (1'h0); (forvar4592 < (2'h2)); forvar4592 = (forvar4592 + (1'h1)))
                    begin
                      reg4593 <= {((8'hb4) ^~ ((~|forvar4602) ?
                              (&(8'ha3)) : {reg4592}))};
                    end
                  reg4594 <= $signed((~&($unsigned(reg4602) ?
                      (forvar4588 != forvar4577) : $unsigned(reg4602))));
                  if (({$signed($unsigned(reg4605))} ?
                      ($unsigned(forvar4608[(3'h7):(3'h4)]) ?
                          forvar4603 : $unsigned($signed(reg4589))) : reg4580[(4'h8):(3'h4)]))
                    begin
                      reg4595 <= {{(~|reg4596[(3'h6):(2'h3)])}};
                      reg4596 <= $signed(({(~^(8'haf))} > $signed((forvar4594 ?
                          (8'hb3) : reg4606))));
                      reg4597 <= {reg4589[(3'h6):(2'h2)]};
                    end
                  else
                    begin
                      reg4595 <= $signed((+({forvar4602} ?
                          forvar4580 : wire4573[(3'h4):(1'h1)])));
                      reg4596 <= reg4606;
                    end
                end
              for (forvar4598 = (1'h0); (forvar4598 < (2'h2)); forvar4598 = (forvar4598 + (1'h1)))
                begin
                  reg4599 <= ((forvar4581 <= reg4593[(2'h2):(2'h2)]) ?
                      forvar4584[(2'h3):(1'h0)] : (~|(reg4582[(1'h0):(1'h0)] + (forvar4598 ?
                          reg4581 : wire4573))));
                  if (($unsigned($signed($signed((8'h9c)))) ?
                      $signed(reg4585) : {(reg4601[(1'h0):(1'h0)] & $signed(forvar4593))}))
                    begin
                      reg4600 <= $signed(forvar4608[(4'hd):(4'hb)]);
                      reg4601 <= {{$unsigned((^~forvar4578))}};
                    end
                  else
                    begin
                      reg4600 <= (+(&(^~$unsigned(forvar4577))));
                      reg4601 <= reg4578[(3'h5):(2'h2)];
                    end
                  for (forvar4602 = (1'h0); (forvar4602 < (2'h3)); forvar4602 = (forvar4602 + (1'h1)))
                    begin
                      reg4603 <= forvar4591[(2'h3):(1'h0)];
                    end
                end
            end
          if (((^~(8'hac)) ? forvar4579[(3'h4):(2'h3)] : reg4603))
            begin
              if ($unsigned($unsigned((forvar4602[(3'h4):(1'h1)] ?
                  $unsigned(wire4576) : {reg4578}))))
                begin
                  for (forvar4604 = (1'h0); (forvar4604 < (2'h2)); forvar4604 = (forvar4604 + (1'h1)))
                    begin
                      reg4605 <= (forvar4579[(1'h1):(1'h0)] >> $signed((+$unsigned(reg4600))));
                      reg4606 <= ($signed(($unsigned(reg4603) ?
                              $unsigned((8'hb2)) : (forvar4598 ^ reg4605))) ?
                          (&$unsigned($unsigned(reg4582))) : (~|$signed($unsigned(forvar4580))));
                      reg4607 <= $signed(reg4581);
                    end
                  if ($signed($signed($signed((&(8'hae))))))
                    begin
                      reg4608 <= $unsigned($signed($signed(wire4575[(1'h1):(1'h0)])));
                      reg4609 <= $signed($unsigned((reg4607 + reg4596[(3'h6):(2'h2)])));
                    end
                  else
                    begin
                      reg4608 <= $unsigned({reg4578});
                      reg4609 <= (($unsigned($unsigned(reg4605)) << $unsigned(reg4582[(1'h1):(1'h0)])) & (-$unsigned((reg4606 ?
                          reg4589 : reg4597))));
                      reg4610 <= ($unsigned(reg4607) ? (!{reg4582}) : reg4583);
                    end
                  for (forvar4611 = (1'h0); (forvar4611 < (2'h2)); forvar4611 = (forvar4611 + (1'h1)))
                    begin
                      reg4612 <= $signed({reg4607});
                      reg4613 <= ($unsigned(reg4580[(3'h4):(2'h2)]) ?
                          (~&{(forvar4577 || forvar4584)}) : $unsigned(($signed(reg4590) << (~|(8'hba)))));
                    end
                  reg4614 <= (-{($unsigned(forvar4578) ^ (reg4586 | reg4592))});
                end
              else
                begin
                  if ((((wire4575 ?
                          $unsigned((8'ha9)) : $signed(reg4594)) ^~ (8'hb8)) ?
                      (~^(forvar4584[(4'ha):(3'h7)] ^~ $signed(reg4595))) : forvar4608))
                    begin
                      reg4604 <= $unsigned({(~^(reg4595 + reg4583))});
                      reg4605 <= (((^((8'ha1) ? forvar4578 : reg4602)) ?
                          $signed($signed(reg4599)) : reg4605[(2'h3):(1'h0)]) || $signed(forvar4592[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg4604 <= $signed({((forvar4598 ? (8'ha1) : (8'hb3)) ?
                              forvar4598[(3'h7):(3'h5)] : $signed(reg4584))});
                      reg4605 <= ((!forvar4602[(3'h6):(3'h6)]) ?
                          reg4603[(4'h8):(3'h6)] : $signed(forvar4608[(1'h0):(1'h0)]));
                    end
                  if (forvar4602)
                    begin
                      reg4606 <= (8'ha7);
                      reg4607 <= (~|($unsigned(reg4606) && (~^(^~reg4603))));
                    end
                  else
                    begin
                      reg4606 <= $signed({reg4598[(3'h6):(3'h6)]});
                      reg4607 <= ((forvar4611[(1'h0):(1'h0)] ?
                              ({reg4587} ?
                                  forvar4584 : (reg4606 <= reg4587)) : $signed({forvar4591})) ?
                          $unsigned({reg4593[(2'h2):(2'h2)]}) : reg4600[(3'h7):(2'h3)]);
                    end
                  for (forvar4608 = (1'h0); (forvar4608 < (2'h2)); forvar4608 = (forvar4608 + (1'h1)))
                    begin
                      reg4609 <= $unsigned(({(8'hb2)} != {reg4610}));
                      reg4610 <= forvar4603[(2'h3):(1'h1)];
                    end
                  for (forvar4611 = (1'h0); (forvar4611 < (1'h0)); forvar4611 = (forvar4611 + (1'h1)))
                    begin
                      reg4612 <= reg4601;
                    end
                end
            end
          else
            begin
              if (forvar4592)
                begin
                  for (forvar4604 = (1'h0); (forvar4604 < (1'h1)); forvar4604 = (forvar4604 + (1'h1)))
                    begin
                      reg4605 <= (8'hb3);
                      reg4606 <= ($signed(forvar4593[(1'h0):(1'h0)]) ?
                          (~|((reg4582 ?
                              wire4574 : forvar4607) || forvar4578[(1'h0):(1'h0)])) : reg4602);
                    end
                  if (reg4596[(1'h1):(1'h1)])
                    begin
                      reg4607 <= (reg4589[(1'h1):(1'h0)] + ($signed(reg4599[(1'h1):(1'h0)]) ?
                          $unsigned($unsigned(wire4576)) : forvar4594));
                      reg4608 <= reg4581[(2'h3):(2'h3)];
                      reg4609 <= $signed(((8'haf) ?
                          $unsigned(forvar4592) : (^~(forvar4592 + forvar4607))));
                    end
                  else
                    begin
                      reg4607 <= reg4601[(3'h7):(1'h0)];
                    end
                  for (forvar4610 = (1'h0); (forvar4610 < (2'h3)); forvar4610 = (forvar4610 + (1'h1)))
                    begin
                      reg4611 <= reg4598[(1'h0):(1'h0)];
                      reg4612 <= $unsigned((&forvar4579));
                    end
                  for (forvar4613 = (1'h0); (forvar4613 < (2'h2)); forvar4613 = (forvar4613 + (1'h1)))
                    begin
                      reg4614 <= reg4597[(2'h3):(2'h3)];
                      reg4615 <= ((~&((~^(8'h9d)) ~^ {reg4584})) <= $signed((reg4590 ?
                          {reg4595} : reg4606[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  for (forvar4604 = (1'h0); (forvar4604 < (2'h3)); forvar4604 = (forvar4604 + (1'h1)))
                    begin
                      reg4605 <= $unsigned(forvar4592);
                      reg4606 <= {((&reg4600[(3'h4):(3'h4)]) ?
                              (forvar4584 ?
                                  (-forvar4591) : $signed((8'hb5))) : (8'ha4))};
                      reg4607 <= $signed(forvar4610);
                      reg4608 <= reg4590[(3'h6):(3'h4)];
                    end
                  for (forvar4609 = (1'h0); (forvar4609 < (1'h0)); forvar4609 = (forvar4609 + (1'h1)))
                    begin
                      reg4610 <= {reg4598};
                    end
                end
              for (forvar4616 = (1'h0); (forvar4616 < (2'h3)); forvar4616 = (forvar4616 + (1'h1)))
                begin
                  for (forvar4617 = (1'h0); (forvar4617 < (1'h1)); forvar4617 = (forvar4617 + (1'h1)))
                    begin
                      reg4618 <= (forvar4609 * (-(~$signed((8'ha5)))));
                      reg4619 <= ($unsigned($unsigned((~|reg4582))) >> reg4612);
                      reg4620 <= reg4609;
                      reg4621 <= (!forvar4594);
                    end
                  if ((~(8'hb6)))
                    begin
                      reg4622 <= forvar4611;
                      reg4623 <= forvar4613[(4'hb):(4'ha)];
                    end
                  else
                    begin
                      reg4622 <= (((8'hb5) ?
                          ((reg4585 ? forvar4579 : (8'had)) ?
                              reg4620[(1'h1):(1'h1)] : (|reg4590)) : (8'h9d)) == {$unsigned($signed(forvar4588))});
                      reg4623 <= (~|$unsigned($signed({wire4575})));
                    end
                end
              if ({((8'ha9) - $unsigned($signed(forvar4591)))})
                begin
                  if (forvar4604[(2'h3):(2'h2)])
                    begin
                      reg4624 <= (8'hb5);
                      reg4625 <= wire4573;
                    end
                  else
                    begin
                      reg4624 <= $unsigned((reg4581 > wire4574));
                    end
                  if (forvar4607[(3'h4):(3'h4)])
                    begin
                      reg4626 <= forvar4580;
                      reg4627 <= $unsigned((^~forvar4591));
                      reg4628 <= ($signed(reg4615[(1'h0):(1'h0)]) ?
                          $signed(reg4611) : ((reg4619[(2'h3):(1'h1)] ?
                                  $signed(reg4604) : (forvar4579 ^ forvar4602)) ?
                              reg4627 : reg4600[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg4626 <= reg4615[(3'h4):(2'h2)];
                      reg4627 <= reg4614[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar4624 = (1'h0); (forvar4624 < (2'h2)); forvar4624 = (forvar4624 + (1'h1)))
                    begin
                      reg4625 <= (reg4589 != $unsigned(($unsigned(reg4592) >>> (reg4606 ?
                          reg4589 : (8'ha5)))));
                      reg4626 <= $signed($signed({$unsigned(forvar4611)}));
                      reg4627 <= $unsigned(($signed($unsigned(reg4595)) ?
                          (forvar4580[(1'h0):(1'h0)] ?
                              (forvar4579 == reg4591) : (~&reg4622)) : $unsigned(((8'hb4) | reg4579))));
                    end
                  if ((forvar4602[(4'ha):(1'h1)] < (~$signed((8'h9e)))))
                    begin
                      reg4628 <= (^(^~((!(8'ha1)) ?
                          (forvar4581 ?
                              forvar4610 : forvar4591) : (^reg4580))));
                    end
                  else
                    begin
                      reg4628 <= $signed((~&$signed((&reg4625))));
                      reg4629 <= {reg4583[(1'h1):(1'h0)]};
                      reg4630 <= reg4594;
                    end
                end
              if (((|wire4575) ?
                  (reg4592 | ({forvar4609} + forvar4593[(3'h4):(2'h3)])) : forvar4611[(3'h7):(2'h2)]))
                begin
                  if ($unsigned($unsigned((((8'hb7) ? reg4624 : reg4620) ?
                      ((8'hba) - (8'haa)) : (reg4591 ? reg4586 : forvar4578)))))
                    begin
                      reg4631 <= forvar4598[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg4631 <= $signed($unsigned($signed($unsigned((8'hac)))));
                    end
                end
              else
                begin
                  reg4631 <= reg4596;
                  reg4632 <= ((-{((8'ha7) - (8'hb8))}) ?
                      (^((reg4596 ^~ forvar4611) || forvar4577[(4'hb):(1'h0)])) : $unsigned((~|$signed((8'ha3)))));
                  if (($unsigned((8'ha8)) ?
                      {reg4579[(4'hf):(4'h8)]} : (~&(reg4606 && $unsigned(reg4579)))))
                    begin
                      reg4633 <= forvar4579;
                      reg4634 <= $signed($unsigned(($signed((8'h9e)) ?
                          ((8'ha8) + forvar4608) : $unsigned(reg4585))));
                    end
                  else
                    begin
                      reg4633 <= forvar4581[(1'h0):(1'h0)];
                      reg4634 <= {forvar4608};
                    end
                end
            end
          if (forvar4577[(4'h9):(1'h0)])
            begin
              reg4635 <= ((($unsigned(reg4630) ?
                      reg4618[(1'h0):(1'h0)] : {reg4607}) & (-reg4602)) ?
                  reg4623 : (~|($signed((8'ha5)) && reg4594)));
              if (((((reg4621 ? reg4614 : reg4621) ?
                      reg4627[(4'h9):(1'h1)] : {reg4612}) ?
                  $signed((|reg4629)) : forvar4592) * reg4618))
                begin
                  if ({reg4583[(3'h4):(1'h1)]})
                    begin
                      reg4636 <= $unsigned((|reg4600));
                      reg4637 <= reg4599[(2'h3):(1'h0)];
                      reg4638 <= reg4621;
                    end
                  else
                    begin
                      reg4636 <= ($signed(forvar4580) ?
                          forvar4591 : reg4635[(4'hb):(3'h5)]);
                      reg4637 <= wire4574[(4'hc):(4'hc)];
                    end
                end
              else
                begin
                  for (forvar4636 = (1'h0); (forvar4636 < (2'h2)); forvar4636 = (forvar4636 + (1'h1)))
                    begin
                      reg4637 <= $signed((((reg4621 ? (8'hb4) : forvar4636) ?
                              {reg4629} : forvar4579[(1'h0):(1'h0)]) ?
                          wire4573[(2'h2):(1'h1)] : ({reg4606} >> {reg4630})));
                      reg4638 <= reg4632[(2'h2):(1'h1)];
                      reg4639 <= (&($signed((reg4600 ?
                          reg4615 : reg4583)) + reg4590));
                    end
                  for (forvar4640 = (1'h0); (forvar4640 < (2'h2)); forvar4640 = (forvar4640 + (1'h1)))
                    begin
                      reg4641 <= $unsigned({($signed(reg4607) ?
                              $unsigned(forvar4593) : $unsigned(reg4628))});
                    end
                end
              if ($unsigned((wire4576 > forvar4578[(1'h1):(1'h1)])))
                begin
                  reg4642 <= reg4609[(3'h7):(2'h2)];
                  for (forvar4643 = (1'h0); (forvar4643 < (2'h3)); forvar4643 = (forvar4643 + (1'h1)))
                    begin
                      reg4644 <= $unsigned(reg4630[(3'h5):(1'h0)]);
                      reg4645 <= forvar4616;
                      reg4646 <= (!(^~$signed((forvar4578 ?
                          (8'ha3) : wire4574))));
                      reg4647 <= (-reg4634);
                    end
                  for (forvar4648 = (1'h0); (forvar4648 < (1'h0)); forvar4648 = (forvar4648 + (1'h1)))
                    begin
                      reg4649 <= (({{reg4644}} ?
                              forvar4588 : ((forvar4608 < forvar4636) + $signed(forvar4616))) ?
                          reg4593[(2'h3):(2'h2)] : (forvar4580 & $unsigned($signed(forvar4579))));
                    end
                  for (forvar4650 = (1'h0); (forvar4650 < (1'h1)); forvar4650 = (forvar4650 + (1'h1)))
                    begin
                      reg4651 <= reg4593[(2'h3):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar4642 = (1'h0); (forvar4642 < (1'h1)); forvar4642 = (forvar4642 + (1'h1)))
                    begin
                      reg4643 <= forvar4648;
                      reg4644 <= reg4629[(3'h5):(3'h4)];
                    end
                  for (forvar4645 = (1'h0); (forvar4645 < (1'h0)); forvar4645 = (forvar4645 + (1'h1)))
                    begin
                      reg4646 <= (reg4605[(3'h5):(2'h2)] ?
                          (({(8'h9c)} ?
                                  reg4577[(3'h6):(3'h4)] : (~&forvar4608)) ?
                              reg4585 : reg4585[(2'h3):(2'h2)]) : $signed(reg4615));
                      reg4647 <= (8'h9c);
                    end
                end
            end
          else
            begin
              reg4635 <= ($unsigned(reg4639) ?
                  reg4639 : (^(wire4575 >>> (forvar4650 ? reg4651 : reg4578))));
            end
        end
      for (forvar4652 = (1'h0); (forvar4652 < (1'h0)); forvar4652 = (forvar4652 + (1'h1)))
        begin
          for (forvar4653 = (1'h0); (forvar4653 < (1'h1)); forvar4653 = (forvar4653 + (1'h1)))
            begin
              if ($unsigned(reg4585[(2'h2):(1'h1)]))
                begin
                  reg4654 <= forvar4603;
                  if (forvar4613)
                    begin
                      reg4655 <= {{(8'hba)}};
                      reg4656 <= (!($signed(reg4619) >= ($signed(reg4628) + reg4596[(1'h1):(1'h0)])));
                      reg4657 <= forvar4652;
                    end
                  else
                    begin
                      reg4655 <= {forvar4577[(3'h5):(1'h1)]};
                      reg4656 <= $unsigned((~$unsigned((reg4619 == (8'ha4)))));
                      reg4657 <= (((+{forvar4580}) ?
                              (reg4647[(3'h5):(2'h3)] + reg4638[(2'h2):(1'h0)]) : $unsigned(reg4604[(2'h3):(1'h1)])) ?
                          (reg4602[(3'h6):(3'h6)] & forvar4594[(1'h1):(1'h0)]) : $signed(($unsigned(forvar4643) == $signed(forvar4648))));
                    end
                  reg4658 <= $unsigned((wire4576 < (forvar4594[(5'h10):(3'h5)] & reg4615[(1'h0):(1'h0)])));
                end
              else
                begin
                  for (forvar4654 = (1'h0); (forvar4654 < (1'h0)); forvar4654 = (forvar4654 + (1'h1)))
                    begin
                      reg4655 <= (($unsigned({wire4574}) ?
                              ((&(8'had)) - reg4609[(3'h6):(3'h6)]) : forvar4608[(4'hd):(4'h8)]) ?
                          reg4642[(1'h1):(1'h0)] : forvar4642);
                    end
                  for (forvar4656 = (1'h0); (forvar4656 < (2'h2)); forvar4656 = (forvar4656 + (1'h1)))
                    begin
                      reg4657 <= reg4655[(3'h6):(3'h6)];
                    end
                end
              for (forvar4659 = (1'h0); (forvar4659 < (2'h3)); forvar4659 = (forvar4659 + (1'h1)))
                begin
                  if ($signed(($signed(forvar4603[(3'h6):(1'h1)]) ?
                      $signed(reg4627) : wire4576[(3'h4):(1'h0)])))
                    begin
                      reg4660 <= $unsigned((-(reg4645[(3'h6):(1'h0)] ?
                          forvar4656[(3'h4):(2'h2)] : (reg4593 ?
                              reg4596 : wire4574))));
                      reg4661 <= $signed((^(+(~&reg4627))));
                      reg4662 <= (wire4575 ?
                          $signed($signed(((8'haf) ?
                              reg4636 : (8'hb6)))) : $signed($signed((+reg4630))));
                    end
                  else
                    begin
                      reg4660 <= {$unsigned($unsigned($unsigned(reg4655)))};
                      reg4661 <= (~$unsigned(forvar4616));
                    end
                  for (forvar4663 = (1'h0); (forvar4663 < (2'h3)); forvar4663 = (forvar4663 + (1'h1)))
                    begin
                      reg4664 <= ($signed(reg4593[(1'h0):(1'h0)]) ?
                          ($unsigned(forvar4608[(1'h0):(1'h0)]) || $signed(wire4574[(2'h2):(1'h0)])) : $unsigned(reg4638[(1'h1):(1'h0)]));
                      reg4665 <= (reg4579[(2'h3):(2'h3)] ?
                          forvar4603 : forvar4611[(4'hb):(4'h9)]);
                      reg4666 <= ($unsigned((~(8'hb2))) <= ($unsigned(reg4606) ?
                          $signed($unsigned(reg4606)) : forvar4593[(3'h4):(1'h0)]));
                    end
                  if ((8'haf))
                    begin
                      reg4667 <= (^~$unsigned($unsigned((reg4579 <<< (8'ha8)))));
                      reg4668 <= $unsigned((~|forvar4584));
                      reg4669 <= reg4662[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg4667 <= wire4573[(4'he):(2'h3)];
                      reg4668 <= $signed({((reg4590 ? (8'ha7) : reg4646) ?
                              (forvar4645 << reg4593) : reg4643[(1'h1):(1'h1)])});
                    end
                  reg4670 <= (|reg4579[(3'h5):(3'h5)]);
                end
              reg4671 <= (~|(~$unsigned(forvar4604)));
            end
        end
      for (forvar4672 = (1'h0); (forvar4672 < (1'h0)); forvar4672 = (forvar4672 + (1'h1)))
        begin
          for (forvar4673 = (1'h0); (forvar4673 < (1'h0)); forvar4673 = (forvar4673 + (1'h1)))
            begin
              if ($unsigned((+((reg4670 ?
                  forvar4613 : (8'hae)) > reg4582[(2'h2):(1'h1)]))))
                begin
                  for (forvar4674 = (1'h0); (forvar4674 < (2'h3)); forvar4674 = (forvar4674 + (1'h1)))
                    begin
                      reg4675 <= (reg4639 > $signed(((forvar4581 * (8'ha6)) - (~&reg4604))));
                    end
                  for (forvar4676 = (1'h0); (forvar4676 < (1'h1)); forvar4676 = (forvar4676 + (1'h1)))
                    begin
                      reg4677 <= (~(+reg4614));
                    end
                  if ($signed((+(reg4607 >= $signed(reg4654)))))
                    begin
                      reg4678 <= (^~forvar4617);
                      reg4679 <= $unsigned($signed((reg4667[(3'h4):(1'h1)] ?
                          (reg4631 == reg4624) : $signed((8'hba)))));
                    end
                  else
                    begin
                      reg4678 <= ((forvar4608 > $signed((forvar4663 ?
                              reg4623 : reg4657))) ?
                          (~^(reg4677[(3'h6):(1'h1)] <<< (forvar4609 ?
                              (8'ha1) : reg4579))) : ((reg4609[(3'h6):(2'h3)] ?
                                  reg4642[(4'ha):(3'h5)] : reg4636) ?
                              $unsigned($unsigned((8'h9f))) : reg4626));
                      reg4679 <= reg4660[(1'h0):(1'h0)];
                      reg4680 <= (^$unsigned(reg4585[(3'h5):(3'h5)]));
                    end
                end
              else
                begin
                  for (forvar4674 = (1'h0); (forvar4674 < (1'h0)); forvar4674 = (forvar4674 + (1'h1)))
                    begin
                      reg4675 <= forvar4598[(1'h1):(1'h1)];
                      reg4676 <= $unsigned(reg4654);
                      reg4677 <= {reg4579};
                    end
                end
              for (forvar4681 = (1'h0); (forvar4681 < (2'h3)); forvar4681 = (forvar4681 + (1'h1)))
                begin
                  if ((((~^reg4626) >> reg4627) >= reg4636))
                    begin
                      reg4682 <= reg4587[(3'h5):(1'h0)];
                      reg4683 <= ($signed($signed(((8'h9d) <= reg4590))) < reg4613[(3'h6):(3'h6)]);
                      reg4684 <= ($signed((^~{reg4578})) ?
                          forvar4624 : (^~reg4582[(2'h2):(2'h2)]));
                      reg4685 <= ((~forvar4659[(3'h4):(1'h1)]) ?
                          forvar4598[(1'h1):(1'h1)] : (~&reg4684));
                    end
                  else
                    begin
                      reg4682 <= $unsigned($signed(forvar4636[(1'h1):(1'h1)]));
                      reg4683 <= ($unsigned(reg4587) ?
                          (8'ha9) : $signed($signed($unsigned((8'ha2)))));
                    end
                end
              reg4686 <= $signed({reg4618[(2'h3):(1'h1)]});
            end
          reg4687 <= (~|$signed(reg4614[(3'h4):(2'h2)]));
          if (forvar4672[(2'h3):(1'h1)])
            begin
              if (((^{(reg4687 ?
                      reg4582 : reg4595)}) == $unsigned((+forvar4613[(4'he):(4'hc)]))))
                begin
                  if ({$unsigned($signed(reg4624[(2'h2):(2'h2)]))})
                    begin
                      reg4688 <= ($signed((forvar4650 ?
                          (~|reg4685) : $signed(reg4679))) > forvar4659);
                    end
                  else
                    begin
                      reg4688 <= $signed($signed(((&reg4680) ?
                          $unsigned(forvar4609) : {reg4584})));
                    end
                  reg4689 <= forvar4648;
                end
              else
                begin
                  for (forvar4688 = (1'h0); (forvar4688 < (1'h1)); forvar4688 = (forvar4688 + (1'h1)))
                    begin
                      reg4689 <= (&$unsigned($signed(reg4590[(1'h0):(1'h0)])));
                      reg4690 <= reg4666[(1'h1):(1'h0)];
                    end
                  reg4691 <= ($unsigned(({reg4602} * (^~reg4587))) || ((~|reg4686) - (reg4577[(3'h4):(3'h4)] ?
                      $unsigned(forvar4579) : ((8'hb7) ~^ reg4609))));
                end
              reg4692 <= (|(((forvar4610 ? (8'haf) : (8'hb9)) ?
                  reg4601[(3'h6):(3'h5)] : (forvar4578 ?
                      (8'h9c) : (8'h9e))) ^ $unsigned(((8'h9f) ?
                  forvar4617 : reg4632))));
            end
          else
            begin
              for (forvar4688 = (1'h0); (forvar4688 < (1'h0)); forvar4688 = (forvar4688 + (1'h1)))
                begin
                  for (forvar4689 = (1'h0); (forvar4689 < (2'h2)); forvar4689 = (forvar4689 + (1'h1)))
                    begin
                      reg4690 <= {reg4631[(2'h3):(2'h3)]};
                      reg4691 <= (reg4642 ?
                          (~^{(reg4628 ? forvar4681 : reg4677)}) : (reg4594 ?
                              reg4668[(1'h1):(1'h1)] : $signed((reg4668 ?
                                  forvar4689 : (8'ha5)))));
                      reg4692 <= (+{reg4684});
                      reg4693 <= (($unsigned($unsigned(reg4609)) * ((reg4597 ?
                                  forvar4579 : forvar4650) ?
                              reg4666[(1'h1):(1'h1)] : (reg4628 ?
                                  forvar4617 : reg4677))) ?
                          $signed($signed($signed(reg4637))) : wire4576);
                    end
                  for (forvar4694 = (1'h0); (forvar4694 < (1'h0)); forvar4694 = (forvar4694 + (1'h1)))
                    begin
                      reg4695 <= forvar4581;
                    end
                  for (forvar4696 = (1'h0); (forvar4696 < (2'h2)); forvar4696 = (forvar4696 + (1'h1)))
                    begin
                      reg4697 <= {(!(^~(~|forvar4604)))};
                    end
                end
              for (forvar4698 = (1'h0); (forvar4698 < (2'h3)); forvar4698 = (forvar4698 + (1'h1)))
                begin
                  if (reg4579[(2'h3):(2'h3)])
                    begin
                      reg4699 <= (((!(^~forvar4609)) >>> reg4581) >>> $unsigned(((reg4688 <= forvar4676) >> $unsigned(forvar4613))));
                      reg4700 <= (reg4699 ?
                          $signed(($signed(reg4656) <<< wire4575)) : forvar4696[(2'h2):(1'h1)]);
                      reg4701 <= reg4625[(3'h6):(3'h5)];
                    end
                  else
                    begin
                      reg4699 <= ((-$signed(reg4701[(2'h3):(1'h0)])) ?
                          forvar4654[(3'h5):(2'h3)] : (&(~|reg4683[(1'h0):(1'h0)])));
                    end
                  if ({$signed($signed((-reg4666)))})
                    begin
                      reg4702 <= ($unsigned(forvar4696) >= forvar4688);
                      reg4703 <= $unsigned(forvar4604[(3'h5):(2'h3)]);
                      reg4704 <= (reg4697 ?
                          reg4686 : {(reg4637[(1'h0):(1'h0)] ?
                                  reg4688 : (reg4627 ? reg4580 : reg4671))});
                    end
                  else
                    begin
                      reg4702 <= reg4643[(2'h2):(1'h1)];
                      reg4703 <= ($unsigned($signed(reg4631)) & (({reg4596} ?
                          (~^(8'hae)) : (forvar4598 | forvar4698)) ~^ (!reg4584)));
                    end
                  for (forvar4705 = (1'h0); (forvar4705 < (1'h1)); forvar4705 = (forvar4705 + (1'h1)))
                    begin
                      reg4706 <= ($unsigned($signed((+reg4680))) <= (8'hb7));
                      reg4707 <= forvar4642[(1'h0):(1'h0)];
                    end
                  if ((&wire4574[(3'h7):(3'h7)]))
                    begin
                      reg4708 <= (((~&$unsigned(forvar4598)) << reg4624) == reg4593);
                      reg4709 <= $signed(forvar4598);
                    end
                  else
                    begin
                      reg4708 <= (!({$signed(reg4599)} & $unsigned((!reg4598))));
                      reg4709 <= ($signed(reg4639[(2'h3):(1'h0)]) + (-forvar4592[(3'h4):(1'h0)]));
                      reg4710 <= $signed($unsigned($unsigned(forvar4592[(2'h2):(1'h1)])));
                      reg4711 <= (~|(8'h9f));
                    end
                end
              if (forvar4611)
                begin
                  for (forvar4712 = (1'h0); (forvar4712 < (1'h0)); forvar4712 = (forvar4712 + (1'h1)))
                    begin
                      reg4713 <= (|(|$signed($signed(reg4600))));
                      reg4714 <= $signed(((|$unsigned(reg4591)) ?
                          (~|$unsigned(reg4693)) : ($signed(reg4632) || (forvar4642 <= reg4702))));
                    end
                  for (forvar4715 = (1'h0); (forvar4715 < (2'h3)); forvar4715 = (forvar4715 + (1'h1)))
                    begin
                      reg4716 <= $signed((~forvar4580[(3'h5):(3'h4)]));
                    end
                  for (forvar4717 = (1'h0); (forvar4717 < (2'h3)); forvar4717 = (forvar4717 + (1'h1)))
                    begin
                      reg4718 <= ((8'h9d) > reg4716[(2'h2):(1'h1)]);
                      reg4719 <= {forvar4617[(2'h3):(1'h1)]};
                      reg4720 <= wire4574;
                    end
                  if ({$unsigned(((~|reg4625) | reg4651))})
                    begin
                      reg4721 <= $unsigned(({$unsigned(reg4622)} ?
                          $signed($unsigned((8'ha1))) : reg4625));
                      reg4722 <= {reg4688[(3'h6):(3'h6)]};
                      reg4723 <= ($signed((^reg4624[(3'h6):(1'h1)])) ?
                          $signed(($signed(reg4622) ?
                              $signed(reg4611) : $unsigned((8'hb5)))) : ({(~reg4670)} ?
                              $signed((reg4646 ?
                                  (8'ha7) : forvar4642)) : ((reg4713 == (8'ha4)) ?
                                  $signed(reg4645) : (forvar4642 ?
                                      reg4609 : forvar4672))));
                      reg4724 <= (reg4577 ?
                          (forvar4696[(2'h2):(2'h2)] ?
                              $unsigned((reg4688 & reg4656)) : reg4677[(2'h2):(2'h2)]) : $signed(reg4687[(3'h5):(2'h2)]));
                    end
                  else
                    begin
                      reg4721 <= (|(($unsigned(reg4632) ? (8'ha3) : reg4655) ?
                          $signed($unsigned(reg4655)) : (^(~|forvar4659))));
                      reg4722 <= ((~&forvar4652[(2'h2):(1'h1)]) ?
                          (reg4623[(3'h4):(2'h2)] ?
                              $signed((reg4604 < reg4624)) : reg4691[(2'h2):(2'h2)]) : {reg4608[(3'h6):(3'h4)]});
                    end
                end
              else
                begin
                  for (forvar4712 = (1'h0); (forvar4712 < (1'h1)); forvar4712 = (forvar4712 + (1'h1)))
                    begin
                      reg4713 <= ($unsigned({reg4623[(4'hb):(4'ha)]}) > (reg4656[(3'h5):(1'h1)] >> (|(^wire4573))));
                      reg4714 <= $unsigned(({reg4600[(2'h2):(1'h1)]} ^ (^~(^forvar4577))));
                      reg4715 <= $signed($unsigned((reg4667 < reg4677)));
                      reg4716 <= ((((~reg4577) | forvar4673[(3'h7):(1'h1)]) * $unsigned(reg4699[(3'h6):(3'h5)])) ?
                          $unsigned(((8'hab) * (|reg4655))) : (reg4722 ?
                              $unsigned(reg4579[(1'h1):(1'h0)]) : $unsigned(reg4693)));
                    end
                  for (forvar4717 = (1'h0); (forvar4717 < (1'h0)); forvar4717 = (forvar4717 + (1'h1)))
                    begin
                      reg4718 <= (8'haa);
                    end
                end
              if (({($unsigned(reg4632) ~^ $unsigned(reg4710))} + ((~^$signed(reg4605)) || reg4626)))
                begin
                  for (forvar4725 = (1'h0); (forvar4725 < (2'h3)); forvar4725 = (forvar4725 + (1'h1)))
                    begin
                      reg4726 <= (~&$unsigned(reg4642));
                    end
                  for (forvar4727 = (1'h0); (forvar4727 < (1'h1)); forvar4727 = (forvar4727 + (1'h1)))
                    begin
                      reg4728 <= forvar4578[(1'h1):(1'h1)];
                      reg4729 <= ($unsigned({(!forvar4579)}) < reg4644);
                    end
                  if ((reg4614[(2'h3):(2'h2)] <<< ((reg4585[(2'h3):(1'h1)] & forvar4604[(1'h1):(1'h0)]) ?
                      forvar4673[(1'h0):(1'h0)] : $unsigned(reg4606))))
                    begin
                      reg4730 <= ((^($signed(forvar4674) ?
                              reg4706 : $signed(reg4657))) ?
                          reg4723 : forvar4672);
                      reg4731 <= (~|(({(8'hb4)} ?
                          (forvar4698 ?
                              forvar4705 : (8'hb2)) : reg4609) ~^ (~&(+reg4729))));
                    end
                  else
                    begin
                      reg4730 <= forvar4654[(3'h5):(2'h2)];
                      reg4731 <= ($signed(((reg4602 ? wire4574 : reg4610) ?
                          $signed(reg4600) : reg4605[(2'h2):(1'h1)])) + ($signed(((8'ha0) ~^ reg4677)) >> $unsigned((reg4641 <= reg4645))));
                      reg4732 <= $signed(forvar4654[(3'h6):(1'h1)]);
                    end
                  for (forvar4733 = (1'h0); (forvar4733 < (2'h3)); forvar4733 = (forvar4733 + (1'h1)))
                    begin
                      reg4734 <= (($signed((reg4713 || reg4685)) ~^ reg4638) * (~reg4685[(2'h3):(1'h0)]));
                      reg4735 <= $signed(reg4619[(3'h4):(2'h3)]);
                      reg4736 <= ($signed(($unsigned(reg4691) ?
                              {(8'hb0)} : reg4704)) ?
                          {(reg4628 ?
                                  forvar4673 : reg4647)} : (wire4573 | (^~(reg4631 >>> forvar4584))));
                    end
                end
              else
                begin
                  if (reg4722)
                    begin
                      reg4725 <= $unsigned({reg4693[(1'h0):(1'h0)]});
                      reg4726 <= (reg4707 >> reg4631);
                    end
                  else
                    begin
                      reg4725 <= reg4584;
                      reg4726 <= (&(reg4642 ^~ $signed($signed(forvar4604))));
                    end
                  if (forvar4603[(1'h1):(1'h0)])
                    begin
                      reg4727 <= ($unsigned(reg4578) ?
                          ($unsigned($signed((8'haf))) ?
                              reg4677[(3'h4):(2'h2)] : $signed({forvar4733})) : (+reg4625[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg4727 <= forvar4689;
                      reg4728 <= reg4664;
                      reg4729 <= ({forvar4656[(4'hd):(4'ha)]} ?
                          {$unsigned((reg4704 << reg4610))} : $signed((-reg4689[(3'h4):(1'h1)])));
                    end
                  reg4730 <= $signed(reg4664);
                  for (forvar4731 = (1'h0); (forvar4731 < (2'h2)); forvar4731 = (forvar4731 + (1'h1)))
                    begin
                      reg4732 <= reg4644[(1'h1):(1'h0)];
                      reg4733 <= (~(~^(8'hb2)));
                      reg4734 <= (-((&(-reg4683)) <<< ({forvar4613} ?
                          ((8'had) ?
                              reg4635 : forvar4642) : $unsigned(reg4693))));
                      reg4735 <= reg4631;
                    end
                end
            end
        end
      if (($unsigned(($signed(reg4632) ^ $signed(wire4574))) >= reg4666))
        begin
          if (reg4641)
            begin
              for (forvar4737 = (1'h0); (forvar4737 < (1'h0)); forvar4737 = (forvar4737 + (1'h1)))
                begin
                  if ((!$signed($unsigned($signed(forvar4616)))))
                    begin
                      reg4738 <= $signed(reg4603[(3'h7):(3'h4)]);
                      reg4739 <= (reg4730[(1'h1):(1'h1)] ?
                          $signed((forvar4591 + {(8'ha4)})) : {reg4598});
                      reg4740 <= (|(!$signed((|reg4585))));
                    end
                  else
                    begin
                      reg4738 <= $signed((^forvar4737));
                      reg4739 <= reg4684[(3'h4):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar4737 = (1'h0); (forvar4737 < (2'h2)); forvar4737 = (forvar4737 + (1'h1)))
                begin
                  for (forvar4738 = (1'h0); (forvar4738 < (1'h0)); forvar4738 = (forvar4738 + (1'h1)))
                    begin
                      reg4739 <= $signed(($unsigned($unsigned(reg4581)) ?
                          (((8'hb1) ? forvar4672 : (8'ha0)) ?
                              $signed(reg4647) : $unsigned(reg4708)) : reg4699[(3'h5):(1'h0)]));
                    end
                  if (reg4684)
                    begin
                      reg4740 <= $unsigned($unsigned(reg4687[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg4740 <= forvar4676;
                      reg4741 <= $signed(((reg4670 ?
                              {reg4635} : $signed(forvar4653)) ?
                          reg4628 : $signed($signed(reg4719))));
                      reg4742 <= $signed((~^($unsigned(reg4579) ?
                          $signed(reg4723) : $unsigned(reg4721))));
                      reg4743 <= $signed((~reg4604[(1'h1):(1'h0)]));
                    end
                end
              reg4744 <= ($unsigned(({reg4636} - ((8'ha8) ?
                      reg4584 : (8'hb4)))) ?
                  (($unsigned(reg4579) ?
                      (reg4591 ?
                          (8'haa) : reg4733) : (reg4625 >= reg4583)) | $unsigned((|forvar4593))) : $signed(($unsigned(reg4683) || (forvar4603 ?
                      (8'hb5) : reg4692))));
            end
          if (((&($unsigned(reg4741) ?
              (reg4720 ?
                  (8'ha1) : (8'ha6)) : reg4700)) ^~ {(((8'ha1) < forvar4738) ?
                  reg4675[(3'h6):(1'h0)] : reg4600)}))
            begin
              for (forvar4745 = (1'h0); (forvar4745 < (2'h3)); forvar4745 = (forvar4745 + (1'h1)))
                begin
                  if ($unsigned(reg4680[(2'h2):(1'h0)]))
                    begin
                      reg4746 <= $unsigned(reg4664);
                      reg4747 <= (reg4719[(1'h1):(1'h1)] || $signed(forvar4588));
                      reg4748 <= (8'ha4);
                    end
                  else
                    begin
                      reg4746 <= (!reg4726[(3'h6):(2'h2)]);
                      reg4747 <= $unsigned(reg4583);
                      reg4748 <= (reg4608 ?
                          {($signed(reg4733) < forvar4610[(3'h4):(3'h4)])} : (8'ha1));
                    end
                  for (forvar4749 = (1'h0); (forvar4749 < (2'h3)); forvar4749 = (forvar4749 + (1'h1)))
                    begin
                      reg4750 <= $unsigned(($unsigned($signed(reg4613)) ?
                          reg4620[(2'h3):(2'h3)] : (~^$unsigned(reg4654))));
                      reg4751 <= $signed($signed(reg4613[(2'h2):(1'h0)]));
                      reg4752 <= ($unsigned(((!forvar4580) <= (!reg4750))) ?
                          ((8'haa) || $signed($unsigned(reg4609))) : (reg4684[(4'hb):(4'h8)] ?
                              (|(reg4668 ?
                                  wire4575 : reg4644)) : (&(+reg4586))));
                      reg4753 <= $unsigned(({(reg4723 ? (8'ha3) : (8'hb2))} ?
                          forvar4616[(4'hd):(2'h2)] : $unsigned((forvar4659 ?
                              reg4593 : forvar4717))));
                    end
                  if (reg4688)
                    begin
                      reg4754 <= $unsigned((^$signed(reg4669)));
                      reg4755 <= reg4726[(3'h7):(2'h3)];
                      reg4756 <= ($unsigned((+$unsigned(forvar4674))) ?
                          ($signed($signed(reg4627)) ?
                              reg4669 : $unsigned((reg4686 ?
                                  reg4669 : reg4595))) : reg4679[(2'h2):(1'h0)]);
                      reg4757 <= forvar4643;
                    end
                  else
                    begin
                      reg4754 <= {(^~reg4710)};
                      reg4755 <= reg4727[(3'h4):(1'h1)];
                      reg4756 <= ((~^reg4644) ?
                          (reg4703[(2'h2):(1'h0)] ?
                              {(^~forvar4659)} : {reg4725}) : $unsigned((~(forvar4738 << forvar4636))));
                    end
                end
              if (reg4586)
                begin
                  reg4758 <= $unsigned((8'hb1));
                  for (forvar4759 = (1'h0); (forvar4759 < (2'h3)); forvar4759 = (forvar4759 + (1'h1)))
                    begin
                      reg4760 <= (wire4574 & (forvar4580[(3'h7):(3'h4)] ?
                          (forvar4694[(1'h1):(1'h1)] | reg4722) : (8'h9d)));
                      reg4761 <= (8'ha9);
                      reg4762 <= reg4590;
                    end
                  for (forvar4763 = (1'h0); (forvar4763 < (1'h1)); forvar4763 = (forvar4763 + (1'h1)))
                    begin
                      reg4764 <= (8'hb3);
                      reg4765 <= forvar4759[(3'h7):(1'h1)];
                      reg4766 <= reg4587;
                    end
                end
              else
                begin
                  for (forvar4758 = (1'h0); (forvar4758 < (2'h3)); forvar4758 = (forvar4758 + (1'h1)))
                    begin
                      reg4759 <= $signed({{$signed(reg4660)}});
                      reg4760 <= (~&{({reg4603} ?
                              (~^forvar4673) : $unsigned(forvar4624))});
                      reg4761 <= ((+{$unsigned(reg4645)}) ?
                          (reg4603[(5'h10):(3'h4)] >= (8'ha7)) : ((&forvar4738[(1'h0):(1'h0)]) - ((~forvar4591) && $signed(reg4750))));
                      reg4762 <= $signed((~^{(reg4644 >= (8'hb8))}));
                    end
                  if ((8'hb3))
                    begin
                      reg4763 <= ((!forvar4727[(3'h4):(1'h1)]) ?
                          (8'hb1) : (!reg4590[(4'h9):(1'h1)]));
                      reg4764 <= (~^(((forvar4745 ^~ reg4595) ?
                          reg4742 : (^~reg4715)) * ($unsigned(reg4724) < $signed(forvar4650))));
                      reg4765 <= {(-reg4718[(1'h1):(1'h0)])};
                      reg4766 <= (8'h9c);
                    end
                  else
                    begin
                      reg4763 <= (!(((8'ha4) ^~ reg4590[(4'h9):(3'h4)]) ?
                          ((reg4693 - forvar4624) == (forvar4578 ?
                              (8'hb3) : reg4606)) : ($unsigned((8'hb0)) & $unsigned(reg4727))));
                      reg4764 <= $signed(((~&$signed(reg4746)) - {$signed(reg4593)}));
                    end
                  if ($signed($signed(forvar4613[(4'ha):(4'h9)])))
                    begin
                      reg4767 <= ($unsigned((|reg4699[(3'h6):(3'h4)])) ?
                          $unsigned(((reg4739 ?
                              reg4675 : reg4676) >> reg4719[(3'h5):(1'h1)])) : (~reg4736));
                    end
                  else
                    begin
                      reg4767 <= (8'hab);
                      reg4768 <= reg4649[(2'h3):(1'h1)];
                      reg4769 <= forvar4593[(2'h3):(2'h2)];
                    end
                  for (forvar4770 = (1'h0); (forvar4770 < (2'h2)); forvar4770 = (forvar4770 + (1'h1)))
                    begin
                      reg4771 <= ($unsigned(((reg4645 + forvar4689) ^ forvar4603)) ^ {reg4740[(2'h2):(2'h2)]});
                      reg4772 <= ({((&reg4707) <= reg4651[(1'h1):(1'h1)])} ?
                          $unsigned(reg4601[(3'h7):(2'h3)]) : $signed((^~(^~forvar4712))));
                    end
                end
              for (forvar4773 = (1'h0); (forvar4773 < (2'h2)); forvar4773 = (forvar4773 + (1'h1)))
                begin
                  reg4774 <= ($unsigned($unsigned(wire4574[(3'h4):(3'h4)])) ^ reg4630);
                end
              for (forvar4775 = (1'h0); (forvar4775 < (2'h3)); forvar4775 = (forvar4775 + (1'h1)))
                begin
                  if (($signed($signed(reg4660)) ?
                      (forvar4579 || ((-(8'hb0)) <<< $signed((8'ha3)))) : ((|$signed((8'ha8))) >= $unsigned(reg4660))))
                    begin
                      reg4776 <= {$unsigned({$signed(reg4686)})};
                      reg4777 <= reg4753[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg4776 <= {forvar4725[(2'h2):(1'h1)]};
                      reg4777 <= ((+(reg4584[(1'h0):(1'h0)] == (~|reg4579))) ?
                          ((!(~|(8'haa))) ?
                              ((reg4661 ? forvar4681 : reg4642) ?
                                  (~reg4583) : reg4670) : (!reg4619)) : reg4630);
                      reg4778 <= ($unsigned(reg4759) ?
                          (($signed(reg4665) && $unsigned(reg4605)) ~^ ((forvar4617 ?
                                  forvar4617 : (8'hb2)) ?
                              forvar4674 : $unsigned(forvar4642))) : (8'hb9));
                    end
                end
            end
          else
            begin
              reg4745 <= (^$unsigned((reg4771 ?
                  (+reg4707) : forvar4715[(3'h6):(3'h6)])));
              if (forvar4607[(2'h2):(2'h2)])
                begin
                  for (forvar4746 = (1'h0); (forvar4746 < (2'h2)); forvar4746 = (forvar4746 + (1'h1)))
                    begin
                      reg4747 <= (~^($signed($unsigned(reg4692)) || reg4760[(4'hb):(4'h8)]));
                      reg4748 <= (((reg4769 ?
                              (+reg4610) : reg4604) | $unsigned((8'ha2))) ?
                          $unsigned($signed((reg4687 ?
                              reg4607 : reg4686))) : reg4765);
                      reg4749 <= reg4733;
                      reg4750 <= $unsigned((!$signed((^~forvar4746))));
                    end
                  reg4751 <= ((^~(8'ha8)) - (^~(~&forvar4717)));
                  reg4752 <= ((reg4691[(3'h7):(3'h6)] >> ((reg4740 ?
                          (8'hb0) : forvar4592) < forvar4584[(2'h2):(2'h2)])) ?
                      $unsigned({$unsigned(reg4635)}) : {$signed((reg4645 ?
                              reg4630 : reg4731))});
                end
              else
                begin
                  if (({reg4579[(4'hb):(4'hb)]} >>> (((reg4680 ?
                          (8'ha6) : reg4612) ?
                      $unsigned(forvar4650) : $signed(reg4702)) * $signed({forvar4676}))))
                    begin
                      reg4746 <= $unsigned($signed($unsigned(forvar4673[(1'h0):(1'h0)])));
                      reg4747 <= (reg4623 ? reg4647 : (8'hb4));
                      reg4748 <= (($signed((&reg4667)) != reg4655) ?
                          (~&wire4575) : ($unsigned(forvar4652[(1'h0):(1'h0)]) ?
                              forvar4581 : $unsigned(((8'hba) * reg4671))));
                    end
                  else
                    begin
                      reg4746 <= $unsigned($signed($unsigned((reg4628 || forvar4616))));
                    end
                  if ((forvar4705 ? {{reg4715}} : reg4589))
                    begin
                      reg4749 <= reg4642;
                    end
                  else
                    begin
                      reg4749 <= (($signed((+reg4691)) ?
                              ($unsigned(reg4749) ?
                                  (reg4615 && (8'ha4)) : (reg4655 ?
                                      reg4716 : reg4735)) : (((8'h9d) >> reg4594) ?
                                  $unsigned(reg4654) : (~|forvar4640))) ?
                          forvar4640[(1'h0):(1'h0)] : $signed($unsigned($unsigned(forvar4594))));
                      reg4750 <= $unsigned(reg4701);
                      reg4751 <= $signed(reg4579);
                    end
                end
              for (forvar4753 = (1'h0); (forvar4753 < (1'h0)); forvar4753 = (forvar4753 + (1'h1)))
                begin
                  reg4754 <= ((~^forvar4737) * {forvar4640});
                  for (forvar4755 = (1'h0); (forvar4755 < (1'h0)); forvar4755 = (forvar4755 + (1'h1)))
                    begin
                      reg4756 <= {reg4678};
                      reg4757 <= $unsigned((((reg4722 << reg4734) ?
                              reg4593[(3'h4):(2'h3)] : (reg4756 ~^ reg4778)) ?
                          ({reg4711} ?
                              (reg4662 ~^ reg4701) : $signed((8'h9e))) : (~|reg4600[(4'h8):(3'h4)])));
                    end
                  for (forvar4758 = (1'h0); (forvar4758 < (1'h0)); forvar4758 = (forvar4758 + (1'h1)))
                    begin
                      reg4759 <= (reg4676 ?
                          $unsigned($signed((+reg4611))) : (8'hac));
                      reg4760 <= ($unsigned(((reg4601 ?
                              reg4602 : (8'h9e)) ^ (reg4655 | reg4777))) ?
                          ($signed((reg4777 ?
                              (8'had) : forvar4636)) && $signed(reg4623)) : $signed(forvar4717[(3'h6):(1'h0)]));
                      reg4761 <= $unsigned(reg4594[(3'h4):(2'h2)]);
                    end
                  if (reg4714)
                    begin
                      reg4762 <= reg4701;
                    end
                  else
                    begin
                      reg4762 <= $signed($unsigned(((reg4583 * (8'hb3)) + {(8'hb7)})));
                      reg4763 <= $signed({((!reg4645) == {reg4596})});
                      reg4764 <= ($unsigned(reg4633[(3'h4):(1'h1)]) ?
                          reg4592[(2'h3):(2'h3)] : (reg4746 ^~ reg4643[(1'h0):(1'h0)]));
                    end
                end
            end
          for (forvar4779 = (1'h0); (forvar4779 < (2'h3)); forvar4779 = (forvar4779 + (1'h1)))
            begin
              for (forvar4780 = (1'h0); (forvar4780 < (2'h3)); forvar4780 = (forvar4780 + (1'h1)))
                begin
                  if (((8'hba) ~^ $signed((~|(reg4651 ? reg4680 : (8'hb3))))))
                    begin
                      reg4781 <= $signed($unsigned($unsigned(reg4631)));
                      reg4782 <= $unsigned($unsigned(forvar4581[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg4781 <= forvar4581;
                      reg4782 <= reg4687[(3'h7):(3'h7)];
                    end
                  reg4783 <= reg4753;
                end
              reg4784 <= {(((forvar4749 ? (8'ha6) : forvar4579) >> forvar4604) ?
                      $unsigned(reg4715[(3'h4):(2'h2)]) : (|(&reg4709)))};
            end
          for (forvar4785 = (1'h0); (forvar4785 < (2'h2)); forvar4785 = (forvar4785 + (1'h1)))
            begin
              if (reg4675)
                begin
                  for (forvar4786 = (1'h0); (forvar4786 < (1'h0)); forvar4786 = (forvar4786 + (1'h1)))
                    begin
                      reg4787 <= (+forvar4636);
                      reg4788 <= $unsigned(($unsigned($signed(reg4733)) ?
                          reg4603[(4'ha):(3'h6)] : reg4732[(3'h6):(3'h6)]));
                      reg4789 <= reg4767[(4'hb):(2'h3)];
                      reg4790 <= reg4752[(4'h9):(3'h4)];
                    end
                end
              else
                begin
                  if ($signed((^forvar4717[(4'hf):(4'he)])))
                    begin
                      reg4786 <= $signed(forvar4727[(3'h5):(2'h2)]);
                      reg4787 <= ((~(8'ha2)) ^~ $unsigned(((~|(8'ha2)) - ((8'hac) ?
                          reg4605 : reg4725))));
                      reg4788 <= (~&forvar4694[(3'h6):(1'h0)]);
                    end
                  else
                    begin
                      reg4786 <= reg4637[(3'h5):(2'h2)];
                      reg4787 <= $signed(((reg4583 >= {forvar4758}) < {$signed(forvar4733)}));
                    end
                  if ($unsigned($unsigned(forvar4738[(1'h1):(1'h1)])))
                    begin
                      reg4789 <= $signed(reg4741[(2'h3):(1'h0)]);
                      reg4790 <= (-((8'h9c) - (~|reg4614)));
                      reg4791 <= ((!wire4574[(4'h9):(2'h3)]) && reg4731[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg4789 <= ($unsigned((((8'ha8) && (8'hb0)) ~^ $signed((8'ha8)))) ?
                          reg4580[(3'h7):(3'h4)] : reg4760[(3'h7):(2'h3)]);
                    end
                  if ((({(^~forvar4717)} | $unsigned((forvar4727 < reg4755))) * $unsigned($unsigned({reg4622}))))
                    begin
                      reg4792 <= $signed({((reg4759 ?
                              reg4755 : reg4747) >> ((8'haf) ?
                              reg4713 : reg4596))});
                      reg4793 <= (reg4603[(4'ha):(4'ha)] ?
                          $signed(($unsigned(forvar4624) ?
                              $unsigned(reg4726) : forvar4654[(2'h3):(2'h3)])) : $unsigned(forvar4698));
                      reg4794 <= (reg4656 <= forvar4676[(4'h8):(1'h1)]);
                    end
                  else
                    begin
                      reg4792 <= $signed((&$signed({reg4600})));
                      reg4793 <= (reg4621[(2'h2):(1'h0)] - $unsigned(((8'hb2) - (reg4777 & forvar4673))));
                    end
                  for (forvar4795 = (1'h0); (forvar4795 < (2'h2)); forvar4795 = (forvar4795 + (1'h1)))
                    begin
                      reg4796 <= $unsigned($signed($unsigned($unsigned(reg4599))));
                      reg4797 <= $signed(($signed($unsigned((8'hb6))) ?
                          $signed((reg4671 ? forvar4581 : reg4658)) : reg4693));
                    end
                end
            end
        end
      else
        begin
          for (forvar4737 = (1'h0); (forvar4737 < (2'h3)); forvar4737 = (forvar4737 + (1'h1)))
            begin
              for (forvar4738 = (1'h0); (forvar4738 < (2'h2)); forvar4738 = (forvar4738 + (1'h1)))
                begin
                  reg4739 <= $unsigned(reg4635[(3'h4):(1'h1)]);
                  reg4740 <= forvar4749;
                  for (forvar4741 = (1'h0); (forvar4741 < (1'h1)); forvar4741 = (forvar4741 + (1'h1)))
                    begin
                      reg4742 <= $unsigned(((~&(reg4636 ?
                          (8'ha9) : reg4707)) | reg4680));
                      reg4743 <= reg4684;
                    end
                end
              for (forvar4744 = (1'h0); (forvar4744 < (2'h2)); forvar4744 = (forvar4744 + (1'h1)))
                begin
                  reg4745 <= $unsigned((^~reg4755));
                end
              for (forvar4746 = (1'h0); (forvar4746 < (2'h3)); forvar4746 = (forvar4746 + (1'h1)))
                begin
                  reg4747 <= {(reg4702 ?
                          reg4667[(4'ha):(4'h9)] : (reg4678 + (reg4695 ?
                              (8'ha0) : forvar4759)))};
                  for (forvar4748 = (1'h0); (forvar4748 < (1'h0)); forvar4748 = (forvar4748 + (1'h1)))
                    begin
                      reg4749 <= {reg4691[(3'h4):(1'h0)]};
                    end
                  for (forvar4750 = (1'h0); (forvar4750 < (2'h3)); forvar4750 = (forvar4750 + (1'h1)))
                    begin
                      reg4751 <= reg4794[(2'h3):(1'h1)];
                      reg4752 <= reg4730[(4'hc):(4'h9)];
                    end
                  for (forvar4753 = (1'h0); (forvar4753 < (2'h3)); forvar4753 = (forvar4753 + (1'h1)))
                    begin
                      reg4754 <= wire4573;
                      reg4755 <= $signed(reg4671);
                      reg4756 <= reg4611[(3'h4):(1'h1)];
                      reg4757 <= (|{((~forvar4603) * {(8'ha1)})});
                    end
                end
              reg4758 <= {(((reg4729 ?
                          forvar4738 : reg4744) > $unsigned(reg4584)) ?
                      reg4734 : reg4600[(1'h0):(1'h0)])};
            end
          if ((~|forvar4610))
            begin
              if ((~|reg4702[(1'h0):(1'h0)]))
                begin
                  if (reg4719[(4'h8):(2'h3)])
                    begin
                      reg4759 <= reg4671[(1'h1):(1'h1)];
                      reg4760 <= $signed($unsigned({reg4794}));
                      reg4761 <= ((($unsigned(reg4592) ?
                          $signed(reg4767) : ((8'hb3) >>> forvar4674)) <<< (~|$signed(reg4718))) - $signed($unsigned($signed(reg4679))));
                      reg4762 <= ($signed(($signed((8'haf)) < $signed(reg4709))) ?
                          ($unsigned(forvar4676) << $signed(((8'h9f) ^~ reg4586))) : $unsigned((~&$signed(reg4604))));
                    end
                  else
                    begin
                      reg4759 <= (8'hac);
                      reg4760 <= (reg4786[(1'h0):(1'h0)] != forvar4592);
                    end
                  if ($unsigned((|reg4714[(4'h9):(3'h6)])))
                    begin
                      reg4763 <= $unsigned(reg4692[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg4763 <= (forvar4727[(3'h4):(3'h4)] ?
                          {$unsigned((reg4690 ?
                                  forvar4663 : reg4586))} : (($signed(reg4735) ?
                              $signed(reg4632) : (8'haf)) <<< $unsigned({(8'hb3)})));
                      reg4764 <= (~&$unsigned(((forvar4643 ?
                              reg4760 : (8'ha9)) ?
                          $signed(reg4786) : (^reg4636))));
                    end
                end
              else
                begin
                  reg4759 <= (({(forvar4593 != forvar4654)} < ((8'hb7) == $signed(forvar4607))) ?
                      (~^$signed($signed((8'hb9)))) : ((8'hb9) << reg4657));
                  if ($unsigned((((reg4720 ?
                      reg4728 : forvar4674) ^~ (|forvar4717)) || reg4701)))
                    begin
                      reg4760 <= (reg4760 ?
                          (((reg4637 ?
                                  (8'hac) : reg4704) >> reg4738[(2'h2):(2'h2)]) ?
                              {$unsigned((8'haa))} : $unsigned(reg4661[(3'h5):(3'h4)])) : (reg4670[(1'h0):(1'h0)] ?
                              {reg4697} : forvar4694));
                      reg4761 <= {((forvar4717[(2'h3):(2'h2)] | (reg4595 - reg4691)) >> forvar4737)};
                      reg4762 <= $unsigned(((8'hb8) >> reg4689));
                    end
                  else
                    begin
                      reg4760 <= $signed($signed((~&reg4627)));
                    end
                end
            end
          else
            begin
              for (forvar4759 = (1'h0); (forvar4759 < (1'h1)); forvar4759 = (forvar4759 + (1'h1)))
                begin
                  for (forvar4760 = (1'h0); (forvar4760 < (2'h3)); forvar4760 = (forvar4760 + (1'h1)))
                    begin
                      reg4761 <= $signed((+reg4766[(1'h0):(1'h0)]));
                      reg4762 <= $unsigned((reg4693[(1'h1):(1'h0)] ?
                          (!$unsigned((8'haf))) : forvar4642[(1'h0):(1'h0)]));
                      reg4763 <= reg4622;
                    end
                  if ($signed(reg4709))
                    begin
                      reg4764 <= ($unsigned({forvar4609[(1'h1):(1'h0)]}) ?
                          $unsigned(reg4662) : ((forvar4659 && $signed(reg4587)) <<< forvar4592));
                    end
                  else
                    begin
                      reg4764 <= (forvar4598[(4'hd):(2'h3)] ?
                          reg4739[(1'h1):(1'h0)] : reg4772);
                      reg4765 <= reg4586;
                    end
                end
            end
          if ($signed($unsigned((forvar4773 * (^reg4730)))))
            begin
              if ((~|$unsigned($unsigned($unsigned(forvar4749)))))
                begin
                  if ($unsigned(reg4645))
                    begin
                      reg4766 <= ({reg4759} ?
                          $signed($unsigned(forvar4608[(3'h4):(1'h1)])) : (-(&((8'hb6) ?
                              reg4742 : reg4739))));
                      reg4767 <= ((~|{$unsigned((8'hb9))}) != $unsigned(($signed(reg4771) | (8'ha9))));
                      reg4768 <= (^(^~forvar4674[(3'h5):(1'h0)]));
                    end
                  else
                    begin
                      reg4766 <= $unsigned(($signed($unsigned(forvar4760)) - $unsigned($signed((8'ha6)))));
                      reg4767 <= $signed((reg4757 ?
                          ((reg4595 ?
                              reg4699 : (8'hb5)) >>> (^forvar4609)) : ((forvar4578 ?
                                  reg4646 : forvar4672) ?
                              forvar4578[(1'h1):(1'h0)] : (reg4601 + (8'hb1)))));
                    end
                  if (reg4665[(3'h6):(3'h4)])
                    begin
                      reg4769 <= reg4765;
                      reg4770 <= forvar4652;
                      reg4771 <= ($signed(($unsigned(reg4654) - {reg4724})) ?
                          wire4576[(2'h3):(2'h2)] : $signed($signed($signed((8'hb4)))));
                      reg4772 <= (|forvar4610[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg4769 <= $signed((((reg4781 ?
                              (8'ha8) : reg4747) ^ reg4599[(3'h7):(1'h1)]) ?
                          $unsigned($signed((8'h9f))) : reg4670));
                      reg4770 <= reg4734[(2'h3):(2'h2)];
                    end
                  for (forvar4773 = (1'h0); (forvar4773 < (1'h0)); forvar4773 = (forvar4773 + (1'h1)))
                    begin
                      reg4774 <= reg4589[(3'h6):(3'h4)];
                      reg4775 <= (($unsigned($signed((8'ha1))) >>> ($signed(forvar4741) || forvar4775[(2'h2):(1'h0)])) ?
                          {$signed(reg4753)} : (|($unsigned((8'ha2)) ?
                              forvar4643[(4'hb):(3'h5)] : forvar4795)));
                      reg4776 <= (forvar4744 ?
                          {((|reg4615) ?
                                  forvar4779 : $signed(forvar4579))} : reg4690);
                    end
                  for (forvar4777 = (1'h0); (forvar4777 < (1'h0)); forvar4777 = (forvar4777 + (1'h1)))
                    begin
                      reg4778 <= forvar4640;
                      reg4779 <= reg4714[(1'h1):(1'h0)];
                      reg4780 <= reg4633[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar4766 = (1'h0); (forvar4766 < (1'h1)); forvar4766 = (forvar4766 + (1'h1)))
                    begin
                      reg4767 <= (^reg4662);
                    end
                  for (forvar4768 = (1'h0); (forvar4768 < (1'h1)); forvar4768 = (forvar4768 + (1'h1)))
                    begin
                      reg4769 <= forvar4694;
                    end
                end
              for (forvar4781 = (1'h0); (forvar4781 < (2'h2)); forvar4781 = (forvar4781 + (1'h1)))
                begin
                  if (({((^~(8'hb8)) ? reg4644 : (~|forvar4636))} ?
                      (8'ha1) : $unsigned((reg4734 ?
                          $signed(reg4682) : $unsigned(reg4632)))))
                    begin
                      reg4782 <= reg4768[(3'h4):(3'h4)];
                      reg4783 <= reg4719[(4'hc):(4'h9)];
                    end
                  else
                    begin
                      reg4782 <= {$signed($unsigned($signed(reg4683)))};
                      reg4783 <= $signed((~&(reg4771 ?
                          (+reg4766) : $signed(reg4624))));
                      reg4784 <= $signed($unsigned($signed(reg4634[(1'h0):(1'h0)])));
                    end
                  for (forvar4785 = (1'h0); (forvar4785 < (2'h3)); forvar4785 = (forvar4785 + (1'h1)))
                    begin
                      reg4786 <= reg4749[(4'hf):(4'hd)];
                      reg4787 <= (~^reg4745[(3'h6):(1'h0)]);
                      reg4788 <= reg4626;
                    end
                  for (forvar4789 = (1'h0); (forvar4789 < (1'h1)); forvar4789 = (forvar4789 + (1'h1)))
                    begin
                      reg4790 <= (&forvar4777[(3'h6):(3'h6)]);
                    end
                  if ($signed((|reg4646)))
                    begin
                      reg4791 <= $unsigned(reg4594);
                      reg4792 <= {($unsigned({(8'ha7)}) && $unsigned({reg4735}))};
                      reg4793 <= ($unsigned((~&(reg4706 ?
                              reg4794 : forvar4609))) ?
                          reg4719[(3'h7):(3'h6)] : (((|(8'ha9)) ^~ (reg4637 + (8'hb1))) >> $unsigned(((8'ha4) ?
                              reg4664 : forvar4705))));
                    end
                  else
                    begin
                      reg4791 <= $signed(reg4780[(3'h4):(1'h0)]);
                      reg4792 <= $unsigned({reg4682[(2'h3):(2'h2)]});
                      reg4793 <= $unsigned(reg4759[(4'hd):(4'h8)]);
                    end
                end
              reg4794 <= reg4580[(4'hc):(1'h0)];
            end
          else
            begin
              for (forvar4766 = (1'h0); (forvar4766 < (2'h2)); forvar4766 = (forvar4766 + (1'h1)))
                begin
                  if (reg4586[(4'h8):(4'h8)])
                    begin
                      reg4767 <= {(((forvar4773 ^~ (8'ha0)) << $unsigned(forvar4610)) > {{reg4763}})};
                    end
                  else
                    begin
                      reg4767 <= ({(-(|reg4655))} ?
                          reg4656 : {reg4791[(3'h5):(2'h2)]});
                    end
                  if (($unsigned(reg4582[(1'h1):(1'h0)]) >>> (+((+(8'hab)) == (reg4757 | forvar4598)))))
                    begin
                      reg4768 <= (forvar4640[(2'h2):(1'h0)] ?
                          $signed({reg4708[(1'h1):(1'h0)]}) : $unsigned($unsigned(reg4787)));
                    end
                  else
                    begin
                      reg4768 <= $signed({$signed($unsigned((8'ha0)))});
                      reg4769 <= $unsigned(($signed($unsigned(reg4719)) != $unsigned($signed(reg4745))));
                      reg4770 <= $unsigned($signed($unsigned(forvar4748[(3'h6):(1'h0)])));
                    end
                end
              if (reg4754)
                begin
                  for (forvar4771 = (1'h0); (forvar4771 < (1'h0)); forvar4771 = (forvar4771 + (1'h1)))
                    begin
                      reg4772 <= (reg4783 ?
                          ((8'ha4) || (~&$unsigned(reg4757))) : $signed(wire4573[(3'h5):(2'h3)]));
                    end
                  reg4773 <= (($unsigned((~(8'h9c))) <= reg4745[(4'h9):(2'h3)]) < ($unsigned({reg4752}) != $unsigned(reg4612)));
                end
              else
                begin
                  if ($unsigned((^~$unsigned($signed(forvar4640)))))
                    begin
                      reg4771 <= (reg4629[(3'h5):(2'h3)] || {$unsigned(reg4727[(1'h0):(1'h0)])});
                      reg4772 <= forvar4759[(3'h7):(1'h1)];
                    end
                  else
                    begin
                      reg4771 <= (8'h9f);
                      reg4772 <= forvar4775;
                      reg4773 <= reg4766;
                      reg4774 <= reg4735;
                    end
                end
              reg4775 <= reg4725[(1'h0):(1'h0)];
            end
        end
    end
  assign wire4798 = $unsigned({(8'had)});
  assign wire4799 = ((~^$signed(reg4589[(1'h1):(1'h1)])) ?
                        ($signed((-reg4732)) ?
                            {(-forvar4715)} : reg4734) : (reg4619[(2'h2):(1'h1)] ?
                            ((~&(8'ha2)) >= (^reg4769)) : (forvar4777[(2'h2):(1'h0)] != (^~reg4624))));
  always
    @(posedge clk) begin
      reg4800 <= ($signed($signed($unsigned(reg4791))) == reg4656);
    end
  always
    @(posedge clk) begin
      for (forvar4801 = (1'h0); (forvar4801 < (2'h2)); forvar4801 = (forvar4801 + (1'h1)))
        begin
          for (forvar4802 = (1'h0); (forvar4802 < (1'h0)); forvar4802 = (forvar4802 + (1'h1)))
            begin
              if ($unsigned($signed(reg4655[(1'h1):(1'h1)])))
                begin
                  if (reg4786[(1'h0):(1'h0)])
                    begin
                      reg4803 <= $signed(($signed((reg4777 ?
                          reg4627 : reg4784)) ~^ (reg4645 <= (8'ha7))));
                      reg4804 <= (|$unsigned($signed(forvar4698[(4'h9):(1'h0)])));
                      reg4805 <= ($signed($signed((reg4726 ?
                              forvar4654 : reg4759))) ?
                          (reg4735 ?
                              $unsigned((!reg4770)) : reg4661[(3'h6):(1'h0)]) : $signed($signed((reg4634 ?
                              reg4608 : (8'haa)))));
                    end
                  else
                    begin
                      reg4803 <= (reg4584 & $unsigned({reg4622[(3'h5):(3'h5)]}));
                      reg4804 <= ((+reg4765) ?
                          forvar4763 : forvar4610[(3'h5):(3'h5)]);
                      reg4805 <= (|reg4746[(3'h6):(1'h1)]);
                    end
                  for (forvar4806 = (1'h0); (forvar4806 < (1'h0)); forvar4806 = (forvar4806 + (1'h1)))
                    begin
                      reg4807 <= (reg4668 ? reg4579 : $signed((-(+reg4658))));
                      reg4808 <= ({reg4606} ~^ reg4701[(2'h2):(1'h0)]);
                    end
                  for (forvar4809 = (1'h0); (forvar4809 < (1'h0)); forvar4809 = (forvar4809 + (1'h1)))
                    begin
                      reg4810 <= (({(reg4762 ?
                                  reg4715 : reg4729)} ^~ {$unsigned((8'hac))}) ?
                          reg4741 : {(^reg4770)});
                      reg4811 <= ({$signed((reg4782 << (8'ha3)))} ?
                          $signed(((|reg4723) ?
                              (reg4768 ?
                                  forvar4694 : reg4775) : (reg4623 & reg4764))) : forvar4748);
                    end
                end
              else
                begin
                  if ((reg4729[(3'h5):(2'h2)] ?
                      (forvar4603[(3'h4):(3'h4)] & (reg4679[(4'hc):(4'hc)] ?
                          $signed(reg4774) : reg4733)) : $unsigned(((reg4724 <<< reg4691) + (reg4701 ?
                          reg4782 : forvar4773)))))
                    begin
                      reg4803 <= reg4789;
                      reg4804 <= (8'ha8);
                    end
                  else
                    begin
                      reg4803 <= $unsigned($signed(reg4637[(3'h7):(1'h0)]));
                    end
                end
              reg4812 <= $unsigned(($signed((^reg4590)) ?
                  reg4682[(1'h0):(1'h0)] : (((8'ha0) ? reg4792 : forvar4760) ?
                      $unsigned(forvar4652) : $signed(reg4726))));
            end
        end
      for (forvar4813 = (1'h0); (forvar4813 < (2'h3)); forvar4813 = (forvar4813 + (1'h1)))
        begin
          for (forvar4814 = (1'h0); (forvar4814 < (1'h1)); forvar4814 = (forvar4814 + (1'h1)))
            begin
              for (forvar4815 = (1'h0); (forvar4815 < (2'h2)); forvar4815 = (forvar4815 + (1'h1)))
                begin
                  reg4816 <= $signed($signed((reg4763 ?
                      {(8'h9d)} : forvar4672)));
                  for (forvar4817 = (1'h0); (forvar4817 < (1'h0)); forvar4817 = (forvar4817 + (1'h1)))
                    begin
                      reg4818 <= reg4769[(2'h2):(2'h2)];
                    end
                  for (forvar4819 = (1'h0); (forvar4819 < (2'h3)); forvar4819 = (forvar4819 + (1'h1)))
                    begin
                      reg4820 <= ($signed(reg4646) ?
                          $signed({reg4638}) : $signed($signed((reg4790 << (8'hb8)))));
                      reg4821 <= (((^~(reg4704 < forvar4731)) ?
                              (8'hb1) : ({(8'hac)} >> $signed((8'ha8)))) ?
                          $signed($signed((reg4750 ?
                              reg4646 : reg4661))) : (~|{(wire4574 ?
                                  (8'ha2) : reg4697)}));
                      reg4822 <= (reg4762[(4'hd):(4'hc)] || reg4585[(3'h7):(3'h4)]);
                      reg4823 <= ((8'ha2) ? (8'hb1) : (~(&forvar4593)));
                    end
                  for (forvar4824 = (1'h0); (forvar4824 < (2'h3)); forvar4824 = (forvar4824 + (1'h1)))
                    begin
                      reg4825 <= ($unsigned((8'hb1)) ?
                          (reg4590 >> ((^reg4660) << reg4647)) : reg4602);
                    end
                end
              for (forvar4826 = (1'h0); (forvar4826 < (2'h3)); forvar4826 = (forvar4826 + (1'h1)))
                begin
                  for (forvar4827 = (1'h0); (forvar4827 < (2'h3)); forvar4827 = (forvar4827 + (1'h1)))
                    begin
                      reg4828 <= (reg4687 >= reg4686);
                    end
                  for (forvar4829 = (1'h0); (forvar4829 < (1'h0)); forvar4829 = (forvar4829 + (1'h1)))
                    begin
                      reg4830 <= reg4601;
                      reg4831 <= (reg4742 ?
                          ($signed((^(8'haa))) ?
                              (~^reg4770[(1'h1):(1'h0)]) : ($signed(forvar4705) ?
                                  (reg4709 ^ reg4761) : reg4626)) : $unsigned($unsigned($signed(reg4702))));
                      reg4832 <= $unsigned($signed(reg4682[(3'h5):(2'h2)]));
                    end
                  if ((reg4711 ?
                      ($signed((~&(8'hb8))) ?
                          (!(+reg4732)) : reg4597[(4'hb):(1'h1)]) : (|forvar4733)))
                    begin
                      reg4833 <= (~^{((8'hb5) ?
                              {reg4590} : $unsigned((8'hba)))});
                      reg4834 <= (!{((reg4595 << forvar4609) << reg4625)});
                      reg4835 <= reg4671;
                      reg4836 <= forvar4610[(3'h4):(3'h4)];
                    end
                  else
                    begin
                      reg4833 <= ($unsigned((8'hae)) ?
                          $unsigned($signed(forvar4815)) : (((!reg4577) ?
                                  reg4742 : {reg4745}) ?
                              (~{reg4821}) : (8'hb9)));
                      reg4834 <= (^$unsigned((-forvar4578)));
                    end
                end
            end
          if ($unsigned($signed(($unsigned((8'h9e)) ^ (+(8'hac))))))
            begin
              reg4837 <= reg4738;
              reg4838 <= (!(8'h9f));
              if ($unsigned($signed(reg4807)))
                begin
                  for (forvar4839 = (1'h0); (forvar4839 < (2'h2)); forvar4839 = (forvar4839 + (1'h1)))
                    begin
                      reg4840 <= (~(8'ha4));
                      reg4841 <= {reg4723[(3'h5):(1'h1)]};
                    end
                  if ({($unsigned(reg4662[(1'h0):(1'h0)]) ?
                          ((reg4654 ?
                              forvar4785 : reg4611) > ((8'ha4) + (8'haf))) : ($unsigned(reg4610) && (~^reg4631)))})
                    begin
                      reg4842 <= $signed($signed($unsigned((reg4577 ^ reg4758))));
                    end
                  else
                    begin
                      reg4842 <= $unsigned(($unsigned($signed(reg4744)) ?
                          reg4679[(3'h6):(3'h5)] : (~^{(8'hb7)})));
                    end
                  for (forvar4843 = (1'h0); (forvar4843 < (2'h3)); forvar4843 = (forvar4843 + (1'h1)))
                    begin
                      reg4844 <= forvar4809;
                    end
                end
              else
                begin
                  for (forvar4839 = (1'h0); (forvar4839 < (2'h2)); forvar4839 = (forvar4839 + (1'h1)))
                    begin
                      reg4840 <= $signed($unsigned((~&(reg4784 >> reg4590))));
                      reg4841 <= reg4837;
                      reg4842 <= reg4721;
                    end
                  for (forvar4843 = (1'h0); (forvar4843 < (1'h1)); forvar4843 = (forvar4843 + (1'h1)))
                    begin
                      reg4844 <= (-(({reg4731} && (reg4784 ?
                              reg4591 : reg4710)) ?
                          forvar4581 : forvar4648[(2'h2):(1'h1)]));
                      reg4845 <= (8'ha9);
                      reg4846 <= reg4581[(3'h4):(1'h1)];
                      reg4847 <= reg4781;
                    end
                  for (forvar4848 = (1'h0); (forvar4848 < (1'h0)); forvar4848 = (forvar4848 + (1'h1)))
                    begin
                      reg4849 <= (&reg4758);
                    end
                end
              for (forvar4850 = (1'h0); (forvar4850 < (2'h3)); forvar4850 = (forvar4850 + (1'h1)))
                begin
                  for (forvar4851 = (1'h0); (forvar4851 < (2'h2)); forvar4851 = (forvar4851 + (1'h1)))
                    begin
                      reg4852 <= reg4647[(1'h1):(1'h1)];
                    end
                  reg4853 <= reg4613[(2'h2):(1'h0)];
                end
            end
          else
            begin
              if (($signed(reg4596) ?
                  ($signed((8'ha6)) ^ (8'hb5)) : (((reg4628 + forvar4753) + (reg4846 < (8'hb4))) & (reg4721 >= reg4703[(1'h0):(1'h0)]))))
                begin
                  for (forvar4837 = (1'h0); (forvar4837 < (1'h0)); forvar4837 = (forvar4837 + (1'h1)))
                    begin
                      reg4838 <= ((forvar4578[(1'h1):(1'h1)] ^ (reg4691 ^~ (wire4798 ?
                          (8'hb2) : reg4676))) + $unsigned((^~{reg4780})));
                    end
                  reg4839 <= {$signed(((|(8'hb8)) ?
                          (~|reg4740) : (forvar4602 & reg4842)))};
                  for (forvar4840 = (1'h0); (forvar4840 < (2'h2)); forvar4840 = (forvar4840 + (1'h1)))
                    begin
                      reg4841 <= reg4847[(1'h0):(1'h0)];
                      reg4842 <= forvar4827[(1'h1):(1'h0)];
                    end
                  if (($unsigned(reg4723[(3'h6):(3'h6)]) ?
                      reg4597[(1'h1):(1'h0)] : $unsigned(reg4805)))
                    begin
                      reg4843 <= $signed((+$signed($signed(reg4593))));
                      reg4844 <= $signed(forvar4748);
                      reg4845 <= reg4804;
                      reg4846 <= (&$unsigned(($unsigned((8'hb2)) ?
                          reg4627 : (forvar4744 & reg4784))));
                    end
                  else
                    begin
                      reg4843 <= forvar4588[(2'h2):(1'h1)];
                      reg4844 <= {reg4770};
                      reg4845 <= ((reg4580 ?
                              ((reg4620 ? reg4750 : forvar4663) ?
                                  (~&forvar4785) : reg4844[(1'h0):(1'h0)]) : ((~|reg4773) ?
                                  (reg4720 == (8'ha9)) : (reg4692 ?
                                      forvar4610 : reg4731))) ?
                          ($unsigned((forvar4781 ?
                              forvar4819 : reg4807)) >> reg4676) : reg4613[(1'h1):(1'h0)]);
                      reg4846 <= $signed(((~|reg4835[(3'h4):(2'h3)]) < ((forvar4652 == forvar4745) ?
                          reg4580[(3'h4):(2'h3)] : (&forvar4598))));
                    end
                end
              else
                begin
                  for (forvar4837 = (1'h0); (forvar4837 < (2'h3)); forvar4837 = (forvar4837 + (1'h1)))
                    begin
                      reg4838 <= reg4831;
                      reg4839 <= (-$signed(((forvar4616 ? reg4846 : reg4701) ?
                          $signed(forvar4763) : (8'haa))));
                      reg4840 <= {(8'ha8)};
                    end
                  if ($signed($signed((forvar4645 ?
                      (8'haf) : reg4841[(3'h7):(3'h7)]))))
                    begin
                      reg4841 <= $unsigned((8'hb1));
                      reg4842 <= $unsigned($unsigned((&reg4647)));
                    end
                  else
                    begin
                      reg4841 <= $signed({reg4740});
                      reg4842 <= forvar4801;
                      reg4843 <= $signed((!$unsigned($unsigned(reg4684))));
                      reg4844 <= forvar4610[(3'h4):(2'h3)];
                    end
                  if ((-forvar4602[(4'h8):(4'h8)]))
                    begin
                      reg4845 <= (~&(~(8'h9f)));
                      reg4846 <= (~($unsigned(forvar4829[(1'h1):(1'h0)]) ?
                          reg4821[(1'h1):(1'h0)] : ($signed((8'haa)) >> $signed(reg4627))));
                      reg4847 <= (!(~^{forvar4843[(4'hb):(3'h5)]}));
                      reg4848 <= $signed(($unsigned(forvar4673) <= ($signed(forvar4594) ?
                          (reg4618 - reg4853) : (&reg4613))));
                    end
                  else
                    begin
                      reg4845 <= reg4669[(2'h2):(1'h1)];
                      reg4846 <= (reg4692 ?
                          forvar4659 : $unsigned($unsigned((~reg4579))));
                    end
                end
              if ((reg4740[(2'h2):(2'h2)] ?
                  $unsigned((!reg4828)) : $signed(((reg4772 ?
                      (8'ha6) : forvar4689) == {wire4574}))))
                begin
                  for (forvar4849 = (1'h0); (forvar4849 < (1'h1)); forvar4849 = (forvar4849 + (1'h1)))
                    begin
                      reg4850 <= {$signed({reg4649})};
                      reg4851 <= (^~((^$unsigned(reg4710)) ?
                          ((&reg4668) * {forvar4696}) : reg4697[(2'h2):(1'h1)]));
                      reg4852 <= $unsigned(forvar4850);
                      reg4853 <= reg4774;
                    end
                  if ({(^~reg4581[(3'h4):(2'h2)])})
                    begin
                      reg4854 <= $signed({((~reg4690) <= $unsigned(forvar4577))});
                      reg4855 <= reg4603;
                      reg4856 <= (reg4581[(4'ha):(4'h9)] && reg4584[(2'h2):(2'h2)]);
                      reg4857 <= (-({forvar4608} >>> {(~reg4611)}));
                    end
                  else
                    begin
                      reg4854 <= $signed($unsigned({{reg4711}}));
                    end
                  for (forvar4858 = (1'h0); (forvar4858 < (1'h1)); forvar4858 = (forvar4858 + (1'h1)))
                    begin
                      reg4859 <= (-{({forvar4654} ?
                              (reg4792 ? (8'ha6) : reg4772) : (|reg4844))});
                      reg4860 <= $unsigned((~^(^$unsigned(reg4610))));
                      reg4861 <= $unsigned(reg4604[(3'h6):(3'h6)]);
                      reg4862 <= (+($signed($unsigned(reg4779)) >> reg4691));
                    end
                  if ($unsigned($unsigned($unsigned((^~reg4735)))))
                    begin
                      reg4863 <= $signed(reg4781[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg4863 <= ((8'ha9) ?
                          {forvar4604[(1'h0):(1'h0)]} : forvar4786);
                    end
                end
              else
                begin
                  if (reg4759)
                    begin
                      reg4849 <= reg4777;
                      reg4850 <= reg4797;
                      reg4851 <= (~&(reg4772[(4'h9):(1'h1)] ?
                          $signed(((8'ha8) ?
                              reg4854 : reg4852)) : forvar4773[(3'h5):(3'h5)]));
                    end
                  else
                    begin
                      reg4849 <= reg4657[(4'hd):(4'ha)];
                      reg4850 <= (~|forvar4839[(3'h5):(2'h3)]);
                      reg4851 <= (((reg4787[(3'h6):(2'h2)] < (~&(8'ha9))) == ((reg4763 ?
                              reg4744 : forvar4763) ?
                          reg4742[(4'hf):(4'he)] : (reg4750 != forvar4604))) >> reg4719);
                    end
                  if (reg4822[(4'he):(4'ha)])
                    begin
                      reg4852 <= (+$signed(((reg4861 ? (8'ha3) : forvar4607) ?
                          reg4658[(3'h6):(1'h1)] : {forvar4604})));
                      reg4853 <= (reg4860[(4'h8):(3'h4)] == $unsigned(reg4762[(3'h5):(2'h3)]));
                    end
                  else
                    begin
                      reg4852 <= ((^forvar4809[(2'h2):(1'h1)]) ?
                          (^forvar4654[(2'h2):(1'h0)]) : {(8'hb7)});
                      reg4853 <= reg4683[(2'h3):(2'h2)];
                    end
                  if ($signed({$signed((forvar4712 ^ reg4787))}))
                    begin
                      reg4854 <= (($unsigned($unsigned(forvar4650)) > (8'haf)) ?
                          forvar4744 : (!reg4605));
                      reg4855 <= $signed({$signed((reg4730 ?
                              reg4638 : forvar4858))});
                    end
                  else
                    begin
                      reg4854 <= ($signed($signed((forvar4607 ^ reg4605))) ?
                          (8'hb0) : (~^forvar4712[(1'h1):(1'h0)]));
                      reg4855 <= $unsigned($signed($signed((~&reg4808))));
                      reg4856 <= forvar4745;
                    end
                end
              if ($signed(forvar4663))
                begin
                  if (({({forvar4593} ? (-reg4646) : reg4702)} ?
                      (reg4710[(2'h3):(1'h1)] ?
                          $signed((|forvar4801)) : reg4744) : forvar4694))
                    begin
                      reg4864 <= reg4734[(4'hb):(2'h3)];
                      reg4865 <= (forvar4824[(2'h2):(2'h2)] - $unsigned(reg4692[(1'h0):(1'h0)]));
                      reg4866 <= {forvar4609[(2'h2):(2'h2)]};
                      reg4867 <= reg4866;
                    end
                  else
                    begin
                      reg4864 <= $signed(reg4752[(4'h8):(2'h3)]);
                      reg4865 <= reg4741;
                    end
                end
              else
                begin
                  for (forvar4864 = (1'h0); (forvar4864 < (1'h1)); forvar4864 = (forvar4864 + (1'h1)))
                    begin
                      reg4865 <= reg4850[(4'hd):(3'h6)];
                      reg4866 <= $signed($signed({(reg4626 ?
                              (8'hb1) : forvar4725)}));
                    end
                end
              if ((((reg4784[(4'hc):(2'h3)] ? (-(8'hba)) : $signed(reg4759)) ?
                      (~^reg4726[(2'h2):(2'h2)]) : (wire4575 >>> (forvar4725 ?
                          reg4609 : reg4791))) ?
                  (~forvar4786) : {reg4709[(3'h6):(1'h1)]}))
                begin
                  reg4868 <= reg4660[(4'h9):(1'h1)];
                  for (forvar4869 = (1'h0); (forvar4869 < (2'h2)); forvar4869 = (forvar4869 + (1'h1)))
                    begin
                      reg4870 <= (~|((forvar4770[(3'h4):(3'h4)] + $signed(reg4670)) ?
                          {forvar4688[(3'h4):(3'h4)]} : $unsigned((|reg4631))));
                      reg4871 <= reg4823[(3'h7):(3'h4)];
                      reg4872 <= (~^forvar4746);
                      reg4873 <= ((-(forvar4603 + (8'h9e))) ?
                          reg4678[(2'h3):(2'h2)] : $signed(($signed(forvar4688) ?
                              {reg4645} : $signed(reg4818))));
                    end
                end
              else
                begin
                  if ({(reg4846 ? (~|$signed(reg4608)) : (8'h9c))})
                    begin
                      reg4868 <= $signed((8'had));
                      reg4869 <= ((reg4703 != $unsigned(wire4574)) ?
                          $signed($unsigned(forvar4795[(4'hc):(2'h2)])) : reg4697[(3'h5):(2'h3)]);
                      reg4870 <= (^~reg4767[(1'h1):(1'h0)]);
                      reg4871 <= (8'hab);
                    end
                  else
                    begin
                      reg4868 <= reg4838;
                      reg4869 <= reg4816;
                      reg4870 <= reg4805;
                      reg4871 <= reg4647[(1'h1):(1'h0)];
                    end
                end
            end
        end
      for (forvar4874 = (1'h0); (forvar4874 < (1'h1)); forvar4874 = (forvar4874 + (1'h1)))
        begin
          reg4875 <= $unsigned({({reg4598} < reg4704)});
          for (forvar4876 = (1'h0); (forvar4876 < (2'h2)); forvar4876 = (forvar4876 + (1'h1)))
            begin
              if (reg4875)
                begin
                  for (forvar4877 = (1'h0); (forvar4877 < (1'h1)); forvar4877 = (forvar4877 + (1'h1)))
                    begin
                      reg4878 <= ($signed(reg4771[(3'h7):(3'h5)]) <<< {{$unsigned(reg4685)}});
                    end
                  for (forvar4879 = (1'h0); (forvar4879 < (1'h0)); forvar4879 = (forvar4879 + (1'h1)))
                    begin
                      reg4880 <= reg4721[(1'h0):(1'h0)];
                      reg4881 <= reg4749[(4'h9):(2'h3)];
                      reg4882 <= forvar4672;
                      reg4883 <= $unsigned((^~$unsigned($signed(forvar4616))));
                    end
                  for (forvar4884 = (1'h0); (forvar4884 < (2'h2)); forvar4884 = (forvar4884 + (1'h1)))
                    begin
                      reg4885 <= ((~reg4654) * forvar4584[(2'h3):(1'h0)]);
                      reg4886 <= $signed((((reg4860 >= forvar4779) ^~ $unsigned(forvar4608)) < {$unsigned(reg4789)}));
                      reg4887 <= $signed($signed((((8'ha1) ?
                              reg4740 : reg4669) ?
                          (reg4651 ? forvar4850 : reg4598) : (~&forvar4817))));
                      reg4888 <= (reg4731 != ((reg4598 | $unsigned(forvar4744)) >> $unsigned(reg4597)));
                    end
                  reg4889 <= $signed((8'hb7));
                end
              else
                begin
                  for (forvar4877 = (1'h0); (forvar4877 < (2'h2)); forvar4877 = (forvar4877 + (1'h1)))
                    begin
                      reg4878 <= {{reg4753[(2'h2):(2'h2)]}};
                      reg4879 <= wire4576;
                      reg4880 <= $unsigned(forvar4848[(2'h2):(2'h2)]);
                    end
                  reg4881 <= reg4747;
                  if ((((&(~|reg4740)) ?
                          ($signed((8'ha2)) >>> (forvar4748 ?
                              reg4859 : reg4835)) : ((forvar4676 < forvar4781) == $signed(reg4702))) ?
                      forvar4645[(1'h0):(1'h0)] : ($signed(((8'h9f) ?
                          (8'hb3) : (8'ha7))) - (8'haf))))
                    begin
                      reg4882 <= {forvar4840};
                    end
                  else
                    begin
                      reg4882 <= {(((forvar4613 ? reg4761 : forvar4779) ?
                                  reg4763[(4'h8):(1'h0)] : $unsigned(reg4606)) ?
                              (^$unsigned(forvar4578)) : reg4782[(1'h0):(1'h0)])};
                      reg4883 <= forvar4824[(4'hb):(3'h7)];
                    end
                end
              for (forvar4890 = (1'h0); (forvar4890 < (1'h0)); forvar4890 = (forvar4890 + (1'h1)))
                begin
                  if ($unsigned($signed($signed(reg4686))))
                    begin
                      reg4891 <= $unsigned((^reg4684[(4'hc):(4'h8)]));
                      reg4892 <= $unsigned(($signed((&reg4578)) == reg4726[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg4891 <= $unsigned($signed(reg4599[(3'h4):(1'h1)]));
                      reg4892 <= ({($unsigned(reg4630) ?
                                  (reg4828 ? (8'ha9) : reg4833) : {reg4706})} ?
                          (reg4644 > ((reg4726 <= forvar4650) ?
                              $signed(forvar4624) : $signed(reg4743))) : (reg4657 ?
                              $signed(reg4658) : ({reg4751} ?
                                  (reg4851 ?
                                      reg4667 : reg4825) : $unsigned((8'hb5)))));
                      reg4893 <= ((-(^{(8'hb6)})) ?
                          (^forvar4789[(1'h0):(1'h0)]) : reg4739[(1'h1):(1'h1)]);
                      reg4894 <= ($unsigned((+(reg4614 ?
                          reg4859 : reg4729))) == (reg4836 ?
                          ((-reg4735) ?
                              (~forvar4642) : (reg4762 && (8'ha4))) : (&$unsigned((8'hae)))));
                    end
                  if ((&(forvar4584[(2'h3):(1'h0)] ?
                      $unsigned((reg4641 <<< (8'hb0))) : {(&forvar4890)})))
                    begin
                      reg4895 <= ((($signed((8'ha4)) > (forvar4593 + reg4893)) == (reg4633[(2'h2):(2'h2)] ?
                              $signed(reg4889) : (forvar4780 ~^ reg4772))) ?
                          (+forvar4851[(1'h0):(1'h0)]) : $signed((|reg4873)));
                      reg4896 <= (&{((reg4579 * reg4738) ?
                              (-reg4781) : (^~reg4655))});
                      reg4897 <= $signed($unsigned((8'hb0)));
                      reg4898 <= (~^(-$signed(reg4853)));
                    end
                  else
                    begin
                      reg4895 <= $unsigned(reg4753);
                    end
                  for (forvar4899 = (1'h0); (forvar4899 < (2'h3)); forvar4899 = (forvar4899 + (1'h1)))
                    begin
                      reg4900 <= forvar4890[(1'h0):(1'h0)];
                      reg4901 <= forvar4869;
                      reg4902 <= $unsigned($unsigned($signed((reg4859 ?
                          reg4676 : reg4604))));
                      reg4903 <= (!($unsigned(reg4893) ^ (8'hb3)));
                    end
                  if (forvar4775[(3'h5):(1'h0)])
                    begin
                      reg4904 <= reg4695;
                      reg4905 <= ($signed((forvar4759[(2'h3):(1'h1)] ?
                              $unsigned(forvar4611) : reg4831[(4'h9):(4'h8)])) ?
                          (8'hb3) : (~$signed((reg4796 ?
                              reg4730 : forvar4840))));
                      reg4906 <= ((forvar4777[(3'h4):(1'h1)] ?
                          $signed(forvar4786) : (+(~|reg4875))) <= $signed(((reg4720 > reg4593) ?
                          {reg4846} : (!reg4703))));
                    end
                  else
                    begin
                      reg4904 <= (8'had);
                    end
                end
              reg4907 <= (((forvar4694 - $unsigned(reg4706)) ?
                  reg4637 : reg4677) < {$unsigned(reg4631)});
            end
        end
      if (reg4720)
        begin
          if (forvar4581)
            begin
              for (forvar4908 = (1'h0); (forvar4908 < (2'h2)); forvar4908 = (forvar4908 + (1'h1)))
                begin
                  for (forvar4909 = (1'h0); (forvar4909 < (2'h3)); forvar4909 = (forvar4909 + (1'h1)))
                    begin
                      reg4910 <= reg4760[(4'h8):(1'h1)];
                    end
                  if (reg4882)
                    begin
                      reg4911 <= $unsigned(forvar4738[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg4911 <= $unsigned((reg4771 != (reg4897[(4'h9):(3'h7)] & $signed((8'haf)))));
                    end
                end
              for (forvar4912 = (1'h0); (forvar4912 < (1'h0)); forvar4912 = (forvar4912 + (1'h1)))
                begin
                  for (forvar4913 = (1'h0); (forvar4913 < (2'h3)); forvar4913 = (forvar4913 + (1'h1)))
                    begin
                      reg4914 <= $signed(forvar4643);
                      reg4915 <= reg4585[(3'h7):(1'h0)];
                      reg4916 <= $unsigned(reg4752[(2'h3):(1'h1)]);
                      reg4917 <= reg4810[(1'h0):(1'h0)];
                    end
                  for (forvar4918 = (1'h0); (forvar4918 < (1'h1)); forvar4918 = (forvar4918 + (1'h1)))
                    begin
                      reg4919 <= forvar4760;
                      reg4920 <= (!$unsigned($signed(reg4844)));
                      reg4921 <= reg4859[(3'h7):(3'h6)];
                      reg4922 <= $unsigned((reg4587 >= reg4636));
                    end
                  for (forvar4923 = (1'h0); (forvar4923 < (2'h2)); forvar4923 = (forvar4923 + (1'h1)))
                    begin
                      reg4924 <= reg4883[(2'h2):(2'h2)];
                      reg4925 <= (-($unsigned((reg4622 + (8'h9d))) ?
                          $unsigned((^forvar4777)) : $signed(reg4878[(3'h6):(3'h4)])));
                      reg4926 <= reg4755;
                      reg4927 <= {(reg4579 | $signed($signed(forvar4839)))};
                    end
                end
              if ((({$unsigned(reg4766)} || ((reg4586 >> (8'ha0)) ?
                      {reg4751} : {reg4895})) ?
                  $unsigned($unsigned($unsigned(forvar4780))) : reg4844[(4'hc):(4'hc)]))
                begin
                  if (($signed(reg4635) ?
                      $unsigned((~$unsigned(reg4656))) : $unsigned((^~{forvar4602}))))
                    begin
                      reg4928 <= {forvar4918[(3'h6):(3'h6)]};
                    end
                  else
                    begin
                      reg4928 <= (8'ha1);
                      reg4929 <= reg4808[(1'h1):(1'h0)];
                    end
                  if (((!$unsigned(forvar4610[(2'h2):(1'h1)])) * (reg4731[(3'h6):(2'h2)] ?
                      (+forvar4913[(1'h0):(1'h0)]) : $unsigned($signed((8'ha2))))))
                    begin
                      reg4930 <= (~^$signed(($unsigned((8'hb5)) ?
                          reg4644 : ((8'ha1) ? reg4774 : reg4811))));
                      reg4931 <= forvar4650;
                      reg4932 <= $unsigned((($signed(reg4682) ?
                              $unsigned(forvar4879) : forvar4681[(1'h1):(1'h1)]) ?
                          (+forvar4912[(4'ha):(4'h9)]) : (8'hb6)));
                      reg4933 <= reg4749;
                    end
                  else
                    begin
                      reg4930 <= reg4836;
                      reg4931 <= (({(forvar4648 ?
                                  forvar4577 : forvar4766)} <= (8'ha0)) ?
                          (reg4727[(1'h1):(1'h1)] | $unsigned($unsigned(reg4927))) : ($unsigned($signed((8'ha6))) == ((&forvar4715) <<< reg4744)));
                      reg4932 <= $signed(forvar4746[(3'h6):(3'h5)]);
                      reg4933 <= (~&(forvar4912 != ((~|reg4750) * (8'h9c))));
                    end
                end
              else
                begin
                  reg4928 <= (~^$unsigned($signed($unsigned(reg4606))));
                  for (forvar4929 = (1'h0); (forvar4929 < (1'h1)); forvar4929 = (forvar4929 + (1'h1)))
                    begin
                      reg4930 <= $unsigned($signed(forvar4584[(3'h7):(2'h3)]));
                      reg4931 <= $unsigned(reg4651[(2'h2):(1'h0)]);
                      reg4932 <= $unsigned(($signed(reg4715[(1'h0):(1'h0)]) && (~&{(8'haa)})));
                      reg4933 <= (({{reg4889}} == (&reg4758)) <<< (((forvar4786 ?
                              (8'hb0) : (8'ha9)) == reg4859[(4'h8):(3'h5)]) ?
                          (+$unsigned(reg4601)) : ($signed((8'ha3)) ?
                              $unsigned(reg4745) : (~|reg4666))));
                    end
                end
            end
          else
            begin
              if (forvar4763)
                begin
                  reg4908 <= reg4881[(2'h3):(1'h1)];
                  for (forvar4909 = (1'h0); (forvar4909 < (1'h1)); forvar4909 = (forvar4909 + (1'h1)))
                    begin
                      reg4910 <= $unsigned(forvar4715);
                    end
                  for (forvar4911 = (1'h0); (forvar4911 < (2'h3)); forvar4911 = (forvar4911 + (1'h1)))
                    begin
                      reg4912 <= reg4875;
                    end
                end
              else
                begin
                  reg4908 <= reg4834;
                end
              for (forvar4913 = (1'h0); (forvar4913 < (2'h2)); forvar4913 = (forvar4913 + (1'h1)))
                begin
                  for (forvar4914 = (1'h0); (forvar4914 < (2'h3)); forvar4914 = (forvar4914 + (1'h1)))
                    begin
                      reg4915 <= $signed($signed(($signed((8'hae)) == forvar4737[(1'h0):(1'h0)])));
                      reg4916 <= reg4842;
                      reg4917 <= (8'ha7);
                      reg4918 <= $unsigned($unsigned($signed((reg4748 ?
                          forvar4913 : reg4916))));
                    end
                  reg4919 <= $unsigned(reg4869[(5'h10):(2'h2)]);
                  for (forvar4920 = (1'h0); (forvar4920 < (1'h1)); forvar4920 = (forvar4920 + (1'h1)))
                    begin
                      reg4921 <= reg4860;
                      reg4922 <= (-$signed({reg4725[(2'h3):(2'h2)]}));
                    end
                end
              if ({forvar4577})
                begin
                  for (forvar4923 = (1'h0); (forvar4923 < (1'h0)); forvar4923 = (forvar4923 + (1'h1)))
                    begin
                      reg4924 <= {$signed($signed($unsigned(reg4747)))};
                      reg4925 <= (8'ha2);
                      reg4926 <= (^($signed(reg4683[(1'h1):(1'h0)]) <= (|reg4816)));
                      reg4927 <= {$unsigned(($unsigned(reg4767) ?
                              (forvar4781 == reg4932) : reg4683))};
                    end
                  if (forvar4850)
                    begin
                      reg4928 <= $unsigned(reg4733);
                      reg4929 <= $unsigned($unsigned($unsigned((~^(8'h9d)))));
                    end
                  else
                    begin
                      reg4928 <= ($unsigned(((reg4638 ? reg4739 : forvar4864) ?
                              (reg4835 | reg4862) : (reg4678 ^~ reg4833))) ?
                          ($unsigned($signed(reg4779)) ?
                              {reg4838[(3'h6):(1'h0)]} : (reg4626[(2'h2):(1'h0)] ?
                                  (forvar4733 ?
                                      forvar4779 : reg4837) : $unsigned(reg4700))) : $signed(forvar4913));
                      reg4929 <= forvar4817[(3'h6):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar4923 = (1'h0); (forvar4923 < (1'h1)); forvar4923 = (forvar4923 + (1'h1)))
                    begin
                      reg4924 <= ({reg4687[(4'ha):(4'ha)]} ?
                          (forvar4775[(1'h0):(1'h0)] ?
                              $signed((~^(8'ha6))) : {$unsigned((8'ha4))}) : (((forvar4581 ?
                                  (8'hb8) : reg4777) == forvar4738) ?
                              reg4684 : (^(reg4816 ?
                                  forvar4696 : forvar4824))));
                      reg4925 <= {(($signed(forvar4698) || (~reg4907)) < ($unsigned((8'ha5)) <= (reg4852 >= reg4719)))};
                    end
                  if ((~&$signed(forvar4681[(2'h2):(1'h1)])))
                    begin
                      reg4926 <= (reg4677 == $unsigned({$unsigned(reg4676)}));
                      reg4927 <= reg4697;
                      reg4928 <= (~|$signed(((~^wire4573) ^~ (reg4636 == (8'hb7)))));
                    end
                  else
                    begin
                      reg4926 <= {(reg4741 ?
                              ($unsigned(reg4916) ?
                                  {reg4714} : reg4630[(3'h7):(2'h2)]) : ((~forvar4676) ?
                                  (~forvar4698) : (-reg4643)))};
                      reg4927 <= $unsigned($signed(($signed(reg4873) ?
                          (reg4844 >> forvar4843) : (reg4903 ?
                              reg4872 : (8'hb7)))));
                      reg4928 <= ((($unsigned(forvar4908) - ((8'haf) ?
                              forvar4760 : reg4731)) ~^ reg4902[(4'hc):(4'hb)]) ?
                          $unsigned($unsigned($signed(reg4699))) : forvar4696[(1'h1):(1'h0)]);
                      reg4929 <= $unsigned({forvar4817});
                    end
                  reg4930 <= forvar4829[(1'h1):(1'h0)];
                  for (forvar4931 = (1'h0); (forvar4931 < (1'h1)); forvar4931 = (forvar4931 + (1'h1)))
                    begin
                      reg4932 <= $unsigned($unsigned(forvar4920[(1'h0):(1'h0)]));
                    end
                end
              for (forvar4933 = (1'h0); (forvar4933 < (1'h0)); forvar4933 = (forvar4933 + (1'h1)))
                begin
                  if (reg4723)
                    begin
                      reg4934 <= $unsigned((&reg4837[(3'h6):(2'h2)]));
                      reg4935 <= $unsigned(reg4738);
                      reg4936 <= {$signed(reg4755)};
                    end
                  else
                    begin
                      reg4934 <= {reg4693};
                      reg4935 <= (8'ha7);
                      reg4936 <= {reg4643};
                    end
                  if ($signed($signed(forvar4840[(4'hd):(4'h8)])))
                    begin
                      reg4937 <= reg4730;
                      reg4938 <= $signed((!((reg4905 ? reg4845 : reg4752) ?
                          forvar4753[(1'h0):(1'h0)] : (reg4805 ?
                              forvar4908 : reg4756))));
                      reg4939 <= (((~{forvar4864}) >> (&$unsigned(reg4604))) - ((8'ha3) | (-(8'hb0))));
                    end
                  else
                    begin
                      reg4937 <= (&(~{((8'hb9) != forvar4814)}));
                      reg4938 <= (forvar4869[(1'h1):(1'h1)] ?
                          reg4666 : ({forvar4608} ?
                              reg4790[(4'hd):(3'h4)] : {(8'hb4)}));
                    end
                end
            end
        end
      else
        begin
          for (forvar4908 = (1'h0); (forvar4908 < (2'h3)); forvar4908 = (forvar4908 + (1'h1)))
            begin
              reg4909 <= reg4590[(4'h9):(3'h4)];
              if (forvar4580)
                begin
                  if (reg4838[(3'h6):(1'h1)])
                    begin
                      reg4910 <= $unsigned(($signed((reg4632 ?
                          reg4820 : reg4865)) ^ reg4605));
                      reg4911 <= reg4654[(2'h3):(2'h3)];
                      reg4912 <= {(($unsigned(reg4688) || (~|reg4736)) > $signed((reg4871 >> forvar4755)))};
                      reg4913 <= $unsigned(reg4834[(2'h2):(1'h1)]);
                    end
                  else
                    begin
                      reg4910 <= $signed((~{$signed(forvar4814)}));
                      reg4911 <= ((((reg4758 ~^ forvar4592) ?
                          (forvar4884 ? forvar4648 : (8'ha3)) : (reg4869 ?
                              (8'ha4) : (8'h9c))) + (~|(reg4584 < reg4578))) | $signed(reg4915));
                      reg4912 <= (~&reg4623[(3'h7):(3'h6)]);
                    end
                end
              else
                begin
                  for (forvar4910 = (1'h0); (forvar4910 < (1'h0)); forvar4910 = (forvar4910 + (1'h1)))
                    begin
                      reg4911 <= (~|reg4682[(1'h0):(1'h0)]);
                      reg4912 <= {{(|(reg4620 ? reg4630 : forvar4755))}};
                      reg4913 <= (~((^$unsigned(reg4728)) ?
                          reg4835[(1'h0):(1'h0)] : (8'hb7)));
                      reg4914 <= ((reg4851 << ($signed(reg4637) ?
                          (reg4893 << reg4868) : (reg4932 << reg4789))) - $signed($signed(reg4893)));
                    end
                  for (forvar4915 = (1'h0); (forvar4915 < (1'h0)); forvar4915 = (forvar4915 + (1'h1)))
                    begin
                      reg4916 <= reg4932;
                    end
                end
            end
        end
    end
  assign wire4940 = $unsigned(forvar4779);
  always
    @(posedge clk) begin
      if (reg4820[(3'h4):(2'h3)])
        begin
          reg4941 <= ($unsigned($unsigned($signed(reg4714))) ~^ {reg4760});
        end
      else
        begin
          if ((|(8'ha2)))
            begin
              if ((&(8'ha4)))
                begin
                  reg4941 <= $unsigned({$unsigned((reg4682 - forvar4705))});
                  if ({($signed(reg4920) ?
                          (!((8'hb8) ?
                              reg4838 : reg4670)) : $signed($signed(reg4796)))})
                    begin
                      reg4942 <= (~&reg4579);
                    end
                  else
                    begin
                      reg4942 <= (~^(reg4794 >> (|forvar4795[(3'h5):(3'h5)])));
                    end
                  reg4943 <= $unsigned(((8'hb7) || reg4762));
                end
              else
                begin
                  if (((~&$signed({reg4907})) ?
                      forvar4694[(4'h9):(2'h2)] : forvar4931[(2'h2):(1'h1)]))
                    begin
                      reg4941 <= ({reg4744[(1'h1):(1'h1)]} ?
                          reg4933 : $signed((8'haa)));
                    end
                  else
                    begin
                      reg4941 <= $unsigned(($unsigned(reg4804[(4'h8):(3'h5)]) ?
                          ({reg4684} | $signed(reg4638)) : (+reg4688[(2'h3):(2'h3)])));
                      reg4942 <= $signed($unsigned($unsigned(wire4940[(1'h1):(1'h0)])));
                      reg4943 <= reg4738;
                    end
                end
              for (forvar4944 = (1'h0); (forvar4944 < (2'h3)); forvar4944 = (forvar4944 + (1'h1)))
                begin
                  reg4945 <= (8'h9e);
                  for (forvar4946 = (1'h0); (forvar4946 < (1'h0)); forvar4946 = (forvar4946 + (1'h1)))
                    begin
                      reg4947 <= reg4771[(4'hc):(4'hb)];
                      reg4948 <= {{$unsigned({reg4745})}};
                      reg4949 <= ((forvar4643[(4'hf):(3'h7)] ?
                              ($signed(forvar4920) > $unsigned(reg4581)) : forvar4908) ?
                          $signed((^reg4855[(4'h8):(2'h2)])) : {(((8'hac) ?
                                      forvar4824 : reg4835) ?
                                  reg4691[(2'h3):(1'h1)] : reg4941)});
                    end
                  if (reg4860[(4'h8):(2'h3)])
                    begin
                      reg4950 <= forvar4908;
                    end
                  else
                    begin
                      reg4950 <= ($unsigned((&$signed(forvar4643))) <<< reg4804[(3'h7):(2'h3)]);
                      reg4951 <= $unsigned($signed({(~|forvar4725)}));
                    end
                  for (forvar4952 = (1'h0); (forvar4952 < (2'h2)); forvar4952 = (forvar4952 + (1'h1)))
                    begin
                      reg4953 <= $unsigned(reg4764[(4'ha):(4'h9)]);
                      reg4954 <= $unsigned($unsigned($unsigned(reg4707)));
                      reg4955 <= (~^reg4638);
                      reg4956 <= ((8'hab) ?
                          (($unsigned(forvar4785) == $signed(wire4575)) ?
                              $unsigned(((8'hb8) < reg4900)) : ($signed(forvar4809) >> $unsigned(reg4602))) : $unsigned(($unsigned(reg4755) << forvar4768[(1'h1):(1'h0)])));
                    end
                end
              for (forvar4957 = (1'h0); (forvar4957 < (2'h2)); forvar4957 = (forvar4957 + (1'h1)))
                begin
                  for (forvar4958 = (1'h0); (forvar4958 < (1'h1)); forvar4958 = (forvar4958 + (1'h1)))
                    begin
                      reg4959 <= ({(reg4907 ?
                              {reg4623} : $signed(forvar4674))} >> ((reg4687[(4'hb):(1'h1)] ?
                          reg4838[(2'h3):(1'h0)] : (reg4835 == reg4848)) << {{wire4799}}));
                      reg4960 <= {((^reg4781[(3'h6):(3'h4)]) ?
                              ((8'ha5) >= reg4761) : (&((8'hba) ?
                                  forvar4688 : reg4580)))};
                      reg4961 <= $unsigned((&reg4665));
                    end
                end
            end
          else
            begin
              for (forvar4941 = (1'h0); (forvar4941 < (1'h1)); forvar4941 = (forvar4941 + (1'h1)))
                begin
                  if ($unsigned((-$unsigned(reg4852))))
                    begin
                      reg4942 <= $unsigned($signed((wire4798[(2'h2):(1'h1)] >= reg4619)));
                      reg4943 <= $signed((~^reg4840));
                    end
                  else
                    begin
                      reg4942 <= reg4586[(2'h2):(1'h1)];
                    end
                  if (((^(((8'hba) ? reg4929 : (8'had)) ?
                          forvar4958 : (reg4941 << reg4775))) ?
                      reg4677[(1'h0):(1'h0)] : $signed($unsigned($signed(forvar4911)))))
                    begin
                      reg4944 <= (+(((reg4808 && forvar4795) ?
                          (-reg4600) : (-reg4601)) > (+(!(8'ha0)))));
                      reg4945 <= $unsigned((reg4657[(2'h3):(1'h0)] == $signed($signed(reg4762))));
                      reg4946 <= {$unsigned((reg4732[(2'h3):(2'h2)] * (reg4892 >> forvar4814)))};
                      reg4947 <= (&{(!forvar4608[(3'h7):(3'h5)])});
                    end
                  else
                    begin
                      reg4944 <= $signed($unsigned({$signed(reg4936)}));
                      reg4945 <= (8'hb8);
                    end
                  if ((^reg4701[(4'h8):(2'h2)]))
                    begin
                      reg4948 <= (&reg4688);
                    end
                  else
                    begin
                      reg4948 <= reg4771[(1'h1):(1'h0)];
                      reg4949 <= $signed(reg4631);
                      reg4950 <= forvar4654;
                      reg4951 <= (reg4821[(3'h7):(1'h1)] > reg4931[(3'h7):(3'h7)]);
                    end
                  if ((&(forvar4712[(1'h1):(1'h1)] != $signed($unsigned((8'h9f))))))
                    begin
                      reg4952 <= $unsigned(((reg4774 == (~reg4913)) ^~ forvar4789));
                      reg4953 <= ((forvar4580 <= reg4707[(4'hc):(4'h8)]) | forvar4760);
                    end
                  else
                    begin
                      reg4952 <= {$unsigned(reg4687[(1'h1):(1'h1)])};
                    end
                end
            end
        end
      if ((forvar4826 ?
          $signed(forvar4941) : $signed(((reg4821 - reg4830) ?
              (reg4790 ~^ forvar4795) : $signed(forvar4915)))))
        begin
          for (forvar4962 = (1'h0); (forvar4962 < (1'h1)); forvar4962 = (forvar4962 + (1'h1)))
            begin
              reg4963 <= (($unsigned({reg4959}) && $signed((8'hae))) ?
                  $signed($signed(reg4660)) : ((~&(forvar4673 ?
                      reg4771 : reg4793)) != (8'ha7)));
            end
          reg4964 <= reg4726[(1'h0):(1'h0)];
        end
      else
        begin
          reg4962 <= $unsigned((!((~reg4757) != reg4771[(4'hd):(3'h6)])));
          reg4963 <= reg4632[(2'h2):(1'h1)];
        end
      if ((~$unsigned($unsigned((reg4585 << reg4583)))))
        begin
          if ((({(8'hb1)} ?
              (^~reg4818[(3'h4):(3'h4)]) : $signed((reg4626 ?
                  (8'hb9) : reg4586))) != ((8'hb3) >>> forvar4689[(4'ha):(4'ha)])))
            begin
              for (forvar4965 = (1'h0); (forvar4965 < (1'h0)); forvar4965 = (forvar4965 + (1'h1)))
                begin
                  for (forvar4966 = (1'h0); (forvar4966 < (1'h1)); forvar4966 = (forvar4966 + (1'h1)))
                    begin
                      reg4967 <= $signed($unsigned({$signed((8'had))}));
                      reg4968 <= {reg4935[(4'h9):(4'h8)]};
                      reg4969 <= $signed($unsigned((reg4894 ?
                          ((8'ha2) || forvar4815) : (~&forvar4755))));
                      reg4970 <= (~^$unsigned(reg4780[(1'h1):(1'h0)]));
                    end
                end
              reg4971 <= $unsigned($unsigned($signed((^reg4822))));
              for (forvar4972 = (1'h0); (forvar4972 < (1'h0)); forvar4972 = (forvar4972 + (1'h1)))
                begin
                  if (reg4577[(3'h5):(3'h5)])
                    begin
                      reg4973 <= $unsigned($unsigned(((~forvar4636) & (forvar4694 ?
                          forvar4594 : reg4680))));
                    end
                  else
                    begin
                      reg4973 <= forvar4768[(2'h2):(1'h1)];
                      reg4974 <= (^~forvar4705[(2'h3):(2'h2)]);
                      reg4975 <= (!$signed(reg4834[(1'h1):(1'h0)]));
                      reg4976 <= (($unsigned($signed(reg4634)) ?
                              forvar4827[(1'h1):(1'h1)] : (wire4574 ?
                                  reg4780 : (reg4867 ? reg4861 : reg4774))) ?
                          ($unsigned((|reg4833)) * reg4631) : reg4707);
                    end
                  for (forvar4977 = (1'h0); (forvar4977 < (2'h2)); forvar4977 = (forvar4977 + (1'h1)))
                    begin
                      reg4978 <= ((~^reg4783) <= $unsigned((|reg4634)));
                      reg4979 <= reg4912;
                    end
                  for (forvar4980 = (1'h0); (forvar4980 < (2'h2)); forvar4980 = (forvar4980 + (1'h1)))
                    begin
                      reg4981 <= (reg4803[(3'h4):(2'h2)] | (|($signed(reg4914) ?
                          (reg4781 * reg4760) : reg4931)));
                      reg4982 <= (~&($signed((reg4888 ? forvar4645 : reg4970)) ?
                          (-{(8'haf)}) : $unsigned((reg4911 <<< forvar4760))));
                      reg4983 <= $unsigned(({$signed(reg4804)} ?
                          {reg4839} : (~(reg4678 >> reg4950))));
                      reg4984 <= forvar4741;
                    end
                  reg4985 <= (forvar4746[(1'h1):(1'h0)] ?
                      {(~|((8'ha4) >> forvar4777))} : forvar4643[(2'h2):(1'h1)]);
                end
            end
          else
            begin
              if (($signed((8'hb2)) >> $signed(({forvar4813} * $signed(reg4955)))))
                begin
                  if ($signed($unsigned((~&reg4677[(3'h7):(2'h3)]))))
                    begin
                      reg4965 <= {(|$signed((!forvar4877)))};
                      reg4966 <= $signed($unsigned(reg4670[(2'h2):(2'h2)]));
                      reg4967 <= {reg4904};
                    end
                  else
                    begin
                      reg4965 <= $unsigned((forvar4775 & reg4683[(2'h2):(1'h0)]));
                      reg4966 <= $signed($signed((wire4940 << reg4842)));
                      reg4967 <= $unsigned($signed($signed($signed(reg4828))));
                      reg4968 <= $unsigned(reg4584[(4'ha):(3'h6)]);
                    end
                end
              else
                begin
                  for (forvar4965 = (1'h0); (forvar4965 < (2'h3)); forvar4965 = (forvar4965 + (1'h1)))
                    begin
                      reg4966 <= $unsigned(reg4760);
                      reg4967 <= reg4837;
                      reg4968 <= (reg4677 <<< reg4724[(1'h1):(1'h1)]);
                    end
                  for (forvar4969 = (1'h0); (forvar4969 < (1'h1)); forvar4969 = (forvar4969 + (1'h1)))
                    begin
                      reg4970 <= reg4834[(2'h2):(1'h1)];
                      reg4971 <= ($unsigned(($unsigned(reg4685) ?
                              ((8'h9d) > (8'hb2)) : (reg4587 ?
                                  reg4633 : (8'h9d)))) ?
                          reg4812 : $signed({(8'h9c)}));
                      reg4972 <= ((((~reg4626) ?
                              (^~reg4766) : (&reg4728)) | ($signed(reg4752) + {forvar4829})) ?
                          (((forvar4654 * reg4768) ?
                                  (reg4835 ^ reg4896) : forvar4876) ?
                              reg4750 : reg4830) : $signed({(|(8'hb1))}));
                    end
                  for (forvar4973 = (1'h0); (forvar4973 < (2'h2)); forvar4973 = (forvar4973 + (1'h1)))
                    begin
                      reg4974 <= (+reg4852);
                    end
                end
              if (reg4761[(2'h2):(1'h1)])
                begin
                  for (forvar4975 = (1'h0); (forvar4975 < (2'h3)); forvar4975 = (forvar4975 + (1'h1)))
                    begin
                      reg4976 <= $unsigned($unsigned({reg4794}));
                      reg4977 <= (forvar4698[(1'h1):(1'h0)] ?
                          reg4731[(1'h0):(1'h0)] : forvar4610[(3'h5):(1'h0)]);
                      reg4978 <= {((~&(!forvar4737)) <= (((8'hb1) << reg4690) && reg4897[(4'h8):(4'h8)]))};
                    end
                  if ({$unsigned(($unsigned(forvar4914) << (^~reg4745)))})
                    begin
                      reg4979 <= $signed(({(reg4812 << reg4973)} == $signed((reg4924 ?
                          reg4651 : reg4891))));
                      reg4980 <= $signed((forvar4913[(1'h0):(1'h0)] <<< $unsigned($signed((8'h9e)))));
                    end
                  else
                    begin
                      reg4979 <= reg4626;
                      reg4980 <= $signed($unsigned(reg4580));
                      reg4981 <= reg4810;
                    end
                  if ($signed(reg4649))
                    begin
                      reg4982 <= (reg4718 - $signed(reg4822));
                      reg4983 <= reg4929;
                      reg4984 <= {(8'ha1)};
                    end
                  else
                    begin
                      reg4982 <= reg4919;
                      reg4983 <= $signed($signed(((forvar4850 ?
                          forvar4688 : reg4577) >= $signed(reg4934))));
                      reg4984 <= ((($signed(forvar4973) ?
                              (forvar4672 ?
                                  reg4597 : reg4796) : (~^reg4901)) < $unsigned($signed(reg4615))) ?
                          reg4898[(2'h3):(2'h2)] : ((reg4897 >> reg4841[(4'hb):(2'h2)]) ?
                              (+(forvar4731 ? reg4697 : wire4575)) : (8'ha1)));
                      reg4985 <= ({reg4686} && $signed(reg4591[(2'h3):(2'h3)]));
                    end
                  for (forvar4986 = (1'h0); (forvar4986 < (1'h1)); forvar4986 = (forvar4986 + (1'h1)))
                    begin
                      reg4987 <= (reg4800[(1'h1):(1'h1)] ?
                          $unsigned((reg4985[(1'h0):(1'h0)] && $unsigned(forvar4884))) : reg4753);
                    end
                end
              else
                begin
                  for (forvar4975 = (1'h0); (forvar4975 < (1'h1)); forvar4975 = (forvar4975 + (1'h1)))
                    begin
                      reg4976 <= reg4693[(2'h3):(1'h1)];
                      reg4977 <= $signed((|reg4762[(2'h2):(1'h0)]));
                      reg4978 <= forvar4884[(3'h5):(1'h0)];
                    end
                  reg4979 <= (($unsigned($signed(reg4662)) ?
                      ($unsigned((8'hb4)) | (reg4621 <<< reg4931)) : reg4984[(3'h4):(2'h3)]) ^ $unsigned((~|(forvar4663 <= (8'hb7)))));
                end
              if ($unsigned((^reg4577[(3'h6):(1'h0)])))
                begin
                  for (forvar4988 = (1'h0); (forvar4988 < (1'h0)); forvar4988 = (forvar4988 + (1'h1)))
                    begin
                      reg4989 <= $signed(forvar4579[(1'h1):(1'h1)]);
                      reg4990 <= reg4908;
                      reg4991 <= {((+(8'ha8)) ?
                              (8'hb5) : $signed(reg4752[(4'h9):(2'h3)]))};
                      reg4992 <= $signed((((reg4745 ? (8'hae) : reg4821) ?
                              (~^forvar4689) : $signed((8'haf))) ?
                          ($signed(reg4707) ?
                              (reg4702 ?
                                  reg4678 : reg4628) : $unsigned(reg4761)) : forvar4914));
                    end
                  reg4993 <= ((($unsigned(reg4634) || forvar4813[(4'hd):(4'hb)]) >>> (~&(8'haf))) ?
                      $signed($unsigned((forvar4588 ?
                          forvar4864 : forvar4616))) : forvar4636);
                  reg4994 <= (~^$unsigned((^(reg4757 ?
                      forvar4848 : forvar4829))));
                end
              else
                begin
                  for (forvar4988 = (1'h0); (forvar4988 < (2'h3)); forvar4988 = (forvar4988 + (1'h1)))
                    begin
                      reg4989 <= $signed($unsigned($unsigned(forvar4745)));
                      reg4990 <= ({$signed(reg4807)} ?
                          forvar4795 : {$signed({forvar4602})});
                    end
                  for (forvar4991 = (1'h0); (forvar4991 < (2'h3)); forvar4991 = (forvar4991 + (1'h1)))
                    begin
                      reg4992 <= reg4864[(4'h9):(2'h3)];
                      reg4993 <= (~^reg4688[(4'h9):(3'h6)]);
                    end
                  reg4994 <= forvar4876[(4'he):(4'ha)];
                end
            end
          if (($signed(($unsigned(reg4761) << (reg4871 < (8'hb1)))) & reg4938[(1'h0):(1'h0)]))
            begin
              if (reg4645)
                begin
                  reg4995 <= $unsigned(reg4794);
                end
              else
                begin
                  if ((&(reg4606 ?
                      (reg4644 != (~|forvar4593)) : (+(reg4932 ~^ reg4581)))))
                    begin
                      reg4995 <= ((($unsigned(reg4873) > (-forvar4676)) - $signed((!forvar4829))) ?
                          $unsigned(($unsigned((8'hab)) ?
                              $unsigned(reg4788) : (reg4880 ?
                                  reg4934 : (8'h9f)))) : forvar4837[(4'hb):(4'h8)]);
                    end
                  else
                    begin
                      reg4995 <= (~(forvar4931[(2'h3):(1'h0)] > reg4885));
                      reg4996 <= {forvar4781[(2'h2):(1'h1)]};
                    end
                  reg4997 <= {reg4747};
                end
              for (forvar4998 = (1'h0); (forvar4998 < (2'h3)); forvar4998 = (forvar4998 + (1'h1)))
                begin
                  for (forvar4999 = (1'h0); (forvar4999 < (2'h2)); forvar4999 = (forvar4999 + (1'h1)))
                    begin
                      reg5000 <= (~|(^~{$unsigned(reg4947)}));
                      reg5001 <= reg4637[(2'h2):(2'h2)];
                      reg5002 <= reg4668[(1'h0):(1'h0)];
                      reg5003 <= $signed(reg4966);
                    end
                  reg5004 <= ((forvar4673[(2'h2):(1'h1)] < $signed((reg4687 ^ forvar4579))) ?
                      reg4715 : reg4808[(1'h0):(1'h0)]);
                  reg5005 <= (($unsigned($unsigned(reg4664)) ?
                      $unsigned(reg4651) : $unsigned((forvar4789 <<< reg4828))) >= ($signed($unsigned(reg4918)) ?
                      (|reg4857[(2'h3):(2'h2)]) : forvar4766[(3'h4):(1'h0)]));
                end
            end
          else
            begin
              for (forvar4995 = (1'h0); (forvar4995 < (2'h3)); forvar4995 = (forvar4995 + (1'h1)))
                begin
                  for (forvar4996 = (1'h0); (forvar4996 < (2'h2)); forvar4996 = (forvar4996 + (1'h1)))
                    begin
                      reg4997 <= (~^forvar4802[(1'h1):(1'h0)]);
                      reg4998 <= (reg4765[(2'h3):(2'h3)] == (($signed((8'hac)) == $signed((8'hb1))) ?
                          $unsigned($unsigned((8'ha7))) : ($unsigned(reg4756) ?
                              (reg4781 ?
                                  forvar4944 : forvar4688) : $unsigned(reg4875))));
                      reg4999 <= ((&reg4612[(2'h2):(2'h2)]) << $unsigned(reg4847));
                    end
                end
              reg5000 <= $signed((($signed(wire4799) ?
                  reg4600[(2'h3):(2'h3)] : $unsigned(forvar4957)) & {$unsigned(reg4675)}));
              if ((forvar4654[(2'h3):(2'h3)] ?
                  {((^(8'h9d)) ?
                          $signed(reg4598) : $unsigned(reg4841))} : $unsigned(reg4979)))
                begin
                  for (forvar5001 = (1'h0); (forvar5001 < (2'h2)); forvar5001 = (forvar5001 + (1'h1)))
                    begin
                      reg5002 <= $unsigned(($unsigned($unsigned(reg4732)) * (8'ha2)));
                    end
                  reg5003 <= reg4963[(3'h5):(3'h5)];
                end
              else
                begin
                  if ({(forvar4848[(1'h1):(1'h0)] ?
                          reg4841 : ((&reg4584) ?
                              (reg4961 << forvar4775) : $signed(reg4840)))})
                    begin
                      reg5001 <= ((^~reg4977[(1'h0):(1'h0)]) ?
                          ((!reg4917[(1'h1):(1'h0)]) ?
                              reg4723[(4'h9):(2'h2)] : ((reg4889 ?
                                  reg4885 : reg4908) | $unsigned(reg4630))) : (-reg4585));
                    end
                  else
                    begin
                      reg5001 <= forvar4973[(4'hc):(4'h8)];
                    end
                end
            end
          if (reg4812[(3'h4):(2'h3)])
            begin
              for (forvar5006 = (1'h0); (forvar5006 < (1'h1)); forvar5006 = (forvar5006 + (1'h1)))
                begin
                  if (((8'hb0) ? (&(8'hb0)) : reg4764[(4'ha):(3'h7)]))
                    begin
                      reg5007 <= $unsigned(((^(8'hb9)) ?
                          $unsigned({reg4949}) : ((+reg4970) >= $unsigned(forvar4941))));
                      reg5008 <= $unsigned(reg4596[(2'h3):(2'h2)]);
                      reg5009 <= (^$unsigned(((forvar4781 < reg4944) ?
                          ((8'hb5) ?
                              reg4991 : reg4938) : $signed(forvar4712))));
                      reg5010 <= ($unsigned($unsigned(forvar4802)) != $signed({$unsigned(forvar4958)}));
                    end
                  else
                    begin
                      reg5007 <= {($unsigned((reg4821 ? reg4935 : forvar4952)) ?
                              (|$unsigned(reg4950)) : ($signed(reg4741) ?
                                  $signed((8'ha6)) : (&reg4925)))};
                    end
                end
            end
          else
            begin
              if ($unsigned(forvar4980))
                begin
                  for (forvar5006 = (1'h0); (forvar5006 < (2'h2)); forvar5006 = (forvar5006 + (1'h1)))
                    begin
                      reg5007 <= (reg4914[(3'h4):(1'h0)] <<< $signed(forvar4840));
                      reg5008 <= wire4574;
                    end
                  for (forvar5009 = (1'h0); (forvar5009 < (1'h0)); forvar5009 = (forvar5009 + (1'h1)))
                    begin
                      reg5010 <= ($unsigned($unsigned(reg4889)) ?
                          $signed(reg4626) : (8'ha6));
                      reg5011 <= reg4703;
                      reg5012 <= forvar4613;
                    end
                  if ((~&$signed($signed(reg4975))))
                    begin
                      reg5013 <= reg4610[(2'h3):(1'h0)];
                      reg5014 <= ((reg5013 ^ $signed((~^forvar4817))) >> (((~&reg4993) ?
                              (forvar5006 - forvar4672) : (~|reg4885)) ?
                          (^~reg4643) : reg4960));
                      reg5015 <= reg4585;
                      reg5016 <= $signed($signed(forvar4915[(3'h7):(2'h3)]));
                    end
                  else
                    begin
                      reg5013 <= {$signed({(reg4959 && forvar5006)})};
                      reg5014 <= reg4708[(3'h6):(3'h6)];
                    end
                end
              else
                begin
                  for (forvar5006 = (1'h0); (forvar5006 < (2'h2)); forvar5006 = (forvar5006 + (1'h1)))
                    begin
                      reg5007 <= forvar4750[(4'hd):(4'hb)];
                    end
                end
              if ($signed((((forvar4771 ? reg4918 : reg4885) | forvar4771) ?
                  ((8'hb0) ^~ forvar4763) : (~(forvar4864 ?
                      (8'had) : reg5002)))))
                begin
                  if ($signed(reg4709))
                    begin
                      reg5017 <= reg4777[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg5017 <= (&($unsigned((forvar4750 ?
                          reg4804 : reg4836)) ~^ (&(reg4898 ?
                          (8'h9c) : reg4765))));
                      reg5018 <= $signed((^~$unsigned({reg5010})));
                    end
                  for (forvar5019 = (1'h0); (forvar5019 < (1'h1)); forvar5019 = (forvar5019 + (1'h1)))
                    begin
                      reg5020 <= $unsigned($unsigned(((reg4820 & reg4772) | {forvar4908})));
                      reg5021 <= reg4675;
                      reg5022 <= {reg4998};
                    end
                  if ($unsigned(reg4695))
                    begin
                      reg5023 <= (!$unsigned((^$signed(reg4782))));
                    end
                  else
                    begin
                      reg5023 <= ($signed($unsigned((!reg4984))) ?
                          forvar4909[(1'h1):(1'h0)] : (((forvar4676 >> forvar4673) >> reg4808[(2'h3):(1'h0)]) < reg4683));
                    end
                end
              else
                begin
                  if ({(-reg4875)})
                    begin
                      reg5017 <= ((~&$unsigned((reg4834 && (8'hb8)))) ?
                          {forvar4914[(1'h1):(1'h1)]} : $unsigned({reg4628[(4'hc):(2'h3)]}));
                    end
                  else
                    begin
                      reg5017 <= ($unsigned($signed($unsigned(reg4879))) ?
                          $signed($signed((|reg4936))) : $unsigned({(8'haf)}));
                    end
                end
              if ((~|$signed($signed(forvar4965[(2'h3):(1'h0)]))))
                begin
                  if (forvar4969[(1'h1):(1'h1)])
                    begin
                      reg5024 <= $unsigned((!($unsigned(reg4869) < (~forvar4975))));
                      reg5025 <= (^~$unsigned(reg4647));
                      reg5026 <= $signed(reg4788);
                    end
                  else
                    begin
                      reg5024 <= (~&forvar4780);
                    end
                  if (({(^~$signed(reg4724))} ^ (+reg4624[(3'h4):(2'h2)])))
                    begin
                      reg5027 <= (-forvar4755);
                    end
                  else
                    begin
                      reg5027 <= reg4861[(2'h3):(2'h3)];
                      reg5028 <= (^~$unsigned($unsigned($unsigned(reg4944))));
                    end
                  for (forvar5029 = (1'h0); (forvar5029 < (2'h3)); forvar5029 = (forvar5029 + (1'h1)))
                    begin
                      reg5030 <= {(!reg4949[(1'h1):(1'h0)])};
                      reg5031 <= ((reg5025 ?
                              (reg4841 ?
                                  reg4657 : reg4891[(3'h4):(1'h1)]) : reg4579) ?
                          (((!(8'h9f)) ?
                              forvar4789[(1'h0):(1'h0)] : reg4937) || forvar4580[(1'h1):(1'h0)]) : ($signed((reg4754 * (8'ha0))) ~^ (reg4749[(1'h0):(1'h0)] ?
                              $signed(reg4711) : reg4834[(1'h1):(1'h0)])));
                      reg5032 <= (&$signed((8'ha4)));
                      reg5033 <= reg4742;
                    end
                  reg5034 <= (({$unsigned(reg4981)} >= $signed(forvar4731[(1'h0):(1'h0)])) ?
                      (($signed(reg4989) ?
                          $unsigned(reg4690) : forvar4640[(2'h2):(1'h0)]) >= (8'h9e)) : $signed(($signed(reg4837) ?
                          reg4768[(1'h0):(1'h0)] : (reg4807 ^~ reg4734))));
                end
              else
                begin
                  if ($unsigned($signed(($signed(reg4613) << reg4996[(3'h4):(2'h3)]))))
                    begin
                      reg5024 <= (({(reg4786 | forvar4941)} >= reg4697) >> $signed(((~(8'hac)) == ((8'hb9) ?
                          forvar4616 : reg4931))));
                      reg5025 <= (8'h9f);
                      reg5026 <= (((reg4747[(2'h3):(2'h2)] ?
                                  (forvar4608 ?
                                      reg4833 : (8'hb6)) : $signed(reg4835)) ?
                              reg4788 : ((reg4651 ? forvar4725 : (8'hb4)) ?
                                  $signed(forvar4733) : (reg4942 ?
                                      reg4975 : reg4985))) ?
                          (forvar4890[(1'h0):(1'h0)] ?
                              ((reg4913 ?
                                  (8'haa) : forvar4584) ^~ ((8'hb7) >= (8'hb8))) : reg4724[(3'h4):(1'h0)]) : ((reg5023 ?
                                  reg5001[(3'h5):(2'h3)] : {reg4722}) ?
                              (((8'had) <<< forvar4858) && (forvar4731 + (8'hb6))) : (forvar4725 ^ $unsigned(reg4928))));
                    end
                  else
                    begin
                      reg5024 <= reg4997;
                      reg5025 <= reg4938;
                      reg5026 <= (~|(^{$signed(reg4807)}));
                    end
                  if ((8'h9f))
                    begin
                      reg5027 <= forvar4813;
                    end
                  else
                    begin
                      reg5027 <= $signed(((+(^reg4907)) ?
                          (reg4854 ?
                              reg4613 : $signed((8'hb4))) : $signed($unsigned(forvar4688))));
                      reg5028 <= (+$signed(({(8'hb5)} ?
                          (|forvar4988) : $unsigned(reg4582))));
                      reg5029 <= {reg4741};
                      reg5030 <= (reg4781[(2'h2):(2'h2)] | reg4907);
                    end
                end
            end
        end
      else
        begin
          reg4965 <= ({(8'ha0)} ?
              (~|({reg5022} >>> $signed((8'ha1)))) : (8'hb1));
          if ($unsigned((reg4782 ?
              $unsigned(reg4643[(1'h0):(1'h0)]) : $unsigned(reg4850[(4'hf):(1'h0)]))))
            begin
              for (forvar4966 = (1'h0); (forvar4966 < (1'h0)); forvar4966 = (forvar4966 + (1'h1)))
                begin
                  if (forvar5009[(3'h5):(3'h4)])
                    begin
                      reg4967 <= $unsigned(forvar4577);
                      reg4968 <= ((($signed(reg4691) ^ (+reg5017)) > $signed((|forvar4591))) ?
                          $unsigned($signed(((8'hab) ?
                              reg4634 : reg4909))) : (reg4868 ?
                              $signed($unsigned((8'ha3))) : reg4660));
                      reg4969 <= forvar4759;
                    end
                  else
                    begin
                      reg4967 <= (reg4803 ?
                          ((forvar4779[(4'hc):(1'h1)] >= $signed(forvar4624)) == reg4945) : ($unsigned((8'hb7)) ?
                              (~$unsigned(reg4626)) : (reg4828 ?
                                  $signed(reg4844) : reg4787[(4'ha):(4'ha)])));
                      reg4968 <= reg4962[(3'h7):(3'h4)];
                      reg4969 <= ({$signed(reg4623[(3'h5):(1'h1)])} ~^ $unsigned(reg4838[(1'h0):(1'h0)]));
                    end
                end
              for (forvar4970 = (1'h0); (forvar4970 < (2'h2)); forvar4970 = (forvar4970 + (1'h1)))
                begin
                  reg4971 <= reg4619[(3'h6):(1'h0)];
                end
              for (forvar4972 = (1'h0); (forvar4972 < (2'h3)); forvar4972 = (forvar4972 + (1'h1)))
                begin
                  reg4973 <= {$unsigned(wire4799)};
                  for (forvar4974 = (1'h0); (forvar4974 < (2'h2)); forvar4974 = (forvar4974 + (1'h1)))
                    begin
                      reg4975 <= (reg4835 <<< (((reg4770 || reg4703) << (forvar4592 ?
                          forvar5006 : forvar4876)) != $unsigned(reg4995[(1'h0):(1'h0)])));
                    end
                  if ((^~$signed(forvar4643)))
                    begin
                      reg4976 <= forvar4750;
                      reg4977 <= reg4761[(2'h3):(2'h3)];
                      reg4978 <= $unsigned(reg4635[(4'hb):(4'ha)]);
                      reg4979 <= {($signed({reg4991}) ?
                              reg4990 : (~^(~&forvar4966)))};
                    end
                  else
                    begin
                      reg4976 <= $unsigned((~^$signed($signed(reg4853))));
                    end
                end
              if (reg4731)
                begin
                  reg4980 <= reg5022;
                  reg4981 <= ($unsigned({$signed(reg4995)}) ?
                      {reg4952} : (~reg4907[(1'h0):(1'h0)]));
                  if ({$signed($signed((~reg4843)))})
                    begin
                      reg4982 <= ($unsigned((&reg4645)) != (8'hae));
                      reg4983 <= reg4738[(1'h1):(1'h0)];
                      reg4984 <= $unsigned((^$unsigned($unsigned((8'hb0)))));
                      reg4985 <= $signed((+(((8'ha1) ^ (8'ha5)) ?
                          {reg4871} : reg4699[(4'h9):(4'h8)])));
                    end
                  else
                    begin
                      reg4982 <= ({((&reg4838) ?
                              (reg4811 ?
                                  forvar4884 : (8'hba)) : reg4977[(1'h0):(1'h0)])} ^~ (^(~^$signed(reg4818))));
                      reg4983 <= {$unsigned($unsigned((+forvar4931)))};
                      reg4984 <= $unsigned({$signed($signed(forvar4731))});
                    end
                  reg4986 <= ({reg4840[(4'hd):(1'h1)]} ?
                      (^~reg4734[(2'h3):(1'h1)]) : (-reg4750));
                end
              else
                begin
                  reg4980 <= reg5015[(4'he):(3'h7)];
                end
            end
          else
            begin
              for (forvar4966 = (1'h0); (forvar4966 < (1'h1)); forvar4966 = (forvar4966 + (1'h1)))
                begin
                  for (forvar4967 = (1'h0); (forvar4967 < (1'h1)); forvar4967 = (forvar4967 + (1'h1)))
                    begin
                      reg4968 <= (reg4695[(2'h2):(2'h2)] ?
                          (~forvar4604[(1'h0):(1'h0)]) : (({reg4610} ?
                              (|(8'hb3)) : (reg4657 ?
                                  (8'hb0) : forvar4603)) ^~ $signed($unsigned(forvar4909))));
                    end
                  for (forvar4969 = (1'h0); (forvar4969 < (1'h1)); forvar4969 = (forvar4969 + (1'h1)))
                    begin
                      reg4970 <= (({$unsigned(reg4978)} <= forvar4995[(2'h2):(2'h2)]) == (^~reg4668));
                      reg4971 <= {reg4645};
                      reg4972 <= {reg5022[(3'h4):(1'h0)]};
                    end
                  for (forvar4973 = (1'h0); (forvar4973 < (2'h2)); forvar4973 = (forvar4973 + (1'h1)))
                    begin
                      reg4974 <= ((|($signed(reg5017) ?
                          (~^forvar4593) : (~&reg4918))) & (!reg4664));
                    end
                end
            end
          reg4987 <= $signed(forvar4775);
          if ($unsigned($unsigned(($signed(reg4636) ^ reg4756))))
            begin
              reg4988 <= $signed($signed(reg4618[(2'h2):(1'h1)]));
              for (forvar4989 = (1'h0); (forvar4989 < (2'h3)); forvar4989 = (forvar4989 + (1'h1)))
                begin
                  if ($signed(reg4855))
                    begin
                      reg4990 <= ($unsigned($signed($unsigned(forvar4771))) <= forvar4988);
                    end
                  else
                    begin
                      reg4990 <= $signed($unsigned(($unsigned((8'ha8)) ?
                          $signed(reg4952) : (reg4740 >= reg4761))));
                      reg4991 <= (($unsigned((reg4688 - reg4668)) < (forvar4869 >= (reg4838 ~^ reg5018))) > (8'hb0));
                      reg4992 <= $signed(reg4821);
                    end
                  if ($signed($signed(reg4750)))
                    begin
                      reg4993 <= forvar4673;
                      reg4994 <= reg4668;
                      reg4995 <= (($signed((+reg4742)) << ((reg4843 == reg4789) ?
                          (reg4779 ?
                              reg5009 : reg4773) : (forvar4962 == (8'hb0)))) & reg4722[(1'h1):(1'h0)]);
                      reg4996 <= $unsigned((~$unsigned((&reg4879))));
                    end
                  else
                    begin
                      reg4993 <= (wire4798[(2'h2):(1'h0)] - ($signed($signed((8'hb9))) ?
                          $signed(reg4812) : reg4675[(4'h8):(3'h4)]));
                      reg4994 <= (~|reg4763[(4'hf):(1'h1)]);
                      reg4995 <= reg4682[(1'h1):(1'h1)];
                    end
                  if (forvar4802[(3'h6):(3'h6)])
                    begin
                      reg4997 <= $unsigned((-forvar4840));
                      reg4998 <= reg4811;
                      reg4999 <= (((reg4823[(3'h5):(1'h0)] & reg4973) ?
                              reg4601 : ($unsigned(reg5013) ?
                                  (forvar4975 >> forvar4640) : $unsigned(forvar4653))) ?
                          reg4961[(2'h2):(1'h0)] : {reg4999});
                    end
                  else
                    begin
                      reg4997 <= reg4578;
                      reg4998 <= $unsigned(($signed(reg4981) <= reg4738));
                    end
                  if ((-(((reg4868 ? reg5027 : reg4840) ?
                          (reg4578 ?
                              reg4856 : (8'ha0)) : reg4873[(1'h0):(1'h0)]) ?
                      reg4600 : reg4933[(4'h8):(2'h3)])))
                    begin
                      reg5000 <= (~&reg4743[(3'h5):(3'h5)]);
                      reg5001 <= reg5023[(2'h2):(1'h1)];
                      reg5002 <= ((^reg4592) ?
                          $signed($signed(forvar4789)) : (~reg4657));
                    end
                  else
                    begin
                      reg5000 <= reg4823;
                      reg5001 <= forvar4972;
                      reg5002 <= {({reg4596[(2'h2):(1'h0)]} ?
                              $signed($unsigned(forvar4869)) : (reg4774[(4'h8):(3'h5)] ?
                                  ((8'h9d) ? reg4596 : reg4845) : (~reg4853)))};
                    end
                end
              if (reg4660[(1'h1):(1'h1)])
                begin
                  for (forvar5003 = (1'h0); (forvar5003 < (2'h2)); forvar5003 = (forvar5003 + (1'h1)))
                    begin
                      reg5004 <= (^~(reg4853[(3'h4):(3'h4)] <<< (-(-reg4729))));
                      reg5005 <= ($unsigned($unsigned($unsigned(forvar4946))) < {$signed((reg4999 & forvar4779))});
                    end
                  for (forvar5006 = (1'h0); (forvar5006 < (1'h1)); forvar5006 = (forvar5006 + (1'h1)))
                    begin
                      reg5007 <= $signed((8'hac));
                      reg5008 <= ($unsigned(reg4787[(4'h9):(4'h8)]) ^ $signed($unsigned({reg4629})));
                      reg5009 <= $signed($signed((~(^reg4857))));
                      reg5010 <= (reg4845[(1'h0):(1'h0)] >> reg4609);
                    end
                end
              else
                begin
                  if ($unsigned(forvar4653[(3'h6):(1'h0)]))
                    begin
                      reg5003 <= ((8'hab) ?
                          $unsigned((8'haf)) : reg4850[(4'hf):(4'h9)]);
                      reg5004 <= {(~^((reg4637 ? reg4882 : reg5017) ?
                              reg5008 : (~|reg5029)))};
                      reg5005 <= (($signed($unsigned(forvar4673)) - $signed(reg4594[(3'h6):(3'h6)])) ?
                          ($unsigned({reg4582}) & {$signed(wire4574)}) : (reg4758 ?
                              ((8'had) ?
                                  $unsigned((8'ha1)) : forvar4755[(1'h1):(1'h1)]) : reg4862));
                      reg5006 <= forvar4849[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg5003 <= (forvar4879[(1'h0):(1'h0)] ?
                          ($signed((~^(8'h9e))) ?
                              (~|forvar4879[(1'h0):(1'h0)]) : forvar4802) : {$signed((~^reg4736))});
                      reg5004 <= (&(($unsigned(forvar4744) ~^ (forvar4848 > reg4590)) ?
                          $signed((~|forvar4581)) : (|$unsigned(reg4607))));
                      reg5005 <= $signed($signed($signed((!reg4945))));
                    end
                end
            end
          else
            begin
              if (reg4865[(1'h1):(1'h0)])
                begin
                  for (forvar4988 = (1'h0); (forvar4988 < (1'h1)); forvar4988 = (forvar4988 + (1'h1)))
                    begin
                      reg4989 <= $signed((~^$unsigned((|reg4789))));
                      reg4990 <= (reg4989 == reg4685[(1'h0):(1'h0)]);
                    end
                  for (forvar4991 = (1'h0); (forvar4991 < (2'h3)); forvar4991 = (forvar4991 + (1'h1)))
                    begin
                      reg4992 <= (+(8'hb8));
                      reg4993 <= (-forvar4581[(1'h1):(1'h1)]);
                      reg4994 <= $unsigned($signed($signed(reg4880[(1'h0):(1'h0)])));
                    end
                  if ($unsigned((reg4808[(1'h0):(1'h0)] != $signed({(8'had)}))))
                    begin
                      reg4995 <= $unsigned((~^((reg4776 ?
                          reg4646 : reg4623) ^ reg4919[(4'h8):(1'h1)])));
                      reg4996 <= (+($signed($unsigned(reg4678)) == (^{forvar4933})));
                      reg4997 <= ((($signed(forvar5009) + {forvar4737}) && reg4955[(1'h0):(1'h0)]) | forvar4946[(4'ha):(3'h5)]);
                      reg4998 <= ($unsigned(reg4635) ?
                          {$signed((reg4709 && (8'ha5)))} : (!$unsigned($signed(reg4683))));
                    end
                  else
                    begin
                      reg4995 <= $signed($signed((-(reg4998 ?
                          reg4823 : forvar4584))));
                    end
                  if (forvar4864)
                    begin
                      reg4999 <= ((-$unsigned((reg4928 ?
                          reg4631 : reg4633))) ^~ ({(-reg4803)} ?
                          ((reg4578 ?
                              reg4869 : reg4730) ^~ $signed(reg4628)) : ($unsigned((8'hae)) ?
                              $unsigned(reg4911) : (reg4598 ?
                                  reg4914 : reg4909))));
                      reg5000 <= (+(({forvar4750} ? {wire4574} : reg4850) ?
                          (~^$signed(forvar4899)) : (((8'hba) ?
                              forvar4753 : forvar4944) <= $signed(reg4584))));
                    end
                  else
                    begin
                      reg4999 <= $signed(($signed(reg4770) ?
                          $unsigned(reg4761) : (~&$unsigned((8'ha5)))));
                      reg5000 <= reg4741[(2'h2):(2'h2)];
                      reg5001 <= {$unsigned(forvar4603)};
                    end
                end
              else
                begin
                  if ((({(forvar4717 || (8'hae))} ?
                          (8'h9c) : (+reg4962[(3'h5):(3'h4)])) ?
                      forvar4642[(2'h2):(1'h0)] : $unsigned(reg5004[(1'h1):(1'h0)])))
                    begin
                      reg4988 <= $signed((8'had));
                      reg4989 <= forvar4910[(3'h4):(2'h2)];
                      reg4990 <= (reg4749 ?
                          (8'hb3) : $unsigned($signed(reg4996[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg4988 <= ((-reg4932) ?
                          {$unsigned($signed((8'h9f)))} : (reg4871 ?
                              $signed((reg4838 ?
                                  forvar4915 : reg4911)) : forvar4972));
                    end
                end
              for (forvar5002 = (1'h0); (forvar5002 < (1'h0)); forvar5002 = (forvar5002 + (1'h1)))
                begin
                  for (forvar5003 = (1'h0); (forvar5003 < (2'h2)); forvar5003 = (forvar5003 + (1'h1)))
                    begin
                      reg5004 <= forvar4877;
                    end
                  for (forvar5005 = (1'h0); (forvar5005 < (1'h1)); forvar5005 = (forvar5005 + (1'h1)))
                    begin
                      reg5006 <= reg4787[(1'h1):(1'h1)];
                      reg5007 <= ((($unsigned(forvar4763) ?
                              reg4901[(2'h3):(2'h2)] : $signed((8'hb8))) << (^(+reg4677))) ?
                          $signed(reg4861) : (((forvar4858 ?
                                  forvar4643 : reg5001) ?
                              $unsigned(reg4715) : $signed(forvar4967)) <<< reg4618));
                    end
                  for (forvar5008 = (1'h0); (forvar5008 < (1'h1)); forvar5008 = (forvar5008 + (1'h1)))
                    begin
                      reg5009 <= (reg4720[(2'h2):(1'h0)] ?
                          $signed({(reg4626 ?
                                  reg4927 : forvar4696)}) : (((&(8'hb5)) < ((8'hb9) ?
                                  (8'ha7) : (8'ha7))) ?
                              (+reg5022[(3'h7):(1'h1)]) : {reg4895}));
                    end
                  reg5010 <= (wire4575 <<< (!((reg4881 ? reg4578 : reg4679) ?
                      forvar4598[(4'hd):(3'h7)] : $unsigned(reg5021))));
                end
              if ({({reg4775[(2'h2):(2'h2)]} <= (forvar4581[(2'h2):(2'h2)] ?
                      reg4654 : reg4976))})
                begin
                  for (forvar5011 = (1'h0); (forvar5011 < (1'h1)); forvar5011 = (forvar5011 + (1'h1)))
                    begin
                      reg5012 <= (((((8'ha2) + forvar4858) ?
                          reg4670[(1'h1):(1'h0)] : $signed(forvar4663)) & (+$unsigned(reg4982))) & reg4933);
                      reg5013 <= $signed((~$unsigned((reg4614 || reg4643))));
                      reg5014 <= reg4837;
                    end
                  for (forvar5015 = (1'h0); (forvar5015 < (2'h3)); forvar5015 = (forvar5015 + (1'h1)))
                    begin
                      reg5016 <= (reg4938[(4'hd):(4'hc)] * reg4747[(4'h8):(4'h8)]);
                    end
                  if (reg4745)
                    begin
                      reg5017 <= reg4915[(3'h5):(1'h0)];
                    end
                  else
                    begin
                      reg5017 <= reg4885;
                      reg5018 <= ((reg5022 <<< $signed(forvar4698)) ?
                          (~&$signed((^reg4764))) : (($unsigned(reg4862) * $signed(reg4835)) <= ({reg4677} >>> $signed(forvar4731))));
                      reg5019 <= $unsigned(forvar4879);
                    end
                end
              else
                begin
                  for (forvar5011 = (1'h0); (forvar5011 < (2'h3)); forvar5011 = (forvar5011 + (1'h1)))
                    begin
                      reg5012 <= ($signed(({reg4913} > {reg4789})) << (~({reg4627} ?
                          $unsigned((8'ha5)) : $unsigned((8'ha6)))));
                      reg5013 <= $signed($unsigned($signed($signed(reg4638))));
                      reg5014 <= reg4760[(1'h1):(1'h1)];
                      reg5015 <= forvar4593;
                    end
                  if ((|$signed(reg4755[(1'h0):(1'h0)])))
                    begin
                      reg5016 <= reg4582[(1'h0):(1'h0)];
                      reg5017 <= reg4828;
                      reg5018 <= ((reg4796 & ((reg4773 ?
                          forvar4613 : forvar4737) * $signed(forvar4770))) >= reg4649[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg5016 <= forvar4962;
                      reg5017 <= $signed((($unsigned(forvar4696) || (forvar5029 * reg4666)) * ((forvar4966 ?
                          reg4633 : reg4783) * reg4637[(4'ha):(1'h0)])));
                      reg5018 <= ((|({wire4940} ?
                              (reg4932 ? forvar4656 : forvar4826) : reg4625)) ?
                          (&({reg5033} ^ reg4701)) : $signed($unsigned((~(8'hb6)))));
                      reg5019 <= $signed((^reg4948));
                    end
                  for (forvar5020 = (1'h0); (forvar5020 < (2'h2)); forvar5020 = (forvar5020 + (1'h1)))
                    begin
                      reg5021 <= $signed((~^$unsigned(forvar4779)));
                      reg5022 <= $signed({$unsigned((forvar4795 ^ reg4892))});
                    end
                end
            end
        end
      if (reg4974[(1'h0):(1'h0)])
        begin
          if ({reg4683[(2'h2):(2'h2)]})
            begin
              reg5035 <= (~$signed(reg4850));
              for (forvar5036 = (1'h0); (forvar5036 < (1'h1)); forvar5036 = (forvar5036 + (1'h1)))
                begin
                  if (forvar4912)
                    begin
                      reg5037 <= $unsigned((((~&reg4727) == reg4733) ^ $signed((|reg5013))));
                      reg5038 <= reg4636;
                    end
                  else
                    begin
                      reg5037 <= forvar4920[(3'h5):(1'h0)];
                      reg5038 <= reg4703;
                      reg5039 <= reg4956[(1'h0):(1'h0)];
                    end
                end
              reg5040 <= (reg4938 ?
                  $unsigned($signed((~reg4981))) : reg4889[(4'h9):(4'h8)]);
            end
          else
            begin
              for (forvar5035 = (1'h0); (forvar5035 < (2'h2)); forvar5035 = (forvar5035 + (1'h1)))
                begin
                  if ({forvar4817[(3'h4):(2'h3)]})
                    begin
                      reg5036 <= $unsigned((-{(~&reg4766)}));
                      reg5037 <= (($signed((reg4870 <= forvar4578)) | {(~^reg4709)}) ?
                          reg5026 : ($unsigned((reg4816 ?
                              forvar4879 : reg4614)) ^~ reg4942));
                      reg5038 <= $signed($signed((((8'had) ?
                          reg4746 : reg5001) <<< (8'ha3))));
                      reg5039 <= reg4913;
                    end
                  else
                    begin
                      reg5036 <= $signed(((reg5027[(1'h1):(1'h1)] ?
                          $signed(reg4642) : reg4793[(4'he):(4'h8)]) & ((reg4583 ?
                              (8'ha0) : reg5006) ?
                          reg4865 : (|(8'had)))));
                    end
                  if (((-(~|$unsigned(forvar4749))) ?
                      ((!(reg4869 ? reg4852 : reg4888)) ?
                          ((~&forvar4829) < wire4940) : {(reg4777 ?
                                  forvar5011 : reg4669)}) : ((forvar4758 ?
                              {reg4831} : (forvar4674 << (8'haf))) ?
                          reg5022[(2'h3):(1'h1)] : $signed((forvar5003 == reg4942)))))
                    begin
                      reg5040 <= {$signed(($unsigned(reg4687) ?
                              (reg4880 >>> (8'hb6)) : (&reg4841)))};
                      reg5041 <= forvar4826;
                    end
                  else
                    begin
                      reg5040 <= ((~^$unsigned((forvar4843 ^ reg4773))) ?
                          (8'had) : $unsigned($unsigned({(8'ha1)})));
                      reg5041 <= reg4638;
                      reg5042 <= $unsigned($signed(((wire4940 <= forvar4972) ?
                          ((8'hb6) ^ reg4766) : (reg4904 >= reg4787))));
                      reg5043 <= $signed((~&$signed((-reg4699))));
                    end
                  if (($signed(reg4768) * (((^~reg4627) ?
                      reg4687[(3'h5):(1'h1)] : $signed(reg4959)) & $signed({reg4682}))))
                    begin
                      reg5044 <= $signed($signed($unsigned($unsigned(reg4753))));
                      reg5045 <= $signed(($unsigned(reg4903) ?
                          $unsigned((reg4952 ?
                              forvar5005 : (8'h9c))) : forvar4766));
                      reg5046 <= (-reg4999);
                    end
                  else
                    begin
                      reg5044 <= $unsigned((reg4883[(2'h2):(1'h0)] >>> {reg4697}));
                      reg5045 <= $signed(reg4781[(3'h4):(1'h1)]);
                      reg5046 <= reg4695[(3'h7):(2'h2)];
                      reg5047 <= ($unsigned((~|reg5018[(3'h7):(2'h3)])) - (|{$unsigned(forvar4727)}));
                    end
                  for (forvar5048 = (1'h0); (forvar5048 < (2'h2)); forvar5048 = (forvar5048 + (1'h1)))
                    begin
                      reg5049 <= ((^$unsigned({forvar4738})) ?
                          (8'ha9) : {$unsigned(reg4766[(1'h1):(1'h1)])});
                      reg5050 <= ({reg4805} ? (^{(!forvar4715)}) : reg4902);
                      reg5051 <= reg4832;
                      reg5052 <= reg4794;
                    end
                end
              for (forvar5053 = (1'h0); (forvar5053 < (1'h1)); forvar5053 = (forvar5053 + (1'h1)))
                begin
                  for (forvar5054 = (1'h0); (forvar5054 < (2'h2)); forvar5054 = (forvar5054 + (1'h1)))
                    begin
                      reg5055 <= $unsigned({($unsigned(forvar4851) ?
                              $unsigned(reg4883) : $signed(forvar4659))});
                      reg5056 <= forvar4617[(2'h2):(1'h0)];
                      reg5057 <= reg5039;
                    end
                  reg5058 <= ($unsigned((wire4798[(4'h8):(3'h6)] - $signed(reg4627))) ?
                      $signed(((forvar4753 < reg4987) ?
                          (reg5006 == reg4642) : (reg5041 * reg4910))) : (forvar4611 < (8'ha2)));
                  for (forvar5059 = (1'h0); (forvar5059 < (1'h1)); forvar5059 = (forvar5059 + (1'h1)))
                    begin
                      reg5060 <= {(+reg4960)};
                    end
                  reg5061 <= reg5023[(4'h8):(2'h2)];
                end
            end
          for (forvar5062 = (1'h0); (forvar5062 < (1'h0)); forvar5062 = (forvar5062 + (1'h1)))
            begin
              for (forvar5063 = (1'h0); (forvar5063 < (1'h0)); forvar5063 = (forvar5063 + (1'h1)))
                begin
                  for (forvar5064 = (1'h0); (forvar5064 < (2'h2)); forvar5064 = (forvar5064 + (1'h1)))
                    begin
                      reg5065 <= $unsigned($unsigned((((8'h9e) ?
                              reg4886 : reg4777) ?
                          (reg4905 <= forvar4996) : (reg4739 >>> (8'ha5)))));
                      reg5066 <= $unsigned($signed(forvar4688));
                      reg5067 <= reg4845[(1'h0):(1'h0)];
                    end
                  for (forvar5068 = (1'h0); (forvar5068 < (2'h3)); forvar5068 = (forvar5068 + (1'h1)))
                    begin
                      reg5069 <= $unsigned($signed({(reg4888 < reg4930)}));
                      reg5070 <= $unsigned(($unsigned($unsigned(forvar4933)) ?
                          (~^(~&forvar4578)) : reg4647));
                      reg5071 <= (~|((+forvar4923) | reg4747[(3'h6):(2'h2)]));
                    end
                  if ($unsigned(reg4912))
                    begin
                      reg5072 <= $signed(forvar4962[(3'h7):(3'h6)]);
                      reg5073 <= reg4782[(2'h3):(1'h1)];
                      reg5074 <= ((reg4770[(3'h4):(1'h0)] ?
                          reg4625[(4'h9):(1'h0)] : $signed($signed((8'haf)))) <<< (!(^~(reg4676 ?
                          reg5067 : forvar4957))));
                    end
                  else
                    begin
                      reg5072 <= {reg4966};
                      reg5073 <= {({$signed(forvar4688)} ?
                              forvar4946[(3'h5):(1'h0)] : ((^~(8'hb2)) ?
                                  forvar4773 : $unsigned(reg4579)))};
                      reg5074 <= ($signed(reg4597) ?
                          {$unsigned(reg4905)} : ($unsigned((reg4692 ?
                                  reg4910 : reg5019)) ?
                              {$unsigned(reg4794)} : {reg4614[(3'h4):(2'h3)]}));
                    end
                end
              for (forvar5075 = (1'h0); (forvar5075 < (2'h3)); forvar5075 = (forvar5075 + (1'h1)))
                begin
                  for (forvar5076 = (1'h0); (forvar5076 < (1'h0)); forvar5076 = (forvar5076 + (1'h1)))
                    begin
                      reg5077 <= (8'hb5);
                      reg5078 <= forvar4766;
                      reg5079 <= $unsigned((~reg4846[(2'h3):(1'h0)]));
                    end
                end
            end
          reg5080 <= ($signed({((8'h9e) >> reg4906)}) <<< $unsigned(($signed(reg4678) ?
              (~|reg4607) : (reg4856 ? reg4725 : reg4660))));
          reg5081 <= $unsigned(reg4611);
        end
      else
        begin
          for (forvar5035 = (1'h0); (forvar5035 < (1'h1)); forvar5035 = (forvar5035 + (1'h1)))
            begin
              if ((((~((8'hac) - reg4688)) | ($unsigned(reg4992) ?
                  reg4723 : (reg4950 ?
                      reg4943 : reg4594))) - (reg4790[(3'h5):(2'h3)] >> (reg5037 != forvar4760))))
                begin
                  for (forvar5036 = (1'h0); (forvar5036 < (1'h0)); forvar5036 = (forvar5036 + (1'h1)))
                    begin
                      reg5037 <= (~|(reg4861[(1'h1):(1'h0)] >> {(&forvar4977)}));
                      reg5038 <= reg4687[(4'hb):(2'h3)];
                      reg5039 <= reg4911[(3'h7):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar5036 = (1'h0); (forvar5036 < (2'h2)); forvar5036 = (forvar5036 + (1'h1)))
                    begin
                      reg5037 <= ($signed(reg5071[(2'h2):(1'h1)]) < $signed(((reg4949 <= forvar4890) == (reg4714 ?
                          reg4670 : reg4796))));
                      reg5038 <= (&(((~|reg4900) ?
                              forvar4766[(1'h0):(1'h0)] : $unsigned(reg5017)) ?
                          reg4928 : {(reg4859 >>> (8'ha9))}));
                    end
                  for (forvar5039 = (1'h0); (forvar5039 < (1'h1)); forvar5039 = (forvar5039 + (1'h1)))
                    begin
                      reg5040 <= ({(~&{reg4767})} || reg4779[(2'h2):(1'h1)]);
                      reg5041 <= $unsigned(reg4695[(4'ha):(2'h2)]);
                      reg5042 <= reg4895;
                    end
                  for (forvar5043 = (1'h0); (forvar5043 < (2'h2)); forvar5043 = (forvar5043 + (1'h1)))
                    begin
                      reg5044 <= {($signed({reg5023}) ?
                              ({reg4839} ?
                                  (reg4975 ?
                                      (8'hb7) : reg5041) : {forvar4946}) : $signed(reg5040))};
                      reg5045 <= reg4904[(1'h0):(1'h0)];
                      reg5046 <= $unsigned($signed((+(~&reg4691))));
                      reg5047 <= $signed((8'ha6));
                    end
                end
              if ($signed(($unsigned($unsigned(reg4847)) ^ {$signed(reg4627)})))
                begin
                  reg5048 <= reg4897[(1'h0):(1'h0)];
                  for (forvar5049 = (1'h0); (forvar5049 < (1'h0)); forvar5049 = (forvar5049 + (1'h1)))
                    begin
                      reg5050 <= ((|$unsigned({forvar4829})) ?
                          $unsigned((~&{reg4993})) : $signed(reg4691));
                      reg5051 <= (reg5004 * {$unsigned($signed((8'ha1)))});
                      reg5052 <= ($signed(forvar5029[(3'h7):(2'h3)]) ?
                          (($signed(reg4870) ?
                                  $signed(reg4804) : (forvar4884 ^ (8'hb3))) ?
                              forvar4653[(1'h1):(1'h0)] : forvar4929[(4'hc):(4'hc)]) : ((~|forvar4737) ?
                              reg4973 : (^~(reg4751 ? reg4692 : reg4808))));
                    end
                  for (forvar5053 = (1'h0); (forvar5053 < (2'h2)); forvar5053 = (forvar5053 + (1'h1)))
                    begin
                      reg5054 <= ($unsigned(((~forvar4689) ?
                              forvar4913[(1'h0):(1'h0)] : {forvar4654})) ?
                          {($unsigned((8'hb6)) <<< $unsigned(reg4989))} : forvar4826);
                      reg5055 <= reg4925[(3'h7):(2'h2)];
                    end
                  if ($unsigned($unsigned(forvar4923[(2'h2):(1'h1)])))
                    begin
                      reg5056 <= (reg4664[(4'h8):(3'h4)] ?
                          {(^(forvar5062 ? reg5057 : reg4987))} : reg4686);
                    end
                  else
                    begin
                      reg5056 <= ($unsigned($unsigned(((8'haa) ?
                              forvar4780 : forvar4824))) ?
                          (~reg4669[(2'h2):(1'h1)]) : (&$signed((reg4854 - reg4912))));
                      reg5057 <= (reg4928 ?
                          forvar5075 : (reg4907 ?
                              reg4914[(3'h5):(1'h0)] : (~^(8'h9f))));
                      reg5058 <= (~reg4774[(4'h9):(4'h9)]);
                      reg5059 <= (8'hab);
                    end
                end
              else
                begin
                  for (forvar5048 = (1'h0); (forvar5048 < (2'h2)); forvar5048 = (forvar5048 + (1'h1)))
                    begin
                      reg5049 <= (forvar4755 * $unsigned(reg4924));
                      reg5050 <= $unsigned((((reg4986 ? reg4746 : reg4649) ?
                          (reg5027 ?
                              reg4744 : reg4926) : (-forvar4911)) >= (8'ha5)));
                    end
                  for (forvar5051 = (1'h0); (forvar5051 < (1'h1)); forvar5051 = (forvar5051 + (1'h1)))
                    begin
                      reg5052 <= (^$unsigned($unsigned((reg4678 ?
                          reg4715 : forvar4970))));
                      reg5053 <= $signed(reg4909[(3'h7):(3'h6)]);
                      reg5054 <= ((!{$unsigned(reg4615)}) > $unsigned(forvar4654[(1'h0):(1'h0)]));
                      reg5055 <= forvar4802;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg4741)
        begin
          if (reg4912[(1'h0):(1'h0)])
            begin
              for (forvar5082 = (1'h0); (forvar5082 < (2'h3)); forvar5082 = (forvar5082 + (1'h1)))
                begin
                  reg5083 <= $unsigned((reg4796 != $unsigned($signed(reg4866))));
                  for (forvar5084 = (1'h0); (forvar5084 < (1'h0)); forvar5084 = (forvar5084 + (1'h1)))
                    begin
                      reg5085 <= ((reg4860 ?
                              $signed($unsigned((8'hb3))) : ($unsigned(reg5046) ?
                                  (reg4830 == forvar4980) : (reg4904 | (8'hab)))) ?
                          {(8'hb7)} : $signed(((reg4882 ?
                                  forvar4604 : reg4977) ?
                              (reg4981 <= forvar5043) : $unsigned(forvar4654))));
                      reg5086 <= {(~^forvar4884)};
                      reg5087 <= reg4836[(2'h2):(1'h0)];
                      reg5088 <= (reg4949 ?
                          $signed(((8'ha3) - (8'h9c))) : reg5045);
                    end
                end
              if (reg4812[(2'h2):(2'h2)])
                begin
                  if (reg5004)
                    begin
                      reg5089 <= (^~$signed($signed($unsigned((8'ha2)))));
                      reg5090 <= {$signed(reg5022[(1'h1):(1'h0)])};
                      reg5091 <= $unsigned((~^forvar4972[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg5089 <= reg4708;
                      reg5090 <= reg4613;
                      reg5091 <= ($unsigned({(forvar5051 ?
                              reg4726 : reg4859)}) || ((^~$signed(reg4954)) ?
                          reg4960 : ((reg5042 ?
                              reg4582 : forvar4616) != (~reg4596))));
                      reg5092 <= $unsigned((($unsigned(forvar4933) << (forvar4908 <<< (8'hae))) <= (reg5053 ^ (forvar4645 ?
                          forvar4727 : forvar4608))));
                    end
                end
              else
                begin
                  for (forvar5089 = (1'h0); (forvar5089 < (1'h0)); forvar5089 = (forvar5089 + (1'h1)))
                    begin
                      reg5090 <= ($unsigned(((reg4937 ?
                              reg4779 : forvar5054) > (|forvar4911))) ?
                          $signed($signed(forvar4611[(3'h7):(3'h6)])) : ((reg5053 - (reg4725 < forvar4598)) < forvar5082[(1'h1):(1'h1)]));
                      reg5091 <= {$unsigned(forvar5036[(3'h4):(2'h3)])};
                    end
                end
              for (forvar5093 = (1'h0); (forvar5093 < (2'h3)); forvar5093 = (forvar5093 + (1'h1)))
                begin
                  if ($unsigned(reg5085))
                    begin
                      reg5094 <= forvar4766;
                      reg5095 <= $unsigned((~|($unsigned(reg4886) - (|forvar4913))));
                    end
                  else
                    begin
                      reg5094 <= wire4798[(3'h5):(2'h2)];
                      reg5095 <= (+(forvar4809[(1'h0):(1'h0)] ?
                          $signed($signed(forvar4607)) : reg4604[(2'h3):(1'h0)]));
                      reg5096 <= (8'hab);
                      reg5097 <= {$unsigned(((reg4745 ? reg4604 : forvar4616) ?
                              (reg4893 ?
                                  reg4585 : reg5095) : $unsigned(reg4583)))};
                    end
                  for (forvar5098 = (1'h0); (forvar5098 < (2'h3)); forvar5098 = (forvar5098 + (1'h1)))
                    begin
                      reg5099 <= reg4786[(2'h2):(1'h1)];
                      reg5100 <= (reg4915 < (reg4580 == reg4738));
                      reg5101 <= reg4953;
                    end
                  for (forvar5102 = (1'h0); (forvar5102 < (1'h1)); forvar5102 = (forvar5102 + (1'h1)))
                    begin
                      reg5103 <= ((~(reg4700 ? reg4907 : {reg4631})) ?
                          (8'hae) : ({reg4979[(1'h0):(1'h0)]} ?
                              reg4934 : reg4602[(3'h4):(1'h1)]));
                    end
                  if (($unsigned($signed($unsigned(reg4885))) - (reg4825[(2'h2):(2'h2)] ^ ((reg4872 | reg4954) && {(8'ha0)}))))
                    begin
                      reg5104 <= forvar5005[(4'h8):(1'h0)];
                      reg5105 <= forvar4817[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg5104 <= reg5048[(2'h2):(2'h2)];
                    end
                end
            end
          else
            begin
              if (reg4701)
                begin
                  reg5082 <= $unsigned($signed(($signed(reg5079) == $signed((8'hb8)))));
                  for (forvar5083 = (1'h0); (forvar5083 < (2'h2)); forvar5083 = (forvar5083 + (1'h1)))
                    begin
                      reg5084 <= reg4769[(3'h4):(1'h1)];
                      reg5085 <= forvar4755;
                      reg5086 <= reg4656[(2'h3):(1'h1)];
                    end
                end
              else
                begin
                  reg5082 <= ((reg4587 ?
                          $signed(((8'hae) ?
                              forvar4989 : reg4636)) : reg4853[(2'h2):(1'h0)]) ?
                      reg4856[(1'h0):(1'h0)] : (8'ha8));
                  if ((forvar4770[(2'h3):(1'h1)] ?
                      {forvar4760} : ($unsigned($unsigned(reg4867)) >>> (forvar4588 ?
                          reg4602[(3'h4):(1'h1)] : reg5007))))
                    begin
                      reg5083 <= $unsigned($signed((forvar5075 ?
                          {reg4932} : {forvar4946})));
                      reg5084 <= (reg4583[(4'hd):(4'hb)] >> (+((&(8'ha0)) >> reg5023[(1'h1):(1'h0)])));
                      reg5085 <= reg4604;
                    end
                  else
                    begin
                      reg5083 <= forvar4698;
                    end
                end
              reg5087 <= {$signed(($unsigned(reg4697) ?
                      $signed(reg5042) : forvar4843[(4'he):(3'h5)]))};
              for (forvar5088 = (1'h0); (forvar5088 < (2'h3)); forvar5088 = (forvar5088 + (1'h1)))
                begin
                  reg5089 <= (8'had);
                end
              for (forvar5090 = (1'h0); (forvar5090 < (2'h3)); forvar5090 = (forvar5090 + (1'h1)))
                begin
                  if ((~^reg4671[(3'h4):(2'h3)]))
                    begin
                      reg5091 <= $unsigned($unsigned(reg4605[(4'hb):(4'h8)]));
                      reg5092 <= ((($signed(reg4853) != $unsigned((8'hb2))) ?
                              (reg4981[(4'h9):(2'h2)] ?
                                  (reg4837 ?
                                      (8'hb5) : (8'ha7)) : {forvar4801}) : $signed((+reg4946))) ?
                          ({reg4968} ?
                              reg4921[(4'h9):(3'h5)] : forvar4781) : (^~$unsigned($signed(reg4776))));
                      reg5093 <= forvar4640;
                    end
                  else
                    begin
                      reg5091 <= $unsigned(forvar4688[(3'h5):(3'h5)]);
                      reg5092 <= (^~(((!reg4907) <= $signed(reg5042)) ?
                          ($signed(reg4991) ?
                              (~|reg4683) : (~reg4646)) : reg4629[(3'h5):(3'h4)]));
                      reg5093 <= $signed((({(8'had)} ?
                              (reg5074 ? reg4756 : reg4840) : (!reg5021)) ?
                          reg5103[(3'h4):(3'h4)] : {reg4695}));
                    end
                end
            end
          for (forvar5106 = (1'h0); (forvar5106 < (2'h3)); forvar5106 = (forvar5106 + (1'h1)))
            begin
              reg5107 <= $signed({$signed((8'ha4))});
              for (forvar5108 = (1'h0); (forvar5108 < (2'h3)); forvar5108 = (forvar5108 + (1'h1)))
                begin
                  for (forvar5109 = (1'h0); (forvar5109 < (2'h3)); forvar5109 = (forvar5109 + (1'h1)))
                    begin
                      reg5110 <= $signed(forvar4653[(4'hc):(4'h8)]);
                      reg5111 <= reg4853[(1'h0):(1'h0)];
                      reg5112 <= (~(($unsigned(reg4997) ?
                              ((8'ha3) ? reg4925 : (8'hb2)) : reg4924) ?
                          $signed(forvar4779[(4'hf):(4'ha)]) : $unsigned(((8'hb3) ?
                              forvar5005 : reg5089))));
                    end
                end
            end
        end
      else
        begin
          if ({reg5091[(4'ha):(3'h4)]})
            begin
              reg5082 <= (reg4629 ~^ reg4733);
            end
          else
            begin
              for (forvar5082 = (1'h0); (forvar5082 < (2'h3)); forvar5082 = (forvar5082 + (1'h1)))
                begin
                  for (forvar5083 = (1'h0); (forvar5083 < (2'h2)); forvar5083 = (forvar5083 + (1'h1)))
                    begin
                      reg5084 <= $unsigned(((8'ha5) ?
                          reg5097 : forvar5019[(1'h1):(1'h0)]));
                    end
                  for (forvar5085 = (1'h0); (forvar5085 < (1'h1)); forvar5085 = (forvar5085 + (1'h1)))
                    begin
                      reg5086 <= (((~$signed((8'h9e))) >> reg4786[(2'h2):(1'h1)]) ?
                          $unsigned($signed($unsigned(reg4904))) : (((8'ha0) ?
                              $unsigned(reg4984) : reg4968[(3'h6):(1'h1)]) && (~|$signed((8'hb7)))));
                      reg5087 <= $unsigned(forvar4824[(1'h0):(1'h0)]);
                      reg5088 <= $unsigned(((forvar4795[(4'hb):(3'h6)] ?
                          {reg5061} : $signed((8'hb7))) ~^ $unsigned($unsigned(reg4577))));
                    end
                  for (forvar5089 = (1'h0); (forvar5089 < (2'h2)); forvar5089 = (forvar5089 + (1'h1)))
                    begin
                      reg5090 <= reg5052[(3'h4):(1'h0)];
                    end
                end
              if ((~forvar4593[(3'h4):(1'h0)]))
                begin
                  for (forvar5091 = (1'h0); (forvar5091 < (2'h3)); forvar5091 = (forvar5091 + (1'h1)))
                    begin
                      reg5092 <= reg4820[(3'h6):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar5091 = (1'h0); (forvar5091 < (1'h0)); forvar5091 = (forvar5091 + (1'h1)))
                    begin
                      reg5092 <= (forvar5002 << reg4731);
                      reg5093 <= (|{(~^{forvar5088})});
                    end
                  if ((({$signed(reg4783)} >= ((!reg4880) | (^~reg4991))) ?
                      reg4839 : {$unsigned(reg4838[(1'h0):(1'h0)])}))
                    begin
                      reg5094 <= (~|(8'ha0));
                      reg5095 <= (^~($signed((8'h9e)) != reg4816));
                      reg5096 <= (8'hb1);
                    end
                  else
                    begin
                      reg5094 <= {$unsigned({(~&(8'h9f))})};
                      reg5095 <= (8'ha1);
                      reg5096 <= {{$signed((wire4799 ^ (8'ha0)))}};
                      reg5097 <= ({{reg4913}} ?
                          ((forvar4577 >>> (forvar4877 + reg4768)) ?
                              $unsigned(reg4956) : $signed(reg4731)) : (reg4643[(1'h0):(1'h0)] >>> $signed((reg4883 >> (8'hba)))));
                    end
                  for (forvar5098 = (1'h0); (forvar5098 < (1'h0)); forvar5098 = (forvar5098 + (1'h1)))
                    begin
                      reg5099 <= {reg4630[(3'h5):(3'h5)]};
                      reg5100 <= wire4798[(2'h3):(2'h3)];
                      reg5101 <= {(|(&forvar4609))};
                    end
                end
              for (forvar5102 = (1'h0); (forvar5102 < (1'h0)); forvar5102 = (forvar5102 + (1'h1)))
                begin
                  reg5103 <= $signed($signed({$unsigned((8'hac))}));
                  for (forvar5104 = (1'h0); (forvar5104 < (2'h2)); forvar5104 = (forvar5104 + (1'h1)))
                    begin
                      reg5105 <= {(reg4695 ?
                              ((&forvar4837) ?
                                  reg4893[(1'h0):(1'h0)] : reg4805) : (reg4693[(3'h4):(1'h1)] ?
                                  (reg4811 ? reg4590 : reg4629) : forvar5064))};
                      reg5106 <= $unsigned($signed(reg4856));
                      reg5107 <= reg5021;
                    end
                end
              reg5108 <= (reg4841[(4'hf):(4'hb)] ?
                  reg4583[(4'h8):(3'h5)] : (reg4915[(4'h8):(1'h0)] != $unsigned((reg5106 > forvar4659))));
            end
          if ({reg5078})
            begin
              for (forvar5109 = (1'h0); (forvar5109 < (2'h2)); forvar5109 = (forvar5109 + (1'h1)))
                begin
                  if (({$signed(reg4933[(4'hc):(1'h0)])} ?
                      (8'ha1) : reg5051[(3'h6):(2'h2)]))
                    begin
                      reg5110 <= $unsigned((forvar4616[(4'hc):(3'h6)] ?
                          reg5041[(4'hc):(2'h3)] : $signed((reg4984 ?
                              forvar5009 : forvar5002))));
                      reg5111 <= reg4854;
                      reg5112 <= $unsigned((reg4869[(4'he):(4'h9)] | reg4887[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg5110 <= $unsigned({($signed(reg4873) ?
                              (forvar5109 ?
                                  (8'hb1) : forvar4806) : reg5091[(1'h1):(1'h1)])});
                      reg5111 <= $unsigned((((reg5013 ? reg4848 : reg5023) ?
                              (8'hb1) : {(8'ha7)}) ?
                          reg4774 : ((forvar4609 <<< reg4856) >>> forvar4973[(4'ha):(3'h7)])));
                      reg5112 <= $unsigned((!forvar4611));
                    end
                  reg5113 <= $signed(($signed({(8'hb2)}) ?
                      {{reg4992}} : reg4781));
                  for (forvar5114 = (1'h0); (forvar5114 < (1'h1)); forvar5114 = (forvar5114 + (1'h1)))
                    begin
                      reg5115 <= (|(reg4601[(1'h0):(1'h0)] ?
                          ((~&reg4938) - (reg4593 ?
                              (8'hab) : reg4735)) : $unsigned({(8'hae)})));
                      reg5116 <= ({forvar4607[(1'h1):(1'h1)]} - ((((8'h9c) | forvar4766) & $signed(reg5069)) && (reg5025 || (reg4782 == reg5002))));
                    end
                end
              if ((forvar4603 ?
                  $unsigned((((8'hac) << forvar4809) ?
                      reg4834 : (~|forvar4689))) : reg4730[(4'ha):(3'h4)]))
                begin
                  if (forvar4988)
                    begin
                      reg5117 <= {reg4850};
                    end
                  else
                    begin
                      reg5117 <= (8'ha6);
                    end
                end
              else
                begin
                  for (forvar5117 = (1'h0); (forvar5117 < (1'h1)); forvar5117 = (forvar5117 + (1'h1)))
                    begin
                      reg5118 <= (8'h9d);
                      reg5119 <= forvar5108[(4'h9):(4'h9)];
                    end
                  reg5120 <= reg5066[(2'h2):(2'h2)];
                end
            end
          else
            begin
              for (forvar5109 = (1'h0); (forvar5109 < (2'h3)); forvar5109 = (forvar5109 + (1'h1)))
                begin
                  reg5110 <= $unsigned((^~((8'ha3) ?
                      (reg5057 ? (8'hb2) : reg4976) : $signed(reg4832))));
                  for (forvar5111 = (1'h0); (forvar5111 < (2'h2)); forvar5111 = (forvar5111 + (1'h1)))
                    begin
                      reg5112 <= reg4724[(4'h8):(3'h4)];
                      reg5113 <= reg4729[(1'h0):(1'h0)];
                      reg5114 <= (^~$signed({(~&reg5001)}));
                      reg5115 <= $signed(reg4656[(3'h5):(3'h5)]);
                    end
                  reg5116 <= reg4947;
                end
              if ((reg4867 > (-reg5084)))
                begin
                  for (forvar5117 = (1'h0); (forvar5117 < (2'h3)); forvar5117 = (forvar5117 + (1'h1)))
                    begin
                      reg5118 <= (8'h9d);
                      reg5119 <= (&{$unsigned((8'ha7))});
                      reg5120 <= {(+$signed($signed((8'ha6))))};
                      reg5121 <= (reg4751[(2'h3):(1'h0)] ~^ {(reg4692[(2'h2):(1'h0)] & (forvar4766 ?
                              reg4848 : (8'h9d)))});
                    end
                  if (reg4842)
                    begin
                      reg5122 <= ((((~&reg4951) ?
                                  (+(8'hab)) : (forvar4759 ?
                                      reg4956 : reg4931)) ?
                              (forvar4694 ?
                                  (forvar4918 * reg4721) : $signed((8'ha9))) : $signed((reg5070 ^~ reg4924))) ?
                          $signed((8'hab)) : ($unsigned(reg4867) || $unsigned($unsigned(forvar4848))));
                      reg5123 <= reg5085;
                      reg5124 <= $signed($signed(($signed(forvar5008) ?
                          reg4702[(1'h1):(1'h1)] : reg4675[(2'h3):(2'h3)])));
                      reg5125 <= {(-$unsigned($unsigned((8'ha9))))};
                    end
                  else
                    begin
                      reg5122 <= (8'hae);
                      reg5123 <= $unsigned({(8'ha6)});
                      reg5124 <= reg5120[(1'h1):(1'h0)];
                    end
                  for (forvar5126 = (1'h0); (forvar5126 < (1'h0)); forvar5126 = (forvar5126 + (1'h1)))
                    begin
                      reg5127 <= (&$signed((^~(forvar5117 ?
                          reg4982 : forvar4640))));
                      reg5128 <= (-(($unsigned(reg4713) ?
                              (reg4840 ^~ forvar4991) : {forvar5011}) ?
                          reg5017 : forvar5011));
                      reg5129 <= {((~^{forvar4858}) ?
                              $signed((|(8'ha5))) : $unsigned({reg4740}))};
                    end
                end
              else
                begin
                  reg5117 <= (|(&$unsigned(reg5000)));
                  reg5118 <= (((&reg5059) << ((reg4927 ?
                          forvar4996 : (8'hb3)) && $unsigned(reg4740))) ?
                      reg5039[(2'h2):(1'h1)] : $signed(($unsigned(reg4593) ?
                          (~reg4585) : (~^reg4944))));
                end
              if (((reg4750[(1'h0):(1'h0)] << $unsigned((+(8'hab)))) ?
                  ((^$signed(reg4837)) == forvar4801[(1'h1):(1'h0)]) : ((forvar5085 ?
                      (&forvar5062) : $unsigned(reg4954)) ~^ $unsigned(reg4623))))
                begin
                  if ((~|$unsigned($unsigned((reg4920 ?
                      reg4646 : forvar5126)))))
                    begin
                      reg5130 <= forvar4659[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg5130 <= {$signed(($unsigned(reg4853) | (reg5079 ?
                              forvar5091 : reg4732)))};
                    end
                end
              else
                begin
                  for (forvar5130 = (1'h0); (forvar5130 < (1'h0)); forvar5130 = (forvar5130 + (1'h1)))
                    begin
                      reg5131 <= {$unsigned(reg5013)};
                      reg5132 <= (+(((|forvar5001) ?
                              reg5024 : reg4928[(2'h3):(1'h0)]) ?
                          ((forvar4884 ?
                              reg5085 : reg4620) * reg4594[(4'ha):(3'h5)]) : $signed((~forvar4688))));
                      reg5133 <= ({reg4825} <= forvar5117);
                      reg5134 <= $unsigned((&$signed($signed(reg4828))));
                    end
                  for (forvar5135 = (1'h0); (forvar5135 < (1'h0)); forvar5135 = (forvar5135 + (1'h1)))
                    begin
                      reg5136 <= (~(&({reg4618} * (^reg4720))));
                      reg5137 <= (~^$unsigned(reg4761[(1'h0):(1'h0)]));
                    end
                end
              if ((|((((8'ha7) ~^ (8'hb8)) >= (reg4823 >= reg5041)) <<< ($unsigned(reg4871) != $signed(reg5014)))))
                begin
                  for (forvar5138 = (1'h0); (forvar5138 < (2'h3)); forvar5138 = (forvar5138 + (1'h1)))
                    begin
                      reg5139 <= reg5008[(3'h6):(3'h4)];
                    end
                  if ($unsigned($signed(((forvar4877 < reg5034) >> reg4869[(4'hd):(4'ha)]))))
                    begin
                      reg5140 <= $unsigned(reg4931);
                    end
                  else
                    begin
                      reg5140 <= $signed($signed(((!reg4733) + (forvar4578 ?
                          (8'hb9) : reg4808))));
                      reg5141 <= ({{{forvar5104}}} * (8'hb7));
                      reg5142 <= {$unsigned(($unsigned(reg4900) >>> {(8'had)}))};
                      reg5143 <= reg4949;
                    end
                  reg5144 <= (reg4955[(2'h2):(1'h1)] & $unsigned((~^forvar4584)));
                  reg5145 <= reg4861;
                end
              else
                begin
                  if (forvar5108[(2'h2):(1'h1)])
                    begin
                      reg5138 <= ((~((~forvar5083) + (~^reg4606))) ?
                          (reg4707[(4'hd):(4'h8)] <<< ($signed(forvar5053) ?
                              {forvar4581} : {reg4797})) : ($signed($signed(reg4842)) ?
                              reg4954[(3'h6):(1'h1)] : $unsigned((forvar5098 ?
                                  reg4967 : forvar5083))));
                      reg5139 <= (($unsigned((|reg4677)) ?
                          (reg4614[(1'h0):(1'h0)] && reg4609) : (+$signed(forvar4824))) < $signed((forvar5093[(2'h3):(1'h0)] ?
                          reg4964 : reg4965)));
                    end
                  else
                    begin
                      reg5138 <= ($unsigned(forvar4876[(4'ha):(3'h5)]) | reg4589);
                      reg5139 <= $unsigned(($signed($signed(forvar4753)) ?
                          $signed(forvar4733) : $signed((reg5048 ?
                              reg4864 : reg4847))));
                      reg5140 <= $signed(((8'haf) ?
                          $unsigned($unsigned((8'hba))) : ($signed(reg4708) & (reg4855 ?
                              wire4576 : reg4837))));
                      reg5141 <= $signed($signed(((forvar4806 >= forvar4663) ?
                          reg4636 : (forvar4785 ^~ (8'haf)))));
                    end
                  reg5142 <= (~$signed(reg5045));
                  for (forvar5143 = (1'h0); (forvar5143 < (2'h2)); forvar5143 = (forvar5143 + (1'h1)))
                    begin
                      reg5144 <= ($signed(reg4783[(2'h2):(1'h0)]) << $signed(reg4600[(2'h3):(1'h1)]));
                      reg5145 <= (~|{reg4723});
                      reg5146 <= ((($signed(forvar5068) ?
                          (!(8'h9d)) : forvar5083) ^ reg4909[(2'h3):(2'h2)]) >> (forvar4840[(4'hb):(4'h8)] ?
                          ($unsigned(reg4871) - (reg4916 || reg5034)) : reg4950));
                    end
                end
            end
        end
      reg5147 <= reg4774;
      if (($signed((^~((8'hab) << forvar4910))) ?
          ($unsigned((reg4581 ? (8'h9e) : reg4807)) ?
              reg4770 : $unsigned((8'hae))) : $signed(($signed(forvar4980) ?
              $signed(reg4591) : (+reg4936)))))
        begin
          reg5148 <= $signed(((+(forvar5064 * reg5058)) << reg4831[(2'h2):(1'h0)]));
          if ($signed(($unsigned(reg4951) ? $signed(reg4995) : reg4791)))
            begin
              reg5149 <= $signed((8'ha7));
              for (forvar5150 = (1'h0); (forvar5150 < (2'h2)); forvar5150 = (forvar5150 + (1'h1)))
                begin
                  if ({(reg4892 >>> $signed(reg4811[(4'h8):(3'h4)]))})
                    begin
                      reg5151 <= $unsigned($unsigned({(reg5026 ?
                              reg4726 : (8'ha2))}));
                      reg5152 <= $unsigned(reg4677[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg5151 <= forvar4689[(1'h0):(1'h0)];
                    end
                  if (forvar4815)
                    begin
                      reg5153 <= (+(^reg4635[(4'ha):(3'h5)]));
                    end
                  else
                    begin
                      reg5153 <= ((~^$signed((reg4770 == reg4789))) == $signed((|$unsigned(forvar4581))));
                    end
                end
            end
          else
            begin
              for (forvar5149 = (1'h0); (forvar5149 < (2'h2)); forvar5149 = (forvar5149 + (1'h1)))
                begin
                  if ($unsigned($signed((-$signed(reg4881)))))
                    begin
                      reg5150 <= reg4703[(1'h1):(1'h1)];
                      reg5151 <= forvar5020[(1'h0):(1'h0)];
                      reg5152 <= ({reg4842} ?
                          (reg5073 != ((reg4766 * reg4723) <<< (^~reg5143))) : reg5144[(4'he):(4'hb)]);
                    end
                  else
                    begin
                      reg5150 <= ({$signed(reg4667[(3'h4):(3'h4)])} >>> $unsigned($unsigned(((8'hb6) ?
                          reg4834 : forvar4913))));
                      reg5151 <= (forvar4777 <= $signed((^(reg4689 ^~ reg5013))));
                    end
                  if ($signed(reg5036[(3'h5):(1'h0)]))
                    begin
                      reg5153 <= $signed(((8'ha4) || (forvar4890[(3'h4):(2'h3)] || (!reg4748))));
                    end
                  else
                    begin
                      reg5153 <= $unsigned((^~forvar5149[(4'h8):(2'h2)]));
                      reg5154 <= (^~$unsigned(reg4883[(2'h2):(1'h0)]));
                      reg5155 <= reg4678[(2'h3):(2'h3)];
                      reg5156 <= $signed(((!(reg4945 ~^ wire4576)) ^ reg5138[(4'hc):(4'ha)]));
                    end
                  for (forvar5157 = (1'h0); (forvar5157 < (1'h1)); forvar5157 = (forvar5157 + (1'h1)))
                    begin
                      reg5158 <= (reg4598[(3'h4):(2'h3)] >= ({((8'hb3) & reg4608)} ?
                          (~^$signed(reg5015)) : {$signed(forvar5111)}));
                      reg5159 <= $unsigned((-(((8'hb8) && (8'hae)) ?
                          (reg4919 && reg5021) : reg4688)));
                      reg5160 <= $signed({(forvar4694[(4'h8):(3'h7)] ?
                              forvar4969 : $unsigned(reg4869))});
                      reg5161 <= $signed($unsigned(($signed(forvar4909) ?
                          (reg5011 && reg4867) : $unsigned(forvar4786))));
                    end
                  for (forvar5162 = (1'h0); (forvar5162 < (2'h3)); forvar5162 = (forvar5162 + (1'h1)))
                    begin
                      reg5163 <= ((($signed(reg4601) ?
                          forvar5093[(1'h1):(1'h1)] : (reg4878 ?
                              reg4938 : reg4841)) != (^~reg4636)) * ({$signed(reg4924)} ?
                          forvar4849 : reg4859));
                      reg5164 <= reg5029[(1'h0):(1'h0)];
                    end
                end
            end
          for (forvar5165 = (1'h0); (forvar5165 < (1'h1)); forvar5165 = (forvar5165 + (1'h1)))
            begin
              for (forvar5166 = (1'h0); (forvar5166 < (2'h3)); forvar5166 = (forvar5166 + (1'h1)))
                begin
                  if ((~|reg4723[(3'h6):(3'h6)]))
                    begin
                      reg5167 <= $unsigned((^~(reg4593[(3'h4):(1'h1)] + {reg4609})));
                      reg5168 <= reg5046[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg5167 <= (-$signed({((8'haa) ? reg4638 : (8'ha1))}));
                      reg5168 <= (forvar5009 >> $unsigned(((reg5057 ^~ reg4684) ?
                          (reg4693 ^~ forvar4609) : $signed((8'ha0)))));
                      reg5169 <= ({reg4912} ~^ forvar4689[(1'h1):(1'h1)]);
                    end
                end
              for (forvar5170 = (1'h0); (forvar5170 < (1'h1)); forvar5170 = (forvar5170 + (1'h1)))
                begin
                  for (forvar5171 = (1'h0); (forvar5171 < (2'h2)); forvar5171 = (forvar5171 + (1'h1)))
                    begin
                      reg5172 <= reg4599[(3'h6):(2'h3)];
                      reg5173 <= $signed(reg5108[(2'h2):(1'h1)]);
                      reg5174 <= (8'hb2);
                    end
                  for (forvar5175 = (1'h0); (forvar5175 < (2'h3)); forvar5175 = (forvar5175 + (1'h1)))
                    begin
                      reg5176 <= {$unsigned($unsigned($unsigned(forvar4958)))};
                    end
                  for (forvar5177 = (1'h0); (forvar5177 < (2'h2)); forvar5177 = (forvar5177 + (1'h1)))
                    begin
                      reg5178 <= reg4715;
                      reg5179 <= $unsigned($unsigned(reg4726[(2'h3):(1'h0)]));
                      reg5180 <= $signed(reg4928[(3'h5):(1'h1)]);
                    end
                  if ((reg4928 ?
                      {$signed({reg4736})} : wire4940[(3'h4):(2'h2)]))
                    begin
                      reg5181 <= (~&reg4954[(3'h7):(3'h6)]);
                    end
                  else
                    begin
                      reg5181 <= $unsigned((reg4731 ~^ $unsigned((forvar4977 ?
                          forvar4915 : forvar4996))));
                      reg5182 <= $unsigned(reg4614[(3'h4):(2'h2)]);
                      reg5183 <= (forvar4785[(4'hb):(3'h6)] ?
                          $signed(reg4871[(2'h2):(1'h0)]) : ($signed((8'hb2)) ?
                              ((8'h9d) >>> {forvar4944}) : {(forvar4717 ~^ reg5113)}));
                      reg5184 <= (~&$signed(($unsigned(forvar4759) <= (~^reg4612))));
                    end
                end
              if ((($unsigned({forvar4967}) | forvar5084[(2'h2):(1'h0)]) >= $unsigned(forvar5084[(1'h0):(1'h0)])))
                begin
                  for (forvar5185 = (1'h0); (forvar5185 < (1'h0)); forvar5185 = (forvar5185 + (1'h1)))
                    begin
                      reg5186 <= $signed((($unsigned(reg4713) <= $unsigned(reg5047)) ?
                          $signed(reg4754[(3'h7):(2'h3)]) : $unsigned(reg4732[(1'h0):(1'h0)])));
                    end
                  for (forvar5187 = (1'h0); (forvar5187 < (1'h1)); forvar5187 = (forvar5187 + (1'h1)))
                    begin
                      reg5188 <= ({$signed((reg5161 ? forvar4915 : (8'hb2)))} ?
                          $unsigned($signed((reg4994 ?
                              reg4666 : reg4921))) : $signed($signed(((8'ha8) | reg4854))));
                    end
                  for (forvar5189 = (1'h0); (forvar5189 < (1'h0)); forvar5189 = (forvar5189 + (1'h1)))
                    begin
                      reg5190 <= (!(-($unsigned((8'hb8)) ?
                          (^~reg4840) : $unsigned((8'ha4)))));
                      reg5191 <= $unsigned($unsigned(forvar4848[(2'h2):(2'h2)]));
                      reg5192 <= reg5149;
                    end
                end
              else
                begin
                  if (((reg4624 && (^reg4729[(1'h0):(1'h0)])) <= ($unsigned($signed(forvar5157)) <<< $signed($unsigned(reg5093)))))
                    begin
                      reg5185 <= $unsigned(({reg4713} ~^ reg4863[(4'hb):(1'h1)]));
                    end
                  else
                    begin
                      reg5185 <= {reg4753};
                    end
                  for (forvar5186 = (1'h0); (forvar5186 < (1'h0)); forvar5186 = (forvar5186 + (1'h1)))
                    begin
                      reg5187 <= {({(~^wire4799)} ?
                              $unsigned($unsigned(reg4679)) : (^((8'ha3) == reg5097)))};
                    end
                  if ({($unsigned({reg5071}) >> ((forvar4909 <= reg4639) ~^ $signed((8'ha8))))})
                    begin
                      reg5188 <= reg4701;
                      reg5189 <= $unsigned($unsigned(reg4999[(3'h4):(2'h3)]));
                      reg5190 <= ((reg4842 & ($unsigned((8'h9e)) - reg5158[(2'h2):(2'h2)])) * {$signed({reg4680})});
                    end
                  else
                    begin
                      reg5188 <= (~$signed(((^reg4860) ?
                          (reg5044 ? reg5082 : forvar4884) : (^(8'hac)))));
                    end
                  if (reg4614)
                    begin
                      reg5191 <= (((reg4755[(1'h1):(1'h1)] ?
                              $unsigned((8'h9f)) : (forvar5165 ?
                                  reg5053 : reg5178)) <<< (!(~(8'h9d)))) ?
                          {(forvar4944 ?
                                  (forvar4957 ?
                                      reg5010 : reg5070) : $signed(reg4912))} : {{(reg4886 ?
                                      forvar4802 : reg4848)}});
                      reg5192 <= {({$signed(forvar4749)} ?
                              ($unsigned(forvar5008) || (^(8'hba))) : ((^~reg4677) ?
                                  $unsigned(reg4965) : (^reg4920)))};
                      reg5193 <= $unsigned($signed(($signed(reg4990) ?
                          forvar4579[(3'h4):(2'h2)] : reg4679)));
                      reg5194 <= $unsigned($signed((8'hb1)));
                    end
                  else
                    begin
                      reg5191 <= ($signed(reg5172) ?
                          (~$signed(forvar4829)) : (^~reg5185[(2'h2):(1'h1)]));
                      reg5192 <= forvar5036[(2'h2):(1'h1)];
                    end
                end
            end
        end
      else
        begin
          for (forvar5148 = (1'h0); (forvar5148 < (2'h2)); forvar5148 = (forvar5148 + (1'h1)))
            begin
              reg5149 <= (^~(~|(reg4728[(3'h6):(1'h0)] ~^ reg4610)));
              if ($signed($unsigned((reg5038[(4'h8):(2'h2)] ?
                  (reg4867 ? reg4774 : reg5118) : (-reg4606)))))
                begin
                  if ($signed(reg4938))
                    begin
                      reg5150 <= (8'h9c);
                      reg5151 <= $signed(forvar4624);
                      reg5152 <= {(forvar4737[(2'h3):(1'h1)] <= ((reg4780 ?
                              reg5000 : forvar4748) && reg5120[(1'h1):(1'h0)]))};
                    end
                  else
                    begin
                      reg5150 <= (!reg4889[(2'h2):(1'h0)]);
                      reg5151 <= (+(~^$signed(reg4645)));
                      reg5152 <= (((-reg5086[(1'h0):(1'h0)]) + reg4660) ?
                          (reg4778[(2'h3):(2'h2)] ?
                              $unsigned($signed(reg4720)) : reg4910) : (($unsigned(reg4754) == reg4845[(1'h1):(1'h0)]) >>> forvar4965[(1'h0):(1'h0)]));
                      reg5153 <= (reg4825 ?
                          {({reg4715} ^ {forvar4694})} : {$signed($unsigned((8'hb1)))});
                    end
                end
              else
                begin
                  if (reg4742[(1'h1):(1'h0)])
                    begin
                      reg5150 <= (reg4687[(4'hb):(3'h7)] - $signed(({reg4924} > forvar4643[(1'h1):(1'h0)])));
                      reg5151 <= reg4983[(2'h3):(2'h2)];
                      reg5152 <= (8'ha7);
                      reg5153 <= $signed((((forvar5102 ?
                          reg5117 : reg4903) << {(8'ha0)}) >> ($unsigned((8'ha0)) & (reg4716 ?
                          forvar5039 : forvar4962))));
                    end
                  else
                    begin
                      reg5150 <= reg4660[(2'h2):(1'h0)];
                    end
                end
            end
        end
    end
  assign wire5195 = ({(reg4596[(3'h5):(1'h1)] ?
                            {(8'h9d)} : ((8'ha8) ?
                                forvar4969 : forvar4931))} ~^ forvar5049);
  assign wire5196 = (reg4676 ?
                        ((^~reg4686[(3'h5):(3'h4)]) != (8'ha5)) : {(^~$signed((8'haa)))});
  assign wire5197 = $unsigned({((~&(8'ha7)) * (8'hb4))});
  always
    @(posedge clk) begin
      for (forvar5198 = (1'h0); (forvar5198 < (2'h2)); forvar5198 = (forvar5198 + (1'h1)))
        begin
          if (((~^(|((8'hb2) == forvar4773))) ~^ ((reg4996[(1'h1):(1'h0)] + (~(8'h9f))) < forvar5170)))
            begin
              if (forvar4813[(4'h8):(1'h0)])
                begin
                  for (forvar5199 = (1'h0); (forvar5199 < (2'h2)); forvar5199 = (forvar5199 + (1'h1)))
                    begin
                      reg5200 <= forvar5062[(1'h1):(1'h0)];
                    end
                  reg5201 <= $unsigned(reg4579[(2'h2):(1'h1)]);
                  reg5202 <= reg4990[(2'h3):(2'h3)];
                end
              else
                begin
                  reg5199 <= {((&$signed(reg4736)) + ((forvar4780 ?
                          forvar5082 : reg5013) || $signed((8'ha4))))};
                  if (((~|$signed((reg4782 <<< (8'ha4)))) == $unsigned($signed((forvar5019 ^ reg4641)))))
                    begin
                      reg5200 <= reg4850[(1'h1):(1'h0)];
                      reg5201 <= reg4953[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg5200 <= ({$unsigned($signed(reg4715))} ?
                          {($unsigned(reg4805) <= reg4867)} : {$unsigned($signed(reg4774))});
                      reg5201 <= forvar4749[(2'h3):(2'h3)];
                    end
                  reg5202 <= forvar4909;
                end
              if (({(^(&reg4605))} > (-reg4639[(2'h3):(2'h2)])))
                begin
                  if ((+forvar5108[(3'h5):(3'h4)]))
                    begin
                      reg5203 <= $signed((^reg4787));
                      reg5204 <= reg4763;
                      reg5205 <= $unsigned((forvar4674[(3'h5):(1'h1)] <<< {{forvar4777}}));
                    end
                  else
                    begin
                      reg5203 <= $signed(reg4701);
                    end
                  for (forvar5206 = (1'h0); (forvar5206 < (1'h0)); forvar5206 = (forvar5206 + (1'h1)))
                    begin
                      reg5207 <= $unsigned($unsigned(((reg4865 != reg4908) | $signed(reg5181))));
                    end
                  for (forvar5208 = (1'h0); (forvar5208 < (2'h3)); forvar5208 = (forvar5208 + (1'h1)))
                    begin
                      reg5209 <= wire5195[(3'h5):(1'h1)];
                      reg5210 <= $unsigned(reg4832[(2'h2):(1'h1)]);
                      reg5211 <= reg5163[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  if (reg5020)
                    begin
                      reg5203 <= reg5125[(2'h2):(1'h1)];
                      reg5204 <= $signed($unsigned((forvar4659[(3'h4):(2'h3)] <<< ((8'ha7) | reg5082))));
                      reg5205 <= $unsigned({{$signed(reg4939)}});
                      reg5206 <= (^forvar4879);
                    end
                  else
                    begin
                      reg5203 <= $unsigned((({forvar5104} && forvar4999[(4'ha):(4'h9)]) ?
                          forvar4952[(1'h0):(1'h0)] : (~{reg4897})));
                    end
                  if (forvar5162)
                    begin
                      reg5207 <= $signed(forvar4581[(1'h0):(1'h0)]);
                      reg5208 <= (8'hb1);
                      reg5209 <= $unsigned({((&reg4579) ?
                              $signed(reg5047) : forvar4858[(3'h4):(2'h2)])});
                    end
                  else
                    begin
                      reg5207 <= (-($signed($unsigned(reg5038)) & $unsigned(forvar4610[(3'h6):(3'h6)])));
                    end
                  if (reg4703[(1'h1):(1'h1)])
                    begin
                      reg5210 <= (reg5138[(4'ha):(4'h8)] ~^ reg4794);
                      reg5211 <= ((!reg5096) ?
                          (-(~&(forvar4717 | reg4954))) : $signed((~&{reg4619})));
                      reg5212 <= (&{(((8'ha7) > reg4683) ?
                              forvar5051 : $unsigned(reg4643))});
                    end
                  else
                    begin
                      reg5210 <= $signed({{(~(8'ha4))}});
                      reg5211 <= reg5100;
                      reg5212 <= reg4722[(1'h0):(1'h0)];
                    end
                  if (($unsigned((8'ha8)) > (^(!((8'ha2) ?
                      forvar5043 : (8'hac))))))
                    begin
                      reg5213 <= {(reg5167[(1'h0):(1'h0)] ?
                              forvar5114 : $unsigned($unsigned(reg4901)))};
                      reg5214 <= (reg4846 == (8'hb2));
                      reg5215 <= {$signed((+((8'hba) && reg4749)))};
                      reg5216 <= $signed((forvar5111 ?
                          $signed((reg4608 < reg4946)) : $unsigned(((8'hb7) ?
                              forvar5109 : reg5097))));
                    end
                  else
                    begin
                      reg5213 <= $signed($signed(((^reg4598) == reg5006)));
                      reg5214 <= forvar5084[(2'h2):(2'h2)];
                    end
                end
              for (forvar5217 = (1'h0); (forvar5217 < (2'h2)); forvar5217 = (forvar5217 + (1'h1)))
                begin
                  for (forvar5218 = (1'h0); (forvar5218 < (1'h1)); forvar5218 = (forvar5218 + (1'h1)))
                    begin
                      reg5219 <= $unsigned($unsigned($signed(reg4628[(2'h2):(2'h2)])));
                    end
                  if (reg4910[(1'h0):(1'h0)])
                    begin
                      reg5220 <= {(((reg4629 ? forvar4758 : reg4849) ?
                                  $signed(reg5073) : (^~reg4928)) ?
                              reg4770 : (reg4969[(2'h3):(2'h3)] - reg4791))};
                      reg5221 <= (~forvar4745);
                      reg5222 <= (~|(~|($signed((8'h9f)) ?
                          (8'hb7) : (reg4797 | forvar4850))));
                      reg5223 <= (($signed($signed(forvar4773)) ?
                              forvar4673[(3'h5):(3'h5)] : $unsigned(reg5012)) ?
                          reg4598[(2'h2):(1'h1)] : reg4857);
                    end
                  else
                    begin
                      reg5220 <= (-$signed(reg4792));
                      reg5221 <= $unsigned(reg4701);
                      reg5222 <= $unsigned(forvar5020);
                      reg5223 <= reg4758;
                    end
                  for (forvar5224 = (1'h0); (forvar5224 < (2'h2)); forvar5224 = (forvar5224 + (1'h1)))
                    begin
                      reg5225 <= $unsigned($signed(reg4893[(1'h0):(1'h0)]));
                    end
                end
              reg5226 <= $unsigned(reg5179);
            end
          else
            begin
              for (forvar5199 = (1'h0); (forvar5199 < (2'h2)); forvar5199 = (forvar5199 + (1'h1)))
                begin
                  for (forvar5200 = (1'h0); (forvar5200 < (2'h2)); forvar5200 = (forvar5200 + (1'h1)))
                    begin
                      reg5201 <= ($signed(((!forvar5108) ~^ forvar4933[(3'h5):(3'h4)])) & $signed((8'hb1)));
                    end
                  reg5202 <= $signed(reg4579[(2'h3):(2'h3)]);
                  reg5203 <= {forvar4991};
                  if ((~|{forvar4785[(1'h1):(1'h0)]}))
                    begin
                      reg5204 <= (~&(({reg5008} ?
                              reg4952 : $unsigned((8'haf))) ?
                          $unsigned(reg4651[(4'ha):(4'h8)]) : (reg5044 ^~ (reg5005 && reg5037))));
                      reg5205 <= forvar4998;
                    end
                  else
                    begin
                      reg5204 <= ((~^({reg5199} ?
                          (+reg4736) : $unsigned(reg5127))) & (reg4820[(3'h7):(2'h2)] ?
                          (|(~forvar4789)) : $unsigned((wire5196 ?
                              reg4635 : reg4789))));
                      reg5205 <= $signed(reg5071[(1'h1):(1'h1)]);
                    end
                end
            end
          reg5227 <= $signed(reg5143);
        end
      if ((reg5183[(4'hb):(4'ha)] ? forvar5109 : (8'hb4)))
        begin
          if (forvar4826)
            begin
              for (forvar5228 = (1'h0); (forvar5228 < (1'h1)); forvar5228 = (forvar5228 + (1'h1)))
                begin
                  reg5229 <= ($unsigned($signed(reg5137)) ?
                      $unsigned(($signed(reg4860) >= $unsigned(reg4601))) : (!((reg4993 ~^ reg5096) - (~^(8'hb1)))));
                  if ($signed(forvar4676))
                    begin
                      reg5230 <= (reg4691[(1'h0):(1'h0)] ?
                          reg5010[(1'h0):(1'h0)] : ((forvar4839 ?
                                  $unsigned(reg5129) : reg5086[(3'h6):(1'h1)]) ?
                              {(forvar4588 ?
                                      reg4816 : reg5100)} : ((forvar4975 ?
                                      reg4907 : reg5172) ?
                                  $signed(reg5057) : forvar4725[(2'h2):(1'h1)])));
                      reg5231 <= (&reg5116);
                      reg5232 <= $signed($signed($unsigned(reg5079)));
                      reg5233 <= $signed((forvar4999[(4'h9):(1'h1)] && (^$unsigned(reg4750))));
                    end
                  else
                    begin
                      reg5230 <= $signed(($unsigned($unsigned(reg4695)) ?
                          ((~^reg4904) ?
                              (~&forvar4579) : $signed((8'hac))) : $unsigned($signed((8'ha9)))));
                      reg5231 <= $signed($signed(((reg5085 ?
                          reg4803 : reg4662) ^ forvar5051)));
                    end
                  for (forvar5234 = (1'h0); (forvar5234 < (2'h3)); forvar5234 = (forvar5234 + (1'h1)))
                    begin
                      reg5235 <= $unsigned((8'hb6));
                      reg5236 <= ($unsigned((reg5013[(2'h2):(1'h1)] | forvar4909[(3'h5):(3'h5)])) < ((~|forvar5068) ?
                          {$unsigned(reg4580)} : reg4852[(4'hd):(4'hd)]));
                      reg5237 <= (~|(!reg4882));
                    end
                  for (forvar5238 = (1'h0); (forvar5238 < (1'h1)); forvar5238 = (forvar5238 + (1'h1)))
                    begin
                      reg5239 <= $unsigned(reg4703[(2'h2):(2'h2)]);
                      reg5240 <= ({((reg4978 + reg5188) ?
                              $signed(forvar4598) : forvar4826[(2'h2):(2'h2)])} >> wire5195);
                      reg5241 <= $unsigned($unsigned($signed((forvar4759 ?
                          (8'haf) : reg4893))));
                      reg5242 <= (~&{{((8'ha2) ? (8'h9d) : (8'hba))}});
                    end
                end
            end
          else
            begin
              if (forvar4970)
                begin
                  for (forvar5228 = (1'h0); (forvar5228 < (2'h3)); forvar5228 = (forvar5228 + (1'h1)))
                    begin
                      reg5229 <= (8'ha9);
                      reg5230 <= reg5085[(2'h2):(1'h1)];
                    end
                  if ((^~$signed((8'hb7))))
                    begin
                      reg5231 <= $signed($signed($unsigned(reg4937)));
                      reg5232 <= (^~((^~$signed(reg5019)) ?
                          reg4885 : {(reg4805 >= forvar4608)}));
                      reg5233 <= $signed(($unsigned($unsigned(forvar5008)) ?
                          ((reg5010 < forvar5106) ?
                              (forvar4755 >= reg4611) : (reg5095 > reg5153)) : ((reg5230 >= (8'hb7)) >> (reg5011 > reg4850))));
                    end
                  else
                    begin
                      reg5231 <= $unsigned(($signed(reg5006) ?
                          $signed((forvar5186 ?
                              reg4966 : reg4627)) : $unsigned(reg5233[(1'h0):(1'h0)])));
                      reg5232 <= $unsigned({$signed(((8'hae) ?
                              forvar4624 : reg4618))});
                      reg5233 <= (forvar4795[(3'h5):(3'h5)] ?
                          reg5043 : reg5057);
                      reg5234 <= ($unsigned((8'hb2)) + forvar5020[(3'h4):(3'h4)]);
                    end
                end
              else
                begin
                  if (forvar5162[(1'h0):(1'h0)])
                    begin
                      reg5228 <= {($signed($signed(forvar4674)) && ((&forvar4998) + (^~reg4684)))};
                      reg5229 <= ((+{(^reg5007)}) ?
                          (($unsigned((8'ha0)) ?
                                  $unsigned(reg4986) : $unsigned(forvar4768)) ?
                              (8'ha6) : $unsigned($unsigned((8'ha9)))) : $signed(((+reg4747) ?
                              reg4893 : {reg5091})));
                      reg5230 <= $unsigned(reg4721);
                    end
                  else
                    begin
                      reg5228 <= (forvar5171 * $signed(((~&reg4868) != (reg5045 ?
                          reg5027 : reg4825))));
                    end
                end
            end
          if (($signed((+(^reg4895))) >>> {(forvar4611 ?
                  (8'ha4) : reg5117[(2'h3):(2'h2)])}))
            begin
              reg5243 <= (($unsigned((~|reg4935)) ?
                      $unsigned({reg5220}) : reg4868) ?
                  reg4746[(1'h1):(1'h0)] : $signed(((8'hab) ?
                      (^~reg5055) : reg4611)));
              reg5244 <= ($unsigned(($unsigned(reg4911) ?
                  (reg4902 >= forvar5138) : forvar5208[(2'h3):(2'h3)])) <<< ($unsigned($signed(reg4664)) >>> reg5017));
              if ($unsigned(($unsigned($unsigned(reg4770)) ?
                  $signed($signed(reg4738)) : reg5169[(2'h3):(1'h1)])))
                begin
                  reg5245 <= $unsigned((reg4929 == $unsigned(forvar4733)));
                end
              else
                begin
                  for (forvar5245 = (1'h0); (forvar5245 < (1'h1)); forvar5245 = (forvar5245 + (1'h1)))
                    begin
                      reg5246 <= forvar4962[(4'h8):(3'h7)];
                      reg5247 <= (reg5107 && ({(8'hac)} ~^ forvar5102[(1'h1):(1'h1)]));
                    end
                  for (forvar5248 = (1'h0); (forvar5248 < (1'h0)); forvar5248 = (forvar5248 + (1'h1)))
                    begin
                      reg5249 <= $signed($signed($unsigned((8'hb9))));
                      reg5250 <= forvar5228;
                      reg5251 <= $signed(($unsigned(reg4594[(3'h5):(1'h0)]) ?
                          ((8'hab) | (reg4609 ?
                              reg5131 : reg4751)) : ((~reg5089) ?
                              (reg4878 > reg4805) : $unsigned(reg4589))));
                    end
                  reg5252 <= reg5012[(1'h1):(1'h0)];
                  if (($unsigned(forvar4731[(1'h1):(1'h1)]) + reg5074[(3'h4):(1'h1)]))
                    begin
                      reg5253 <= (^~((reg4810[(1'h1):(1'h0)] ?
                          $unsigned(forvar5170) : $signed(reg5183)) <= (8'ha3)));
                      reg5254 <= reg5138;
                    end
                  else
                    begin
                      reg5253 <= ($signed(reg4955[(3'h7):(2'h2)]) ?
                          reg4927 : (forvar4588[(4'h8):(3'h6)] || ((reg4679 ?
                              reg4740 : reg5057) | (reg5011 ?
                              reg4911 : reg4883))));
                      reg5254 <= ($signed(reg4732) << ((~^(+reg5042)) ?
                          ((reg5052 ?
                              reg5169 : reg4768) * $unsigned(forvar4848)) : $unsigned((|forvar5075))));
                    end
                end
            end
          else
            begin
              if (((~&$unsigned($unsigned((8'h9f)))) ?
                  $unsigned($unsigned((reg4779 ?
                      forvar5218 : (8'hac)))) : (^~forvar5238[(2'h2):(2'h2)])))
                begin
                  for (forvar5243 = (1'h0); (forvar5243 < (2'h2)); forvar5243 = (forvar5243 + (1'h1)))
                    begin
                      reg5244 <= $signed(({reg5251} || reg5146));
                      reg5245 <= ($signed($signed((reg4878 ?
                              reg5053 : reg5110))) ?
                          $signed((^(reg4830 ?
                              forvar4577 : reg4756))) : ((-$unsigned(reg4741)) ^ ($unsigned(forvar4768) ?
                              (forvar5171 ?
                                  reg4715 : reg4680) : $unsigned(reg4604))));
                      reg5246 <= (((((8'hb1) ?
                          forvar5218 : (8'hba)) && {reg4990}) <<< {$unsigned(reg5129)}) <= {$unsigned((8'had))});
                    end
                  for (forvar5247 = (1'h0); (forvar5247 < (2'h2)); forvar5247 = (forvar5247 + (1'h1)))
                    begin
                      reg5248 <= ({($signed(reg4928) & forvar5189[(3'h7):(3'h5)])} ?
                          forvar4580 : reg4800);
                      reg5249 <= (reg4999[(2'h2):(1'h1)] ?
                          ({reg4780} ?
                              forvar4758[(1'h0):(1'h0)] : ($signed(reg5071) >= $unsigned((8'hb1)))) : (((^~forvar4929) ?
                              (reg4805 ?
                                  reg4628 : reg4768) : reg4767) == reg5143[(3'h6):(3'h6)]));
                      reg5250 <= reg4666[(2'h2):(1'h1)];
                      reg5251 <= $unsigned($signed((!forvar4579[(1'h0):(1'h0)])));
                    end
                  for (forvar5252 = (1'h0); (forvar5252 < (1'h1)); forvar5252 = (forvar5252 + (1'h1)))
                    begin
                      reg5253 <= $signed(($signed({reg5128}) >> $signed((8'ha2))));
                      reg5254 <= $signed((!({reg5032} & (reg5247 | reg5128))));
                      reg5255 <= ($signed($signed((forvar4996 | reg5145))) ?
                          $signed(reg4861) : (&forvar5171[(1'h1):(1'h1)]));
                      reg5256 <= ($signed($unsigned((8'h9c))) ?
                          $unsigned({{forvar4594}}) : (($signed(reg4998) >> (~|reg4595)) <= $signed(reg4835)));
                    end
                end
              else
                begin
                  for (forvar5243 = (1'h0); (forvar5243 < (2'h3)); forvar5243 = (forvar5243 + (1'h1)))
                    begin
                      reg5244 <= ((~^$unsigned(forvar5162[(1'h1):(1'h0)])) ?
                          reg4742[(4'hf):(3'h6)] : ($unsigned(reg5219) ?
                              reg5125 : $unsigned(forvar5029)));
                    end
                  if ($unsigned(reg4621[(2'h3):(1'h1)]))
                    begin
                      reg5245 <= (reg4749 ?
                          {$signed(reg5116[(3'h4):(3'h4)])} : ($unsigned($signed(forvar4616)) << forvar5224));
                      reg5246 <= ({$signed($unsigned(reg4793))} ?
                          (((forvar4766 ? reg5240 : reg4930) ?
                                  forvar5019 : forvar5002) ?
                              reg4755 : reg4761) : $signed($signed((8'had))));
                      reg5247 <= $signed($signed(reg4639));
                    end
                  else
                    begin
                      reg5245 <= $signed((reg4677 ?
                          $signed($signed(reg4847)) : forvar4770[(3'h6):(1'h1)]));
                      reg5246 <= (reg4740[(1'h1):(1'h1)] == (!reg4582[(1'h1):(1'h0)]));
                      reg5247 <= ((reg5045[(1'h1):(1'h0)] ?
                          forvar4909 : (reg4599[(1'h1):(1'h1)] >= reg4837[(3'h4):(1'h1)])) * $signed(forvar4738));
                    end
                end
              for (forvar5257 = (1'h0); (forvar5257 < (2'h3)); forvar5257 = (forvar5257 + (1'h1)))
                begin
                  if (({($unsigned((8'ha4)) ? reg4792 : reg5136)} | {reg5079}))
                    begin
                      reg5258 <= ({$signed((8'hb2))} ?
                          $unsigned($signed((reg4929 ?
                              forvar4610 : reg5252))) : (($signed(reg4612) & {forvar4995}) ?
                              wire5197[(4'h8):(3'h7)] : (8'h9f)));
                      reg5259 <= reg4766;
                    end
                  else
                    begin
                      reg5258 <= $signed((((reg4724 && forvar4801) == forvar5091) >= ((reg4872 ?
                          reg4822 : reg5037) <= (reg5207 & (8'hb2)))));
                      reg5259 <= $signed(($unsigned($unsigned(reg5207)) ?
                          (~|$unsigned(reg4954)) : $unsigned((8'ha7))));
                    end
                  reg5260 <= $signed($unsigned($unsigned($unsigned(reg4803))));
                  for (forvar5261 = (1'h0); (forvar5261 < (1'h0)); forvar5261 = (forvar5261 + (1'h1)))
                    begin
                      reg5262 <= ((+(((8'hb0) ? reg5259 : reg4638) ?
                              forvar4674[(3'h5):(1'h1)] : $unsigned(reg4846))) ?
                          (|(reg4583 ?
                              (reg5143 ?
                                  (8'hb0) : forvar5029) : (reg4789 > reg5235))) : $signed(reg4596[(1'h0):(1'h0)]));
                      reg5263 <= {((8'h9f) ?
                              $signed((reg5211 ?
                                  wire4576 : reg4959)) : $signed((-reg5117)))};
                      reg5264 <= reg4704[(4'hc):(3'h6)];
                      reg5265 <= $signed((reg5118[(1'h1):(1'h1)] ?
                          (-{reg5234}) : (-forvar5217[(1'h1):(1'h0)])));
                    end
                  for (forvar5266 = (1'h0); (forvar5266 < (2'h2)); forvar5266 = (forvar5266 + (1'h1)))
                    begin
                      reg5267 <= reg4789[(1'h0):(1'h0)];
                      reg5268 <= ((-(~|forvar5091)) & (+{{reg5263}}));
                    end
                end
            end
          reg5269 <= forvar4877;
        end
      else
        begin
          for (forvar5228 = (1'h0); (forvar5228 < (2'h2)); forvar5228 = (forvar5228 + (1'h1)))
            begin
              for (forvar5229 = (1'h0); (forvar5229 < (1'h0)); forvar5229 = (forvar5229 + (1'h1)))
                begin
                  if ({reg4679[(3'h4):(1'h1)]})
                    begin
                      reg5230 <= forvar5064;
                    end
                  else
                    begin
                      reg5230 <= {(((forvar4851 & reg5108) || {forvar5108}) ?
                              ((reg4719 != forvar5247) ?
                                  (~^(8'ha4)) : (reg4667 ?
                                      reg4780 : reg4679)) : (|(forvar4694 ?
                                  (8'ha9) : forvar5148)))};
                    end
                end
              for (forvar5231 = (1'h0); (forvar5231 < (2'h3)); forvar5231 = (forvar5231 + (1'h1)))
                begin
                  if ($signed(reg4722[(1'h1):(1'h0)]))
                    begin
                      reg5232 <= $unsigned((&forvar4989));
                      reg5233 <= ($signed(reg4726[(3'h4):(1'h1)]) ?
                          {(~&(reg4687 ?
                                  (8'ha8) : reg5028))} : (reg4660 >>> $unsigned($signed((8'hb8)))));
                      reg5234 <= (~|(8'ha9));
                      reg5235 <= $unsigned(($signed(reg5136) + $signed((~reg4658))));
                    end
                  else
                    begin
                      reg5232 <= reg5048[(3'h4):(2'h2)];
                      reg5233 <= $signed($unsigned((~^$unsigned(reg5054))));
                    end
                  if (reg5226[(3'h4):(1'h0)])
                    begin
                      reg5236 <= reg5169;
                      reg5237 <= $unsigned((-(reg4950[(3'h6):(2'h2)] < (reg5087 ?
                          reg5192 : reg5172))));
                    end
                  else
                    begin
                      reg5236 <= {reg4775};
                      reg5237 <= (-$unsigned(forvar4977[(2'h2):(1'h1)]));
                      reg5238 <= reg4594[(3'h5):(3'h4)];
                    end
                end
            end
        end
      for (forvar5270 = (1'h0); (forvar5270 < (1'h0)); forvar5270 = (forvar5270 + (1'h1)))
        begin
          reg5271 <= reg4888[(2'h2):(1'h0)];
          if (($unsigned((((8'ha8) & reg4710) || reg5037[(2'h2):(1'h1)])) < forvar4616))
            begin
              for (forvar5272 = (1'h0); (forvar5272 < (2'h3)); forvar5272 = (forvar5272 + (1'h1)))
                begin
                  reg5273 <= (($signed((-reg4776)) ?
                      $signed((reg4985 - reg4914)) : (^reg4770)) & reg5140);
                  for (forvar5274 = (1'h0); (forvar5274 < (1'h0)); forvar5274 = (forvar5274 + (1'h1)))
                    begin
                      reg5275 <= $signed($signed(forvar4663));
                      reg5276 <= {reg4934};
                      reg5277 <= ((~reg5072[(4'hc):(4'h9)]) ?
                          ((8'hb9) - forvar4813) : forvar4910[(3'h7):(2'h2)]);
                      reg5278 <= forvar4617;
                    end
                  reg5279 <= reg4984;
                end
              for (forvar5280 = (1'h0); (forvar5280 < (2'h2)); forvar5280 = (forvar5280 + (1'h1)))
                begin
                  for (forvar5281 = (1'h0); (forvar5281 < (2'h2)); forvar5281 = (forvar5281 + (1'h1)))
                    begin
                      reg5282 <= {{reg4741[(3'h4):(2'h2)]}};
                      reg5283 <= {reg5163[(3'h5):(2'h3)]};
                      reg5284 <= ($unsigned(reg5263) <= forvar5062[(2'h3):(1'h1)]);
                    end
                  for (forvar5285 = (1'h0); (forvar5285 < (2'h3)); forvar5285 = (forvar5285 + (1'h1)))
                    begin
                      reg5286 <= (!$signed($unsigned((8'hb0))));
                      reg5287 <= $signed($signed($signed((reg5216 << reg5273))));
                      reg5288 <= $signed($unsigned((reg4852 > $signed(reg4926))));
                      reg5289 <= (($signed((reg5237 & (8'hb1))) ?
                          reg4866[(3'h4):(3'h4)] : reg4676) ^ $signed($signed($unsigned(reg4871))));
                    end
                  if (($signed((~{reg4880})) <<< (~&((reg5242 << reg4861) ?
                      reg5013[(1'h1):(1'h0)] : reg4928))))
                    begin
                      reg5290 <= (-(((8'ha6) + (reg4680 ?
                              reg5030 : forvar4689)) ?
                          (reg5021[(2'h2):(1'h1)] >> $unsigned(forvar4969)) : $unsigned((|reg4793))));
                      reg5291 <= reg5164[(4'hc):(4'ha)];
                    end
                  else
                    begin
                      reg5290 <= (reg5127[(2'h2):(2'h2)] ?
                          ({$signed(reg5144)} ?
                              $signed($unsigned((8'h9d))) : (((8'h9d) <= reg4701) ?
                                  reg5081[(3'h5):(1'h0)] : (-(8'haa)))) : $signed({forvar5076}));
                    end
                end
              if (((reg4690[(1'h1):(1'h0)] != $signed(((8'hb0) ?
                  forvar5238 : reg4793))) <<< (|$signed(forvar5088))))
                begin
                  if (reg4638)
                    begin
                      reg5292 <= (^{$unsigned((reg5245 || forvar5234))});
                    end
                  else
                    begin
                      reg5292 <= {$signed((8'hba))};
                      reg5293 <= (reg4921 >> (reg4909 == $unsigned($unsigned(reg4741))));
                      reg5294 <= ((~^(forvar5088[(2'h3):(2'h2)] ?
                              (reg5249 ? forvar5093 : reg4883) : reg4895)) ?
                          reg5032[(2'h3):(1'h1)] : ($signed((forvar5185 ?
                                  reg4901 : wire4574)) ?
                              (|{reg4883}) : ((reg5055 ? forvar4839 : (8'hb1)) ?
                                  forvar4909 : forvar4795[(4'hc):(1'h1)])));
                      reg5295 <= (~|$signed(reg4627));
                    end
                  if ({reg4727[(1'h1):(1'h0)]})
                    begin
                      reg5296 <= (reg5199 ?
                          $signed(($unsigned(reg4584) ?
                              reg5080 : ((8'ha8) <= (8'hab)))) : $signed(($unsigned(forvar4806) <= (reg5192 ?
                              forvar5084 : reg5086))));
                    end
                  else
                    begin
                      reg5296 <= (8'hb0);
                      reg5297 <= forvar4663[(1'h1):(1'h0)];
                    end
                  for (forvar5298 = (1'h0); (forvar5298 < (1'h1)); forvar5298 = (forvar5298 + (1'h1)))
                    begin
                      reg5299 <= (~|(|($unsigned((8'ha2)) ?
                          {forvar5090} : forvar5083)));
                      reg5300 <= (reg4636 || ($signed((reg5297 ?
                              reg4969 : reg4794)) ?
                          reg4778[(3'h4):(1'h1)] : (8'hb2)));
                    end
                end
              else
                begin
                  for (forvar5292 = (1'h0); (forvar5292 < (1'h0)); forvar5292 = (forvar5292 + (1'h1)))
                    begin
                      reg5293 <= {{{$unsigned((8'hb2))}}};
                      reg5294 <= ((&reg4961) && $unsigned(reg5293[(3'h4):(1'h0)]));
                      reg5295 <= (((8'hb8) ?
                          forvar4705[(1'h1):(1'h1)] : reg4913[(1'h1):(1'h0)]) - reg4784);
                    end
                  reg5296 <= {{((^~reg5037) ?
                              $signed(reg4932) : (forvar5280 ?
                                  forvar4801 : reg5253))}};
                  for (forvar5297 = (1'h0); (forvar5297 < (2'h3)); forvar5297 = (forvar5297 + (1'h1)))
                    begin
                      reg5298 <= $unsigned($unsigned(((reg5023 ?
                          reg4773 : forvar4624) ~^ (reg4600 ?
                          reg5069 : reg4959))));
                      reg5299 <= (&reg4719);
                      reg5300 <= ($unsigned(reg5024) < (forvar4591[(1'h0):(1'h0)] ^~ $unsigned((reg5220 || forvar5064))));
                      reg5301 <= $signed($unsigned(reg5103));
                    end
                  if (((~^reg5014[(1'h1):(1'h0)]) >>> ((reg4914[(1'h1):(1'h0)] ?
                      (+forvar5049) : (reg5133 ?
                          reg4967 : forvar5157)) << $unsigned({reg4587}))))
                    begin
                      reg5302 <= $unsigned(({reg4903} ?
                          (~|(forvar5076 < (8'h9d))) : {reg5144}));
                    end
                  else
                    begin
                      reg5302 <= ($signed(reg5214[(3'h5):(3'h4)]) ?
                          (^(-(reg5084 | reg5271))) : reg5039[(1'h0):(1'h0)]);
                    end
                end
            end
          else
            begin
              if (reg5254)
                begin
                  reg5272 <= $unsigned((~&(~|(reg5215 ?
                      reg5042 : forvar5063))));
                  if (reg5260)
                    begin
                      reg5273 <= ((reg4708[(2'h3):(1'h0)] * (+reg5256[(4'hd):(4'h9)])) ?
                          $unsigned($unsigned((~^forvar4941))) : (~|$unsigned((reg4700 ?
                              (8'hab) : forvar5157))));
                      reg5274 <= ($signed({reg4784}) ?
                          reg5089 : ($unsigned(reg4996[(3'h6):(2'h2)]) ?
                              {$unsigned(forvar4933)} : ({forvar4974} ?
                                  (forvar4839 ?
                                      reg5227 : forvar4652) : $signed(forvar5068))));
                      reg5275 <= reg4738[(1'h0):(1'h0)];
                      reg5276 <= {{($signed(reg4808) <= (reg4939 >= reg4845))}};
                    end
                  else
                    begin
                      reg5273 <= {(&{{reg4794}})};
                      reg5274 <= $unsigned($unsigned($unsigned($signed(forvar4944))));
                      reg5275 <= $unsigned(reg4784);
                    end
                  for (forvar5277 = (1'h0); (forvar5277 < (2'h3)); forvar5277 = (forvar5277 + (1'h1)))
                    begin
                      reg5278 <= forvar5035[(2'h2):(2'h2)];
                      reg5279 <= {(^$unsigned(forvar5084[(1'h0):(1'h0)]))};
                      reg5280 <= (~$signed(forvar4777));
                    end
                end
              else
                begin
                  for (forvar5272 = (1'h0); (forvar5272 < (1'h1)); forvar5272 = (forvar5272 + (1'h1)))
                    begin
                      reg5273 <= $signed($unsigned(((forvar4826 ?
                          reg4750 : forvar5008) >= $unsigned(reg5027))));
                    end
                  for (forvar5274 = (1'h0); (forvar5274 < (2'h2)); forvar5274 = (forvar5274 + (1'h1)))
                    begin
                      reg5275 <= reg4857;
                      reg5276 <= ($signed(reg5201) ?
                          $signed((~&(reg5154 + reg4748))) : ($signed(reg4655[(1'h1):(1'h0)]) >> ($signed(reg5184) ?
                              (~|reg5011) : (!(8'hb1)))));
                    end
                  for (forvar5277 = (1'h0); (forvar5277 < (2'h2)); forvar5277 = (forvar5277 + (1'h1)))
                    begin
                      reg5278 <= ($unsigned($unsigned($signed(reg4885))) ~^ ($unsigned({reg4607}) ?
                          $unsigned((reg5077 ?
                              reg5022 : forvar5243)) : $unsigned($unsigned(forvar5150))));
                    end
                  if ($signed(reg4851))
                    begin
                      reg5279 <= {((-$unsigned(forvar5198)) << $signed((!reg5077)))};
                      reg5280 <= (~&$unsigned({reg4680}));
                    end
                  else
                    begin
                      reg5279 <= reg4872[(1'h1):(1'h0)];
                    end
                end
              if (forvar4758)
                begin
                  if ((^~($signed(forvar4609) ?
                      ($signed(forvar4745) ?
                          (reg4847 ?
                              reg5112 : reg5054) : forvar4654[(1'h1):(1'h0)]) : (((8'ha1) * (8'ha4)) ?
                          (8'haa) : $unsigned(reg5053)))))
                    begin
                      reg5281 <= $unsigned(reg5056[(3'h7):(3'h7)]);
                      reg5282 <= forvar5039[(3'h4):(3'h4)];
                      reg5283 <= ($unsigned((&(reg5122 ? (8'ha6) : reg4729))) ?
                          {(-reg4908)} : (8'hb3));
                      reg5284 <= reg4632;
                    end
                  else
                    begin
                      reg5281 <= $unsigned($unsigned(reg5007[(2'h2):(1'h0)]));
                      reg5282 <= $signed((~&(~&forvar5270[(2'h3):(2'h3)])));
                    end
                end
              else
                begin
                  for (forvar5281 = (1'h0); (forvar5281 < (1'h1)); forvar5281 = (forvar5281 + (1'h1)))
                    begin
                      reg5282 <= $unsigned((reg4862 ?
                          reg5159[(1'h0):(1'h0)] : $signed({reg4735})));
                      reg5283 <= $signed(forvar5114[(1'h1):(1'h0)]);
                    end
                  for (forvar5284 = (1'h0); (forvar5284 < (1'h1)); forvar5284 = (forvar5284 + (1'h1)))
                    begin
                      reg5285 <= forvar4858[(2'h2):(2'h2)];
                      reg5286 <= $signed({reg4602});
                      reg5287 <= reg5131;
                    end
                  if (($signed(($signed(reg4654) <= reg4591[(1'h0):(1'h0)])) ?
                      (+($signed(forvar5114) ?
                          (^forvar4801) : $unsigned(forvar4760))) : reg5158))
                    begin
                      reg5288 <= (({reg4969} ?
                          (-$signed((8'hba))) : reg4590) || (+$unsigned($unsigned(reg4660))));
                    end
                  else
                    begin
                      reg5288 <= $signed((8'ha9));
                      reg5289 <= (((reg4969[(2'h2):(1'h1)] ?
                                  $unsigned(reg4709) : (+reg5035)) ?
                              reg4692 : forvar5114) ?
                          $unsigned({(~^reg4633)}) : wire5196[(2'h3):(1'h0)]);
                    end
                  if (((-reg5199[(2'h2):(1'h0)]) ?
                      ($signed({forvar4815}) ?
                          $signed((reg5139 ?
                              reg5289 : reg4949)) : ((~&(8'hab)) ?
                              reg4779[(2'h2):(2'h2)] : (reg4670 ?
                                  reg5118 : reg5252))) : ((reg5036 <= $unsigned(forvar5162)) & $signed((~reg4646)))))
                    begin
                      reg5290 <= forvar4610[(3'h5):(1'h1)];
                      reg5291 <= $signed(((8'h9f) != $signed(reg5228)));
                      reg5292 <= ($signed((reg4994 ?
                          (-reg4591) : {reg5080})) >= reg4986);
                      reg5293 <= ($unsigned(reg4925) || {(~^reg4853)});
                    end
                  else
                    begin
                      reg5290 <= ($unsigned($unsigned(reg4822[(4'h9):(3'h4)])) ?
                          ((reg5016 ?
                              {reg5011} : (~|reg4762)) && reg4728) : (~^reg4607[(3'h6):(3'h5)]));
                      reg5291 <= reg4952;
                      reg5292 <= {reg5023};
                    end
                end
              if ((reg5103[(2'h3):(1'h1)] ^ forvar4689[(4'hd):(4'hd)]))
                begin
                  if ($signed(reg4646[(2'h3):(2'h3)]))
                    begin
                      reg5294 <= (!reg4645[(2'h3):(2'h3)]);
                      reg5295 <= reg4790;
                      reg5296 <= reg4689[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg5294 <= $unsigned($unsigned(((+forvar4914) >> {reg4709})));
                      reg5295 <= (~((reg4581 ?
                          forvar4640 : {(8'haa)}) != ($signed((8'ha7)) <= (forvar5104 != reg5143))));
                      reg5296 <= ((($signed(reg4780) ~^ $unsigned(reg4729)) | forvar4759) ?
                          ($signed((~^forvar4584)) ?
                              $unsigned(forvar4837[(4'hc):(3'h7)]) : ({reg4752} ?
                                  reg4948[(2'h2):(1'h1)] : forvar4763)) : (($signed(reg4838) ?
                                  (reg5254 ? forvar4694 : reg5186) : reg4992) ?
                              ((forvar5284 ? reg4622 : forvar4594) ?
                                  {reg4615} : $unsigned(reg5049)) : {$signed(reg5032)}));
                      reg5297 <= (!((&$signed(reg5131)) ?
                          $unsigned((forvar5234 ^~ reg4942)) : ((~|(8'ha0)) ?
                              reg4642[(3'h6):(3'h4)] : (^reg4614))));
                    end
                  if (reg5192)
                    begin
                      reg5298 <= reg5227[(1'h1):(1'h0)];
                      reg5299 <= (8'ha6);
                    end
                  else
                    begin
                      reg5298 <= reg4906[(3'h6):(1'h0)];
                      reg5299 <= reg4708;
                      reg5300 <= $signed(wire5196[(2'h3):(1'h0)]);
                    end
                  for (forvar5301 = (1'h0); (forvar5301 < (1'h1)); forvar5301 = (forvar5301 + (1'h1)))
                    begin
                      reg5302 <= forvar5248[(2'h3):(1'h0)];
                      reg5303 <= ({reg5037} ?
                          (!((reg4999 ?
                              forvar4584 : forvar5252) << (8'ha2))) : (^($signed(forvar4944) >> $signed(reg4935))));
                      reg5304 <= ($signed($signed($unsigned((8'ha5)))) > (~^$unsigned(((8'hae) ?
                          reg5297 : forvar4656))));
                    end
                  reg5305 <= (reg4912[(3'h4):(2'h2)] ?
                      (^(8'hb7)) : $unsigned($signed($signed(reg5011))));
                end
              else
                begin
                  if ($signed(((reg5249[(4'hb):(2'h2)] ?
                      {reg4767} : (reg5033 ?
                          reg5245 : forvar4745)) || (+$signed(forvar4827)))))
                    begin
                      reg5294 <= reg5003[(1'h0):(1'h0)];
                      reg5295 <= reg4680[(3'h7):(3'h5)];
                    end
                  else
                    begin
                      reg5294 <= ((reg4996[(3'h6):(3'h5)] ?
                          (8'hba) : reg4791) == reg4988[(1'h1):(1'h1)]);
                      reg5295 <= ((-{{forvar4819}}) || forvar4786[(3'h6):(3'h4)]);
                      reg5296 <= (reg5069[(4'hb):(4'h8)] ?
                          (((|reg4996) ?
                              $signed((8'hb7)) : (reg5093 ?
                                  reg5296 : reg5258)) + reg4702[(3'h5):(1'h0)]) : ($unsigned((reg4720 - reg4605)) > (8'hb1)));
                    end
                  for (forvar5297 = (1'h0); (forvar5297 < (2'h3)); forvar5297 = (forvar5297 + (1'h1)))
                    begin
                      reg5298 <= forvar5083;
                      reg5299 <= $unsigned(reg5152[(4'hb):(3'h7)]);
                      reg5300 <= reg4584;
                      reg5301 <= reg5027[(1'h0):(1'h0)];
                    end
                  for (forvar5302 = (1'h0); (forvar5302 < (2'h2)); forvar5302 = (forvar5302 + (1'h1)))
                    begin
                      reg5303 <= (({$unsigned((8'hae))} < {{reg5268}}) * reg4855[(2'h2):(1'h1)]);
                      reg5304 <= $signed((forvar4602[(3'h6):(2'h3)] + (^~$unsigned((8'h9c)))));
                      reg5305 <= (forvar5002 ?
                          $signed($signed((reg4834 ?
                              reg5143 : forvar5198))) : $signed(($unsigned(reg5241) ?
                              reg4857 : reg5174[(4'h8):(3'h5)])));
                    end
                end
            end
        end
      for (forvar5306 = (1'h0); (forvar5306 < (2'h3)); forvar5306 = (forvar5306 + (1'h1)))
        begin
          for (forvar5307 = (1'h0); (forvar5307 < (1'h1)); forvar5307 = (forvar5307 + (1'h1)))
            begin
              if ($signed((-(reg5185 ?
                  reg4873[(2'h2):(1'h1)] : reg5107[(2'h2):(1'h1)]))))
                begin
                  if (reg4895)
                    begin
                      reg5308 <= $unsigned($signed(($signed(reg4584) ?
                          $signed(reg4612) : {(8'had)})));
                      reg5309 <= (|reg4880[(3'h7):(2'h3)]);
                    end
                  else
                    begin
                      reg5308 <= reg4888;
                      reg5309 <= reg5210[(3'h4):(3'h4)];
                    end
                  reg5310 <= (-(forvar4688 ?
                      forvar5186 : (~^reg4686[(3'h6):(2'h3)])));
                end
              else
                begin
                  reg5308 <= reg4624[(3'h5):(3'h5)];
                  reg5309 <= (forvar5117[(3'h4):(1'h1)] >>> ($unsigned((forvar5149 ?
                          reg5002 : reg4961)) ?
                      forvar4672[(2'h2):(1'h0)] : $signed(((8'hb4) <<< reg4850))));
                  if (reg4740)
                    begin
                      reg5310 <= reg5121[(4'h8):(4'h8)];
                      reg5311 <= (((8'haf) ?
                              ($signed(wire4576) <= reg5243[(3'h4):(2'h3)]) : (forvar4698 <<< $signed(reg5119))) ?
                          (8'ha1) : (&reg4622[(1'h0):(1'h0)]));
                      reg5312 <= reg5262[(3'h4):(2'h2)];
                      reg5313 <= ((((!reg5247) > forvar5068[(2'h3):(1'h0)]) << (^~(8'haf))) <<< (reg4715[(1'h1):(1'h0)] * (reg5142 ?
                          $signed(reg5094) : $unsigned(reg5227))));
                    end
                  else
                    begin
                      reg5310 <= $signed(forvar4912);
                      reg5311 <= reg5023;
                    end
                end
              if ({reg4605[(3'h5):(3'h5)]})
                begin
                  for (forvar5314 = (1'h0); (forvar5314 < (1'h1)); forvar5314 = (forvar5314 + (1'h1)))
                    begin
                      reg5315 <= (~reg4636);
                      reg5316 <= $signed($signed(((reg5023 ?
                          reg4791 : wire4575) ^~ (reg4930 ?
                          reg4623 : reg4723))));
                      reg5317 <= (8'ha5);
                      reg5318 <= ($signed(reg4745[(3'h7):(3'h6)]) != $signed(((reg4825 ?
                          reg5061 : forvar4744) && reg4630[(3'h5):(3'h4)])));
                    end
                  if ($unsigned($unsigned($signed($unsigned(reg5183)))))
                    begin
                      reg5319 <= $unsigned(reg5090[(2'h3):(2'h3)]);
                      reg5320 <= $unsigned((~reg5299[(3'h5):(3'h4)]));
                    end
                  else
                    begin
                      reg5319 <= $signed({reg4935});
                      reg5320 <= (^~reg5038[(3'h5):(3'h5)]);
                      reg5321 <= (forvar5138[(1'h0):(1'h0)] & forvar4648[(3'h4):(1'h1)]);
                      reg5322 <= forvar4577;
                    end
                end
              else
                begin
                  if ((forvar5280 ?
                      reg5042[(1'h1):(1'h1)] : forvar4698[(4'h9):(1'h1)]))
                    begin
                      reg5314 <= ($unsigned(((reg5020 >> reg4955) | ((8'hb1) ?
                              reg4860 : reg5209))) ?
                          reg4988 : (^(!(~^reg4909))));
                      reg5315 <= $signed(($signed(reg4771) && reg5243[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg5314 <= $unsigned($unsigned($signed((forvar4663 ?
                          reg5029 : (8'had)))));
                    end
                end
              for (forvar5323 = (1'h0); (forvar5323 < (2'h2)); forvar5323 = (forvar5323 + (1'h1)))
                begin
                  if (reg4707[(4'hd):(3'h6)])
                    begin
                      reg5324 <= $signed(((~^$signed(reg4912)) ?
                          $signed({(8'hba)}) : $unsigned($unsigned(forvar5298))));
                    end
                  else
                    begin
                      reg5324 <= (8'hb5);
                      reg5325 <= (($signed({reg4936}) ?
                              reg4586[(2'h3):(1'h0)] : ((+forvar4972) & forvar4738[(1'h1):(1'h1)])) ?
                          ((^(reg4611 <= reg5305)) ?
                              (reg5121 ?
                                  (reg5161 ?
                                      reg5069 : forvar5106) : reg4846) : {$unsigned(forvar4603)}) : {$signed((reg5085 && forvar4593))});
                    end
                  for (forvar5326 = (1'h0); (forvar5326 < (1'h1)); forvar5326 = (forvar5326 + (1'h1)))
                    begin
                      reg5327 <= ((|forvar4850[(3'h6):(3'h6)]) ?
                          ((&reg5095[(3'h4):(3'h4)]) - ($signed(forvar5261) ?
                              (~|(8'ha8)) : reg4816[(4'hc):(4'h9)])) : (~^($unsigned(reg4609) ?
                              {reg4951} : $unsigned(reg4742))));
                    end
                end
              for (forvar5328 = (1'h0); (forvar5328 < (1'h0)); forvar5328 = (forvar5328 + (1'h1)))
                begin
                  if (($unsigned($signed(reg5258[(2'h3):(1'h1)])) && (forvar4986[(2'h3):(2'h2)] <= ((reg4859 - reg4997) * reg5114[(1'h0):(1'h0)]))))
                    begin
                      reg5329 <= forvar4694[(4'hc):(1'h1)];
                      reg5330 <= $signed(({(reg5194 ? reg5208 : forvar5006)} ?
                          ((^~(8'hb9)) << {reg4748}) : $signed((reg4692 ?
                              reg4993 : wire4940))));
                      reg5331 <= ((+(reg5033 ? (^(8'haa)) : reg4948)) ?
                          reg4697 : forvar4877[(4'hc):(3'h7)]);
                    end
                  else
                    begin
                      reg5329 <= reg5145[(2'h3):(2'h3)];
                      reg5330 <= $signed($signed((reg4751[(2'h2):(1'h1)] ?
                          (forvar5208 ?
                              reg4658 : (8'ha9)) : (forvar4986 || reg5304))));
                      reg5331 <= forvar5082;
                      reg5332 <= ((8'hae) ?
                          $unsigned(reg4828[(3'h6):(1'h0)]) : ($signed((reg5072 ?
                                  forvar5234 : (8'h9f))) ?
                              {$unsigned(forvar4915)} : ((~reg4697) ?
                                  (reg4832 ? reg5312 : reg4714) : {reg4999})));
                    end
                  if ({{$unsigned((reg5287 ? forvar4712 : reg5073))}})
                    begin
                      reg5333 <= (~|$unsigned(reg5254));
                      reg5334 <= (~^wire4798[(3'h6):(1'h0)]);
                      reg5335 <= ({(reg4635[(3'h5):(3'h5)] ?
                                  $unsigned(reg4727) : (forvar4814 >>> reg4647))} ?
                          ((^(reg5154 ?
                              reg4786 : reg4775)) + reg5303) : (8'hae));
                    end
                  else
                    begin
                      reg5333 <= (~|$signed(({forvar5088} ?
                          ((8'ha6) != reg4603) : forvar4694[(2'h2):(1'h0)])));
                      reg5334 <= ($unsigned((~^reg4684)) * reg5085[(3'h6):(2'h2)]);
                      reg5335 <= forvar4969;
                    end
                  if ((!reg4803[(1'h1):(1'h1)]))
                    begin
                      reg5336 <= reg4844;
                      reg5337 <= $unsigned((+$unsigned((forvar4819 ?
                          reg4810 : reg4728))));
                    end
                  else
                    begin
                      reg5336 <= reg5125;
                      reg5337 <= forvar5186;
                      reg5338 <= $unsigned($unsigned((-(reg5191 ?
                          reg5290 : (8'hb0)))));
                      reg5339 <= $unsigned((~^$unsigned($unsigned(reg4743))));
                    end
                end
            end
          for (forvar5340 = (1'h0); (forvar5340 < (2'h3)); forvar5340 = (forvar5340 + (1'h1)))
            begin
              for (forvar5341 = (1'h0); (forvar5341 < (2'h3)); forvar5341 = (forvar5341 + (1'h1)))
                begin
                  if ($signed((reg5022 ?
                      reg4907[(3'h5):(1'h0)] : $unsigned(((8'hb4) ?
                          forvar5165 : forvar5217)))))
                    begin
                      reg5342 <= ({reg5057[(2'h3):(2'h2)]} * ((8'h9f) * reg5189[(2'h3):(2'h2)]));
                      reg5343 <= (~reg4882);
                      reg5344 <= $signed({(-(!reg4928))});
                    end
                  else
                    begin
                      reg5342 <= reg5053[(1'h1):(1'h0)];
                      reg5343 <= reg5309;
                      reg5344 <= reg5014[(1'h1):(1'h0)];
                    end
                  if ($signed(reg5344))
                    begin
                      reg5345 <= ((((!forvar4749) || $signed((8'h9d))) & forvar5005) || reg4766[(1'h1):(1'h1)]);
                      reg5346 <= ($signed(forvar4929) <<< $signed(forvar4840[(4'h9):(1'h1)]));
                      reg5347 <= forvar5229[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg5345 <= ({reg5236} <= {forvar5198});
                      reg5346 <= (reg4613 ?
                          (|(-$unsigned((8'hb8)))) : (reg4807[(3'h5):(1'h1)] ?
                              $signed($signed(forvar4913)) : ($signed(reg4997) ?
                                  (~|wire4576) : reg4976[(3'h4):(1'h0)])));
                      reg5347 <= $signed({forvar4636});
                      reg5348 <= $unsigned((|reg4742[(2'h3):(1'h1)]));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ((reg4655[(3'h6):(3'h6)] ?
          reg4682[(1'h0):(1'h0)] : $unsigned($signed((8'ha3)))))
        begin
          for (forvar5349 = (1'h0); (forvar5349 < (1'h1)); forvar5349 = (forvar5349 + (1'h1)))
            begin
              for (forvar5350 = (1'h0); (forvar5350 < (2'h2)); forvar5350 = (forvar5350 + (1'h1)))
                begin
                  if (forvar4933)
                    begin
                      reg5351 <= (reg5011[(3'h4):(2'h3)] ~^ $unsigned((+(reg4744 != reg4989))));
                    end
                  else
                    begin
                      reg5351 <= forvar4877;
                      reg5352 <= forvar4749[(2'h2):(1'h1)];
                      reg5353 <= ($signed(forvar4777) >> reg4656[(2'h2):(2'h2)]);
                    end
                  reg5354 <= (reg4970[(2'h3):(1'h0)] ?
                      (~&$unsigned((reg5054 ?
                          reg4893 : reg4916))) : ($signed(((8'hb6) >>> reg5342)) - (reg5325[(4'h8):(2'h2)] ?
                          reg5074 : (reg4928 ? reg4687 : reg5072))));
                end
              if ((($unsigned((^~forvar4578)) ~^ {reg4744[(1'h1):(1'h0)]}) & $signed($signed($unsigned((8'hb3))))))
                begin
                  for (forvar5355 = (1'h0); (forvar5355 < (2'h3)); forvar5355 = (forvar5355 + (1'h1)))
                    begin
                      reg5356 <= ((~|$signed($signed((8'hba)))) || (((forvar4642 ?
                              forvar4988 : reg4579) ?
                          $unsigned(reg5025) : {reg5236}) >> reg4789));
                      reg5357 <= (~^reg4598);
                      reg5358 <= reg4627[(2'h2):(2'h2)];
                    end
                  if ((&reg4834[(2'h2):(1'h1)]))
                    begin
                      reg5359 <= (~^{reg4986[(2'h3):(1'h0)]});
                    end
                  else
                    begin
                      reg5359 <= (8'ha5);
                      reg5360 <= (~|reg4662);
                      reg5361 <= $unsigned(($signed((~&forvar4815)) & ($signed(reg4880) != (~reg4589))));
                      reg5362 <= ((!reg5201) << $unsigned($unsigned((8'hab))));
                    end
                end
              else
                begin
                  reg5355 <= reg5130;
                end
              for (forvar5363 = (1'h0); (forvar5363 < (2'h2)); forvar5363 = (forvar5363 + (1'h1)))
                begin
                  if ($signed($signed($unsigned($signed(forvar5135)))))
                    begin
                      reg5364 <= (8'hb2);
                      reg5365 <= ($signed(reg5249[(1'h0):(1'h0)]) - reg4581[(3'h5):(3'h5)]);
                      reg5366 <= ((~&$signed(reg5181)) ?
                          (&forvar5208[(1'h1):(1'h0)]) : forvar5297[(1'h0):(1'h0)]);
                      reg5367 <= reg5353;
                    end
                  else
                    begin
                      reg5364 <= $unsigned({($unsigned(forvar5148) + $unsigned(reg4900))});
                      reg5365 <= {{($unsigned(reg5238) * ((8'ha6) ?
                                  reg4631 : (8'ha3)))}};
                      reg5366 <= $signed((+reg5240));
                    end
                end
              for (forvar5368 = (1'h0); (forvar5368 < (2'h2)); forvar5368 = (forvar5368 + (1'h1)))
                begin
                  if ($unsigned($signed((forvar4611 << (~|reg5318)))))
                    begin
                      reg5369 <= reg4744[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg5369 <= reg5156;
                    end
                  for (forvar5370 = (1'h0); (forvar5370 < (2'h2)); forvar5370 = (forvar5370 + (1'h1)))
                    begin
                      reg5371 <= {((reg4765 >= (forvar5006 ?
                              forvar5111 : reg4954)) < (((8'ha5) ~^ reg5263) ?
                              $signed(reg5295) : $signed(reg4839)))};
                    end
                  for (forvar5372 = (1'h0); (forvar5372 < (2'h2)); forvar5372 = (forvar5372 + (1'h1)))
                    begin
                      reg5373 <= $signed({$unsigned((^reg5121))});
                      reg5374 <= ($signed(forvar5284[(2'h3):(2'h3)]) ?
                          (~^(8'hab)) : (reg4932[(4'he):(4'h9)] ~^ reg4741));
                    end
                end
            end
          if ($unsigned((reg5255 | $unsigned(reg4683))))
            begin
              for (forvar5375 = (1'h0); (forvar5375 < (1'h0)); forvar5375 = (forvar5375 + (1'h1)))
                begin
                  reg5376 <= $signed($unsigned($unsigned((-reg5080))));
                end
              for (forvar5377 = (1'h0); (forvar5377 < (2'h3)); forvar5377 = (forvar5377 + (1'h1)))
                begin
                  reg5378 <= $signed((reg5074[(1'h0):(1'h0)] && ($signed((8'ha3)) * {reg4590})));
                  reg5379 <= (-(~reg4930));
                  for (forvar5380 = (1'h0); (forvar5380 < (2'h2)); forvar5380 = (forvar5380 + (1'h1)))
                    begin
                      reg5381 <= $signed($unsigned(forvar4745[(3'h6):(3'h6)]));
                      reg5382 <= ((forvar4643[(4'hd):(2'h3)] ?
                          (~^(!(8'hac))) : ({forvar4910} < (forvar4819 ?
                              reg4902 : forvar4598))) ^ (!((~reg4931) || (reg5204 ?
                          reg4864 : reg4719))));
                      reg5383 <= (((~&(forvar4843 ?
                          reg4897 : (8'ha7))) >>> $signed(reg4942)) | {$signed((reg5009 && forvar5020))});
                      reg5384 <= {$signed({((8'ha4) ? reg5366 : reg4910)})};
                    end
                end
              reg5385 <= $unsigned((forvar4914[(1'h0):(1'h0)] * $unsigned((~&reg4910))));
            end
          else
            begin
              for (forvar5375 = (1'h0); (forvar5375 < (1'h1)); forvar5375 = (forvar5375 + (1'h1)))
                begin
                  for (forvar5376 = (1'h0); (forvar5376 < (1'h0)); forvar5376 = (forvar5376 + (1'h1)))
                    begin
                      reg5377 <= (reg5285 ?
                          (reg4711 ^~ (~^reg5019)) : $signed($unsigned((forvar4815 ?
                              reg5018 : (8'ha1)))));
                      reg5378 <= forvar4864;
                    end
                  reg5379 <= (+(($unsigned(reg4591) != $unsigned(reg4639)) ?
                      forvar5372 : $unsigned((reg5208 < (8'hb8)))));
                end
              if ((reg5142[(2'h3):(2'h3)] <<< $unsigned(forvar4986)))
                begin
                  if ((-forvar4909))
                    begin
                      reg5380 <= ($signed($unsigned((~&(8'ha3)))) ?
                          $unsigned(($unsigned(forvar4874) ?
                              {(8'ha5)} : (-reg4948))) : (((forvar4636 ?
                              reg5273 : reg4757) || $signed(forvar4673)) >> (reg5237[(3'h6):(2'h3)] >> (reg4660 ^~ reg5029))));
                      reg5381 <= forvar5370;
                      reg5382 <= ($unsigned(reg4664[(2'h3):(1'h0)]) == {reg5140[(1'h0):(1'h0)]});
                      reg5383 <= $unsigned($signed($unsigned(((8'hb4) ?
                          reg5163 : reg4788))));
                    end
                  else
                    begin
                      reg5380 <= (~&(reg4771[(4'h8):(3'h4)] >>> reg4907));
                      reg5381 <= {$signed((8'ha0))};
                      reg5382 <= {$signed(({reg4903} - $unsigned(reg4818)))};
                    end
                  if (reg5351)
                    begin
                      reg5384 <= ($unsigned($unsigned((forvar4688 ?
                              reg4695 : reg5211))) ?
                          $unsigned($signed((^reg4776))) : reg4765);
                    end
                  else
                    begin
                      reg5384 <= $unsigned((reg4635 ?
                          reg4677[(1'h0):(1'h0)] : (^(reg4999 ?
                              forvar4749 : reg4736))));
                      reg5385 <= ($unsigned(reg4985) ?
                          (forvar4727[(4'h8):(3'h7)] ?
                              wire4940 : ((!reg4782) + (forvar5117 < reg4726))) : (reg5085[(3'h5):(1'h1)] ?
                              (reg5278[(3'h4):(2'h2)] ^~ (reg5105 ~^ reg5117)) : reg4686[(2'h3):(1'h1)]));
                      reg5386 <= ($unsigned(((+reg4689) ?
                          reg5120[(1'h0):(1'h0)] : $signed(reg5301))) > (reg4788[(2'h2):(1'h0)] * (~(forvar5175 ?
                          (8'ha3) : reg5320))));
                    end
                end
              else
                begin
                  if (reg5315[(3'h4):(2'h3)])
                    begin
                      reg5380 <= reg4905[(4'ha):(1'h0)];
                    end
                  else
                    begin
                      reg5380 <= reg4632[(2'h3):(1'h0)];
                      reg5381 <= (8'hb8);
                    end
                  for (forvar5382 = (1'h0); (forvar5382 < (2'h3)); forvar5382 = (forvar5382 + (1'h1)))
                    begin
                      reg5383 <= $unsigned($unsigned(reg5347[(4'h9):(3'h4)]));
                      reg5384 <= reg4778;
                    end
                end
              for (forvar5387 = (1'h0); (forvar5387 < (2'h3)); forvar5387 = (forvar5387 + (1'h1)))
                begin
                  for (forvar5388 = (1'h0); (forvar5388 < (1'h0)); forvar5388 = (forvar5388 + (1'h1)))
                    begin
                      reg5389 <= (+$signed(forvar5084[(2'h2):(1'h1)]));
                      reg5390 <= (^$unsigned((~reg5191[(1'h0):(1'h0)])));
                      reg5391 <= $unsigned((reg4946 - ((|reg5096) < $signed((8'hb8)))));
                      reg5392 <= reg5114;
                    end
                  for (forvar5393 = (1'h0); (forvar5393 < (2'h3)); forvar5393 = (forvar5393 + (1'h1)))
                    begin
                      reg5394 <= (($unsigned((^forvar5098)) > (|$signed(reg4910))) ?
                          (8'hac) : reg5116);
                    end
                  for (forvar5395 = (1'h0); (forvar5395 < (2'h2)); forvar5395 = (forvar5395 + (1'h1)))
                    begin
                      reg5396 <= (forvar4809 == $unsigned((!(reg4769 >> reg4656))));
                      reg5397 <= wire4575[(1'h1):(1'h1)];
                      reg5398 <= reg4911[(3'h6):(3'h6)];
                    end
                  if (reg5229)
                    begin
                      reg5399 <= $unsigned((((|(8'h9f)) ^~ reg4991[(2'h2):(1'h0)]) ?
                          (|(8'hb4)) : ($unsigned(reg5080) < forvar4689[(1'h1):(1'h1)])));
                      reg5400 <= reg5242[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg5399 <= wire4576[(2'h2):(2'h2)];
                      reg5400 <= $signed($unsigned(($signed(reg5356) ?
                          (~forvar5083) : reg5356)));
                      reg5401 <= (-({(~|reg5147)} ?
                          ((reg5345 && reg5055) ?
                              forvar5001[(2'h3):(2'h2)] : $unsigned(forvar4851)) : (~reg5269)));
                      reg5402 <= {($unsigned(forvar4848[(2'h2):(2'h2)]) ?
                              {(+reg5002)} : ((reg5223 << forvar5307) ?
                                  (|forvar4988) : (|reg4973)))};
                    end
                end
            end
          for (forvar5403 = (1'h0); (forvar5403 < (2'h2)); forvar5403 = (forvar5403 + (1'h1)))
            begin
              for (forvar5404 = (1'h0); (forvar5404 < (2'h3)); forvar5404 = (forvar5404 + (1'h1)))
                begin
                  for (forvar5405 = (1'h0); (forvar5405 < (2'h3)); forvar5405 = (forvar5405 + (1'h1)))
                    begin
                      reg5406 <= {$unsigned($unsigned((reg5069 ?
                              reg5048 : reg5232)))};
                      reg5407 <= (((!$signed(reg4960)) ?
                          (reg5325[(3'h5):(3'h5)] <<< $unsigned((8'hb9))) : forvar4988) >>> reg4735);
                      reg5408 <= (~|reg4989[(4'h9):(4'h9)]);
                    end
                  for (forvar5409 = (1'h0); (forvar5409 < (2'h2)); forvar5409 = (forvar5409 + (1'h1)))
                    begin
                      reg5410 <= forvar5001[(3'h7):(1'h0)];
                    end
                  if ((forvar5198 << (~|reg4818[(1'h0):(1'h0)])))
                    begin
                      reg5411 <= forvar4840;
                      reg5412 <= (~^$unsigned(forvar4694[(4'he):(4'ha)]));
                      reg5413 <= $signed((^$unsigned(reg4946[(2'h2):(1'h0)])));
                      reg5414 <= $signed($unsigned(((8'h9c) ?
                          ((8'ha9) << forvar4613) : reg4803[(3'h4):(2'h2)])));
                    end
                  else
                    begin
                      reg5411 <= $signed(reg4725[(1'h0):(1'h0)]);
                    end
                  reg5415 <= $unsigned(reg5214);
                end
              for (forvar5416 = (1'h0); (forvar5416 < (1'h1)); forvar5416 = (forvar5416 + (1'h1)))
                begin
                  if ({reg4888})
                    begin
                      reg5417 <= $unsigned(forvar4899[(1'h0):(1'h0)]);
                      reg5418 <= $signed(({(reg4796 >>> (8'hba))} ?
                          $unsigned({(8'hab)}) : ($unsigned(forvar5297) ?
                              (8'hab) : $unsigned(reg5286))));
                      reg5419 <= {(&reg4839[(2'h2):(1'h1)])};
                    end
                  else
                    begin
                      reg5417 <= ((8'hae) << $signed((!$unsigned(reg4669))));
                      reg5418 <= ((~^(^reg4843[(4'h9):(3'h5)])) ~^ ((reg5362 >> (reg4722 ?
                              reg4835 : reg5332)) ?
                          ($unsigned(reg5211) ?
                              forvar4624[(3'h5):(3'h4)] : $unsigned(reg5386)) : (wire5196 ?
                              $signed(reg5332) : (^reg5277))));
                      reg5419 <= (&$signed((~|(8'ha6))));
                    end
                end
              for (forvar5420 = (1'h0); (forvar5420 < (2'h3)); forvar5420 = (forvar5420 + (1'h1)))
                begin
                  if (reg4676)
                    begin
                      reg5421 <= (reg5352 ?
                          {{$signed((8'ha6))}} : (((reg5319 ?
                                      forvar4890 : wire5197) ?
                                  $unsigned(reg4722) : $unsigned(forvar5395)) ?
                              {{reg4763}} : $signed((reg4853 ?
                                  forvar5098 : reg4656))));
                    end
                  else
                    begin
                      reg5421 <= $unsigned(forvar4920[(2'h3):(1'h0)]);
                      reg5422 <= reg4689[(1'h1):(1'h1)];
                    end
                end
            end
          if (reg5160[(1'h1):(1'h0)])
            begin
              reg5423 <= (($signed((-reg4733)) ?
                  $signed({reg5081}) : $signed(reg4680)) <<< (-$signed((reg4831 <<< reg4807))));
              for (forvar5424 = (1'h0); (forvar5424 < (1'h0)); forvar5424 = (forvar5424 + (1'h1)))
                begin
                  if (reg5327[(1'h1):(1'h1)])
                    begin
                      reg5425 <= forvar4806;
                      reg5426 <= $unsigned($signed($unsigned(reg4664[(3'h5):(2'h2)])));
                    end
                  else
                    begin
                      reg5425 <= forvar4789[(2'h3):(1'h1)];
                      reg5426 <= (reg5413 + wire5196[(3'h4):(3'h4)]);
                      reg5427 <= (((~^{forvar4749}) <<< $unsigned(reg5006[(1'h0):(1'h0)])) ?
                          (((reg5410 != reg4658) - {(8'ha7)}) ?
                              (forvar5285 ^ forvar4996) : (^$unsigned((8'haa)))) : $unsigned(reg4838));
                    end
                end
            end
          else
            begin
              for (forvar5423 = (1'h0); (forvar5423 < (2'h3)); forvar5423 = (forvar5423 + (1'h1)))
                begin
                  for (forvar5424 = (1'h0); (forvar5424 < (1'h0)); forvar5424 = (forvar5424 + (1'h1)))
                    begin
                      reg5425 <= ((!(reg4900[(2'h2):(1'h0)] << $unsigned((8'hb8)))) ?
                          reg5276[(2'h2):(1'h0)] : (reg5264[(2'h2):(1'h0)] ?
                              (reg5184 ?
                                  $unsigned(forvar4912) : {reg5178}) : reg4654[(4'hd):(1'h1)]));
                      reg5426 <= $signed({$signed(reg4972[(3'h6):(3'h4)])});
                    end
                  for (forvar5427 = (1'h0); (forvar5427 < (1'h0)); forvar5427 = (forvar5427 + (1'h1)))
                    begin
                      reg5428 <= (~forvar4681);
                      reg5429 <= (forvar4640[(2'h2):(1'h1)] < (forvar4579[(3'h4):(2'h2)] ?
                          reg5359[(3'h5):(1'h1)] : reg5337[(1'h0):(1'h0)]));
                      reg5430 <= reg5026[(1'h1):(1'h1)];
                    end
                  if ($signed(reg4966))
                    begin
                      reg5431 <= $unsigned(((reg4924[(3'h6):(1'h0)] ^~ reg5415[(2'h3):(1'h0)]) + $signed((forvar5297 | reg5054))));
                      reg5432 <= $signed(reg4778);
                      reg5433 <= reg5088[(3'h6):(1'h1)];
                      reg5434 <= (forvar4744[(1'h1):(1'h1)] == reg4864);
                    end
                  else
                    begin
                      reg5431 <= {$signed($unsigned($unsigned(reg5336)))};
                      reg5432 <= (forvar5130 > $signed($unsigned((~|reg5226))));
                      reg5433 <= $signed((reg5337 ?
                          {(reg5297 <<< (8'hb9))} : forvar5186[(3'h5):(2'h3)]));
                    end
                end
              for (forvar5435 = (1'h0); (forvar5435 < (2'h2)); forvar5435 = (forvar5435 + (1'h1)))
                begin
                  for (forvar5436 = (1'h0); (forvar5436 < (1'h0)); forvar5436 = (forvar5436 + (1'h1)))
                    begin
                      reg5437 <= (reg5212 ^ $unsigned(forvar4727[(4'h8):(3'h7)]));
                    end
                  for (forvar5438 = (1'h0); (forvar5438 < (1'h1)); forvar5438 = (forvar5438 + (1'h1)))
                    begin
                      reg5439 <= reg5256[(4'h9):(1'h0)];
                    end
                  for (forvar5440 = (1'h0); (forvar5440 < (2'h2)); forvar5440 = (forvar5440 + (1'h1)))
                    begin
                      reg5441 <= reg4836[(1'h1):(1'h0)];
                    end
                end
              for (forvar5442 = (1'h0); (forvar5442 < (2'h3)); forvar5442 = (forvar5442 + (1'h1)))
                begin
                  if (((-$unsigned((!(8'haa)))) != $signed((reg5286 ^~ (reg5094 != forvar4929)))))
                    begin
                      reg5443 <= (~^($unsigned($signed(reg4763)) ?
                          reg5297 : $unsigned((^forvar4952))));
                      reg5444 <= (!{(reg5214[(2'h3):(2'h3)] & forvar5093[(2'h2):(2'h2)])});
                      reg5445 <= reg5312;
                    end
                  else
                    begin
                      reg5443 <= $signed((reg5112[(4'hd):(3'h5)] == forvar5247));
                      reg5444 <= (^~reg4646[(4'ha):(3'h5)]);
                      reg5445 <= reg5163[(1'h0):(1'h0)];
                    end
                end
              if ((reg5141 && (reg4928 ? reg5179 : (|(reg5347 < reg5015)))))
                begin
                  reg5446 <= ((forvar4688 ?
                      (|(reg4979 ?
                          reg5422 : forvar4899)) : {(forvar4580 == reg4915)}) > (~^((reg5288 - reg4600) << (reg4852 ?
                      forvar4773 : forvar5165))));
                end
              else
                begin
                  if (reg4830)
                    begin
                      reg5446 <= $unsigned(($unsigned(reg4849[(2'h2):(1'h0)]) ?
                          $unsigned((reg4841 <<< reg4577)) : $signed(reg5026)));
                      reg5447 <= $signed(forvar4910);
                      reg5448 <= reg5107[(4'h8):(3'h6)];
                    end
                  else
                    begin
                      reg5446 <= (reg4978[(4'h8):(3'h6)] ?
                          ({{reg5364}} - $signed(forvar5376)) : $signed(((!reg4700) ^ reg5168[(1'h1):(1'h0)])));
                      reg5447 <= $signed($signed($signed((forvar5106 > reg5343))));
                    end
                  reg5449 <= $signed((((reg4879 == forvar5314) << reg4589[(2'h2):(2'h2)]) ?
                      ((reg4599 != reg5223) + $signed(reg4964)) : (^~$signed((8'ha7)))));
                  for (forvar5450 = (1'h0); (forvar5450 < (1'h0)); forvar5450 = (forvar5450 + (1'h1)))
                    begin
                      reg5451 <= reg5181[(3'h4):(3'h4)];
                    end
                  reg5452 <= $signed((~$unsigned($unsigned(reg5253))));
                end
            end
        end
      else
        begin
          if ((^{{(forvar4604 ? reg5276 : reg4618)}}))
            begin
              if ($signed(reg4963[(1'h1):(1'h1)]))
                begin
                  for (forvar5349 = (1'h0); (forvar5349 < (2'h3)); forvar5349 = (forvar5349 + (1'h1)))
                    begin
                      reg5350 <= reg5160[(2'h2):(2'h2)];
                    end
                  reg5351 <= (!forvar5088);
                end
              else
                begin
                  if ({({(forvar5064 ? (8'ha7) : reg4577)} >> $signed((reg5014 ?
                          reg5354 : forvar5054)))})
                    begin
                      reg5349 <= ((forvar4781[(3'h6):(2'h3)] >= $signed((-reg4718))) - $signed($unsigned((~&reg4639))));
                      reg5350 <= $unsigned(((reg4793 ? {reg5086} : forvar4806) ?
                          ((8'ha1) <<< $unsigned(reg4871)) : (~^(reg4896 & (8'hae)))));
                    end
                  else
                    begin
                      reg5349 <= reg4622;
                      reg5350 <= reg5362[(1'h0):(1'h0)];
                      reg5351 <= reg4651;
                      reg5352 <= $signed($unsigned({((8'hb2) || reg4973)}));
                    end
                  for (forvar5353 = (1'h0); (forvar5353 < (1'h1)); forvar5353 = (forvar5353 + (1'h1)))
                    begin
                      reg5354 <= (8'haa);
                      reg5355 <= (reg5400[(4'hb):(4'hb)] == $unsigned((-(|(8'ha1)))));
                      reg5356 <= $signed(reg5070[(3'h4):(3'h4)]);
                      reg5357 <= forvar4914;
                    end
                end
            end
          else
            begin
              if ({reg4723[(4'ha):(4'ha)]})
                begin
                  for (forvar5349 = (1'h0); (forvar5349 < (2'h3)); forvar5349 = (forvar5349 + (1'h1)))
                    begin
                      reg5350 <= {$unsigned(reg5321)};
                    end
                  if ($signed(reg4782[(2'h3):(2'h2)]))
                    begin
                      reg5351 <= reg5400;
                      reg5352 <= ({$unsigned((-reg5392))} & ((+(reg4836 ?
                          reg4623 : (8'hb0))) ^ (~&(reg5303 ?
                          reg5447 : reg5025))));
                    end
                  else
                    begin
                      reg5351 <= (+reg5256[(3'h6):(3'h5)]);
                    end
                  for (forvar5353 = (1'h0); (forvar5353 < (1'h1)); forvar5353 = (forvar5353 + (1'h1)))
                    begin
                      reg5354 <= ($signed($unsigned((~|reg4796))) ?
                          (reg4657 ?
                              (~$signed(forvar4645)) : $unsigned((reg5110 ?
                                  (8'h9e) : forvar4636))) : (($unsigned(reg4675) >= (reg4762 ?
                              reg5083 : reg5333)) - $signed((reg5222 - forvar5440))));
                      reg5355 <= $unsigned((|{(reg4780 ? (8'hb3) : reg4666)}));
                      reg5356 <= forvar4607;
                    end
                end
              else
                begin
                  reg5349 <= (forvar4848[(1'h1):(1'h1)] - $unsigned(((forvar4705 <<< reg4930) <= $signed(reg4608))));
                  for (forvar5350 = (1'h0); (forvar5350 < (1'h0)); forvar5350 = (forvar5350 + (1'h1)))
                    begin
                      reg5351 <= ($signed($unsigned($signed(reg5352))) >= (-reg5263));
                      reg5352 <= (~&$signed((~reg4796[(2'h3):(1'h0)])));
                    end
                  for (forvar5353 = (1'h0); (forvar5353 < (2'h2)); forvar5353 = (forvar5353 + (1'h1)))
                    begin
                      reg5354 <= ((reg5158[(1'h0):(1'h0)] - reg4852) - $signed(((~&reg5145) ?
                          $signed(reg5210) : forvar5423)));
                      reg5355 <= (~^reg5258[(2'h3):(2'h2)]);
                      reg5356 <= reg4854;
                      reg5357 <= ($signed($signed((^reg4724))) ?
                          ($signed($unsigned(reg4897)) ?
                              (&reg5213[(3'h4):(1'h1)]) : $signed((forvar4837 ?
                                  (8'ha4) : (8'ha9)))) : reg5111[(2'h2):(1'h0)]);
                    end
                end
              reg5358 <= $unsigned((~^$signed((^~forvar5084))));
              if (((forvar5380 <= ((reg4688 >>> forvar5143) < ((8'ha1) <= reg5200))) == (((^~reg5129) ?
                      $signed(forvar4717) : (~^reg5106)) ?
                  reg4779 : {(reg4767 ? reg5047 : forvar4915)})))
                begin
                  if (({reg4936[(1'h0):(1'h0)]} ?
                      (!$unsigned($unsigned((8'ha1)))) : reg4700))
                    begin
                      reg5359 <= reg5183;
                      reg5360 <= ($unsigned($unsigned($signed(forvar5165))) ?
                          {reg4926} : forvar5350);
                    end
                  else
                    begin
                      reg5359 <= forvar5006;
                      reg5360 <= (forvar4929[(1'h1):(1'h1)] ?
                          reg5156[(4'hc):(1'h1)] : (($unsigned(reg5140) ?
                              (+reg5037) : (8'hba)) ^ ($signed(reg5252) ?
                              (forvar5440 & reg4723) : forvar4777[(2'h2):(1'h0)])));
                      reg5361 <= reg5091;
                      reg5362 <= $signed($signed($unsigned(reg5364)));
                    end
                end
              else
                begin
                  reg5359 <= reg4974[(2'h3):(1'h0)];
                  for (forvar5360 = (1'h0); (forvar5360 < (2'h2)); forvar5360 = (forvar5360 + (1'h1)))
                    begin
                      reg5361 <= {$signed({(-reg5302)})};
                    end
                  for (forvar5362 = (1'h0); (forvar5362 < (2'h3)); forvar5362 = (forvar5362 + (1'h1)))
                    begin
                      reg5363 <= (~^(^~(forvar4849[(3'h5):(3'h4)] <<< reg4964)));
                    end
                end
              for (forvar5364 = (1'h0); (forvar5364 < (1'h1)); forvar5364 = (forvar5364 + (1'h1)))
                begin
                  reg5365 <= {$unsigned((~^wire4798))};
                end
            end
          if ($unsigned((^~reg4850)))
            begin
              if (($unsigned($unsigned((forvar4642 ? reg4748 : reg5008))) ?
                  forvar4962[(2'h2):(2'h2)] : {reg4966}))
                begin
                  for (forvar5366 = (1'h0); (forvar5366 < (1'h0)); forvar5366 = (forvar5366 + (1'h1)))
                    begin
                      reg5367 <= $signed((8'ha1));
                      reg5368 <= reg4613[(3'h4):(2'h2)];
                      reg5369 <= {reg4820};
                    end
                  if ($signed($signed(reg4845)))
                    begin
                      reg5370 <= (reg4853[(3'h5):(2'h2)] ?
                          {((reg4907 ?
                                  forvar4967 : forvar5011) ^ (8'hb7))} : (~&((reg4584 > reg4780) && (reg4933 << reg4670))));
                    end
                  else
                    begin
                      reg5370 <= $unsigned((&{forvar5091}));
                      reg5371 <= reg5033;
                    end
                  if (($unsigned($signed((reg5133 < reg5339))) ?
                      {(8'hb4)} : ((^(8'ha6)) ?
                          $signed((reg4768 >= reg5373)) : ((reg4881 <= (8'h9d)) ?
                              $unsigned((8'h9c)) : $signed(reg4788)))))
                    begin
                      reg5372 <= ((forvar5217[(2'h3):(2'h2)] < (+$signed(reg5430))) ?
                          $signed(reg4614[(2'h3):(2'h3)]) : $unsigned($signed(forvar4741[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg5372 <= $signed((($unsigned(reg5317) ?
                          ((8'ha3) ?
                              reg5378 : forvar4588) : forvar5350[(1'h0):(1'h0)]) >> reg4607[(2'h3):(1'h0)]));
                      reg5373 <= reg4902;
                      reg5374 <= (((^~(reg4844 ? forvar4755 : reg4905)) ?
                          (((8'hb3) >= wire4574) < (~^forvar4989)) : forvar4789) & (reg5000[(3'h5):(1'h0)] & (8'hb3)));
                    end
                end
              else
                begin
                  if ($unsigned(reg4848))
                    begin
                      reg5366 <= ($signed(((+forvar5171) ?
                          $signed((8'ha8)) : reg4927)) * (~&$signed({reg5319})));
                      reg5367 <= reg4998;
                      reg5368 <= $signed($signed(reg5150[(4'ha):(2'h3)]));
                    end
                  else
                    begin
                      reg5366 <= ((($signed((8'hb1)) ?
                          ((8'hb3) ? forvar4815 : forvar4779) : (forvar5270 ?
                              reg4875 : reg5202)) != ($signed((8'hb7)) ?
                          reg5188 : reg4626[(2'h2):(2'h2)])) ~^ ($signed($signed(reg5301)) ?
                          ((reg4885 != forvar5143) ?
                              reg5168 : $signed((8'ha0))) : (reg4749 >> {reg4629})));
                    end
                  for (forvar5369 = (1'h0); (forvar5369 < (2'h3)); forvar5369 = (forvar5369 + (1'h1)))
                    begin
                      reg5370 <= $signed((reg5112 ~^ reg4718[(3'h7):(3'h4)]));
                      reg5371 <= (($signed((reg5184 ?
                          (8'ha7) : forvar5011)) < ((|forvar4876) < (-(8'hae)))) >= reg5020[(2'h2):(1'h0)]);
                    end
                  for (forvar5372 = (1'h0); (forvar5372 < (2'h3)); forvar5372 = (forvar5372 + (1'h1)))
                    begin
                      reg5373 <= (!(({reg5264} ?
                              $signed(reg5042) : (wire5195 != (8'hac))) ?
                          reg4584 : reg4936[(1'h0):(1'h0)]));
                      reg5374 <= $unsigned((&$signed((~|(8'ha1)))));
                      reg5375 <= forvar4579[(3'h4):(1'h0)];
                      reg5376 <= $unsigned($unsigned((~^(reg4948 + reg4922))));
                    end
                end
              reg5377 <= {{$unsigned((forvar5270 ? forvar4879 : reg5375))}};
              for (forvar5378 = (1'h0); (forvar5378 < (1'h0)); forvar5378 = (forvar5378 + (1'h1)))
                begin
                  for (forvar5379 = (1'h0); (forvar5379 < (2'h2)); forvar5379 = (forvar5379 + (1'h1)))
                    begin
                      reg5380 <= $signed(reg5120[(1'h0):(1'h0)]);
                      reg5381 <= $signed((~^forvar4592[(3'h5):(3'h5)]));
                    end
                end
              for (forvar5382 = (1'h0); (forvar5382 < (2'h2)); forvar5382 = (forvar5382 + (1'h1)))
                begin
                  for (forvar5383 = (1'h0); (forvar5383 < (1'h0)); forvar5383 = (forvar5383 + (1'h1)))
                    begin
                      reg5384 <= $signed((+$unsigned({(8'had)})));
                      reg5385 <= reg4861;
                    end
                  reg5386 <= ($signed((~(8'hb9))) ?
                      (~$signed((^(8'ha5)))) : $signed((8'hb2)));
                  for (forvar5387 = (1'h0); (forvar5387 < (1'h0)); forvar5387 = (forvar5387 + (1'h1)))
                    begin
                      reg5388 <= $signed((reg5430[(2'h2):(2'h2)] * wire4799));
                      reg5389 <= (|((-(reg5142 - (8'haa))) ?
                          $signed($unsigned(reg4997)) : wire5195[(4'hb):(2'h2)]));
                      reg5390 <= (reg4973[(2'h2):(1'h1)] & (($unsigned(forvar5157) ?
                              (reg4630 >= forvar5165) : (~forvar5189)) ?
                          (~forvar5064) : (|forvar4766)));
                    end
                  for (forvar5391 = (1'h0); (forvar5391 < (2'h2)); forvar5391 = (forvar5391 + (1'h1)))
                    begin
                      reg5392 <= {$unsigned(reg5011)};
                      reg5393 <= (~|$signed($signed(reg4800)));
                      reg5394 <= $unsigned(((8'hba) ?
                          reg5445[(2'h3):(1'h0)] : (8'h9e)));
                      reg5395 <= reg5096;
                    end
                end
            end
          else
            begin
              for (forvar5366 = (1'h0); (forvar5366 < (2'h3)); forvar5366 = (forvar5366 + (1'h1)))
                begin
                  if ($signed(reg4753[(4'hc):(3'h4)]))
                    begin
                      reg5367 <= {((~|{(8'haf)}) ?
                              (reg4973[(2'h2):(2'h2)] ?
                                  (forvar4712 ^ reg4739) : (forvar4779 ?
                                      reg4600 : reg5263)) : reg5287)};
                      reg5368 <= ($signed(reg4912) ?
                          $signed((+(8'ha8))) : ($signed((reg4725 ?
                                  reg4946 : reg5017)) ?
                              reg5055 : $unsigned(reg4685[(1'h0):(1'h0)])));
                      reg5369 <= ((^((+forvar5435) ? (8'h9f) : (+reg5303))) ?
                          (forvar5435[(2'h2):(1'h1)] <= forvar5148) : $signed(reg4642[(4'ha):(4'h8)]));
                    end
                  else
                    begin
                      reg5367 <= reg4892[(1'h0):(1'h0)];
                    end
                  if ($signed(reg4645[(3'h7):(2'h3)]))
                    begin
                      reg5370 <= reg5023;
                      reg5371 <= (|reg4715);
                      reg5372 <= ((-$signed($unsigned(reg5023))) ^ reg5159[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg5370 <= (8'ha9);
                    end
                  for (forvar5373 = (1'h0); (forvar5373 < (1'h1)); forvar5373 = (forvar5373 + (1'h1)))
                    begin
                      reg5374 <= (($unsigned($signed(reg5443)) ?
                          $unsigned({reg4825}) : reg4609[(3'h7):(2'h3)]) >>> forvar4911[(1'h0):(1'h0)]);
                    end
                end
              for (forvar5375 = (1'h0); (forvar5375 < (1'h0)); forvar5375 = (forvar5375 + (1'h1)))
                begin
                  if ((&(reg4581[(2'h3):(2'h2)] ?
                      $signed($signed(reg4597)) : reg4783)))
                    begin
                      reg5376 <= $unsigned((!(reg4965[(3'h4):(1'h0)] ?
                          {(8'ha0)} : (reg4912 ? reg4713 : reg5074))));
                      reg5377 <= reg5299;
                      reg5378 <= ((({reg4757} | (8'ha5)) ?
                          $signed(reg5390) : ((reg4863 ? (8'hb2) : forvar4578) ?
                              (~^forvar5029) : (|forvar5005))) <= ({{forvar5362}} & {(reg5103 == reg4767)}));
                      reg5379 <= {(($unsigned(reg5369) != reg4834[(2'h2):(2'h2)]) >= ($unsigned(reg5040) ?
                              (^reg5187) : reg4905[(1'h1):(1'h1)]))};
                    end
                  else
                    begin
                      reg5376 <= (($signed({reg5040}) ?
                          ($signed(reg4600) ?
                              reg4745[(3'h5):(3'h4)] : reg4664[(4'hf):(4'hb)]) : reg5241[(4'hd):(4'hb)]) != (reg4729 - ((&forvar4864) - reg5397[(1'h0):(1'h0)])));
                      reg5377 <= $signed((8'hb7));
                    end
                  for (forvar5380 = (1'h0); (forvar5380 < (2'h2)); forvar5380 = (forvar5380 + (1'h1)))
                    begin
                      reg5381 <= reg5342;
                      reg5382 <= $unsigned((&$signed(forvar5048)));
                      reg5383 <= $unsigned($signed($signed(((8'hb5) - forvar5285))));
                    end
                  reg5384 <= $unsigned($unsigned(((+reg4928) >= (^reg4859))));
                  reg5385 <= ($unsigned($signed((forvar5068 < forvar5423))) - ({reg5145} ?
                      $unsigned((reg5249 != (8'ha3))) : $signed((reg5179 ^~ reg5439))));
                end
            end
          if ((($signed($signed(forvar5307)) ?
                  {(~reg4989)} : ((reg5209 ? forvar5114 : reg5009) + (reg5349 ?
                      forvar4617 : reg4942))) ?
              reg4679 : ($signed((reg5367 ?
                  reg4848 : forvar4609)) <= forvar5341[(2'h2):(1'h1)])))
            begin
              for (forvar5396 = (1'h0); (forvar5396 < (2'h2)); forvar5396 = (forvar5396 + (1'h1)))
                begin
                  reg5397 <= reg4728[(1'h0):(1'h0)];
                  for (forvar5398 = (1'h0); (forvar5398 < (2'h3)); forvar5398 = (forvar5398 + (1'h1)))
                    begin
                      reg5399 <= reg4768;
                    end
                end
            end
          else
            begin
              for (forvar5396 = (1'h0); (forvar5396 < (2'h3)); forvar5396 = (forvar5396 + (1'h1)))
                begin
                  reg5397 <= reg4871[(4'h8):(2'h3)];
                end
            end
        end
      for (forvar5453 = (1'h0); (forvar5453 < (2'h3)); forvar5453 = (forvar5453 + (1'h1)))
        begin
          for (forvar5454 = (1'h0); (forvar5454 < (2'h3)); forvar5454 = (forvar5454 + (1'h1)))
            begin
              for (forvar5455 = (1'h0); (forvar5455 < (1'h0)); forvar5455 = (forvar5455 + (1'h1)))
                begin
                  if ({$signed(reg4709[(4'hd):(3'h7)])})
                    begin
                      reg5456 <= (reg5269 ?
                          $signed($unsigned((forvar5396 ?
                              forvar4923 : reg5021))) : (!((reg4912 + reg4830) ?
                              (8'ha3) : reg5209[(2'h3):(2'h3)])));
                      reg5457 <= {(^$signed($signed(reg5018)))};
                    end
                  else
                    begin
                      reg5456 <= (|reg5321[(3'h5):(2'h2)]);
                    end
                  for (forvar5458 = (1'h0); (forvar5458 < (1'h0)); forvar5458 = (forvar5458 + (1'h1)))
                    begin
                      reg5459 <= forvar5301[(4'hb):(2'h2)];
                    end
                  for (forvar5460 = (1'h0); (forvar5460 < (2'h3)); forvar5460 = (forvar5460 + (1'h1)))
                    begin
                      reg5461 <= $signed({{$unsigned(reg4746)}});
                      reg5462 <= reg4910[(2'h2):(1'h1)];
                      reg5463 <= (reg4954 || $unsigned((reg4774 << (~|forvar5187))));
                    end
                  reg5464 <= reg4691[(1'h0):(1'h0)];
                end
              reg5465 <= ((~reg5311) ?
                  $unsigned($unsigned(reg5317)) : $unsigned({$signed((8'hb3))}));
              if (((forvar5341 ^~ (~|(~|reg5447))) >= ((&forvar4819[(2'h3):(1'h1)]) ?
                  $unsigned((reg5136 ~^ reg4790)) : ($signed(reg5058) <<< (reg5167 ?
                      (8'h9e) : forvar5353)))))
                begin
                  for (forvar5466 = (1'h0); (forvar5466 < (1'h1)); forvar5466 = (forvar5466 + (1'h1)))
                    begin
                      reg5467 <= ((reg5429 > $signed({reg5037})) ?
                          $unsigned(($unsigned((8'haf)) ?
                              (reg4812 ?
                                  (8'hab) : reg5020) : reg5280)) : reg4982);
                      reg5468 <= $signed((reg4769[(2'h3):(1'h1)] < ($signed(reg5446) ?
                          $unsigned(reg5377) : (!(8'hb3)))));
                    end
                end
              else
                begin
                  reg5466 <= forvar4616;
                  for (forvar5467 = (1'h0); (forvar5467 < (2'h2)); forvar5467 = (forvar5467 + (1'h1)))
                    begin
                      reg5468 <= (&$signed((~&(forvar5171 ?
                          reg5259 : reg4822))));
                      reg5469 <= ($signed(($unsigned(reg5283) >= $unsigned(forvar5398))) | reg4868);
                      reg5470 <= reg5205[(3'h7):(3'h4)];
                      reg5471 <= reg5384;
                    end
                  for (forvar5472 = (1'h0); (forvar5472 < (1'h1)); forvar5472 = (forvar5472 + (1'h1)))
                    begin
                      reg5473 <= $unsigned((($signed(reg4928) && (forvar4802 ?
                              reg5159 : forvar4584)) ?
                          $unsigned((reg4942 ^ reg5202)) : (~|$signed(reg4722))));
                    end
                end
            end
          for (forvar5474 = (1'h0); (forvar5474 < (2'h2)); forvar5474 = (forvar5474 + (1'h1)))
            begin
              if (reg5174[(4'hb):(3'h6)])
                begin
                  reg5475 <= $unsigned(forvar5245[(3'h5):(2'h2)]);
                  for (forvar5476 = (1'h0); (forvar5476 < (2'h3)); forvar5476 = (forvar5476 + (1'h1)))
                    begin
                      reg5477 <= {(forvar4763 ?
                              (^(reg4861 ?
                                  reg5411 : (8'h9d))) : $unsigned((~&reg4926)))};
                      reg5478 <= reg4741;
                      reg5479 <= {$unsigned({$unsigned(reg5125)})};
                    end
                end
              else
                begin
                  reg5475 <= $unsigned(({((8'hb9) ? (8'ha1) : reg5104)} ?
                      {((8'haa) ? reg4621 : reg5391)} : forvar5231));
                  for (forvar5476 = (1'h0); (forvar5476 < (1'h0)); forvar5476 = (forvar5476 + (1'h1)))
                    begin
                      reg5477 <= forvar5117[(2'h3):(2'h3)];
                    end
                end
              if (reg5250)
                begin
                  for (forvar5480 = (1'h0); (forvar5480 < (1'h0)); forvar5480 = (forvar5480 + (1'h1)))
                    begin
                      reg5481 <= reg5122[(1'h1):(1'h0)];
                      reg5482 <= $signed((((~reg4929) ?
                          (forvar5423 ^~ reg5427) : (reg4658 - reg5250)) < (~|reg4753[(1'h0):(1'h0)])));
                      reg5483 <= reg4847[(1'h1):(1'h0)];
                    end
                  if ({((&$unsigned(reg4901)) >> $unsigned($unsigned(reg4854)))})
                    begin
                      reg5484 <= (~&(!(^(forvar4910 ? (8'hb4) : reg5478))));
                      reg5485 <= reg5141;
                    end
                  else
                    begin
                      reg5484 <= forvar4674[(3'h7):(3'h6)];
                      reg5485 <= $unsigned({(^(reg5029 ^~ reg4920))});
                    end
                  if ($signed(((((8'hb1) != forvar4581) ?
                          reg5317[(4'hb):(4'ha)] : ((8'hb8) & reg5305)) ?
                      forvar4696 : (reg4955 >= (reg5412 >= (8'ha1))))))
                    begin
                      reg5486 <= (reg5152[(4'he):(3'h4)] ?
                          $signed(reg4742) : (reg5357 ^~ (~|reg4997[(1'h0):(1'h0)])));
                      reg5487 <= (($unsigned(forvar4737) ?
                          (forvar4610 ?
                              reg5324[(1'h1):(1'h1)] : (&reg5060)) : $unsigned((forvar5404 ?
                              reg5231 : reg4894))) < reg5208);
                      reg5488 <= $unsigned((^(~|$signed(forvar4840))));
                      reg5489 <= $unsigned(($signed((forvar5369 ?
                          reg4869 : reg4832)) ^~ reg4870));
                    end
                  else
                    begin
                      reg5486 <= (reg5002 ?
                          $signed(($signed(reg4909) ?
                              reg4903 : (reg5287 ?
                                  reg4908 : forvar4840))) : $unsigned((~^forvar5008[(4'h8):(3'h7)])));
                      reg5487 <= (reg4896[(4'h9):(3'h5)] << reg5004);
                      reg5488 <= (8'ha6);
                    end
                  if ($signed(($unsigned((forvar4745 | reg4656)) && $unsigned(reg5360[(4'hc):(3'h4)]))))
                    begin
                      reg5490 <= {$unsigned(reg5213[(3'h7):(3'h4)])};
                      reg5491 <= $unsigned((forvar5171 ?
                          reg5355 : $signed(reg5324)));
                      reg5492 <= (((!$unsigned((8'hb0))) >>> (~&$unsigned((8'hac)))) ?
                          forvar5467[(1'h0):(1'h0)] : (((reg4761 ?
                                  reg4915 : reg5466) ?
                              reg4699[(3'h5):(2'h3)] : reg4863) <<< (reg4730 ?
                              (reg5365 * (8'h9d)) : (reg5122 ?
                                  (8'ha7) : (8'hb7)))));
                    end
                  else
                    begin
                      reg5490 <= $signed((~&((forvar5049 | (8'hba)) & $unsigned(reg4836))));
                    end
                end
              else
                begin
                  if ($unsigned(reg4934))
                    begin
                      reg5480 <= ((reg4860[(3'h7):(3'h4)] ?
                              ((reg5252 ^~ reg5337) != $unsigned(forvar5039)) : (^~(^~reg5115))) ?
                          {reg5287} : ((8'ha9) ?
                              ({forvar4952} * (reg5142 ?
                                  forvar4659 : reg4834)) : $unsigned($unsigned(forvar4970))));
                      reg5481 <= wire4798[(1'h0):(1'h0)];
                      reg5482 <= reg5152[(3'h5):(1'h0)];
                      reg5483 <= reg4744;
                    end
                  else
                    begin
                      reg5480 <= reg5233[(4'hb):(4'h8)];
                      reg5481 <= $signed((((forvar4604 || reg4869) <<< {forvar4712}) ?
                          $unsigned($unsigned(forvar4996)) : reg5351));
                      reg5482 <= (-reg4721[(1'h1):(1'h0)]);
                    end
                  for (forvar5484 = (1'h0); (forvar5484 < (1'h1)); forvar5484 = (forvar5484 + (1'h1)))
                    begin
                      reg5485 <= $signed((forvar5350 << (forvar5126[(4'h9):(3'h7)] <= (!reg5079))));
                    end
                  reg5486 <= $signed($unsigned((forvar4795 ~^ ((8'haa) >> (8'hb9)))));
                end
            end
          for (forvar5493 = (1'h0); (forvar5493 < (2'h2)); forvar5493 = (forvar5493 + (1'h1)))
            begin
              reg5494 <= (reg4701[(3'h7):(3'h7)] ?
                  $signed(forvar5387) : $signed($unsigned(forvar5109)));
              if (($unsigned($unsigned({(8'h9d)})) ?
                  reg4983 : $unsigned(reg4634)))
                begin
                  if ((reg5184[(3'h7):(3'h5)] ?
                      $unsigned({reg5194}) : forvar4593[(1'h1):(1'h0)]))
                    begin
                      reg5495 <= ((+(~(&reg4852))) ?
                          reg4752[(4'h8):(2'h3)] : ($unsigned($signed(reg4952)) >= $unsigned((reg4691 ?
                              forvar4759 : reg5219))));
                    end
                  else
                    begin
                      reg5495 <= (!$unsigned(((~&reg4611) ^~ (&forvar4759))));
                      reg5496 <= reg5206[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  if ((!$unsigned(((^forvar4975) >>> reg5394))))
                    begin
                      reg5495 <= (((reg5347[(1'h1):(1'h1)] >> reg5301[(2'h3):(2'h2)]) < reg4960[(2'h2):(1'h1)]) < forvar5051[(4'h8):(4'h8)]);
                      reg5496 <= ((~&$unsigned($signed(reg4947))) >>> reg5286[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg5495 <= ($unsigned({(forvar4815 ?
                                  forvar5051 : reg5412)}) ?
                          reg5238[(2'h2):(1'h0)] : (((^~reg4667) ~^ (reg5187 + reg4916)) ?
                              {reg4848[(1'h1):(1'h1)]} : $signed({reg4850})));
                    end
                  for (forvar5497 = (1'h0); (forvar5497 < (2'h2)); forvar5497 = (forvar5497 + (1'h1)))
                    begin
                      reg5498 <= forvar5284;
                      reg5499 <= ($signed($unsigned(reg5263)) ?
                          {(^~(forvar5355 ?
                                  reg4658 : reg4678))} : (($signed(reg5223) - {reg5365}) >> (forvar4640[(3'h4):(1'h1)] ?
                              (8'ha8) : (forvar4577 * (8'hb9)))));
                      reg5500 <= (reg5357[(2'h3):(1'h1)] ?
                          {($unsigned(reg5494) ^ reg5150)} : ($unsigned((8'ha1)) ?
                              ((forvar5297 <<< (8'h9c)) && reg4929) : {(reg4937 ?
                                      reg5055 : reg4861)}));
                      reg5501 <= forvar5148;
                    end
                  reg5502 <= (|(^{(forvar4988 ? reg4907 : reg4707)}));
                end
              for (forvar5503 = (1'h0); (forvar5503 < (2'h3)); forvar5503 = (forvar5503 + (1'h1)))
                begin
                  if ($signed((^~$signed((^~(8'ha5))))))
                    begin
                      reg5504 <= reg5167;
                    end
                  else
                    begin
                      reg5504 <= (-$signed({(reg5365 ? reg5377 : reg4980)}));
                    end
                end
            end
        end
    end
  module5505 modinst6863 (.wire5507(forvar5454), .clk(clk), .wire5509(reg4993), .wire5506(forvar5231), .wire5508(reg4668), .wire5510(reg4747), .y(wire6862));
  assign wire6864 = {((forvar5231[(2'h3):(1'h0)] & (forvar5054 <= reg5149)) >> reg5329[(1'h1):(1'h0)])};
  assign wire6865 = (reg5239 != reg5269);
  assign wire6866 = (({{reg4917}} && $signed(reg5448[(3'h7):(3'h7)])) ?
                        $signed(((forvar4578 <<< forvar4824) * reg4680[(4'h9):(3'h6)])) : (reg4670[(2'h2):(1'h1)] * (reg5219 ?
                            $unsigned((8'had)) : reg5378)));
  always
    @(posedge clk) begin
      for (forvar6867 = (1'h0); (forvar6867 < (1'h0)); forvar6867 = (forvar6867 + (1'h1)))
        begin
          reg6868 <= reg4580;
          if ((((~&{reg4863}) ?
              reg4909[(3'h6):(2'h3)] : ($unsigned(reg5378) * $signed((8'hb6)))) * $signed((((8'ha5) ?
              (8'hb3) : forvar5117) >> (reg4700 ? reg4757 : (8'hb6))))))
            begin
              if (reg4960[(1'h1):(1'h1)])
                begin
                  for (forvar6869 = (1'h0); (forvar6869 < (2'h2)); forvar6869 = (forvar6869 + (1'h1)))
                    begin
                      reg6870 <= ($signed(($signed(reg4639) ?
                              $unsigned((8'hb4)) : ((8'h9e) ?
                                  reg4638 : reg4903))) ?
                          $signed(((~|(8'haa)) == (reg4733 ?
                              wire4799 : forvar4624))) : $signed({forvar5108}));
                      reg6871 <= (^~{(~&reg5463[(2'h3):(1'h1)])});
                      reg6872 <= $signed($unsigned($unsigned((~|forvar5043))));
                      reg6873 <= $signed(({$signed(reg5325)} ^ ((reg4895 >>> reg4985) ?
                          reg5192[(1'h0):(1'h0)] : forvar4848)));
                    end
                  for (forvar6874 = (1'h0); (forvar6874 < (2'h3)); forvar6874 = (forvar6874 + (1'h1)))
                    begin
                      reg6875 <= (reg5114 == $unsigned($signed(reg5089[(2'h2):(1'h1)])));
                      reg6876 <= $signed({reg5244});
                      reg6877 <= (forvar5062[(1'h0):(1'h0)] <= $signed((|(reg4932 ?
                          reg5275 : wire5197))));
                    end
                end
              else
                begin
                  for (forvar6869 = (1'h0); (forvar6869 < (2'h3)); forvar6869 = (forvar6869 + (1'h1)))
                    begin
                      reg6870 <= (!reg4630[(1'h1):(1'h0)]);
                      reg6871 <= $unsigned((+reg5159[(3'h7):(3'h4)]));
                      reg6872 <= (8'hb9);
                    end
                  reg6873 <= (reg5181[(1'h0):(1'h0)] <= (+$signed((reg5373 * reg5180))));
                end
              reg6878 <= forvar4715[(3'h5):(3'h4)];
              if (($unsigned($unsigned(reg4946)) || $unsigned((8'hae))))
                begin
                  reg6879 <= reg4831[(3'h6):(2'h2)];
                  for (forvar6880 = (1'h0); (forvar6880 < (1'h0)); forvar6880 = (forvar6880 + (1'h1)))
                    begin
                      reg6881 <= reg4909[(2'h2):(1'h0)];
                    end
                  for (forvar6882 = (1'h0); (forvar6882 < (2'h2)); forvar6882 = (forvar6882 + (1'h1)))
                    begin
                      reg6883 <= reg5155[(3'h4):(1'h0)];
                      reg6884 <= (({(~|reg5444)} ~^ forvar5440[(3'h6):(2'h3)]) ?
                          {reg4794} : (reg4830 ?
                              ((^reg5029) ?
                                  (8'hab) : reg5106[(1'h1):(1'h0)]) : $signed(reg5379)));
                    end
                end
              else
                begin
                  if ((8'h9e))
                    begin
                      reg6879 <= $unsigned((|$unsigned($unsigned((8'h9c)))));
                      reg6880 <= (reg5448[(3'h4):(1'h1)] ?
                          ((+(-forvar5363)) ?
                              $signed((reg5345 || forvar5472)) : $signed($unsigned(forvar4795))) : forvar4839);
                      reg6881 <= (^$signed(((reg4604 >= reg4591) ?
                          (reg4719 ? reg5118 : (8'hb9)) : $signed(reg4887))));
                      reg6882 <= (reg5299[(3'h5):(1'h1)] ?
                          $unsigned($unsigned((~&reg5176))) : $signed(reg4974));
                    end
                  else
                    begin
                      reg6879 <= $unsigned($unsigned((+(-reg4786))));
                      reg6880 <= ({$unsigned(reg4771)} ?
                          $signed(forvar4977[(3'h4):(3'h4)]) : reg4775);
                    end
                end
              if (reg5495[(1'h1):(1'h1)])
                begin
                  for (forvar6885 = (1'h0); (forvar6885 < (2'h3)); forvar6885 = (forvar6885 + (1'h1)))
                    begin
                      reg6886 <= reg4964[(2'h2):(2'h2)];
                      reg6887 <= (reg5496 - ((8'h9c) < $signed((^~forvar5460))));
                    end
                  if ((8'hb2))
                    begin
                      reg6888 <= (8'hba);
                      reg6889 <= ((~&((!reg4879) ?
                          (reg5215 == (8'ha1)) : (|forvar4755))) | reg4964[(2'h3):(2'h2)]);
                      reg6890 <= {$signed(($unsigned(reg4760) ?
                              (-reg4664) : (forvar4962 ? reg5465 : reg5486)))};
                      reg6891 <= ((8'ha4) ?
                          (reg4818[(3'h4):(3'h4)] ?
                              ((wire6864 ? forvar4843 : forvar4610) ?
                                  $unsigned(reg4781) : (&(8'hb4))) : reg4989[(3'h7):(3'h7)]) : (($unsigned(reg4820) > (reg5237 <= reg4903)) & $unsigned((-reg5298))));
                    end
                  else
                    begin
                      reg6888 <= reg5488;
                    end
                  for (forvar6892 = (1'h0); (forvar6892 < (2'h2)); forvar6892 = (forvar6892 + (1'h1)))
                    begin
                      reg6893 <= (({(8'h9f)} ?
                          (8'hb7) : $unsigned(((8'hb2) ?
                              reg5118 : (8'hab)))) < {forvar4694[(4'h8):(3'h4)]});
                      reg6894 <= forvar5048[(2'h3):(1'h0)];
                    end
                end
              else
                begin
                  reg6885 <= $unsigned(({$signed((8'hb3))} - ((|forvar4591) <<< (reg4774 || (8'ha9)))));
                  for (forvar6886 = (1'h0); (forvar6886 < (1'h1)); forvar6886 = (forvar6886 + (1'h1)))
                    begin
                      reg6887 <= wire4799;
                      reg6888 <= forvar5266[(2'h3):(1'h0)];
                      reg6889 <= $unsigned($signed({$unsigned(forvar5143)}));
                    end
                  for (forvar6890 = (1'h0); (forvar6890 < (2'h3)); forvar6890 = (forvar6890 + (1'h1)))
                    begin
                      reg6891 <= {$unsigned(forvar5403[(1'h0):(1'h0)])};
                    end
                  for (forvar6892 = (1'h0); (forvar6892 < (1'h1)); forvar6892 = (forvar6892 + (1'h1)))
                    begin
                      reg6893 <= $unsigned(($unsigned((8'ha1)) ?
                          {(&reg4985)} : $signed((8'h9f))));
                      reg6894 <= reg4642;
                      reg6895 <= $unsigned($signed({$unsigned(reg5080)}));
                    end
                end
            end
          else
            begin
              for (forvar6869 = (1'h0); (forvar6869 < (1'h1)); forvar6869 = (forvar6869 + (1'h1)))
                begin
                  reg6870 <= reg5346[(1'h0):(1'h0)];
                end
              for (forvar6871 = (1'h0); (forvar6871 < (2'h2)); forvar6871 = (forvar6871 + (1'h1)))
                begin
                  if ((~^(reg4904 ~^ {(~&reg4973)})))
                    begin
                      reg6872 <= $signed(($unsigned((reg5208 ?
                              forvar4965 : reg5483)) ?
                          reg5164 : (~reg4933[(4'h8):(2'h2)])));
                      reg6873 <= (~|reg5116[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg6872 <= {(~&reg5074[(4'ha):(3'h4)])};
                      reg6873 <= reg4972;
                    end
                  if ((~&(-reg4779[(1'h0):(1'h0)])))
                    begin
                      reg6874 <= (~reg4983);
                      reg6875 <= reg4864[(4'hd):(3'h7)];
                      reg6876 <= reg5078;
                    end
                  else
                    begin
                      reg6874 <= (reg4852[(4'ha):(4'h9)] ?
                          $unsigned(((forvar5440 | reg4999) > $unsigned(reg4586))) : reg4810);
                      reg6875 <= (~^(forvar4908 ^ {forvar4698}));
                    end
                  for (forvar6877 = (1'h0); (forvar6877 < (2'h3)); forvar6877 = (forvar6877 + (1'h1)))
                    begin
                      reg6878 <= reg5305;
                    end
                end
              if ((((-reg5189[(4'h9):(4'h9)]) ?
                      {{reg5345}} : {(forvar4727 ? (8'h9c) : reg5216)}) ?
                  forvar4869 : forvar4850))
                begin
                  reg6879 <= reg4986;
                  reg6880 <= (~$unsigned($unsigned({reg4608})));
                  if ((reg4755[(1'h1):(1'h0)] ? (~|reg6868) : (~reg4907)))
                    begin
                      reg6881 <= $signed((~|$signed({reg5359})));
                    end
                  else
                    begin
                      reg6881 <= reg4927[(1'h1):(1'h1)];
                      reg6882 <= (+$unsigned(($unsigned(reg4937) ?
                          (reg5278 ?
                              reg4608 : forvar5048) : $unsigned((8'hb8)))));
                    end
                  if (forvar5059[(1'h0):(1'h0)])
                    begin
                      reg6883 <= reg5303;
                    end
                  else
                    begin
                      reg6883 <= (&($unsigned(forvar4642) ?
                          {(reg4822 ? (8'hb0) : reg5107)} : {forvar5340}));
                      reg6884 <= (|(forvar6892[(1'h1):(1'h0)] ?
                          (~^$signed(reg4885)) : (reg5019[(4'he):(1'h0)] ?
                              reg5499[(2'h3):(2'h3)] : (forvar5020 < reg5259))));
                      reg6885 <= $unsigned(({(forvar5423 && forvar5206)} & ($unsigned(reg4736) - (forvar5326 + reg5080))));
                      reg6886 <= {$signed(reg5421)};
                    end
                end
              else
                begin
                  if (reg4950)
                    begin
                      reg6879 <= $unsigned(forvar4918);
                      reg6880 <= $signed(($unsigned($unsigned(reg4803)) ?
                          $signed({(8'ha3)}) : reg4607));
                      reg6881 <= ({reg5287} ?
                          $unsigned((~^$unsigned(forvar4640))) : $signed((forvar5011 ?
                              reg5311[(3'h7):(3'h4)] : (^~reg5329))));
                    end
                  else
                    begin
                      reg6879 <= {(reg5130[(3'h7):(3'h7)] < (~{reg4755}))};
                    end
                end
              if (reg5124)
                begin
                  reg6887 <= (($signed((reg4772 && forvar4698)) <= reg4641[(4'h8):(1'h0)]) ?
                      (!$signed((reg5083 ?
                          forvar4674 : reg5142))) : $unsigned((+$signed((8'ha4)))));
                  if (reg5189[(4'ha):(2'h2)])
                    begin
                      reg6888 <= ($unsigned($signed({reg4821})) ?
                          (+reg4637[(1'h0):(1'h0)]) : (forvar4652[(2'h2):(2'h2)] ~^ (((8'hb2) <<< (8'hb3)) ?
                              $unsigned(reg4840) : $unsigned(forvar5292))));
                      reg6889 <= {(!((reg5291 != reg5209) ?
                              forvar4929 : reg4757))};
                      reg6890 <= (reg4848[(2'h2):(2'h2)] || $unsigned(($signed(forvar5387) ?
                          reg5291 : $unsigned(reg5437))));
                    end
                  else
                    begin
                      reg6888 <= (&$unsigned(($unsigned((8'hae)) ?
                          (forvar5420 ~^ reg5342) : $unsigned(forvar4696))));
                      reg6889 <= forvar4869;
                      reg6890 <= forvar4738;
                      reg6891 <= (reg4684[(4'h8):(3'h5)] || reg6895[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  reg6887 <= (^(~|(~&(&reg4715))));
                end
            end
        end
      reg6896 <= reg5385[(4'hd):(4'h8)];
      if ($unsigned(reg5023[(4'ha):(4'h9)]))
        begin
          for (forvar6897 = (1'h0); (forvar6897 < (2'h3)); forvar6897 = (forvar6897 + (1'h1)))
            begin
              reg6898 <= (~&reg5267[(4'hd):(4'hd)]);
            end
        end
      else
        begin
          for (forvar6897 = (1'h0); (forvar6897 < (1'h1)); forvar6897 = (forvar6897 + (1'h1)))
            begin
              for (forvar6898 = (1'h0); (forvar6898 < (2'h2)); forvar6898 = (forvar6898 + (1'h1)))
                begin
                  for (forvar6899 = (1'h0); (forvar6899 < (2'h2)); forvar6899 = (forvar6899 + (1'h1)))
                    begin
                      reg6900 <= {$unsigned($unsigned($signed(forvar5075)))};
                      reg6901 <= forvar4763[(4'hb):(1'h0)];
                      reg6902 <= $unsigned({((forvar4604 ? reg5444 : reg5042) ?
                              $signed(reg5038) : (reg5156 | (8'hb6)))});
                    end
                  reg6903 <= $signed((&(forvar5068 ?
                      (reg4782 ? forvar4801 : reg5267) : $signed(reg4942))));
                  reg6904 <= $unsigned($unsigned(reg5258));
                  for (forvar6905 = (1'h0); (forvar6905 < (1'h0)); forvar6905 = (forvar6905 + (1'h1)))
                    begin
                      reg6906 <= ($signed((forvar4996 ?
                              (wire5196 ? reg4699 : reg4726) : {forvar5472})) ?
                          $signed(reg4840[(4'ha):(3'h7)]) : reg5146[(2'h3):(1'h1)]);
                      reg6907 <= reg5410;
                      reg6908 <= (8'ha4);
                    end
                end
              for (forvar6909 = (1'h0); (forvar6909 < (2'h3)); forvar6909 = (forvar6909 + (1'h1)))
                begin
                  for (forvar6910 = (1'h0); (forvar6910 < (1'h0)); forvar6910 = (forvar6910 + (1'h1)))
                    begin
                      reg6911 <= $unsigned(reg4834);
                      reg6912 <= $unsigned((8'ha9));
                    end
                  for (forvar6913 = (1'h0); (forvar6913 < (2'h3)); forvar6913 = (forvar6913 + (1'h1)))
                    begin
                      reg6914 <= $signed($unsigned({(8'had)}));
                      reg6915 <= forvar5466;
                      reg6916 <= $unsigned(reg5410[(4'h8):(2'h2)]);
                    end
                end
              reg6917 <= {forvar4819};
              reg6918 <= ((8'ha0) ^ forvar5458);
            end
          for (forvar6919 = (1'h0); (forvar6919 < (2'h2)); forvar6919 = (forvar6919 + (1'h1)))
            begin
              if ((((~|$unsigned(reg4818)) ?
                      reg5057 : $unsigned(forvar5177[(1'h0):(1'h0)])) ?
                  $signed((~^reg5125[(1'h0):(1'h0)])) : $unsigned($unsigned((reg4872 ?
                      forvar4986 : reg4839)))))
                begin
                  for (forvar6920 = (1'h0); (forvar6920 < (2'h2)); forvar6920 = (forvar6920 + (1'h1)))
                    begin
                      reg6921 <= reg5113;
                      reg6922 <= reg4992[(2'h2):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar6920 = (1'h0); (forvar6920 < (1'h0)); forvar6920 = (forvar6920 + (1'h1)))
                    begin
                      reg6921 <= $unsigned(($signed($unsigned(forvar4712)) ?
                          $signed((reg4821 < forvar5043)) : (~(forvar4858 < reg4678))));
                      reg6922 <= $signed((8'hb1));
                      reg6923 <= {($unsigned(reg4961[(3'h6):(1'h1)]) << $unsigned(forvar5398[(1'h1):(1'h1)]))};
                      reg6924 <= reg5325[(2'h3):(2'h3)];
                    end
                  for (forvar6925 = (1'h0); (forvar6925 < (1'h1)); forvar6925 = (forvar6925 + (1'h1)))
                    begin
                      reg6926 <= $signed((8'haf));
                      reg6927 <= (&(((reg4633 ^ forvar5011) <<< {reg5013}) ?
                          (8'hb1) : $signed(reg5053)));
                    end
                end
              for (forvar6928 = (1'h0); (forvar6928 < (1'h1)); forvar6928 = (forvar6928 + (1'h1)))
                begin
                  if (forvar5165)
                    begin
                      reg6929 <= {$signed(forvar5206)};
                      reg6930 <= {(reg4730[(3'h5):(2'h3)] > (~reg4704[(2'h3):(2'h2)]))};
                      reg6931 <= {forvar5085[(4'hb):(3'h5)]};
                    end
                  else
                    begin
                      reg6929 <= ($signed($signed((reg5421 >= reg4684))) < $signed(($signed(reg4883) < reg5111[(4'hc):(3'h7)])));
                      reg6930 <= (($signed($signed(forvar4676)) ?
                          reg5204 : {$unsigned(forvar5270)}) >>> reg5273);
                    end
                end
            end
        end
      for (forvar6932 = (1'h0); (forvar6932 < (1'h0)); forvar6932 = (forvar6932 + (1'h1)))
        begin
          if ($unsigned(wire4799[(1'h0):(1'h0)]))
            begin
              reg6933 <= $unsigned({((forvar4607 == (8'ha5)) < reg5014)});
              for (forvar6934 = (1'h0); (forvar6934 < (2'h3)); forvar6934 = (forvar6934 + (1'h1)))
                begin
                  if ((reg4976[(4'he):(4'he)] ?
                      (reg5434 >> ({reg5083} >= (reg4916 & reg5087))) : $signed(((reg4988 ?
                          forvar5003 : reg4970) < (-reg4822)))))
                    begin
                      reg6935 <= (reg4974[(2'h2):(1'h0)] | (forvar5109 ?
                          (|reg4797) : (~&forvar5398[(3'h4):(3'h4)])));
                      reg6936 <= (+(&$signed((8'ha1))));
                      reg6937 <= $signed((reg5259[(4'h8):(3'h4)] ?
                          $unsigned(reg5001[(4'ha):(3'h6)]) : forvar4694[(4'h8):(3'h4)]));
                    end
                  else
                    begin
                      reg6935 <= reg4784;
                      reg6936 <= reg5365[(4'hb):(4'h9)];
                      reg6937 <= {(~^(+reg5423))};
                    end
                  for (forvar6938 = (1'h0); (forvar6938 < (2'h3)); forvar6938 = (forvar6938 + (1'h1)))
                    begin
                      reg6939 <= $unsigned(forvar4806[(1'h1):(1'h0)]);
                      reg6940 <= reg4746[(3'h4):(1'h0)];
                    end
                end
            end
          else
            begin
              reg6933 <= {(8'ha3)};
              for (forvar6934 = (1'h0); (forvar6934 < (1'h0)); forvar6934 = (forvar6934 + (1'h1)))
                begin
                  reg6935 <= $unsigned(((forvar5059[(2'h2):(2'h2)] ?
                      (reg4764 ? reg6927 : (8'hb2)) : reg5417) - (reg5028 ?
                      ((8'hae) * (8'hb6)) : $unsigned(reg4679))));
                  for (forvar6936 = (1'h0); (forvar6936 < (1'h1)); forvar6936 = (forvar6936 + (1'h1)))
                    begin
                      reg6937 <= ($signed($signed((reg6891 ?
                          reg4973 : reg5296))) ^ ({$unsigned(reg5349)} + ((~|reg5264) ~^ $signed(reg5019))));
                      reg6938 <= ($unsigned((~|(+reg5414))) <= (^($unsigned(reg5161) ~^ (forvar4923 >>> reg5463))));
                      reg6939 <= (|reg5146);
                      reg6940 <= $unsigned((reg4759[(2'h3):(2'h2)] <= (~|(reg4859 ?
                          forvar5200 : reg5093))));
                    end
                  if ($signed((^~(reg5067 ?
                      $signed(reg5277) : (~&forvar5420)))))
                    begin
                      reg6941 <= $signed(reg5096[(3'h4):(2'h2)]);
                      reg6942 <= (((forvar5234 ?
                              ((8'hb5) ?
                                  reg5056 : (8'hb3)) : (reg4898 == reg5444)) ?
                          ($unsigned(reg5359) >> (reg4738 + (8'h9e))) : $unsigned($unsigned(reg4919))) <<< {($unsigned(reg4857) ?
                              reg5364 : ((8'haa) ? reg4718 : reg5134))});
                      reg6943 <= ((^~((reg5012 < reg4912) && reg4950[(3'h6):(3'h4)])) ?
                          (+(&$unsigned(forvar4594))) : ($signed($signed(forvar5248)) ?
                              ((~&reg4770) ?
                                  $signed((8'hb9)) : $signed(forvar5270)) : reg6896[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg6941 <= $signed({$unsigned((~^(8'hb5)))});
                      reg6942 <= (&({(~&reg5457)} ?
                          (wire6866[(2'h2):(2'h2)] == reg4671[(1'h1):(1'h0)]) : ((forvar5019 ?
                              reg5394 : reg5346) != $signed(reg4631))));
                      reg6943 <= reg4767;
                    end
                end
              if ($signed({{((8'ha1) < forvar5360)}}))
                begin
                  for (forvar6944 = (1'h0); (forvar6944 < (1'h0)); forvar6944 = (forvar6944 + (1'h1)))
                    begin
                      reg6945 <= ($signed((~(8'hb2))) ?
                          (~reg4594[(1'h1):(1'h1)]) : ({reg5407} ?
                              $signed((forvar4973 == forvar5376)) : (|((8'hab) * (8'ha5)))));
                      reg6946 <= $unsigned($signed((((8'hb2) >= forvar4995) ?
                          (reg5034 ?
                              reg5129 : forvar5171) : reg5070[(4'h8):(3'h6)])));
                    end
                  if ($unsigned($unsigned(($unsigned((8'hba)) != reg6943))))
                    begin
                      reg6947 <= reg5127[(3'h6):(1'h0)];
                      reg6948 <= (forvar5247 > (-reg5238));
                    end
                  else
                    begin
                      reg6947 <= $signed(reg5329);
                      reg6948 <= $unsigned((-reg5105));
                      reg6949 <= {(($signed(wire4940) ?
                              $signed(reg5152) : $signed(reg6876)) < reg5406)};
                      reg6950 <= reg5110;
                    end
                end
              else
                begin
                  reg6944 <= reg6888;
                end
              reg6951 <= reg5073[(3'h4):(3'h4)];
            end
          for (forvar6952 = (1'h0); (forvar6952 < (1'h0)); forvar6952 = (forvar6952 + (1'h1)))
            begin
              for (forvar6953 = (1'h0); (forvar6953 < (2'h3)); forvar6953 = (forvar6953 + (1'h1)))
                begin
                  for (forvar6954 = (1'h0); (forvar6954 < (2'h3)); forvar6954 = (forvar6954 + (1'h1)))
                    begin
                      reg6955 <= (($unsigned(reg5264[(1'h0):(1'h0)]) < $unsigned({forvar5089})) ~^ (+$unsigned((^reg4688))));
                      reg6956 <= forvar4809[(2'h2):(1'h1)];
                      reg6957 <= (reg6870[(2'h2):(1'h0)] ? reg5055 : reg5316);
                    end
                  for (forvar6958 = (1'h0); (forvar6958 < (2'h2)); forvar6958 = (forvar6958 + (1'h1)))
                    begin
                      reg6959 <= {($unsigned((-reg5092)) == ({reg6918} ?
                              (reg4833 | reg6881) : (reg5357 ?
                                  forvar5001 : wire5195)))};
                      reg6960 <= $unsigned($signed((!reg4892[(3'h4):(2'h2)])));
                      reg6961 <= (reg5429 ?
                          reg4597[(1'h0):(1'h0)] : (((~^forvar5217) ?
                                  $unsigned(reg5154) : (~reg4715)) ?
                              (!((8'hb3) ?
                                  forvar6874 : forvar5261)) : (~&$signed(reg5408))));
                    end
                  if ($signed($unsigned($unsigned({forvar4879}))))
                    begin
                      reg6962 <= $unsigned(reg5445);
                    end
                  else
                    begin
                      reg6962 <= ($unsigned($signed((~^reg4736))) <= {{(forvar4642 ?
                                  reg4769 : forvar4988)}});
                      reg6963 <= forvar5458;
                    end
                end
              for (forvar6964 = (1'h0); (forvar6964 < (1'h0)); forvar6964 = (forvar6964 + (1'h1)))
                begin
                  reg6965 <= $unsigned($unsigned(($unsigned(reg4711) ?
                      (reg5304 >= reg4879) : (~^reg6940))));
                  for (forvar6966 = (1'h0); (forvar6966 < (1'h1)); forvar6966 = (forvar6966 + (1'h1)))
                    begin
                      reg6967 <= forvar5104[(3'h5):(2'h3)];
                      reg6968 <= $signed((-((reg4975 >= reg4846) ?
                          $signed(reg5495) : $unsigned((8'hb4)))));
                      reg6969 <= (^~$signed(reg4955));
                    end
                end
              reg6970 <= reg5413[(4'ha):(3'h4)];
              for (forvar6971 = (1'h0); (forvar6971 < (1'h1)); forvar6971 = (forvar6971 + (1'h1)))
                begin
                  for (forvar6972 = (1'h0); (forvar6972 < (2'h2)); forvar6972 = (forvar6972 + (1'h1)))
                    begin
                      reg6973 <= $signed(($unsigned(forvar4843) <<< $signed((reg4589 ?
                          forvar5165 : reg6876))));
                      reg6974 <= $unsigned(forvar4827);
                      reg6975 <= $signed((-$unsigned(reg6937[(2'h3):(2'h3)])));
                      reg6976 <= $signed((~^$signed(forvar4850)));
                    end
                  for (forvar6977 = (1'h0); (forvar6977 < (1'h1)); forvar6977 = (forvar6977 + (1'h1)))
                    begin
                      reg6978 <= $signed($signed((-$signed(reg5139))));
                      reg6979 <= reg5212;
                      reg6980 <= reg5445;
                    end
                end
            end
          if ((reg4975[(2'h3):(1'h1)] || $signed((8'ha0))))
            begin
              reg6981 <= reg5241[(4'h8):(3'h7)];
            end
          else
            begin
              if ((reg5099 ?
                  $signed($unsigned((~&reg5449))) : reg5093[(4'hf):(1'h0)]))
                begin
                  reg6981 <= reg4594[(4'ha):(2'h2)];
                end
              else
                begin
                  reg6981 <= ((reg5250 ?
                          (reg4722 ?
                              (+(8'had)) : forvar4577[(2'h2):(2'h2)]) : $signed($unsigned(forvar4727))) ?
                      (8'hb6) : reg5268[(1'h1):(1'h0)]);
                  if (($unsigned(({reg5280} ?
                      (reg4739 != reg5441) : $unsigned(forvar5064))) <<< (((reg5299 ?
                              reg5047 : reg4902) ?
                          (forvar5247 & reg5134) : {reg5339}) ?
                      (~|((8'hac) ^ reg6900)) : reg4894[(3'h6):(1'h0)])))
                    begin
                      reg6982 <= ((($unsigned(reg5501) ?
                                  $unsigned(forvar5314) : $signed(reg5187)) ?
                              reg5032[(4'ha):(3'h6)] : ((reg5385 - reg4692) ?
                                  (forvar4908 >>> reg5106) : reg4992[(1'h1):(1'h0)])) ?
                          $unsigned($unsigned(forvar4588[(4'h8):(3'h5)])) : (reg4908 ^~ ((~&reg5034) << (reg5078 ?
                              reg4856 : reg4740))));
                      reg6983 <= $signed($unsigned($signed($signed(forvar5165))));
                      reg6984 <= $signed(reg5227[(3'h5):(3'h5)]);
                    end
                  else
                    begin
                      reg6982 <= (forvar4958[(1'h0):(1'h0)] <<< (reg6868 + ($unsigned(forvar4578) ?
                          forvar4843 : (^(8'hb2)))));
                      reg6983 <= (^~$signed(forvar5036[(4'hc):(3'h5)]));
                      reg6984 <= ({$unsigned(reg5016[(3'h4):(2'h3)])} ?
                          reg5333[(1'h1):(1'h1)] : reg6885[(2'h3):(2'h3)]);
                    end
                end
              if ((reg4702 ^ (~|$signed(((8'ha5) ? forvar4819 : (8'haf))))))
                begin
                  for (forvar6985 = (1'h0); (forvar6985 < (1'h0)); forvar6985 = (forvar6985 + (1'h1)))
                    begin
                      reg6986 <= (reg5369 ~^ $signed((!reg5199)));
                      reg6987 <= (($signed((|reg4746)) * reg5136) > $signed($unsigned((+forvar5150))));
                      reg6988 <= ({(reg5427[(4'ha):(3'h6)] >>> $signed(forvar4814))} ?
                          {{(|reg6948)}} : (forvar6952 ?
                              $unsigned((^~reg4624)) : reg5254));
                    end
                end
              else
                begin
                  for (forvar6985 = (1'h0); (forvar6985 < (1'h1)); forvar6985 = (forvar6985 + (1'h1)))
                    begin
                      reg6986 <= {reg6982};
                      reg6987 <= forvar5208[(3'h6):(3'h5)];
                    end
                  if ((reg5033 == $signed(reg6906)))
                    begin
                      reg6988 <= {(~^reg4693)};
                    end
                  else
                    begin
                      reg6988 <= (reg5043[(3'h7):(1'h0)] ~^ ({reg5390} ?
                          {forvar5148[(1'h0):(1'h0)]} : (~|$unsigned(reg6881))));
                      reg6989 <= $unsigned(forvar5111[(1'h0):(1'h0)]);
                    end
                  if (reg5358)
                    begin
                      reg6990 <= forvar4819[(1'h0):(1'h0)];
                      reg6991 <= (((~reg6986) ?
                              $signed((reg5411 <<< reg5388)) : $signed((reg4582 - (8'ha7)))) ?
                          forvar4840[(2'h3):(2'h3)] : (((&forvar5252) ?
                                  forvar5382[(3'h5):(1'h1)] : ((8'hb3) ~^ reg5496)) ?
                              forvar5102 : {reg4719[(4'ha):(2'h3)]}));
                      reg6992 <= forvar5453;
                    end
                  else
                    begin
                      reg6990 <= (8'hb1);
                      reg6991 <= (reg5429[(3'h4):(2'h3)] ^ (($unsigned(forvar5416) >>> $signed(forvar4952)) - $unsigned(reg5129)));
                      reg6992 <= $unsigned((forvar4609[(1'h1):(1'h0)] != {forvar5130}));
                    end
                end
              if ($signed((~^reg4791[(4'h8):(4'h8)])))
                begin
                  if ($unsigned($signed(($unsigned(forvar4789) <= forvar4759[(3'h4):(2'h2)]))))
                    begin
                      reg6993 <= (~^reg5464[(2'h2):(2'h2)]);
                      reg6994 <= {$unsigned($unsigned($signed(reg5189)))};
                      reg6995 <= (~forvar6897);
                    end
                  else
                    begin
                      reg6993 <= forvar5165;
                      reg6994 <= (~^($signed((~|forvar4715)) == forvar4760[(3'h5):(3'h4)]));
                      reg6995 <= {(!{((8'hb9) ^~ forvar4777)})};
                      reg6996 <= reg5330[(4'hc):(3'h7)];
                    end
                end
              else
                begin
                  if (reg5149)
                    begin
                      reg6993 <= {$signed($signed($signed(forvar5379)))};
                      reg6994 <= (|(($signed(reg5482) < reg6933[(3'h5):(2'h2)]) ?
                          (^~{reg4900}) : ($signed(forvar4602) ?
                              (^forvar5368) : reg4975[(1'h0):(1'h0)])));
                      reg6995 <= reg4793;
                      reg6996 <= reg4843[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg6993 <= (reg5038 ?
                          forvar4648[(2'h3):(2'h2)] : $unsigned((&(reg5199 >> (8'hb7)))));
                    end
                end
              for (forvar6997 = (1'h0); (forvar6997 < (1'h0)); forvar6997 = (forvar6997 + (1'h1)))
                begin
                  reg6998 <= ($unsigned((~^$signed(reg5430))) ?
                      (~reg5374[(2'h3):(1'h0)]) : $unsigned(((forvar4738 ?
                          reg4687 : reg4867) >> $signed(reg4859))));
                  if ((!$unsigned($signed((reg5004 ? reg5136 : reg5343)))))
                    begin
                      reg6999 <= reg4836;
                      reg7000 <= (|$signed(($unsigned(forvar4913) ?
                          reg5025[(3'h4):(1'h0)] : ((8'hb5) ?
                              forvar5427 : forvar4768))));
                      reg7001 <= ((($signed(reg4688) - reg5030) >>> (~&$signed(reg6961))) ?
                          ((forvar6909[(3'h7):(1'h0)] ?
                              reg4613 : $signed(reg4836)) >>> (!reg4869)) : reg5448[(2'h2):(1'h0)]);
                      reg7002 <= (&reg5268);
                    end
                  else
                    begin
                      reg6999 <= (!{reg4941[(3'h6):(3'h5)]});
                      reg7000 <= $unsigned(reg4755[(1'h0):(1'h0)]);
                      reg7001 <= $signed(reg5319[(4'h8):(3'h6)]);
                    end
                  if ((((~&(&(8'ha9))) ?
                      {(reg5313 == reg5187)} : $signed((reg4590 << forvar5175))) & $unsigned({(~^forvar5380)})))
                    begin
                      reg7003 <= (^((~&(reg4959 ? forvar4952 : (8'ha9))) ?
                          forvar4977[(3'h5):(2'h3)] : (forvar5307 ?
                              (reg5496 ?
                                  forvar4929 : reg5169) : $signed(reg4970))));
                      reg7004 <= forvar4749;
                    end
                  else
                    begin
                      reg7003 <= (~|(8'hab));
                    end
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5505  (y, clk, wire5510, wire5509, wire5508, wire5507, wire5506);
  output wire [(32'h22da):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire5510;
  input wire [(4'hd):(1'h0)] wire5509;
  input wire [(4'hb):(1'h0)] wire5508;
  input wire signed [(4'ha):(1'h0)] wire5507;
  input wire signed [(4'h8):(1'h0)] wire5506;
  wire [(3'h6):(1'h0)] wire6861;
  reg [(3'h7):(1'h0)] reg6860 = (1'h0);
  reg [(4'hc):(1'h0)] reg6859 = (1'h0);
  reg [(5'h10):(1'h0)] reg6858 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6857 = (1'h0);
  reg [(3'h5):(1'h0)] reg6856 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6855 = (1'h0);
  reg [(4'hf):(1'h0)] reg6854 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6853 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6852 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6851 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar6850 = (1'h0);
  reg [(4'he):(1'h0)] forvar6849 = (1'h0);
  reg [(4'h8):(1'h0)] reg6848 = (1'h0);
  reg [(2'h2):(1'h0)] reg6847 = (1'h0);
  reg [(3'h4):(1'h0)] reg6846 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6845 = (1'h0);
  reg [(4'he):(1'h0)] reg6844 = (1'h0);
  reg [(4'he):(1'h0)] reg6843 = (1'h0);
  reg [(4'hb):(1'h0)] reg6842 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6841 = (1'h0);
  reg [(4'hb):(1'h0)] forvar6840 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6839 = (1'h0);
  reg [(2'h2):(1'h0)] forvar6838 = (1'h0);
  reg [(5'h10):(1'h0)] reg6837 = (1'h0);
  reg [(2'h3):(1'h0)] reg6836 = (1'h0);
  reg [(4'he):(1'h0)] reg6835 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6834 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6833 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6832 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6831 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6830 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6829 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6828 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6827 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6826 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6825 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6824 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6823 = (1'h0);
  reg [(4'h9):(1'h0)] reg6822 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6821 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6820 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6819 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6818 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6810 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6817 = (1'h0);
  reg [(4'h8):(1'h0)] reg6816 = (1'h0);
  reg [(3'h4):(1'h0)] reg6815 = (1'h0);
  reg [(4'h9):(1'h0)] reg6814 = (1'h0);
  reg [(4'hb):(1'h0)] reg6813 = (1'h0);
  reg [(4'h8):(1'h0)] reg6812 = (1'h0);
  reg [(3'h5):(1'h0)] reg6811 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar6810 = (1'h0);
  reg [(2'h3):(1'h0)] reg6809 = (1'h0);
  reg [(2'h2):(1'h0)] forvar6808 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6807 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6784 = (1'h0);
  reg [(3'h4):(1'h0)] reg6783 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6775 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6773 = (1'h0);
  reg [(3'h7):(1'h0)] reg6806 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6805 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6804 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6803 = (1'h0);
  reg [(4'hd):(1'h0)] reg6802 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6801 = (1'h0);
  reg [(4'h8):(1'h0)] reg6800 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6799 = (1'h0);
  reg [(5'h10):(1'h0)] reg6798 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6797 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6796 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6795 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6794 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6793 = (1'h0);
  reg [(3'h7):(1'h0)] reg6792 = (1'h0);
  reg [(3'h6):(1'h0)] reg6791 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6790 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6789 = (1'h0);
  reg [(4'h9):(1'h0)] reg6788 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6787 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6786 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6785 = (1'h0);
  reg [(3'h4):(1'h0)] reg6784 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6783 = (1'h0);
  reg [(4'he):(1'h0)] forvar6779 = (1'h0);
  reg [(4'he):(1'h0)] forvar6774 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6782 = (1'h0);
  reg [(4'hf):(1'h0)] reg6781 = (1'h0);
  reg [(4'hb):(1'h0)] reg6780 = (1'h0);
  reg [(4'h8):(1'h0)] reg6779 = (1'h0);
  reg [(4'hb):(1'h0)] reg6778 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6777 = (1'h0);
  reg [(5'h10):(1'h0)] reg6776 = (1'h0);
  reg [(2'h2):(1'h0)] reg6775 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6774 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6773 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6772 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6763 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6769 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6764 = (1'h0);
  reg [(3'h7):(1'h0)] reg6762 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6760 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6759 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar6753 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6749 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6744 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6752 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6740 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6739 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6734 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6733 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6732 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6771 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6770 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6769 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6768 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6767 = (1'h0);
  reg [(4'h8):(1'h0)] reg6766 = (1'h0);
  reg [(5'h10):(1'h0)] reg6765 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6764 = (1'h0);
  reg [(4'ha):(1'h0)] reg6763 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6762 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6761 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6760 = (1'h0);
  reg [(2'h2):(1'h0)] reg6759 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6756 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6755 = (1'h0);
  reg [(4'he):(1'h0)] reg6758 = (1'h0);
  reg [(5'h10):(1'h0)] reg6757 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6756 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6755 = (1'h0);
  reg [(4'hd):(1'h0)] reg6754 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6750 = (1'h0);
  reg [(4'h9):(1'h0)] reg6746 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6745 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6753 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6752 = (1'h0);
  reg [(3'h5):(1'h0)] reg6751 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6750 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6749 = (1'h0);
  reg [(4'he):(1'h0)] reg6748 = (1'h0);
  reg [(3'h6):(1'h0)] reg6747 = (1'h0);
  reg [(4'he):(1'h0)] forvar6746 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6745 = (1'h0);
  reg [(3'h4):(1'h0)] reg6744 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6743 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6742 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6741 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6740 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6739 = (1'h0);
  reg [(3'h4):(1'h0)] reg6738 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6737 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6736 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6735 = (1'h0);
  reg [(4'he):(1'h0)] forvar6734 = (1'h0);
  reg [(2'h2):(1'h0)] reg6733 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6732 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6731 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6726 = (1'h0);
  reg [(5'h10):(1'h0)] reg6730 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6729 = (1'h0);
  reg [(2'h3):(1'h0)] reg6728 = (1'h0);
  reg [(2'h3):(1'h0)] reg6727 = (1'h0);
  reg [(3'h4):(1'h0)] reg6726 = (1'h0);
  reg [(3'h7):(1'h0)] reg6725 = (1'h0);
  reg [(3'h6):(1'h0)] reg6724 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6723 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6722 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6721 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6720 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6719 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6718 = (1'h0);
  reg [(4'hb):(1'h0)] reg6717 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6716 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6715 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6714 = (1'h0);
  reg [(4'hb):(1'h0)] reg6713 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6712 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6711 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6710 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6709 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6708 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6707 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6706 = (1'h0);
  reg [(4'h8):(1'h0)] reg6705 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6704 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6703 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6702 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6701 = (1'h0);
  reg [(3'h6):(1'h0)] reg6700 = (1'h0);
  reg [(4'hc):(1'h0)] reg6699 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6697 = (1'h0);
  reg [(4'he):(1'h0)] reg6698 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6697 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6696 = (1'h0);
  reg [(2'h3):(1'h0)] reg6695 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6694 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6693 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6692 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6691 = (1'h0);
  reg [(4'h8):(1'h0)] reg6690 = (1'h0);
  reg [(4'ha):(1'h0)] reg6689 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6688 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6687 = (1'h0);
  reg [(4'hd):(1'h0)] reg6686 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar6685 = (1'h0);
  reg [(5'h10):(1'h0)] reg6684 = (1'h0);
  reg [(4'h9):(1'h0)] reg6683 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar6682 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6681 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6680 = (1'h0);
  reg [(4'h8):(1'h0)] reg6679 = (1'h0);
  reg [(4'hb):(1'h0)] reg6678 = (1'h0);
  reg [(4'h8):(1'h0)] reg6677 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6676 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6675 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6674 = (1'h0);
  reg [(4'hd):(1'h0)] reg6673 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6672 = (1'h0);
  reg [(3'h5):(1'h0)] reg6671 = (1'h0);
  reg [(3'h5):(1'h0)] reg6670 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6669 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6668 = (1'h0);
  reg [(4'ha):(1'h0)] reg6667 = (1'h0);
  reg [(3'h6):(1'h0)] reg6666 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6665 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6664 = (1'h0);
  reg [(5'h10):(1'h0)] reg6663 = (1'h0);
  reg [(2'h3):(1'h0)] reg6662 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar6661 = (1'h0);
  reg [(4'hd):(1'h0)] reg6660 = (1'h0);
  reg [(4'hd):(1'h0)] reg6659 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6658 = (1'h0);
  reg [(4'hf):(1'h0)] reg6657 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6656 = (1'h0);
  reg [(3'h6):(1'h0)] reg6655 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6654 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6653 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6652 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6651 = (1'h0);
  reg [(2'h2):(1'h0)] reg6650 = (1'h0);
  reg [(4'hb):(1'h0)] forvar6649 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6649 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6639 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar6637 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar6636 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6624 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6623 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6621 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6646 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6645 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6644 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6641 = (1'h0);
  reg [(4'hc):(1'h0)] reg6648 = (1'h0);
  reg [(4'hd):(1'h0)] reg6647 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6646 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6645 = (1'h0);
  reg [(5'h10):(1'h0)] reg6644 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6643 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6642 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6641 = (1'h0);
  reg [(4'hd):(1'h0)] reg6640 = (1'h0);
  reg [(3'h4):(1'h0)] reg6639 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6638 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6637 = (1'h0);
  reg [(3'h6):(1'h0)] reg6636 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6635 = (1'h0);
  reg [(3'h4):(1'h0)] reg6634 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6633 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6632 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6631 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6629 = (1'h0);
  reg [(3'h7):(1'h0)] reg6630 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6629 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6628 = (1'h0);
  reg [(5'h10):(1'h0)] reg6627 = (1'h0);
  reg [(4'hc):(1'h0)] reg6626 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6625 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6624 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6623 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6622 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6621 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar6620 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6619 = (1'h0);
  wire [(2'h3):(1'h0)] wire6618;
  wire [(4'ha):(1'h0)] wire6617;
  wire signed [(4'hc):(1'h0)] wire6616;
  reg [(3'h6):(1'h0)] forvar6609 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6615 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6614 = (1'h0);
  reg [(3'h4):(1'h0)] reg6613 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6612 = (1'h0);
  reg [(4'hf):(1'h0)] reg6611 = (1'h0);
  reg [(4'hf):(1'h0)] reg6610 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6609 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6608 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6607 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6606 = (1'h0);
  reg [(4'hf):(1'h0)] reg6605 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6603 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6602 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6601 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6597 = (1'h0);
  reg [(4'ha):(1'h0)] reg6604 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6603 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6602 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6601 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6600 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6599 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6598 = (1'h0);
  reg [(3'h7):(1'h0)] reg6597 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6596 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6595 = (1'h0);
  reg [(4'hb):(1'h0)] reg6594 = (1'h0);
  reg [(4'h8):(1'h0)] reg6593 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6592 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6591 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6590 = (1'h0);
  reg [(3'h4):(1'h0)] reg6589 = (1'h0);
  reg [(4'he):(1'h0)] forvar6588 = (1'h0);
  reg [(3'h6):(1'h0)] reg6587 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6586 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6585 = (1'h0);
  reg [(4'he):(1'h0)] reg6584 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar6583 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6582 = (1'h0);
  reg [(4'he):(1'h0)] reg6581 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6580 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6579 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6578 = (1'h0);
  reg [(4'he):(1'h0)] reg6577 = (1'h0);
  reg [(4'he):(1'h0)] forvar6576 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6575 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6574 = (1'h0);
  reg [(3'h4):(1'h0)] reg6546 = (1'h0);
  reg [(2'h2):(1'h0)] reg6573 = (1'h0);
  reg [(2'h2):(1'h0)] reg6571 = (1'h0);
  reg [(3'h7):(1'h0)] reg6572 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6571 = (1'h0);
  reg [(4'hd):(1'h0)] reg6570 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6564 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6562 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6559 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6557 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6555 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6554 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6549 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar6548 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6569 = (1'h0);
  reg [(3'h5):(1'h0)] reg6568 = (1'h0);
  reg [(4'hb):(1'h0)] reg6567 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6566 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6565 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6564 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6563 = (1'h0);
  reg [(4'hd):(1'h0)] reg6562 = (1'h0);
  reg [(4'hc):(1'h0)] reg6561 = (1'h0);
  reg [(2'h3):(1'h0)] reg6560 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6559 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6558 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6557 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6556 = (1'h0);
  reg [(4'he):(1'h0)] reg6555 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6554 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6553 = (1'h0);
  reg [(4'h9):(1'h0)] reg6552 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6551 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6550 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6549 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6548 = (1'h0);
  reg [(4'hc):(1'h0)] reg6547 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6546 = (1'h0);
  wire [(4'hd):(1'h0)] wire6545;
  reg [(4'hb):(1'h0)] reg6544 = (1'h0);
  reg [(2'h3):(1'h0)] reg6543 = (1'h0);
  reg [(4'hb):(1'h0)] reg6542 = (1'h0);
  reg [(2'h2):(1'h0)] reg6541 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6540 = (1'h0);
  reg [(4'h9):(1'h0)] reg6539 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6538 = (1'h0);
  reg [(2'h2):(1'h0)] reg6537 = (1'h0);
  reg [(4'h9):(1'h0)] reg6536 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6535 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6534 = (1'h0);
  reg [(4'hd):(1'h0)] reg6533 = (1'h0);
  reg [(4'hc):(1'h0)] reg6532 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6531 = (1'h0);
  reg [(3'h7):(1'h0)] reg6530 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6529 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6528 = (1'h0);
  reg [(4'ha):(1'h0)] reg6525 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6522 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6521 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6527 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6526 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6525 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6524 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6523 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6522 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6521 = (1'h0);
  reg [(5'h10):(1'h0)] reg6520 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6519 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6517 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6514 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6513 = (1'h0);
  reg [(4'h9):(1'h0)] reg6512 = (1'h0);
  reg [(5'h10):(1'h0)] reg6518 = (1'h0);
  reg [(4'hb):(1'h0)] reg6517 = (1'h0);
  reg [(4'hd):(1'h0)] reg6516 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6515 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6514 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6513 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6512 = (1'h0);
  reg [(3'h6):(1'h0)] reg6511 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6510 = (1'h0);
  reg [(4'hb):(1'h0)] reg6509 = (1'h0);
  reg [(5'h10):(1'h0)] reg6508 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6507 = (1'h0);
  reg [(4'h8):(1'h0)] reg6506 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6505 = (1'h0);
  reg [(4'he):(1'h0)] reg6504 = (1'h0);
  reg [(4'hc):(1'h0)] reg6503 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6502 = (1'h0);
  reg [(4'hd):(1'h0)] reg6501 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6500 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6499 = (1'h0);
  reg [(4'hb):(1'h0)] forvar6498 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6497 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6496 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6495 = (1'h0);
  reg [(5'h10):(1'h0)] reg6494 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6493 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6492 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6491 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6490 = (1'h0);
  reg [(4'hc):(1'h0)] reg6489 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6488 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6487 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6486 = (1'h0);
  reg [(3'h6):(1'h0)] reg6485 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6484 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6483 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6482 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6470 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6469 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6465 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6481 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6480 = (1'h0);
  reg [(4'ha):(1'h0)] reg6479 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6478 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6477 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6476 = (1'h0);
  reg [(4'h9):(1'h0)] reg6475 = (1'h0);
  reg [(4'h8):(1'h0)] reg6474 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6473 = (1'h0);
  reg [(5'h10):(1'h0)] reg6472 = (1'h0);
  reg [(4'hc):(1'h0)] reg6471 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6470 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6469 = (1'h0);
  reg [(4'hf):(1'h0)] reg6468 = (1'h0);
  reg [(4'hd):(1'h0)] reg6467 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6466 = (1'h0);
  reg [(2'h3):(1'h0)] reg6465 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6464 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar6463 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6462 = (1'h0);
  reg [(4'hd):(1'h0)] reg6461 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6460 = (1'h0);
  reg [(3'h5):(1'h0)] reg6459 = (1'h0);
  reg [(2'h2):(1'h0)] reg6458 = (1'h0);
  reg [(2'h3):(1'h0)] reg6457 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6456 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6455 = (1'h0);
  reg [(4'hd):(1'h0)] reg6454 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6453 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6452 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6451 = (1'h0);
  reg [(4'hb):(1'h0)] reg6450 = (1'h0);
  reg [(4'hd):(1'h0)] reg6449 = (1'h0);
  reg [(3'h4):(1'h0)] reg6448 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6447 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6446 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6445 = (1'h0);
  wire [(2'h2):(1'h0)] wire6444;
  wire [(4'hb):(1'h0)] wire6443;
  reg signed [(4'he):(1'h0)] reg6442 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6441 = (1'h0);
  reg [(3'h6):(1'h0)] reg6440 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6439 = (1'h0);
  reg [(4'hc):(1'h0)] reg6438 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6437 = (1'h0);
  reg [(4'hc):(1'h0)] reg6436 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6435 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6434 = (1'h0);
  reg [(4'hc):(1'h0)] reg6433 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6432 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6431 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6430 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6429 = (1'h0);
  reg [(2'h3):(1'h0)] reg6428 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6427 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6426 = (1'h0);
  reg [(4'hf):(1'h0)] reg6425 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6424 = (1'h0);
  reg [(4'h9):(1'h0)] reg6423 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6422 = (1'h0);
  reg [(4'he):(1'h0)] reg6421 = (1'h0);
  reg [(3'h6):(1'h0)] reg6420 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6419 = (1'h0);
  reg [(3'h6):(1'h0)] reg6418 = (1'h0);
  reg [(4'he):(1'h0)] forvar6417 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6416 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6415 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6414 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6413 = (1'h0);
  reg [(4'h9):(1'h0)] reg6412 = (1'h0);
  reg [(4'he):(1'h0)] forvar6411 = (1'h0);
  reg [(2'h2):(1'h0)] reg6410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6409 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6407 = (1'h0);
  reg [(2'h3):(1'h0)] reg6406 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6408 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6407 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6406 = (1'h0);
  reg [(4'hb):(1'h0)] forvar6405 = (1'h0);
  reg [(3'h5):(1'h0)] reg6404 = (1'h0);
  reg [(3'h7):(1'h0)] reg6403 = (1'h0);
  reg [(4'h8):(1'h0)] reg6402 = (1'h0);
  reg [(3'h6):(1'h0)] reg6401 = (1'h0);
  reg [(4'ha):(1'h0)] reg6400 = (1'h0);
  reg [(4'ha):(1'h0)] reg6399 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6398 = (1'h0);
  reg [(4'hb):(1'h0)] reg6397 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6394 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6393 = (1'h0);
  reg [(4'he):(1'h0)] forvar6384 = (1'h0);
  reg [(4'ha):(1'h0)] reg6381 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6379 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6377 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6375 = (1'h0);
  reg [(4'h8):(1'h0)] reg6396 = (1'h0);
  reg [(2'h3):(1'h0)] reg6392 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6387 = (1'h0);
  reg [(4'hf):(1'h0)] reg6395 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6394 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6393 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6392 = (1'h0);
  reg [(4'hf):(1'h0)] reg6391 = (1'h0);
  reg [(2'h2):(1'h0)] reg6390 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6389 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6388 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6387 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6386 = (1'h0);
  reg [(3'h6):(1'h0)] reg6385 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6384 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6383 = (1'h0);
  reg [(4'hf):(1'h0)] reg6382 = (1'h0);
  reg [(4'he):(1'h0)] forvar6381 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6380 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6379 = (1'h0);
  reg [(3'h5):(1'h0)] reg6378 = (1'h0);
  reg [(4'ha):(1'h0)] reg6377 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6376 = (1'h0);
  reg [(4'hb):(1'h0)] reg6375 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6374 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6373 = (1'h0);
  reg [(2'h2):(1'h0)] reg6361 = (1'h0);
  reg [(4'hc):(1'h0)] reg6372 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar6371 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6370 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6369 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6368 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6367 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6366 = (1'h0);
  reg [(2'h3):(1'h0)] reg6365 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6364 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6363 = (1'h0);
  reg [(4'hb):(1'h0)] reg6362 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6361 = (1'h0);
  reg [(4'hb):(1'h0)] reg6352 = (1'h0);
  reg [(4'hf):(1'h0)] reg6360 = (1'h0);
  reg [(5'h10):(1'h0)] reg6359 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6358 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6357 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6356 = (1'h0);
  reg [(3'h7):(1'h0)] reg6355 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6354 = (1'h0);
  reg [(3'h5):(1'h0)] reg6353 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6352 = (1'h0);
  reg [(4'hf):(1'h0)] reg6351 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6350 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6349 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6348 = (1'h0);
  reg [(2'h2):(1'h0)] forvar6347 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6346 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6345 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6344 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6343 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6342 = (1'h0);
  reg [(4'he):(1'h0)] reg6341 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6340 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6339 = (1'h0);
  reg [(4'hb):(1'h0)] reg6339 = (1'h0);
  reg [(4'h8):(1'h0)] reg6338 = (1'h0);
  reg [(4'he):(1'h0)] reg6337 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6336 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6335 = (1'h0);
  reg [(2'h2):(1'h0)] reg6334 = (1'h0);
  reg [(4'hc):(1'h0)] reg6333 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6332 = (1'h0);
  reg [(3'h5):(1'h0)] reg6331 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6330 = (1'h0);
  reg [(4'hb):(1'h0)] reg6329 = (1'h0);
  reg [(3'h5):(1'h0)] reg6328 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6327 = (1'h0);
  reg [(2'h3):(1'h0)] reg6326 = (1'h0);
  reg [(4'he):(1'h0)] forvar6325 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6324 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6317 = (1'h0);
  reg [(3'h5):(1'h0)] forvar6316 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6312 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6323 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6322 = (1'h0);
  reg [(3'h4):(1'h0)] reg6321 = (1'h0);
  reg [(4'hd):(1'h0)] reg6320 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar6319 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6318 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6317 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6316 = (1'h0);
  reg [(4'hb):(1'h0)] reg6315 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6314 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6313 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6312 = (1'h0);
  reg [(3'h4):(1'h0)] reg6311 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6310 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6309 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6308 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6307 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6306 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6305 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6304 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6303 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6302 = (1'h0);
  reg [(2'h2):(1'h0)] reg6301 = (1'h0);
  reg [(4'ha):(1'h0)] reg6300 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6299 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6298 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6297 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6296 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6295 = (1'h0);
  reg [(2'h2):(1'h0)] reg6294 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6293 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6292 = (1'h0);
  reg [(4'ha):(1'h0)] reg6291 = (1'h0);
  reg [(2'h3):(1'h0)] reg6290 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6289 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6288 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6287 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6286 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6285 = (1'h0);
  reg [(2'h3):(1'h0)] reg6284 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6283 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6282 = (1'h0);
  reg [(2'h2):(1'h0)] reg6281 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6280 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6279 = (1'h0);
  reg [(4'hd):(1'h0)] reg6278 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6277 = (1'h0);
  reg [(3'h7):(1'h0)] reg6276 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6275 = (1'h0);
  reg [(4'h9):(1'h0)] reg6274 = (1'h0);
  reg [(3'h4):(1'h0)] reg6273 = (1'h0);
  reg [(3'h6):(1'h0)] reg6272 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6271 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6270 = (1'h0);
  reg [(4'hb):(1'h0)] forvar6269 = (1'h0);
  reg [(4'he):(1'h0)] reg6268 = (1'h0);
  reg [(4'hd):(1'h0)] reg6267 = (1'h0);
  reg [(3'h4):(1'h0)] reg6266 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6265 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6264 = (1'h0);
  reg [(4'ha):(1'h0)] reg6263 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6262 = (1'h0);
  reg [(4'he):(1'h0)] reg6261 = (1'h0);
  reg [(4'hd):(1'h0)] reg6260 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6257 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6259 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6258 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6257 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6244 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6243 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6256 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6255 = (1'h0);
  reg [(2'h2):(1'h0)] reg6254 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6253 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6252 = (1'h0);
  reg [(4'hc):(1'h0)] reg6251 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6250 = (1'h0);
  reg [(4'he):(1'h0)] reg6249 = (1'h0);
  reg [(4'h8):(1'h0)] reg6248 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6247 = (1'h0);
  reg [(3'h7):(1'h0)] reg6246 = (1'h0);
  reg [(4'h9):(1'h0)] reg6245 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6244 = (1'h0);
  reg [(4'h9):(1'h0)] reg6243 = (1'h0);
  reg [(3'h4):(1'h0)] reg6242 = (1'h0);
  reg [(4'hb):(1'h0)] reg6241 = (1'h0);
  reg [(2'h2):(1'h0)] reg6240 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6239 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6238 = (1'h0);
  reg [(3'h6):(1'h0)] reg6237 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6236 = (1'h0);
  reg [(4'hb):(1'h0)] reg6235 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6234 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6233 = (1'h0);
  reg [(4'he):(1'h0)] forvar6232 = (1'h0);
  reg [(4'hd):(1'h0)] reg6231 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6230 = (1'h0);
  reg [(4'hf):(1'h0)] reg6229 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6228 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6227 = (1'h0);
  reg [(3'h4):(1'h0)] reg6226 = (1'h0);
  reg [(4'h8):(1'h0)] reg6225 = (1'h0);
  reg [(4'h8):(1'h0)] reg6224 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6223 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6222 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6221 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6220 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar6219 = (1'h0);
  wire [(5'h10):(1'h0)] wire6218;
  reg [(2'h3):(1'h0)] reg6217 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6216 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6215 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6214 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6213 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6212 = (1'h0);
  reg [(3'h7):(1'h0)] reg6211 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6210 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6209 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6208 = (1'h0);
  reg [(4'hc):(1'h0)] reg6207 = (1'h0);
  reg [(4'he):(1'h0)] forvar6139 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6134 = (1'h0);
  reg [(3'h7):(1'h0)] reg6127 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6122 = (1'h0);
  reg [(4'hb):(1'h0)] reg6131 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6129 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar6126 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6123 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6120 = (1'h0);
  reg [(4'ha):(1'h0)] reg6116 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6106 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6105 = (1'h0);
  reg [(3'h5):(1'h0)] reg6206 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6195 = (1'h0);
  reg [(2'h3):(1'h0)] reg6191 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6205 = (1'h0);
  reg [(4'h9):(1'h0)] reg6204 = (1'h0);
  reg [(3'h5):(1'h0)] reg6203 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar6202 = (1'h0);
  reg [(4'hb):(1'h0)] reg6201 = (1'h0);
  reg [(5'h10):(1'h0)] reg6200 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6199 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6198 = (1'h0);
  reg [(4'h9):(1'h0)] reg6197 = (1'h0);
  reg [(3'h6):(1'h0)] reg6196 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6195 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6194 = (1'h0);
  reg [(2'h3):(1'h0)] reg6193 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6192 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6191 = (1'h0);
  reg [(4'hc):(1'h0)] reg6190 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6189 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6188 = (1'h0);
  reg [(3'h5):(1'h0)] reg6187 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6186 = (1'h0);
  reg [(4'hf):(1'h0)] reg6185 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6184 = (1'h0);
  reg [(3'h4):(1'h0)] reg6183 = (1'h0);
  reg [(2'h2):(1'h0)] reg6182 = (1'h0);
  reg [(2'h3):(1'h0)] reg6181 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6180 = (1'h0);
  reg [(3'h6):(1'h0)] forvar6179 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6178 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6177 = (1'h0);
  reg [(4'hb):(1'h0)] reg6176 = (1'h0);
  reg [(2'h3):(1'h0)] reg6175 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6174 = (1'h0);
  reg [(4'hf):(1'h0)] reg6173 = (1'h0);
  reg [(4'h9):(1'h0)] reg6172 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6171 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6170 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6168 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6166 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6165 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6164 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6161 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6159 = (1'h0);
  reg [(4'hf):(1'h0)] reg6171 = (1'h0);
  reg [(3'h5):(1'h0)] reg6170 = (1'h0);
  reg [(3'h6):(1'h0)] reg6169 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6168 = (1'h0);
  reg [(3'h5):(1'h0)] reg6167 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6166 = (1'h0);
  reg [(3'h4):(1'h0)] reg6165 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6164 = (1'h0);
  reg [(4'he):(1'h0)] reg6163 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6162 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6161 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6160 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6159 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6158 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6157 = (1'h0);
  reg [(4'he):(1'h0)] forvar6156 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6155 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6154 = (1'h0);
  reg [(3'h6):(1'h0)] reg6153 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6152 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6151 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6150 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6149 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6148 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6147 = (1'h0);
  reg [(4'he):(1'h0)] forvar6145 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6146 = (1'h0);
  reg [(3'h7):(1'h0)] reg6145 = (1'h0);
  reg [(4'ha):(1'h0)] reg6144 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar6143 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6142 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6141 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6140 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6139 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6137 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6136 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar6135 = (1'h0);
  reg [(5'h10):(1'h0)] reg6138 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6137 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6136 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6135 = (1'h0);
  reg [(3'h7):(1'h0)] reg6134 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6133 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6132 = (1'h0);
  reg [(4'h8):(1'h0)] forvar6131 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6121 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar6117 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6130 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6129 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6128 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar6127 = (1'h0);
  reg [(3'h5):(1'h0)] reg6126 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6125 = (1'h0);
  reg [(3'h4):(1'h0)] reg6124 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6123 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6122 = (1'h0);
  reg [(4'hd):(1'h0)] forvar6121 = (1'h0);
  reg [(4'hc):(1'h0)] reg6120 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6119 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6118 = (1'h0);
  reg [(4'hf):(1'h0)] reg6117 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6116 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6099 = (1'h0);
  reg [(3'h6):(1'h0)] reg6100 = (1'h0);
  reg [(4'hb):(1'h0)] reg6115 = (1'h0);
  reg [(4'hd):(1'h0)] reg6114 = (1'h0);
  reg [(3'h5):(1'h0)] reg6113 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6111 = (1'h0);
  reg [(3'h7):(1'h0)] reg6110 = (1'h0);
  reg [(4'hb):(1'h0)] reg6104 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6112 = (1'h0);
  reg [(3'h4):(1'h0)] reg6111 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6110 = (1'h0);
  reg [(3'h5):(1'h0)] reg6109 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6108 = (1'h0);
  reg [(2'h3):(1'h0)] reg6107 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6106 = (1'h0);
  reg [(4'h8):(1'h0)] reg6105 = (1'h0);
  reg [(4'hf):(1'h0)] forvar6104 = (1'h0);
  reg [(2'h2):(1'h0)] reg6103 = (1'h0);
  reg [(4'he):(1'h0)] reg6102 = (1'h0);
  reg [(4'hb):(1'h0)] reg6101 = (1'h0);
  reg [(4'h9):(1'h0)] forvar6100 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6099 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6098 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6097 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6091 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6096 = (1'h0);
  reg [(4'hc):(1'h0)] reg6095 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6094 = (1'h0);
  reg [(3'h7):(1'h0)] reg6093 = (1'h0);
  reg [(3'h4):(1'h0)] reg6092 = (1'h0);
  reg [(4'hf):(1'h0)] reg6091 = (1'h0);
  reg [(4'he):(1'h0)] reg6090 = (1'h0);
  reg [(4'hc):(1'h0)] reg6089 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6088 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6087 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6086 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6085 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6084 = (1'h0);
  reg [(4'h8):(1'h0)] reg6083 = (1'h0);
  reg [(4'hd):(1'h0)] reg6082 = (1'h0);
  reg [(2'h2):(1'h0)] forvar6081 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6080 = (1'h0);
  reg [(4'ha):(1'h0)] forvar6079 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar6078 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6077 = (1'h0);
  reg [(4'hf):(1'h0)] reg6076 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6075 = (1'h0);
  reg [(4'he):(1'h0)] reg6074 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6073 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6072 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg6071 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6070 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6069 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6068 = (1'h0);
  reg [(4'hb):(1'h0)] reg6067 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6066 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6065 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6064 = (1'h0);
  reg [(5'h10):(1'h0)] reg6063 = (1'h0);
  reg [(4'hd):(1'h0)] reg6062 = (1'h0);
  reg [(4'hb):(1'h0)] forvar6061 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6060 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg6059 = (1'h0);
  reg [(4'hf):(1'h0)] reg6058 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar6050 = (1'h0);
  reg [(4'h8):(1'h0)] reg6044 = (1'h0);
  reg [(4'hd):(1'h0)] reg6057 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar6049 = (1'h0);
  reg [(4'hb):(1'h0)] reg6045 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6056 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar6055 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6054 = (1'h0);
  reg [(4'hd):(1'h0)] reg6053 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6052 = (1'h0);
  reg signed [(4'he):(1'h0)] reg6051 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg6050 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6049 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6048 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6047 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6046 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar6045 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6044 = (1'h0);
  reg [(4'hd):(1'h0)] reg6043 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6042 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg6041 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6040 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6039 = (1'h0);
  reg [(4'h9):(1'h0)] reg6038 = (1'h0);
  reg [(4'hd):(1'h0)] reg6037 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6036 = (1'h0);
  reg [(3'h4):(1'h0)] forvar6035 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6034 = (1'h0);
  reg [(4'h8):(1'h0)] reg6033 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg6032 = (1'h0);
  reg [(4'h9):(1'h0)] reg6031 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6030 = (1'h0);
  reg [(5'h10):(1'h0)] reg6029 = (1'h0);
  reg [(3'h7):(1'h0)] reg6028 = (1'h0);
  reg [(4'hd):(1'h0)] reg6027 = (1'h0);
  reg [(4'hc):(1'h0)] forvar6026 = (1'h0);
  reg [(2'h2):(1'h0)] reg6025 = (1'h0);
  reg [(3'h6):(1'h0)] reg6024 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg6023 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg6022 = (1'h0);
  reg [(3'h7):(1'h0)] forvar6021 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6020 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar6019 = (1'h0);
  reg [(5'h10):(1'h0)] forvar6018 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire6016;
  assign y = {wire6861,
                 reg6860,
                 reg6859,
                 reg6858,
                 reg6857,
                 reg6856,
                 reg6855,
                 reg6854,
                 forvar6853,
                 reg6852,
                 forvar6851,
                 forvar6850,
                 forvar6849,
                 reg6848,
                 reg6847,
                 reg6846,
                 forvar6845,
                 reg6844,
                 reg6843,
                 reg6842,
                 reg6841,
                 forvar6840,
                 forvar6839,
                 forvar6838,
                 reg6837,
                 reg6836,
                 reg6835,
                 reg6834,
                 forvar6833,
                 reg6832,
                 reg6831,
                 reg6830,
                 forvar6829,
                 reg6828,
                 reg6827,
                 forvar6826,
                 forvar6825,
                 forvar6824,
                 reg6823,
                 reg6822,
                 reg6821,
                 reg6820,
                 forvar6819,
                 reg6818,
                 reg6810,
                 reg6817,
                 reg6816,
                 reg6815,
                 reg6814,
                 reg6813,
                 reg6812,
                 reg6811,
                 forvar6810,
                 reg6809,
                 forvar6808,
                 forvar6807,
                 forvar6784,
                 reg6783,
                 forvar6775,
                 forvar6773,
                 reg6806,
                 reg6805,
                 reg6804,
                 reg6803,
                 reg6802,
                 forvar6801,
                 reg6800,
                 reg6799,
                 reg6798,
                 reg6797,
                 forvar6796,
                 forvar6795,
                 reg6794,
                 forvar6793,
                 reg6792,
                 reg6791,
                 reg6790,
                 reg6789,
                 reg6788,
                 reg6787,
                 reg6786,
                 reg6785,
                 reg6784,
                 forvar6783,
                 forvar6779,
                 forvar6774,
                 reg6782,
                 reg6781,
                 reg6780,
                 reg6779,
                 reg6778,
                 reg6777,
                 reg6776,
                 reg6775,
                 reg6774,
                 reg6773,
                 forvar6772,
                 forvar6763,
                 reg6769,
                 reg6764,
                 reg6762,
                 forvar6760,
                 forvar6759,
                 forvar6753,
                 forvar6749,
                 forvar6744,
                 forvar6752,
                 reg6740,
                 reg6739,
                 reg6734,
                 forvar6733,
                 forvar6732,
                 reg6771,
                 reg6770,
                 forvar6769,
                 reg6768,
                 reg6767,
                 reg6766,
                 reg6765,
                 forvar6764,
                 reg6763,
                 forvar6762,
                 reg6761,
                 reg6760,
                 reg6759,
                 forvar6756,
                 forvar6755,
                 reg6758,
                 reg6757,
                 reg6756,
                 reg6755,
                 reg6754,
                 reg6750,
                 reg6746,
                 forvar6745,
                 reg6753,
                 reg6752,
                 reg6751,
                 forvar6750,
                 reg6749,
                 reg6748,
                 reg6747,
                 forvar6746,
                 reg6745,
                 reg6744,
                 reg6743,
                 reg6742,
                 reg6741,
                 forvar6740,
                 forvar6739,
                 reg6738,
                 reg6737,
                 reg6736,
                 reg6735,
                 forvar6734,
                 reg6733,
                 reg6732,
                 forvar6731,
                 forvar6726,
                 reg6730,
                 reg6729,
                 reg6728,
                 reg6727,
                 reg6726,
                 reg6725,
                 reg6724,
                 forvar6723,
                 forvar6722,
                 reg6721,
                 reg6720,
                 reg6719,
                 reg6718,
                 reg6717,
                 forvar6716,
                 reg6715,
                 reg6714,
                 reg6713,
                 forvar6712,
                 reg6711,
                 reg6710,
                 reg6709,
                 reg6708,
                 reg6707,
                 forvar6706,
                 reg6705,
                 reg6704,
                 reg6703,
                 reg6702,
                 forvar6701,
                 reg6700,
                 reg6699,
                 forvar6697,
                 reg6698,
                 reg6697,
                 reg6696,
                 reg6695,
                 reg6694,
                 reg6693,
                 reg6692,
                 forvar6691,
                 reg6690,
                 reg6689,
                 reg6688,
                 forvar6687,
                 reg6686,
                 forvar6685,
                 reg6684,
                 reg6683,
                 forvar6682,
                 forvar6681,
                 forvar6680,
                 reg6679,
                 reg6678,
                 reg6677,
                 forvar6676,
                 forvar6675,
                 reg6674,
                 reg6673,
                 reg6672,
                 reg6671,
                 reg6670,
                 forvar6669,
                 reg6668,
                 reg6667,
                 reg6666,
                 reg6665,
                 reg6664,
                 reg6663,
                 reg6662,
                 forvar6661,
                 reg6660,
                 reg6659,
                 forvar6658,
                 reg6657,
                 reg6656,
                 reg6655,
                 reg6654,
                 reg6653,
                 reg6652,
                 reg6651,
                 reg6650,
                 forvar6649,
                 reg6649,
                 forvar6639,
                 forvar6637,
                 forvar6636,
                 forvar6624,
                 forvar6623,
                 forvar6621,
                 forvar6646,
                 reg6645,
                 forvar6644,
                 reg6641,
                 reg6648,
                 reg6647,
                 reg6646,
                 forvar6645,
                 reg6644,
                 reg6643,
                 reg6642,
                 forvar6641,
                 reg6640,
                 reg6639,
                 reg6638,
                 reg6637,
                 reg6636,
                 reg6635,
                 reg6634,
                 reg6633,
                 reg6632,
                 reg6631,
                 forvar6629,
                 reg6630,
                 reg6629,
                 reg6628,
                 reg6627,
                 reg6626,
                 reg6625,
                 reg6624,
                 reg6623,
                 reg6622,
                 reg6621,
                 forvar6620,
                 forvar6619,
                 wire6618,
                 wire6617,
                 wire6616,
                 forvar6609,
                 reg6615,
                 reg6614,
                 reg6613,
                 reg6612,
                 reg6611,
                 reg6610,
                 reg6609,
                 reg6608,
                 reg6607,
                 forvar6606,
                 reg6605,
                 forvar6603,
                 reg6602,
                 forvar6601,
                 forvar6597,
                 reg6604,
                 reg6603,
                 forvar6602,
                 reg6601,
                 reg6600,
                 reg6599,
                 reg6598,
                 reg6597,
                 reg6596,
                 forvar6595,
                 reg6594,
                 reg6593,
                 forvar6592,
                 forvar6591,
                 reg6590,
                 reg6589,
                 forvar6588,
                 reg6587,
                 forvar6586,
                 reg6585,
                 reg6584,
                 forvar6583,
                 reg6582,
                 reg6581,
                 reg6580,
                 forvar6579,
                 reg6578,
                 reg6577,
                 forvar6576,
                 reg6575,
                 forvar6574,
                 reg6546,
                 reg6573,
                 reg6571,
                 reg6572,
                 forvar6571,
                 reg6570,
                 reg6564,
                 forvar6562,
                 reg6559,
                 reg6557,
                 forvar6555,
                 reg6554,
                 reg6549,
                 forvar6548,
                 reg6569,
                 reg6568,
                 reg6567,
                 reg6566,
                 reg6565,
                 forvar6564,
                 reg6563,
                 reg6562,
                 reg6561,
                 reg6560,
                 forvar6559,
                 reg6558,
                 forvar6557,
                 reg6556,
                 reg6555,
                 forvar6554,
                 reg6553,
                 reg6552,
                 reg6551,
                 reg6550,
                 forvar6549,
                 reg6548,
                 reg6547,
                 forvar6546,
                 wire6545,
                 reg6544,
                 reg6543,
                 reg6542,
                 reg6541,
                 forvar6540,
                 reg6539,
                 reg6538,
                 reg6537,
                 reg6536,
                 reg6535,
                 forvar6534,
                 reg6533,
                 reg6532,
                 reg6531,
                 reg6530,
                 forvar6529,
                 forvar6528,
                 reg6525,
                 forvar6522,
                 reg6521,
                 reg6527,
                 reg6526,
                 forvar6525,
                 reg6524,
                 reg6523,
                 reg6522,
                 forvar6521,
                 reg6520,
                 forvar6519,
                 forvar6517,
                 reg6514,
                 forvar6513,
                 reg6512,
                 reg6518,
                 reg6517,
                 reg6516,
                 reg6515,
                 forvar6514,
                 reg6513,
                 forvar6512,
                 reg6511,
                 reg6510,
                 reg6509,
                 reg6508,
                 forvar6507,
                 reg6506,
                 reg6505,
                 reg6504,
                 reg6503,
                 forvar6502,
                 reg6501,
                 reg6500,
                 reg6499,
                 forvar6498,
                 reg6497,
                 forvar6496,
                 reg6495,
                 reg6494,
                 reg6493,
                 forvar6492,
                 forvar6491,
                 reg6490,
                 reg6489,
                 forvar6488,
                 forvar6487,
                 reg6486,
                 reg6485,
                 forvar6484,
                 forvar6483,
                 forvar6482,
                 forvar6470,
                 reg6469,
                 forvar6465,
                 reg6481,
                 reg6480,
                 reg6479,
                 reg6478,
                 forvar6477,
                 reg6476,
                 reg6475,
                 reg6474,
                 reg6473,
                 reg6472,
                 reg6471,
                 reg6470,
                 forvar6469,
                 reg6468,
                 reg6467,
                 reg6466,
                 reg6465,
                 forvar6464,
                 forvar6463,
                 reg6462,
                 reg6461,
                 reg6460,
                 reg6459,
                 reg6458,
                 reg6457,
                 reg6456,
                 reg6455,
                 reg6454,
                 forvar6453,
                 forvar6452,
                 reg6451,
                 reg6450,
                 reg6449,
                 reg6448,
                 forvar6447,
                 forvar6446,
                 forvar6445,
                 wire6444,
                 wire6443,
                 reg6442,
                 reg6441,
                 reg6440,
                 reg6439,
                 reg6438,
                 reg6437,
                 reg6436,
                 forvar6435,
                 reg6434,
                 reg6433,
                 forvar6432,
                 forvar6431,
                 forvar6430,
                 reg6429,
                 reg6428,
                 reg6427,
                 forvar6426,
                 reg6425,
                 reg6424,
                 reg6423,
                 reg6422,
                 reg6421,
                 reg6420,
                 reg6419,
                 reg6418,
                 forvar6417,
                 reg6416,
                 reg6415,
                 reg6414,
                 reg6413,
                 reg6412,
                 forvar6411,
                 reg6410,
                 reg6409,
                 forvar6407,
                 reg6406,
                 reg6408,
                 reg6407,
                 forvar6406,
                 forvar6405,
                 reg6404,
                 reg6403,
                 reg6402,
                 reg6401,
                 reg6400,
                 reg6399,
                 forvar6398,
                 reg6397,
                 forvar6394,
                 forvar6393,
                 forvar6384,
                 reg6381,
                 reg6379,
                 forvar6377,
                 forvar6375,
                 reg6396,
                 reg6392,
                 reg6387,
                 reg6395,
                 reg6394,
                 reg6393,
                 forvar6392,
                 reg6391,
                 reg6390,
                 reg6389,
                 reg6388,
                 forvar6387,
                 reg6386,
                 reg6385,
                 reg6384,
                 reg6383,
                 reg6382,
                 forvar6381,
                 reg6380,
                 forvar6379,
                 reg6378,
                 reg6377,
                 reg6376,
                 reg6375,
                 forvar6374,
                 forvar6373,
                 reg6361,
                 reg6372,
                 forvar6371,
                 reg6370,
                 reg6369,
                 reg6368,
                 reg6367,
                 forvar6366,
                 reg6365,
                 reg6364,
                 reg6363,
                 reg6362,
                 forvar6361,
                 reg6352,
                 reg6360,
                 reg6359,
                 reg6358,
                 forvar6357,
                 reg6356,
                 reg6355,
                 reg6354,
                 reg6353,
                 forvar6352,
                 reg6351,
                 reg6350,
                 forvar6349,
                 reg6348,
                 forvar6347,
                 reg6346,
                 reg6345,
                 reg6344,
                 reg6343,
                 reg6342,
                 reg6341,
                 reg6340,
                 forvar6339,
                 reg6339,
                 reg6338,
                 reg6337,
                 forvar6336,
                 forvar6335,
                 reg6334,
                 reg6333,
                 forvar6332,
                 reg6331,
                 reg6330,
                 reg6329,
                 reg6328,
                 forvar6327,
                 reg6326,
                 forvar6325,
                 forvar6324,
                 reg6317,
                 forvar6316,
                 reg6312,
                 reg6323,
                 forvar6322,
                 reg6321,
                 reg6320,
                 forvar6319,
                 reg6318,
                 forvar6317,
                 reg6316,
                 reg6315,
                 reg6314,
                 reg6313,
                 forvar6312,
                 reg6311,
                 reg6310,
                 reg6309,
                 reg6308,
                 forvar6307,
                 forvar6306,
                 reg6305,
                 reg6304,
                 forvar6303,
                 forvar6302,
                 reg6301,
                 reg6300,
                 reg6299,
                 forvar6298,
                 forvar6297,
                 forvar6296,
                 forvar6295,
                 reg6294,
                 forvar6293,
                 reg6292,
                 reg6291,
                 reg6290,
                 reg6289,
                 forvar6288,
                 reg6287,
                 forvar6286,
                 reg6285,
                 reg6284,
                 forvar6283,
                 forvar6282,
                 reg6281,
                 reg6280,
                 reg6279,
                 reg6278,
                 forvar6277,
                 reg6276,
                 reg6275,
                 reg6274,
                 reg6273,
                 reg6272,
                 reg6271,
                 forvar6270,
                 forvar6269,
                 reg6268,
                 reg6267,
                 reg6266,
                 reg6265,
                 reg6264,
                 reg6263,
                 reg6262,
                 reg6261,
                 reg6260,
                 reg6257,
                 reg6259,
                 reg6258,
                 forvar6257,
                 reg6244,
                 forvar6243,
                 reg6256,
                 reg6255,
                 reg6254,
                 forvar6253,
                 reg6252,
                 reg6251,
                 reg6250,
                 reg6249,
                 reg6248,
                 reg6247,
                 reg6246,
                 reg6245,
                 forvar6244,
                 reg6243,
                 reg6242,
                 reg6241,
                 reg6240,
                 reg6239,
                 reg6238,
                 reg6237,
                 reg6236,
                 reg6235,
                 forvar6234,
                 reg6233,
                 forvar6232,
                 reg6231,
                 reg6230,
                 reg6229,
                 forvar6228,
                 reg6227,
                 reg6226,
                 reg6225,
                 reg6224,
                 reg6223,
                 reg6222,
                 forvar6221,
                 forvar6220,
                 forvar6219,
                 wire6218,
                 reg6217,
                 reg6216,
                 reg6215,
                 reg6214,
                 reg6213,
                 forvar6212,
                 reg6211,
                 forvar6210,
                 forvar6209,
                 forvar6208,
                 reg6207,
                 forvar6139,
                 forvar6134,
                 reg6127,
                 forvar6122,
                 reg6131,
                 forvar6129,
                 forvar6126,
                 forvar6123,
                 forvar6120,
                 reg6116,
                 forvar6106,
                 forvar6105,
                 reg6206,
                 reg6195,
                 reg6191,
                 reg6205,
                 reg6204,
                 reg6203,
                 forvar6202,
                 reg6201,
                 reg6200,
                 reg6199,
                 forvar6198,
                 reg6197,
                 reg6196,
                 forvar6195,
                 reg6194,
                 reg6193,
                 reg6192,
                 forvar6191,
                 reg6190,
                 reg6189,
                 reg6188,
                 reg6187,
                 forvar6186,
                 reg6185,
                 reg6184,
                 reg6183,
                 reg6182,
                 reg6181,
                 reg6180,
                 forvar6179,
                 forvar6178,
                 forvar6177,
                 reg6176,
                 reg6175,
                 reg6174,
                 reg6173,
                 reg6172,
                 forvar6171,
                 forvar6170,
                 reg6168,
                 forvar6166,
                 forvar6165,
                 reg6164,
                 forvar6161,
                 reg6159,
                 reg6171,
                 reg6170,
                 reg6169,
                 forvar6168,
                 reg6167,
                 reg6166,
                 reg6165,
                 forvar6164,
                 reg6163,
                 reg6162,
                 reg6161,
                 reg6160,
                 forvar6159,
                 reg6158,
                 reg6157,
                 forvar6156,
                 forvar6155,
                 reg6154,
                 reg6153,
                 reg6152,
                 reg6151,
                 reg6150,
                 forvar6149,
                 reg6148,
                 reg6147,
                 forvar6145,
                 reg6146,
                 reg6145,
                 reg6144,
                 forvar6143,
                 reg6142,
                 reg6141,
                 reg6140,
                 reg6139,
                 forvar6137,
                 reg6136,
                 forvar6135,
                 reg6138,
                 reg6137,
                 forvar6136,
                 reg6135,
                 reg6134,
                 reg6133,
                 reg6132,
                 forvar6131,
                 reg6121,
                 forvar6117,
                 reg6130,
                 reg6129,
                 reg6128,
                 forvar6127,
                 reg6126,
                 reg6125,
                 reg6124,
                 reg6123,
                 reg6122,
                 forvar6121,
                 reg6120,
                 reg6119,
                 reg6118,
                 reg6117,
                 forvar6116,
                 reg6099,
                 reg6100,
                 reg6115,
                 reg6114,
                 reg6113,
                 forvar6111,
                 reg6110,
                 reg6104,
                 reg6112,
                 reg6111,
                 forvar6110,
                 reg6109,
                 reg6108,
                 reg6107,
                 reg6106,
                 reg6105,
                 forvar6104,
                 reg6103,
                 reg6102,
                 reg6101,
                 forvar6100,
                 forvar6099,
                 reg6098,
                 forvar6097,
                 forvar6091,
                 reg6096,
                 reg6095,
                 forvar6094,
                 reg6093,
                 reg6092,
                 reg6091,
                 reg6090,
                 reg6089,
                 forvar6088,
                 forvar6087,
                 reg6086,
                 reg6085,
                 reg6084,
                 reg6083,
                 reg6082,
                 forvar6081,
                 reg6080,
                 forvar6079,
                 forvar6078,
                 reg6077,
                 reg6076,
                 reg6075,
                 reg6074,
                 forvar6073,
                 reg6072,
                 reg6071,
                 reg6070,
                 reg6069,
                 reg6068,
                 reg6067,
                 reg6066,
                 forvar6065,
                 reg6064,
                 reg6063,
                 reg6062,
                 forvar6061,
                 forvar6060,
                 reg6059,
                 reg6058,
                 forvar6050,
                 reg6044,
                 reg6057,
                 forvar6049,
                 reg6045,
                 reg6056,
                 forvar6055,
                 reg6054,
                 reg6053,
                 reg6052,
                 reg6051,
                 reg6050,
                 reg6049,
                 reg6048,
                 reg6047,
                 reg6046,
                 forvar6045,
                 forvar6044,
                 reg6043,
                 reg6042,
                 reg6041,
                 reg6040,
                 reg6039,
                 reg6038,
                 reg6037,
                 forvar6036,
                 forvar6035,
                 reg6034,
                 reg6033,
                 reg6032,
                 reg6031,
                 reg6030,
                 reg6029,
                 reg6028,
                 reg6027,
                 forvar6026,
                 reg6025,
                 reg6024,
                 reg6023,
                 reg6022,
                 forvar6021,
                 forvar6020,
                 forvar6019,
                 forvar6018,
                 wire6016,
                 (1'h0)};
  module5511 modinst6017 (.wire5515(wire5509), .clk(clk), .wire5514(wire5508), .wire5513(wire5506), .y(wire6016), .wire5512(wire5510));
  always
    @(posedge clk) begin
      for (forvar6018 = (1'h0); (forvar6018 < (2'h3)); forvar6018 = (forvar6018 + (1'h1)))
        begin
          for (forvar6019 = (1'h0); (forvar6019 < (1'h0)); forvar6019 = (forvar6019 + (1'h1)))
            begin
              for (forvar6020 = (1'h0); (forvar6020 < (2'h3)); forvar6020 = (forvar6020 + (1'h1)))
                begin
                  for (forvar6021 = (1'h0); (forvar6021 < (2'h2)); forvar6021 = (forvar6021 + (1'h1)))
                    begin
                      reg6022 <= {forvar6019};
                      reg6023 <= wire5506;
                      reg6024 <= reg6022;
                      reg6025 <= ((|{wire5508}) < $signed(reg6022[(3'h5):(3'h5)]));
                    end
                  for (forvar6026 = (1'h0); (forvar6026 < (1'h1)); forvar6026 = (forvar6026 + (1'h1)))
                    begin
                      reg6027 <= $signed(forvar6020);
                      reg6028 <= {$unsigned($signed($unsigned(wire5508)))};
                      reg6029 <= (reg6022 << reg6023);
                      reg6030 <= $signed((reg6029 ?
                          ((!forvar6018) ?
                              $signed(reg6024) : (wire5506 & reg6024)) : $signed(reg6023[(3'h7):(1'h0)])));
                    end
                  if (reg6030)
                    begin
                      reg6031 <= forvar6020;
                      reg6032 <= {($unsigned($unsigned((8'hb8))) == ((forvar6020 ?
                              forvar6019 : (8'h9e)) << $unsigned(reg6028)))};
                    end
                  else
                    begin
                      reg6031 <= $unsigned(reg6031[(1'h0):(1'h0)]);
                      reg6032 <= $unsigned($signed({(~^wire5508)}));
                      reg6033 <= reg6027[(4'hd):(3'h5)];
                      reg6034 <= (~|(wire5509[(4'h9):(1'h0)] ?
                          reg6031[(2'h3):(1'h1)] : reg6027[(3'h7):(3'h5)]));
                    end
                end
              for (forvar6035 = (1'h0); (forvar6035 < (2'h3)); forvar6035 = (forvar6035 + (1'h1)))
                begin
                  for (forvar6036 = (1'h0); (forvar6036 < (1'h0)); forvar6036 = (forvar6036 + (1'h1)))
                    begin
                      reg6037 <= $unsigned(wire5507);
                      reg6038 <= {(8'hb2)};
                    end
                end
              if ((-$signed((8'ha4))))
                begin
                  reg6039 <= wire6016;
                  reg6040 <= (~($unsigned($signed((8'ha6))) ?
                      (8'hae) : (~&wire5507[(2'h2):(1'h0)])));
                end
              else
                begin
                  if ($unsigned($signed($unsigned(wire5507[(4'h8):(1'h0)]))))
                    begin
                      reg6039 <= ($unsigned((-{wire5509})) >= reg6032[(2'h3):(2'h2)]);
                      reg6040 <= ($signed($unsigned((8'hb1))) ?
                          reg6032 : ({$unsigned(forvar6018)} ?
                              $signed((reg6027 ?
                                  reg6033 : reg6029)) : {$unsigned(forvar6021)}));
                    end
                  else
                    begin
                      reg6039 <= $unsigned(reg6034[(3'h4):(1'h0)]);
                    end
                  reg6041 <= ((reg6037[(4'hb):(4'ha)] >= ($unsigned(wire5509) ?
                          (reg6028 * reg6034) : (wire6016 & reg6022))) ?
                      reg6038 : $unsigned($unsigned(reg6028[(2'h3):(2'h3)])));
                end
            end
        end
      reg6042 <= ({((wire6016 ?
              forvar6019 : wire5508) <= reg6027[(2'h3):(1'h0)])} - {reg6041});
      reg6043 <= ($unsigned($unsigned({(8'h9d)})) <<< (($unsigned(forvar6036) << reg6027) ?
          forvar6019[(1'h0):(1'h0)] : (^((8'ha5) > wire5506))));
      if ((~wire5506))
        begin
          for (forvar6044 = (1'h0); (forvar6044 < (1'h1)); forvar6044 = (forvar6044 + (1'h1)))
            begin
              if ({$signed(wire5510[(4'h8):(3'h4)])})
                begin
                  for (forvar6045 = (1'h0); (forvar6045 < (2'h2)); forvar6045 = (forvar6045 + (1'h1)))
                    begin
                      reg6046 <= (!($signed($unsigned(forvar6019)) + ($signed(reg6029) ?
                          reg6034[(2'h2):(1'h0)] : (forvar6026 && (8'haa)))));
                      reg6047 <= $unsigned($signed((^~reg6032[(3'h6):(3'h5)])));
                    end
                  if ((reg6029[(4'ha):(4'h9)] >>> $unsigned($signed($unsigned(reg6025)))))
                    begin
                      reg6048 <= ($unsigned(((forvar6045 ?
                                  forvar6019 : reg6023) ?
                              (wire5509 ? wire5509 : reg6025) : {reg6038})) ?
                          $signed(((reg6039 ? (8'hb6) : reg6029) ?
                              (8'h9e) : $signed((8'h9f)))) : $signed(((forvar6019 * wire5510) ?
                              reg6030[(1'h1):(1'h0)] : $unsigned(wire5508))));
                      reg6049 <= forvar6044;
                      reg6050 <= wire5510[(4'h8):(1'h1)];
                      reg6051 <= ($unsigned($unsigned({wire5507})) ?
                          $signed((~$unsigned(wire5509))) : ($unsigned($signed((8'ha8))) ?
                              (((8'ha1) == reg6050) ?
                                  {(8'h9d)} : forvar6045[(1'h1):(1'h0)]) : ($unsigned(reg6048) ?
                                  (!reg6033) : (reg6030 ?
                                      reg6039 : forvar6036))));
                    end
                  else
                    begin
                      reg6048 <= ($unsigned({(forvar6026 ?
                              reg6024 : forvar6036)}) <= reg6032[(1'h1):(1'h0)]);
                      reg6049 <= (~&((reg6033 ? reg6033 : (8'hb9)) ^ reg6023));
                      reg6050 <= (((~^(reg6050 ^~ reg6027)) ?
                              $signed((reg6046 ?
                                  reg6029 : (8'h9f))) : $unsigned({reg6033})) ?
                          $signed((((8'ha4) ? forvar6035 : wire6016) ?
                              reg6032 : (forvar6035 ?
                                  reg6022 : reg6038))) : $signed($signed((8'hac))));
                    end
                  if ({(($signed(forvar6036) ?
                              reg6051[(2'h3):(2'h3)] : $signed((8'hb6))) ?
                          wire6016 : {reg6041})})
                    begin
                      reg6052 <= ($unsigned($unsigned(forvar6021[(3'h7):(3'h4)])) ?
                          ((reg6048[(1'h1):(1'h0)] ?
                                  $signed((8'hab)) : reg6046[(3'h4):(1'h1)]) ?
                              (reg6033 <= (reg6023 ?
                                  reg6049 : forvar6035)) : reg6028) : {((+reg6043) ?
                                  forvar6018[(4'hf):(4'h8)] : ((8'hab) ?
                                      forvar6019 : reg6041))});
                    end
                  else
                    begin
                      reg6052 <= ($signed($signed((reg6043 < reg6043))) ?
                          $unsigned((~&reg6041)) : $signed((|reg6038[(3'h6):(1'h1)])));
                      reg6053 <= (reg6051[(4'h8):(1'h0)] ?
                          (reg6034 ?
                              $unsigned((+reg6041)) : (-forvar6044)) : ({(~^reg6027)} == reg6037[(4'hd):(4'hc)]));
                      reg6054 <= (((wire5510[(1'h0):(1'h0)] ?
                                  (~^(8'hb1)) : $signed((8'hb1))) ?
                              $signed((^~reg6048)) : $unsigned($signed((8'ha8)))) ?
                          $signed({$unsigned(reg6024)}) : (8'ha5));
                    end
                  for (forvar6055 = (1'h0); (forvar6055 < (1'h0)); forvar6055 = (forvar6055 + (1'h1)))
                    begin
                      reg6056 <= $signed($unsigned($unsigned($unsigned(forvar6019))));
                    end
                end
              else
                begin
                  if ($unsigned($unsigned($unsigned((|reg6041)))))
                    begin
                      reg6045 <= (reg6029[(4'hd):(3'h6)] || (~^reg6034));
                      reg6046 <= (+$unsigned((~&((8'hae) ?
                          forvar6044 : forvar6045))));
                      reg6047 <= ((~(reg6056[(3'h5):(1'h1)] && forvar6021)) ?
                          $signed(((8'h9e) <= (forvar6035 ?
                              reg6037 : reg6049))) : (~|$unsigned((~|(8'hb8)))));
                      reg6048 <= (wire5506 <<< (8'h9e));
                    end
                  else
                    begin
                      reg6045 <= (~|reg6047);
                      reg6046 <= $unsigned((($unsigned(forvar6045) < (reg6027 <= reg6041)) || reg6041));
                      reg6047 <= {(^~(^~(reg6032 <= reg6031)))};
                    end
                  for (forvar6049 = (1'h0); (forvar6049 < (2'h2)); forvar6049 = (forvar6049 + (1'h1)))
                    begin
                      reg6050 <= $signed(reg6048[(1'h0):(1'h0)]);
                      reg6051 <= reg6052[(3'h5):(1'h1)];
                      reg6052 <= ($signed(forvar6035) ?
                          $signed(reg6040[(4'he):(3'h5)]) : (~|$signed(forvar6049[(1'h1):(1'h1)])));
                    end
                end
              reg6057 <= reg6029[(4'he):(4'hb)];
            end
        end
      else
        begin
          if ((!$unsigned((-(forvar6035 ? reg6027 : reg6032)))))
            begin
              if (((forvar6036 ?
                  $signed($unsigned(reg6045)) : (+(reg6025 ?
                      reg6057 : wire5506))) << $unsigned({forvar6035})))
                begin
                  if (wire6016)
                    begin
                      reg6044 <= wire5510;
                      reg6045 <= $signed($unsigned($unsigned($unsigned(reg6044))));
                    end
                  else
                    begin
                      reg6044 <= reg6057[(4'hc):(4'ha)];
                      reg6045 <= ((&$signed($signed(reg6044))) > (~&forvar6021[(2'h2):(1'h0)]));
                    end
                end
              else
                begin
                  for (forvar6044 = (1'h0); (forvar6044 < (1'h1)); forvar6044 = (forvar6044 + (1'h1)))
                    begin
                      reg6045 <= reg6039;
                      reg6046 <= reg6038;
                    end
                end
            end
          else
            begin
              for (forvar6044 = (1'h0); (forvar6044 < (1'h1)); forvar6044 = (forvar6044 + (1'h1)))
                begin
                  for (forvar6045 = (1'h0); (forvar6045 < (1'h0)); forvar6045 = (forvar6045 + (1'h1)))
                    begin
                      reg6046 <= $signed($signed((reg6034 | (reg6050 ?
                          reg6025 : reg6042))));
                      reg6047 <= $signed((^~(((8'hb9) >= reg6029) ?
                          $signed(wire5507) : (~|reg6032))));
                      reg6048 <= (forvar6018[(3'h5):(3'h5)] ?
                          (+(^~$signed(reg6048))) : reg6041[(2'h2):(1'h1)]);
                      reg6049 <= reg6034;
                    end
                end
              for (forvar6050 = (1'h0); (forvar6050 < (1'h1)); forvar6050 = (forvar6050 + (1'h1)))
                begin
                  if (((~&(~|(reg6039 ^ (8'ha5)))) > $signed((reg6030[(3'h4):(2'h3)] || (8'ha4)))))
                    begin
                      reg6051 <= reg6053;
                      reg6052 <= {$unsigned(($unsigned(reg6032) * (~|(8'ha7))))};
                      reg6053 <= ($unsigned(((wire5510 ? (8'haf) : reg6033) ?
                          $unsigned((8'hb9)) : (reg6043 == reg6028))) + $unsigned(reg6033[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg6051 <= $signed(forvar6020);
                      reg6052 <= reg6045[(2'h2):(2'h2)];
                      reg6053 <= {$signed({reg6028[(2'h3):(2'h2)]})};
                    end
                  if ($unsigned(($signed(((8'hb5) ? reg6031 : forvar6021)) ?
                      (~^forvar6050) : $signed($unsigned(reg6039)))))
                    begin
                      reg6054 <= $unsigned(reg6044[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg6054 <= $unsigned(($signed((reg6043 || reg6047)) <<< ($unsigned((8'ha4)) == $signed(reg6044))));
                    end
                  for (forvar6055 = (1'h0); (forvar6055 < (2'h3)); forvar6055 = (forvar6055 + (1'h1)))
                    begin
                      reg6056 <= wire5510[(4'h8):(2'h2)];
                      reg6057 <= (8'hb2);
                      reg6058 <= $signed((^~({reg6047} ?
                          (forvar6055 ? reg6047 : reg6056) : (wire6016 ?
                              forvar6018 : reg6028))));
                      reg6059 <= $signed($unsigned(reg6024));
                    end
                end
              for (forvar6060 = (1'h0); (forvar6060 < (1'h1)); forvar6060 = (forvar6060 + (1'h1)))
                begin
                  for (forvar6061 = (1'h0); (forvar6061 < (1'h1)); forvar6061 = (forvar6061 + (1'h1)))
                    begin
                      reg6062 <= reg6053;
                      reg6063 <= $signed((((8'hb3) ?
                              $signed((8'hb1)) : reg6057) ?
                          ((~&(8'hb0)) ?
                              $unsigned(reg6058) : (~reg6044)) : $unsigned((~&(8'hba)))));
                      reg6064 <= (8'hb0);
                    end
                  for (forvar6065 = (1'h0); (forvar6065 < (1'h0)); forvar6065 = (forvar6065 + (1'h1)))
                    begin
                      reg6066 <= (^$signed(((forvar6060 >= reg6034) ?
                          {forvar6035} : (~&reg6051))));
                      reg6067 <= ((reg6042[(1'h0):(1'h0)] ?
                              $signed($signed(reg6045)) : (~((8'hab) <= reg6048))) ?
                          $unsigned(forvar6050) : $unsigned(forvar6036));
                      reg6068 <= wire5510;
                    end
                  if ($signed({((8'hb3) == wire5506[(3'h7):(1'h1)])}))
                    begin
                      reg6069 <= $signed((+(reg6024[(3'h4):(1'h1)] ?
                          (reg6037 * forvar6049) : (reg6038 ?
                              reg6048 : forvar6045))));
                      reg6070 <= (^~$signed(reg6039[(4'ha):(3'h4)]));
                      reg6071 <= reg6049[(1'h1):(1'h1)];
                      reg6072 <= $unsigned((($signed((8'hb0)) * reg6032[(3'h5):(3'h5)]) ?
                          wire5506[(3'h5):(3'h5)] : $unsigned($unsigned(reg6071))));
                    end
                  else
                    begin
                      reg6069 <= (reg6052[(3'h5):(3'h5)] ?
                          reg6045[(2'h2):(1'h1)] : $unsigned(reg6042));
                      reg6070 <= $unsigned((8'hac));
                      reg6071 <= ({$unsigned($unsigned(forvar6035))} > (~{((8'ha8) ?
                              wire5508 : reg6029)}));
                    end
                  for (forvar6073 = (1'h0); (forvar6073 < (2'h2)); forvar6073 = (forvar6073 + (1'h1)))
                    begin
                      reg6074 <= (($signed((reg6048 <= reg6071)) && reg6051[(3'h7):(1'h0)]) != (~|reg6066[(4'hb):(4'h9)]));
                      reg6075 <= reg6032;
                      reg6076 <= (reg6037 ?
                          (({reg6022} ? reg6072 : {reg6071}) ?
                              ($signed(forvar6036) >= $unsigned(reg6071)) : ($signed((8'ha9)) << (8'hb3))) : reg6044[(3'h7):(3'h7)]);
                      reg6077 <= $unsigned($unsigned(((reg6046 ?
                          reg6044 : reg6053) == (8'h9c))));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar6078 = (1'h0); (forvar6078 < (1'h1)); forvar6078 = (forvar6078 + (1'h1)))
        begin
          for (forvar6079 = (1'h0); (forvar6079 < (2'h2)); forvar6079 = (forvar6079 + (1'h1)))
            begin
              reg6080 <= (8'ha8);
              for (forvar6081 = (1'h0); (forvar6081 < (2'h2)); forvar6081 = (forvar6081 + (1'h1)))
                begin
                  if (reg6044)
                    begin
                      reg6082 <= $signed($signed($unsigned($unsigned(reg6059))));
                      reg6083 <= (~|(+reg6058));
                    end
                  else
                    begin
                      reg6082 <= reg6049[(2'h3):(2'h3)];
                      reg6083 <= (|$signed($signed($unsigned(reg6022))));
                      reg6084 <= (reg6033[(3'h6):(3'h6)] ~^ $unsigned(reg6025[(2'h2):(2'h2)]));
                    end
                  if ((($unsigned((reg6049 ?
                          (8'hab) : reg6062)) < reg6071[(3'h5):(2'h3)]) ?
                      reg6053[(1'h1):(1'h1)] : reg6041[(2'h3):(2'h3)]))
                    begin
                      reg6085 <= (($signed(reg6076[(4'hd):(4'h9)]) << reg6031) ~^ (($unsigned(reg6070) ?
                              (reg6053 ? reg6031 : reg6028) : (!(8'hb3))) ?
                          forvar6065 : ({reg6054} <<< reg6053)));
                    end
                  else
                    begin
                      reg6085 <= reg6077[(3'h4):(1'h1)];
                    end
                  reg6086 <= {{$signed((~^forvar6018))}};
                end
            end
          for (forvar6087 = (1'h0); (forvar6087 < (2'h3)); forvar6087 = (forvar6087 + (1'h1)))
            begin
              if ((({(wire5507 + (8'h9f))} <= reg6045) ?
                  (&{reg6049[(2'h2):(1'h0)]}) : (forvar6036[(2'h3):(2'h3)] ?
                      (|$signed(reg6045)) : reg6054)))
                begin
                  for (forvar6088 = (1'h0); (forvar6088 < (1'h1)); forvar6088 = (forvar6088 + (1'h1)))
                    begin
                      reg6089 <= ($unsigned($unsigned($unsigned(reg6084))) ?
                          $signed($signed((reg6041 || forvar6065))) : ($unsigned({forvar6055}) ?
                              reg6025 : $signed($signed(reg6054))));
                    end
                  if (forvar6078)
                    begin
                      reg6090 <= ((reg6082 != $unsigned((reg6027 >= reg6072))) ?
                          $signed(forvar6050[(3'h7):(1'h1)]) : reg6053);
                      reg6091 <= reg6044[(4'h8):(4'h8)];
                      reg6092 <= ((^~((!reg6033) ?
                          $unsigned(reg6090) : $signed(reg6047))) << (~|reg6076[(1'h1):(1'h0)]));
                      reg6093 <= ({reg6089[(4'hb):(4'h9)]} * $signed(({reg6039} + wire5507[(3'h4):(1'h1)])));
                    end
                  else
                    begin
                      reg6090 <= (forvar6021[(3'h5):(1'h0)] ~^ (+$signed((reg6082 ~^ reg6042))));
                      reg6091 <= reg6071;
                      reg6092 <= {$unsigned(($unsigned(reg6064) || $unsigned(reg6083)))};
                      reg6093 <= (reg6069[(1'h1):(1'h0)] >>> $unsigned((reg6082[(4'hb):(2'h2)] ?
                          {reg6051} : forvar6073)));
                    end
                  for (forvar6094 = (1'h0); (forvar6094 < (1'h0)); forvar6094 = (forvar6094 + (1'h1)))
                    begin
                      reg6095 <= (~&(reg6028[(3'h5):(3'h5)] ?
                          forvar6049[(1'h0):(1'h0)] : ((-reg6033) ?
                              $signed(reg6025) : (^~(8'haa)))));
                      reg6096 <= forvar6021[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  for (forvar6088 = (1'h0); (forvar6088 < (2'h3)); forvar6088 = (forvar6088 + (1'h1)))
                    begin
                      reg6089 <= $signed((^($unsigned(wire5506) && $signed((8'hb4)))));
                      reg6090 <= (&($unsigned((reg6093 > reg6030)) ?
                          ($signed(forvar6073) ?
                              forvar6078[(1'h1):(1'h0)] : {(8'hb4)}) : $signed(reg6047)));
                    end
                  for (forvar6091 = (1'h0); (forvar6091 < (1'h0)); forvar6091 = (forvar6091 + (1'h1)))
                    begin
                      reg6092 <= ((($signed(reg6032) ?
                              reg6039[(4'h9):(4'h8)] : reg6050) == ((wire6016 >> forvar6026) == (+forvar6055))) ?
                          (~&{(|reg6095)}) : wire6016[(2'h3):(1'h1)]);
                      reg6093 <= {$signed($signed((&reg6046)))};
                    end
                end
            end
          for (forvar6097 = (1'h0); (forvar6097 < (2'h2)); forvar6097 = (forvar6097 + (1'h1)))
            begin
              reg6098 <= forvar6044;
            end
        end
      if ((^(reg6033 > reg6033[(3'h6):(1'h1)])))
        begin
          if (({$unsigned($signed(forvar6018))} ?
              $unsigned(wire5507[(4'ha):(2'h3)]) : reg6090[(1'h0):(1'h0)]))
            begin
              for (forvar6099 = (1'h0); (forvar6099 < (2'h2)); forvar6099 = (forvar6099 + (1'h1)))
                begin
                  for (forvar6100 = (1'h0); (forvar6100 < (1'h1)); forvar6100 = (forvar6100 + (1'h1)))
                    begin
                      reg6101 <= $unsigned((reg6089[(3'h6):(3'h6)] ?
                          ((-reg6075) != forvar6073) : reg6041[(2'h2):(2'h2)]));
                      reg6102 <= (forvar6061 && $signed(forvar6094));
                      reg6103 <= reg6034[(2'h3):(1'h0)];
                    end
                end
              if ($unsigned((((forvar6045 == (8'haa)) | reg6101) != (-(reg6080 ?
                  reg6074 : wire5509)))))
                begin
                  for (forvar6104 = (1'h0); (forvar6104 < (2'h2)); forvar6104 = (forvar6104 + (1'h1)))
                    begin
                      reg6105 <= $signed((($unsigned(reg6068) ?
                          (reg6098 - reg6029) : ((8'hb1) ?
                              reg6062 : forvar6026)) ~^ ((&forvar6078) ?
                          wire5510 : (reg6086 ? forvar6097 : forvar6026))));
                      reg6106 <= $unsigned(reg6098);
                      reg6107 <= $unsigned((~&{$unsigned(reg6046)}));
                    end
                  if ($unsigned($signed((reg6085[(4'h9):(4'h8)] ?
                      (reg6103 + reg6064) : $signed(reg6041)))))
                    begin
                      reg6108 <= ($unsigned((|(reg6052 - forvar6091))) >>> (reg6038[(4'h8):(2'h3)] ?
                          ($signed(reg6076) ?
                              (reg6051 ?
                                  forvar6060 : (8'ha9)) : wire5510) : reg6024[(2'h3):(1'h0)]));
                      reg6109 <= forvar6094[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg6108 <= {((~^{reg6043}) + ((~reg6075) ?
                              (|reg6034) : (reg6105 ? (8'hb6) : reg6049)))};
                      reg6109 <= (~&(~^reg6058));
                    end
                  for (forvar6110 = (1'h0); (forvar6110 < (2'h2)); forvar6110 = (forvar6110 + (1'h1)))
                    begin
                      reg6111 <= $signed($unsigned($signed(forvar6087)));
                      reg6112 <= reg6064;
                    end
                end
              else
                begin
                  if (forvar6099[(2'h2):(1'h0)])
                    begin
                      reg6104 <= (~reg6048[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg6104 <= (^~reg6090[(1'h1):(1'h1)]);
                      reg6105 <= {({((8'hba) ? reg6045 : (8'h9d))} ?
                              reg6062 : reg6024)};
                      reg6106 <= (((~&{reg6045}) || (reg6068[(4'h8):(2'h2)] <= (^~reg6032))) ?
                          reg6040[(4'hb):(4'h8)] : forvar6100);
                    end
                  if (((^~{(~&wire5510)}) ?
                      reg6049 : $signed(((reg6048 >= reg6039) ?
                          $signed(forvar6100) : reg6083[(3'h6):(1'h1)]))))
                    begin
                      reg6107 <= reg6057[(4'hd):(2'h3)];
                    end
                  else
                    begin
                      reg6107 <= $unsigned({reg6068});
                      reg6108 <= $unsigned((|(&(~|(8'hb5)))));
                      reg6109 <= ($unsigned($unsigned((reg6082 ?
                              reg6054 : forvar6100))) ?
                          reg6049[(2'h3):(2'h3)] : $signed($signed($unsigned(wire5509))));
                      reg6110 <= forvar6097[(2'h2):(2'h2)];
                    end
                  for (forvar6111 = (1'h0); (forvar6111 < (1'h1)); forvar6111 = (forvar6111 + (1'h1)))
                    begin
                      reg6112 <= forvar6073;
                      reg6113 <= ((reg6046[(1'h1):(1'h0)] ?
                              reg6095 : $signed($unsigned(wire6016))) ?
                          reg6044 : $signed($signed((reg6069 <<< forvar6079))));
                      reg6114 <= reg6063;
                    end
                  reg6115 <= (reg6022[(3'h5):(2'h3)] | reg6093[(1'h1):(1'h1)]);
                end
            end
          else
            begin
              if ($signed(forvar6094[(1'h1):(1'h0)]))
                begin
                  for (forvar6099 = (1'h0); (forvar6099 < (2'h3)); forvar6099 = (forvar6099 + (1'h1)))
                    begin
                      reg6100 <= ((+reg6047) ?
                          reg6098 : {({(8'hb5)} ?
                                  reg6086 : forvar6111[(3'h4):(2'h2)])});
                      reg6101 <= $signed(($signed(forvar6026[(3'h6):(2'h2)]) > (!(8'h9e))));
                    end
                  if ((&($unsigned(reg6039[(4'h9):(4'h8)]) ?
                      $signed((reg6114 == reg6043)) : (forvar6018[(5'h10):(1'h0)] ?
                          (^reg6070) : (reg6108 == reg6040)))))
                    begin
                      reg6102 <= $signed($signed($unsigned(forvar6061)));
                      reg6103 <= (wire5510[(3'h5):(2'h2)] * $unsigned(reg6096[(2'h2):(2'h2)]));
                      reg6104 <= $unsigned(reg6086[(3'h5):(2'h2)]);
                    end
                  else
                    begin
                      reg6102 <= (($signed(reg6113[(1'h0):(1'h0)]) ?
                          reg6072[(2'h3):(1'h1)] : $unsigned(forvar6065[(4'ha):(1'h1)])) ^ $signed((8'ha4)));
                      reg6103 <= (!({(reg6080 & reg6067)} != ($unsigned(reg6059) <<< (wire5507 ?
                          forvar6055 : wire5507))));
                      reg6104 <= {(~^($signed(reg6022) ?
                              (reg6033 ? reg6105 : reg6067) : (+(8'hb2))))};
                    end
                end
              else
                begin
                  if ({$unsigned($unsigned(forvar6018))})
                    begin
                      reg6099 <= reg6063[(4'hc):(1'h1)];
                      reg6100 <= forvar6104;
                      reg6101 <= $signed((~&$signed(reg6115[(3'h5):(1'h0)])));
                    end
                  else
                    begin
                      reg6099 <= $unsigned(forvar6097);
                      reg6100 <= (-((((8'hb5) ^~ wire5509) < $unsigned(forvar6035)) ?
                          reg6098 : (8'hac)));
                      reg6101 <= forvar6049[(2'h2):(1'h1)];
                      reg6102 <= ((reg6050[(2'h2):(1'h1)] ?
                              forvar6050 : (~^$unsigned(forvar6035))) ?
                          $unsigned(wire5506) : (+$unsigned($unsigned(reg6022))));
                    end
                  if (reg6025)
                    begin
                      reg6103 <= (forvar6049 ^ $signed((~^(!wire5509))));
                      reg6104 <= (&$unsigned(reg6114));
                      reg6105 <= ($signed((8'h9d)) > $unsigned((reg6110 ?
                          reg6114[(2'h3):(1'h1)] : reg6092[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg6103 <= (~|(~&$unsigned((|reg6052))));
                      reg6104 <= reg6106[(3'h5):(3'h4)];
                      reg6105 <= (&reg6030[(3'h5):(2'h3)]);
                      reg6106 <= reg6022;
                    end
                  if ($signed((~^(reg6022[(3'h7):(3'h5)] == $unsigned(reg6032)))))
                    begin
                      reg6107 <= ({$unsigned({(8'ha6)})} ?
                          $unsigned($signed(reg6030[(2'h3):(1'h0)])) : forvar6097[(3'h7):(3'h5)]);
                      reg6108 <= reg6032;
                      reg6109 <= forvar6078;
                      reg6110 <= $unsigned($signed(reg6027[(4'h9):(3'h4)]));
                    end
                  else
                    begin
                      reg6107 <= reg6114[(3'h5):(1'h1)];
                    end
                  if (forvar6100)
                    begin
                      reg6111 <= ((8'hae) ?
                          (&((forvar6088 << forvar6044) >>> $unsigned((8'hac)))) : (reg6101[(4'h9):(3'h7)] ?
                              ((|reg6051) < $signed(forvar6091)) : $signed(forvar6079[(4'ha):(4'h9)])));
                      reg6112 <= $unsigned($unsigned(reg6033));
                      reg6113 <= (!{(^~(~^reg6032))});
                      reg6114 <= $signed(reg6024);
                    end
                  else
                    begin
                      reg6111 <= ($signed(forvar6094[(1'h0):(1'h0)]) ?
                          reg6031 : {forvar6035});
                      reg6112 <= (-(($signed((8'hb7)) << (~reg6068)) ?
                          $signed((forvar6110 ?
                              forvar6055 : wire5509)) : ($unsigned(reg6052) ?
                              (reg6044 ? forvar6020 : forvar6036) : (reg6033 ?
                                  reg6100 : forvar6087))));
                      reg6113 <= wire5509;
                    end
                end
            end
          for (forvar6116 = (1'h0); (forvar6116 < (2'h3)); forvar6116 = (forvar6116 + (1'h1)))
            begin
              if ($unsigned($unsigned(((|reg6072) ?
                  (forvar6091 - reg6093) : reg6100[(1'h1):(1'h1)]))))
                begin
                  if (((-((reg6077 == reg6058) * ((8'ha2) && reg6077))) ?
                      ((~|$unsigned(reg6028)) != ({(8'hb8)} ?
                          ((8'ha8) | reg6093) : $unsigned(reg6084))) : ((reg6031[(2'h2):(2'h2)] <= reg6083[(3'h4):(2'h3)]) ?
                          reg6023 : reg6037)))
                    begin
                      reg6117 <= (+(&(~{forvar6045})));
                      reg6118 <= reg6024[(1'h0):(1'h0)];
                      reg6119 <= $unsigned({$unsigned($unsigned(forvar6035))});
                      reg6120 <= (^($unsigned($signed((8'h9c))) || (^(~^forvar6055))));
                    end
                  else
                    begin
                      reg6117 <= $unsigned(reg6069);
                      reg6118 <= $signed(((|(&reg6098)) ?
                          (^~$unsigned(reg6112)) : $unsigned($signed((8'haf)))));
                    end
                  for (forvar6121 = (1'h0); (forvar6121 < (2'h2)); forvar6121 = (forvar6121 + (1'h1)))
                    begin
                      reg6122 <= (8'ha7);
                      reg6123 <= $signed(reg6032[(3'h4):(1'h1)]);
                      reg6124 <= ($signed($unsigned({(8'hb4)})) ?
                          reg6111[(2'h2):(1'h1)] : ($unsigned(reg6023[(2'h3):(2'h3)]) ?
                              $signed((reg6098 ?
                                  reg6023 : forvar6104)) : $signed(reg6066[(3'h6):(2'h2)])));
                      reg6125 <= (-$unsigned((reg6066[(4'h9):(3'h4)] ?
                          (forvar6060 <= reg6074) : ((8'hae) ~^ forvar6081))));
                    end
                  reg6126 <= (&(8'ha4));
                  for (forvar6127 = (1'h0); (forvar6127 < (2'h3)); forvar6127 = (forvar6127 + (1'h1)))
                    begin
                      reg6128 <= ($signed({(reg6029 ? (8'hab) : reg6054)}) ?
                          ({reg6054[(3'h6):(1'h0)]} ~^ ((~&forvar6097) + {reg6045})) : (+forvar6116[(2'h2):(1'h1)]));
                      reg6129 <= (~reg6076);
                      reg6130 <= reg6069;
                    end
                end
              else
                begin
                  for (forvar6117 = (1'h0); (forvar6117 < (1'h0)); forvar6117 = (forvar6117 + (1'h1)))
                    begin
                      reg6118 <= reg6042;
                      reg6119 <= forvar6073;
                      reg6120 <= forvar6036;
                    end
                  if ((reg6102[(4'hc):(4'hb)] ?
                      {forvar6078} : $signed($unsigned(forvar6091))))
                    begin
                      reg6121 <= (|reg6025);
                      reg6122 <= ((^((reg6074 - (8'ha3)) < $signed(forvar6060))) ?
                          reg6057[(2'h3):(2'h2)] : forvar6026);
                      reg6123 <= $signed((((forvar6036 ? reg6031 : forvar6020) ?
                              (~|reg6096) : (reg6115 ? reg6068 : (8'ha7))) ?
                          (~|(forvar6078 ?
                              reg6067 : reg6076)) : ({reg6066} * $unsigned(reg6051))));
                      reg6124 <= (reg6130[(2'h3):(2'h2)] < $unsigned(($signed((8'hac)) || reg6028[(3'h4):(1'h1)])));
                    end
                  else
                    begin
                      reg6121 <= (reg6106 == (reg6071 ? reg6052 : reg6075));
                      reg6122 <= (&reg6022[(3'h4):(3'h4)]);
                    end
                end
              if ((|(reg6025[(2'h2):(1'h1)] | ((reg6064 ?
                  reg6080 : forvar6088) <= ((8'hab) ? reg6054 : (8'hb0))))))
                begin
                  for (forvar6131 = (1'h0); (forvar6131 < (2'h3)); forvar6131 = (forvar6131 + (1'h1)))
                    begin
                      reg6132 <= reg6115;
                    end
                  if (forvar6116[(3'h5):(2'h3)])
                    begin
                      reg6133 <= reg6098;
                      reg6134 <= ($signed(reg6091) | (8'hab));
                      reg6135 <= (&$signed((-(reg6063 < forvar6091))));
                    end
                  else
                    begin
                      reg6133 <= forvar6091;
                    end
                  for (forvar6136 = (1'h0); (forvar6136 < (1'h1)); forvar6136 = (forvar6136 + (1'h1)))
                    begin
                      reg6137 <= ((wire5506[(2'h3):(2'h3)] >= $signed($unsigned(reg6134))) >= (!reg6102[(2'h3):(1'h0)]));
                      reg6138 <= reg6029[(4'he):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar6131 = (1'h0); (forvar6131 < (2'h2)); forvar6131 = (forvar6131 + (1'h1)))
                    begin
                      reg6132 <= forvar6065[(2'h2):(1'h0)];
                      reg6133 <= (~&{$signed(((8'hb2) + reg6048))});
                      reg6134 <= (reg6105[(1'h1):(1'h1)] ?
                          reg6068[(4'hf):(3'h5)] : (reg6107 ?
                              {(-forvar6045)} : forvar6019[(1'h0):(1'h0)]));
                    end
                  for (forvar6135 = (1'h0); (forvar6135 < (2'h3)); forvar6135 = (forvar6135 + (1'h1)))
                    begin
                      reg6136 <= reg6121;
                    end
                  for (forvar6137 = (1'h0); (forvar6137 < (2'h2)); forvar6137 = (forvar6137 + (1'h1)))
                    begin
                      reg6138 <= wire6016[(3'h5):(1'h1)];
                    end
                  if ($unsigned($signed((+(+reg6037)))))
                    begin
                      reg6139 <= $unsigned(reg6101);
                      reg6140 <= reg6034[(3'h5):(1'h0)];
                      reg6141 <= $unsigned(reg6040);
                      reg6142 <= reg6063;
                    end
                  else
                    begin
                      reg6139 <= reg6098[(4'ha):(3'h6)];
                      reg6140 <= $signed(reg6135);
                      reg6141 <= reg6076[(3'h7):(2'h2)];
                      reg6142 <= $signed(reg6077[(2'h2):(1'h0)]);
                    end
                end
              if (((~|((~reg6112) ?
                  reg6076 : reg6092[(1'h1):(1'h1)])) >> (|((8'ha2) ?
                  reg6077 : (reg6104 ? reg6071 : (8'had))))))
                begin
                  for (forvar6143 = (1'h0); (forvar6143 < (2'h3)); forvar6143 = (forvar6143 + (1'h1)))
                    begin
                      reg6144 <= (wire6016 ?
                          $unsigned($unsigned((8'hb4))) : forvar6019[(1'h0):(1'h0)]);
                      reg6145 <= $unsigned((!(forvar6018[(4'hf):(4'he)] || ((8'h9f) ?
                          reg6047 : forvar6079))));
                      reg6146 <= {(reg6052 ?
                              (~^$unsigned(forvar6121)) : (~reg6034))};
                    end
                end
              else
                begin
                  for (forvar6143 = (1'h0); (forvar6143 < (1'h0)); forvar6143 = (forvar6143 + (1'h1)))
                    begin
                      reg6144 <= {reg6108};
                    end
                  for (forvar6145 = (1'h0); (forvar6145 < (2'h2)); forvar6145 = (forvar6145 + (1'h1)))
                    begin
                      reg6146 <= forvar6117[(1'h1):(1'h1)];
                      reg6147 <= ((^forvar6020[(2'h2):(1'h0)]) ?
                          $signed(($unsigned(forvar6111) ?
                              $unsigned(reg6041) : (!forvar6121))) : (((!(8'hb8)) - wire5508[(1'h1):(1'h1)]) >> ({(8'hb5)} >>> $signed(forvar6137))));
                      reg6148 <= ({(!(reg6032 >>> reg6106))} ?
                          forvar6117[(3'h5):(2'h2)] : reg6100);
                    end
                  for (forvar6149 = (1'h0); (forvar6149 < (1'h1)); forvar6149 = (forvar6149 + (1'h1)))
                    begin
                      reg6150 <= {forvar6079};
                      reg6151 <= $unsigned($unsigned((^~(reg6126 ?
                          reg6071 : reg6121))));
                      reg6152 <= $signed(($signed((forvar6127 + reg6058)) ?
                          $unsigned((^reg6054)) : forvar6061));
                      reg6153 <= {reg6108[(2'h2):(1'h1)]};
                    end
                end
              reg6154 <= ((reg6108 - (~^reg6098[(5'h10):(1'h1)])) <<< (~^((reg6123 ?
                      reg6101 : reg6141) ?
                  (reg6068 & reg6029) : $unsigned(reg6114))));
            end
          if ($signed({($unsigned(forvar6078) ?
                  $signed(forvar6021) : reg6128[(4'hc):(3'h5)])}))
            begin
              for (forvar6155 = (1'h0); (forvar6155 < (1'h0)); forvar6155 = (forvar6155 + (1'h1)))
                begin
                  for (forvar6156 = (1'h0); (forvar6156 < (1'h1)); forvar6156 = (forvar6156 + (1'h1)))
                    begin
                      reg6157 <= $signed((|((^reg6066) ?
                          (forvar6094 ? forvar6060 : reg6052) : (reg6151 ?
                              reg6076 : reg6044))));
                      reg6158 <= (~^(forvar6094 ?
                          $signed($unsigned(reg6098)) : reg6058[(3'h5):(3'h4)]));
                    end
                  for (forvar6159 = (1'h0); (forvar6159 < (2'h2)); forvar6159 = (forvar6159 + (1'h1)))
                    begin
                      reg6160 <= reg6066[(1'h1):(1'h0)];
                      reg6161 <= $unsigned(($unsigned(reg6122) >> $signed((forvar6143 ?
                          reg6128 : reg6108))));
                      reg6162 <= $signed($unsigned({$signed(reg6102)}));
                      reg6163 <= reg6071;
                    end
                  for (forvar6164 = (1'h0); (forvar6164 < (2'h2)); forvar6164 = (forvar6164 + (1'h1)))
                    begin
                      reg6165 <= reg6120;
                      reg6166 <= reg6029;
                      reg6167 <= ($unsigned(reg6023) != reg6044[(2'h2):(1'h1)]);
                    end
                  for (forvar6168 = (1'h0); (forvar6168 < (1'h0)); forvar6168 = (forvar6168 + (1'h1)))
                    begin
                      reg6169 <= (reg6033 ?
                          ($unsigned((reg6062 && reg6142)) > reg6084) : (8'h9c));
                      reg6170 <= forvar6079;
                      reg6171 <= forvar6087;
                    end
                end
            end
          else
            begin
              for (forvar6155 = (1'h0); (forvar6155 < (1'h0)); forvar6155 = (forvar6155 + (1'h1)))
                begin
                  for (forvar6156 = (1'h0); (forvar6156 < (2'h3)); forvar6156 = (forvar6156 + (1'h1)))
                    begin
                      reg6157 <= (forvar6099[(2'h2):(2'h2)] ?
                          ((8'ha5) * $unsigned(reg6118)) : $signed((~(reg6115 >> reg6132))));
                      reg6158 <= (&($unsigned($unsigned(forvar6156)) < ((reg6030 ?
                              reg6139 : reg6082) ?
                          forvar6049[(1'h1):(1'h1)] : reg6123)));
                      reg6159 <= (^reg6160);
                      reg6160 <= $unsigned({reg6030});
                    end
                  for (forvar6161 = (1'h0); (forvar6161 < (1'h0)); forvar6161 = (forvar6161 + (1'h1)))
                    begin
                      reg6162 <= (!reg6024);
                      reg6163 <= {$unsigned(reg6135[(1'h1):(1'h1)])};
                      reg6164 <= ((+($signed(forvar6018) >= (~|forvar6099))) <<< (~|(^{reg6089})));
                    end
                end
              for (forvar6165 = (1'h0); (forvar6165 < (1'h0)); forvar6165 = (forvar6165 + (1'h1)))
                begin
                  for (forvar6166 = (1'h0); (forvar6166 < (2'h2)); forvar6166 = (forvar6166 + (1'h1)))
                    begin
                      reg6167 <= ({{reg6110}} ?
                          (~^(((8'hb3) != reg6099) > reg6123)) : $signed(forvar6091[(4'hd):(4'hb)]));
                      reg6168 <= ($unsigned($signed($signed((8'hb8)))) ?
                          (forvar6073 ?
                              $unsigned(((8'hb1) <<< reg6076)) : $signed((reg6147 <= forvar6155))) : reg6062);
                    end
                end
              reg6169 <= $signed($unsigned(reg6165[(3'h4):(2'h3)]));
              for (forvar6170 = (1'h0); (forvar6170 < (1'h1)); forvar6170 = (forvar6170 + (1'h1)))
                begin
                  for (forvar6171 = (1'h0); (forvar6171 < (2'h3)); forvar6171 = (forvar6171 + (1'h1)))
                    begin
                      reg6172 <= forvar6079;
                      reg6173 <= forvar6121;
                      reg6174 <= reg6148;
                      reg6175 <= ({(+reg6076[(4'hd):(4'ha)])} >> $unsigned(($unsigned(reg6030) | (^~forvar6091))));
                    end
                  reg6176 <= $unsigned(reg6129);
                end
            end
          for (forvar6177 = (1'h0); (forvar6177 < (1'h1)); forvar6177 = (forvar6177 + (1'h1)))
            begin
              for (forvar6178 = (1'h0); (forvar6178 < (2'h2)); forvar6178 = (forvar6178 + (1'h1)))
                begin
                  for (forvar6179 = (1'h0); (forvar6179 < (1'h0)); forvar6179 = (forvar6179 + (1'h1)))
                    begin
                      reg6180 <= (reg6159 ?
                          reg6115 : $unsigned(((reg6041 ? reg6080 : reg6135) ?
                              $signed((8'h9c)) : (~reg6138))));
                      reg6181 <= reg6090;
                      reg6182 <= $unsigned($signed(((reg6086 || forvar6116) == forvar6060[(3'h6):(3'h5)])));
                    end
                  if ($unsigned(({reg6037[(4'hc):(3'h5)]} ?
                      $signed(forvar6099[(1'h1):(1'h1)]) : $unsigned(forvar6117))))
                    begin
                      reg6183 <= $unsigned(reg6117);
                      reg6184 <= (reg6075 ?
                          forvar6166[(1'h1):(1'h0)] : $unsigned(((|forvar6159) << (^reg6092))));
                      reg6185 <= (~&{((+reg6181) >> (reg6068 ?
                              reg6053 : reg6165))});
                    end
                  else
                    begin
                      reg6183 <= $signed((forvar6131 ?
                          ($unsigned(reg6105) | (~reg6031)) : (reg6095[(4'hb):(4'h8)] << (-reg6110))));
                    end
                  for (forvar6186 = (1'h0); (forvar6186 < (1'h1)); forvar6186 = (forvar6186 + (1'h1)))
                    begin
                      reg6187 <= forvar6061;
                      reg6188 <= reg6140;
                      reg6189 <= reg6033;
                    end
                end
              reg6190 <= (!reg6147);
              if ((reg6063[(4'h9):(1'h0)] >= $signed($signed((forvar6137 * reg6106)))))
                begin
                  for (forvar6191 = (1'h0); (forvar6191 < (2'h3)); forvar6191 = (forvar6191 + (1'h1)))
                    begin
                      reg6192 <= $signed(reg6089);
                      reg6193 <= (+($signed((forvar6165 ?
                          reg6172 : (8'h9e))) << ((reg6046 ^~ reg6189) ?
                          (forvar6019 ~^ forvar6136) : ((8'ha5) && forvar6050))));
                      reg6194 <= forvar6104[(1'h0):(1'h0)];
                    end
                  for (forvar6195 = (1'h0); (forvar6195 < (2'h2)); forvar6195 = (forvar6195 + (1'h1)))
                    begin
                      reg6196 <= (~&(($signed(reg6039) >= ((8'had) ?
                          forvar6104 : forvar6121)) >= ((reg6027 ?
                              (8'hb0) : forvar6116) ?
                          $signed((8'h9e)) : (^reg6042))));
                      reg6197 <= {reg6164};
                    end
                  for (forvar6198 = (1'h0); (forvar6198 < (1'h1)); forvar6198 = (forvar6198 + (1'h1)))
                    begin
                      reg6199 <= $signed($unsigned({(-(8'h9e))}));
                      reg6200 <= reg6032[(3'h4):(2'h2)];
                      reg6201 <= (((reg6096[(3'h5):(3'h4)] * {reg6091}) < $signed({forvar6156})) ?
                          (8'ha6) : reg6058);
                    end
                  for (forvar6202 = (1'h0); (forvar6202 < (2'h3)); forvar6202 = (forvar6202 + (1'h1)))
                    begin
                      reg6203 <= (reg6125[(1'h0):(1'h0)] ?
                          (-forvar6020) : $signed((!$signed(reg6083))));
                      reg6204 <= reg6043;
                      reg6205 <= ($signed($signed((^(8'haa)))) < reg6158);
                    end
                end
              else
                begin
                  if ($signed($signed(reg6022)))
                    begin
                      reg6191 <= ((reg6071 == $unsigned((|reg6110))) ?
                          (~^(&(^(8'ha6)))) : forvar6060[(3'h7):(3'h7)]);
                      reg6192 <= (($signed((reg6032 ?
                          (8'ha2) : reg6172)) && (~|reg6163)) == reg6205[(3'h4):(1'h0)]);
                      reg6193 <= $unsigned({reg6033[(1'h1):(1'h0)]});
                    end
                  else
                    begin
                      reg6191 <= ({(forvar6177 && $signed(reg6151))} ?
                          (8'hb4) : ($signed((wire5509 + reg6046)) * ((+reg6204) != (reg6100 ?
                              reg6185 : reg6067))));
                    end
                  if ((^~{(+(reg6114 ? reg6134 : reg6057))}))
                    begin
                      reg6194 <= $unsigned(forvar6137[(1'h0):(1'h0)]);
                      reg6195 <= {($unsigned((reg6105 ?
                              (8'hba) : reg6189)) & $unsigned((~(8'hb3))))};
                      reg6196 <= (~^reg6182[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg6194 <= (reg6092 ?
                          (forvar6179[(1'h1):(1'h0)] ?
                              reg6175 : ($signed(forvar6168) ?
                                  reg6091[(1'h1):(1'h0)] : (forvar6100 >= forvar6159))) : ((reg6040[(1'h0):(1'h0)] ?
                              {forvar6045} : (reg6112 ?
                                  reg6129 : reg6196)) ^ reg6071[(1'h0):(1'h0)]));
                    end
                end
              reg6206 <= forvar6020[(2'h3):(1'h1)];
            end
        end
      else
        begin
          if ({reg6192})
            begin
              if ((8'haa))
                begin
                  if (reg6114)
                    begin
                      reg6099 <= (~|((forvar6019 && (reg6163 ?
                          forvar6136 : forvar6191)) + $unsigned($signed(reg6199))));
                      reg6100 <= (8'hb0);
                      reg6101 <= (reg6180[(1'h1):(1'h0)] ?
                          ($signed(reg6075) ?
                              {(forvar6161 && reg6123)} : $unsigned((^~(8'ha6)))) : reg6067);
                    end
                  else
                    begin
                      reg6099 <= reg6140[(2'h2):(2'h2)];
                      reg6100 <= (forvar6060 ^ (^reg6062[(4'h9):(3'h4)]));
                    end
                end
              else
                begin
                  for (forvar6099 = (1'h0); (forvar6099 < (1'h1)); forvar6099 = (forvar6099 + (1'h1)))
                    begin
                      reg6100 <= reg6070;
                      reg6101 <= $signed($signed((|((8'h9c) ?
                          reg6075 : reg6153))));
                    end
                end
              if (((&((reg6197 || reg6080) > {(8'ha9)})) ?
                  forvar6050 : (8'haa)))
                begin
                  if ($signed(($signed((&reg6106)) * reg6069[(3'h6):(1'h1)])))
                    begin
                      reg6102 <= ({({wire5508} - (reg6067 - reg6069))} ?
                          reg6057[(4'hc):(3'h6)] : $signed((|((8'h9e) ?
                              reg6203 : (8'ha0)))));
                    end
                  else
                    begin
                      reg6102 <= $signed((~|reg6174[(2'h2):(1'h0)]));
                      reg6103 <= wire5510;
                    end
                end
              else
                begin
                  if ($unsigned($signed($unsigned((^reg6206)))))
                    begin
                      reg6102 <= forvar6161[(3'h6):(3'h6)];
                      reg6103 <= {{$signed((reg6191 < reg6059))}};
                    end
                  else
                    begin
                      reg6102 <= (^$signed(($signed(forvar6078) ?
                          {reg6203} : {reg6091})));
                    end
                end
            end
          else
            begin
              for (forvar6099 = (1'h0); (forvar6099 < (1'h1)); forvar6099 = (forvar6099 + (1'h1)))
                begin
                  for (forvar6100 = (1'h0); (forvar6100 < (2'h2)); forvar6100 = (forvar6100 + (1'h1)))
                    begin
                      reg6101 <= $unsigned($signed(($unsigned(forvar6164) - reg6030[(2'h3):(2'h2)])));
                      reg6102 <= reg6030;
                      reg6103 <= $signed((|(8'hb4)));
                      reg6104 <= $unsigned(reg6080);
                    end
                end
              for (forvar6105 = (1'h0); (forvar6105 < (2'h2)); forvar6105 = (forvar6105 + (1'h1)))
                begin
                  for (forvar6106 = (1'h0); (forvar6106 < (1'h1)); forvar6106 = (forvar6106 + (1'h1)))
                    begin
                      reg6107 <= $unsigned(($signed(forvar6195) ?
                          reg6053 : (~$unsigned(reg6175))));
                      reg6108 <= $signed((forvar6094 << (^$signed(reg6130))));
                      reg6109 <= ((!({reg6132} ?
                              (~|reg6047) : (reg6206 ? wire5508 : (8'ha1)))) ?
                          (reg6059 ?
                              forvar6161 : $signed(reg6128)) : $unsigned(reg6101));
                    end
                end
            end
          reg6110 <= {reg6040[(3'h5):(1'h0)]};
          for (forvar6111 = (1'h0); (forvar6111 < (2'h3)); forvar6111 = (forvar6111 + (1'h1)))
            begin
              if ((forvar6020[(3'h4):(1'h0)] - $unsigned(((8'ha0) & (reg6022 ^~ reg6041)))))
                begin
                  if ($unsigned($signed(reg6108)))
                    begin
                      reg6112 <= ((((reg6111 ? reg6051 : reg6190) ?
                              (-reg6206) : (|forvar6019)) | ((^~(8'ha5)) ?
                              (forvar6170 ^~ reg6133) : ((8'ha5) ^ reg6038))) ?
                          $signed(forvar6065[(4'hd):(4'h9)]) : forvar6018[(3'h5):(1'h0)]);
                      reg6113 <= ($signed(($signed(forvar6145) ~^ (reg6139 <<< reg6159))) ?
                          $signed(reg6194[(4'hb):(4'hb)]) : reg6104[(2'h3):(2'h2)]);
                      reg6114 <= ($signed(forvar6137[(2'h3):(1'h1)]) ^ $signed((~^$signed((8'hac)))));
                      reg6115 <= (reg6067[(4'h9):(4'h8)] ?
                          forvar6094[(3'h5):(2'h3)] : (8'h9e));
                    end
                  else
                    begin
                      reg6112 <= (reg6034 ?
                          forvar6136[(4'h8):(1'h0)] : {forvar6155});
                      reg6113 <= ((8'ha1) ? forvar6159 : (8'h9d));
                      reg6114 <= $signed(reg6135[(4'h8):(2'h3)]);
                    end
                  if (reg6203)
                    begin
                      reg6116 <= (forvar6168 ?
                          $unsigned($unsigned((forvar6104 <<< forvar6106))) : ($signed((~&reg6173)) || $signed((forvar6186 ?
                              reg6028 : reg6095))));
                      reg6117 <= reg6072[(3'h6):(3'h4)];
                      reg6118 <= $unsigned((forvar6161 ?
                          ((+wire5507) <= (~^forvar6117)) : ($signed(reg6038) ?
                              $signed(reg6072) : reg6205)));
                      reg6119 <= $signed((~|reg6199));
                    end
                  else
                    begin
                      reg6116 <= (((&(reg6025 ?
                              (8'ha8) : reg6111)) + (reg6034[(3'h7):(1'h1)] ?
                              (reg6101 + forvar6061) : ((8'hb4) ?
                                  (8'haf) : reg6157))) ?
                          reg6192[(3'h4):(2'h3)] : wire5508[(4'h8):(3'h7)]);
                      reg6117 <= ($signed($signed($unsigned(reg6092))) ?
                          (&(~|reg6053)) : ((~^reg6096[(2'h2):(2'h2)]) ?
                              reg6132 : (forvar6171[(4'h9):(2'h2)] ?
                                  reg6051 : $unsigned(forvar6143))));
                      reg6118 <= reg6031[(4'h8):(1'h1)];
                    end
                  for (forvar6120 = (1'h0); (forvar6120 < (1'h0)); forvar6120 = (forvar6120 + (1'h1)))
                    begin
                      reg6121 <= ((reg6167[(2'h3):(1'h1)] ?
                          reg6053 : {(reg6051 ?
                                  reg6107 : reg6191)}) ~^ $signed((8'ha2)));
                    end
                end
              else
                begin
                  reg6112 <= forvar6050;
                end
            end
          if ($signed(reg6106[(1'h0):(1'h0)]))
            begin
              if ((-reg6175[(2'h3):(2'h3)]))
                begin
                  reg6122 <= $unsigned(wire5509[(4'ha):(3'h6)]);
                  for (forvar6123 = (1'h0); (forvar6123 < (2'h2)); forvar6123 = (forvar6123 + (1'h1)))
                    begin
                      reg6124 <= reg6185[(4'he):(2'h2)];
                      reg6125 <= {$signed(($unsigned(reg6161) >= $unsigned(reg6041)))};
                    end
                end
              else
                begin
                  if ((~|{forvar6159}))
                    begin
                      reg6122 <= forvar6137[(4'hb):(2'h3)];
                      reg6123 <= (~|reg6112[(3'h5):(3'h5)]);
                      reg6124 <= forvar6079[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg6122 <= {forvar6127[(3'h6):(2'h2)]};
                      reg6123 <= {$signed(($signed(reg6125) ?
                              reg6189[(1'h1):(1'h1)] : (reg6029 & (8'h9e))))};
                      reg6124 <= $unsigned((($signed((8'h9f)) ?
                          $unsigned(forvar6178) : reg6066) < (reg6095 ?
                          (wire5510 != reg6151) : forvar6050)));
                      reg6125 <= $signed(reg6164);
                    end
                end
              for (forvar6126 = (1'h0); (forvar6126 < (2'h3)); forvar6126 = (forvar6126 + (1'h1)))
                begin
                  for (forvar6127 = (1'h0); (forvar6127 < (1'h1)); forvar6127 = (forvar6127 + (1'h1)))
                    begin
                      reg6128 <= ($unsigned($signed($signed(reg6130))) && $unsigned((|(forvar6155 | (8'ha0)))));
                    end
                  for (forvar6129 = (1'h0); (forvar6129 < (2'h3)); forvar6129 = (forvar6129 + (1'h1)))
                    begin
                      reg6130 <= (&($signed(reg6150) & ($signed((8'h9f)) ?
                          reg6135 : reg6153)));
                    end
                end
              reg6131 <= reg6154[(4'hd):(4'h9)];
            end
          else
            begin
              if ((reg6058 ?
                  $signed({(~|(8'ha9))}) : (reg6187 ^~ {(forvar6111 == reg6159)})))
                begin
                  for (forvar6122 = (1'h0); (forvar6122 < (1'h0)); forvar6122 = (forvar6122 + (1'h1)))
                    begin
                      reg6123 <= $unsigned((reg6115[(4'ha):(3'h7)] ?
                          $unsigned($signed(reg6158)) : $unsigned($unsigned(reg6190))));
                      reg6124 <= forvar6165[(2'h3):(1'h0)];
                      reg6125 <= reg6074[(4'he):(4'ha)];
                      reg6126 <= $unsigned(((|$signed(reg6090)) ?
                          $signed($signed(reg6033)) : (~(reg6050 ?
                              forvar6143 : reg6141))));
                    end
                end
              else
                begin
                  for (forvar6122 = (1'h0); (forvar6122 < (2'h2)); forvar6122 = (forvar6122 + (1'h1)))
                    begin
                      reg6123 <= reg6192;
                      reg6124 <= $unsigned($signed({{reg6023}}));
                      reg6125 <= $unsigned((8'ha6));
                    end
                  if (reg6201)
                    begin
                      reg6126 <= reg6199[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg6126 <= (8'hb5);
                      reg6127 <= reg6170[(2'h3):(1'h0)];
                      reg6128 <= (reg6201[(4'ha):(1'h0)] >> (8'haa));
                    end
                  if (reg6160[(3'h4):(1'h1)])
                    begin
                      reg6129 <= $unsigned(reg6190[(4'h9):(2'h2)]);
                      reg6130 <= ($signed((+(forvar6161 ?
                              (8'hb0) : forvar6186))) ?
                          reg6044[(2'h3):(1'h0)] : ((^(reg6057 ~^ (8'h9c))) == $signed($signed(reg6106))));
                      reg6131 <= $unsigned((^reg6076[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg6129 <= $unsigned((~^{$unsigned((8'hb2))}));
                      reg6130 <= (~^reg6192[(3'h5):(3'h5)]);
                    end
                  if (reg6151)
                    begin
                      reg6132 <= $signed(($unsigned($signed(forvar6060)) && reg6068[(3'h7):(1'h0)]));
                      reg6133 <= $unsigned($signed(reg6168[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg6132 <= reg6175[(1'h0):(1'h0)];
                    end
                end
              for (forvar6134 = (1'h0); (forvar6134 < (2'h2)); forvar6134 = (forvar6134 + (1'h1)))
                begin
                  for (forvar6135 = (1'h0); (forvar6135 < (1'h0)); forvar6135 = (forvar6135 + (1'h1)))
                    begin
                      reg6136 <= (~|wire5508);
                      reg6137 <= reg6136;
                      reg6138 <= $signed(reg6052);
                    end
                end
              if ($signed((~$unsigned({(8'hb8)}))))
                begin
                  for (forvar6139 = (1'h0); (forvar6139 < (1'h1)); forvar6139 = (forvar6139 + (1'h1)))
                    begin
                      reg6140 <= reg6199;
                      reg6141 <= reg6152;
                      reg6142 <= $unsigned(reg6159);
                    end
                end
              else
                begin
                  for (forvar6139 = (1'h0); (forvar6139 < (2'h3)); forvar6139 = (forvar6139 + (1'h1)))
                    begin
                      reg6140 <= (({(^reg6030)} ?
                          forvar6079 : (~&(reg6049 + reg6181))) >= reg6163);
                      reg6141 <= ({{$unsigned(reg6166)}} ?
                          $unsigned(($unsigned(reg6199) || reg6022)) : forvar6136);
                    end
                end
            end
        end
      reg6207 <= (-($signed(reg6024[(3'h4):(2'h3)]) && $signed(reg6106)));
      for (forvar6208 = (1'h0); (forvar6208 < (1'h1)); forvar6208 = (forvar6208 + (1'h1)))
        begin
          for (forvar6209 = (1'h0); (forvar6209 < (2'h3)); forvar6209 = (forvar6209 + (1'h1)))
            begin
              for (forvar6210 = (1'h0); (forvar6210 < (1'h1)); forvar6210 = (forvar6210 + (1'h1)))
                begin
                  reg6211 <= $unsigned(reg6069[(3'h4):(3'h4)]);
                end
              for (forvar6212 = (1'h0); (forvar6212 < (1'h0)); forvar6212 = (forvar6212 + (1'h1)))
                begin
                  if ($signed(reg6105[(3'h4):(2'h2)]))
                    begin
                      reg6213 <= reg6096;
                      reg6214 <= forvar6035;
                      reg6215 <= $signed(reg6114);
                      reg6216 <= reg6194[(3'h6):(2'h3)];
                    end
                  else
                    begin
                      reg6213 <= (8'hb1);
                      reg6214 <= reg6189[(2'h2):(1'h0)];
                      reg6215 <= $unsigned((8'ha8));
                    end
                  reg6217 <= {$signed(((-reg6050) ?
                          {(8'hae)} : $unsigned(reg6080)))};
                end
            end
        end
    end
  assign wire6218 = $signed($unsigned((~&reg6172[(2'h3):(2'h2)])));
  always
    @(posedge clk) begin
      for (forvar6219 = (1'h0); (forvar6219 < (2'h2)); forvar6219 = (forvar6219 + (1'h1)))
        begin
          for (forvar6220 = (1'h0); (forvar6220 < (2'h2)); forvar6220 = (forvar6220 + (1'h1)))
            begin
              if ((reg6189[(2'h2):(1'h1)] > ($unsigned(wire5506) ?
                  ({forvar6155} ?
                      (^~reg6130) : (reg6118 ?
                          forvar6049 : (8'hb3))) : ($unsigned(forvar6045) || reg6089[(4'h9):(3'h4)]))))
                begin
                  for (forvar6221 = (1'h0); (forvar6221 < (2'h3)); forvar6221 = (forvar6221 + (1'h1)))
                    begin
                      reg6222 <= $unsigned((8'hb1));
                      reg6223 <= reg6139[(4'h9):(3'h5)];
                    end
                  if (((($signed(reg6024) ?
                          $signed(reg6103) : $unsigned(forvar6065)) <= (reg6222[(4'h9):(3'h6)] + (^reg6128))) ?
                      (((forvar6208 ? reg6167 : forvar6104) ?
                          $signed(reg6110) : {(8'h9c)}) < ({forvar6178} ~^ ((8'ha5) <= reg6146))) : $unsigned(forvar6145[(3'h4):(1'h0)])))
                    begin
                      reg6224 <= reg6091;
                      reg6225 <= reg6023;
                      reg6226 <= forvar6131;
                      reg6227 <= forvar6198[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg6224 <= (~(~&$unsigned((forvar6019 ^ reg6130))));
                    end
                  for (forvar6228 = (1'h0); (forvar6228 < (1'h0)); forvar6228 = (forvar6228 + (1'h1)))
                    begin
                      reg6229 <= (~&(|((8'hac) > (wire6218 & reg6136))));
                      reg6230 <= (~^reg6223[(1'h1):(1'h1)]);
                      reg6231 <= $signed(((8'hab) ?
                          (reg6123[(4'hb):(4'ha)] ?
                              (forvar6055 < (8'hae)) : $signed(reg6184)) : ((-reg6122) ?
                              (8'hab) : $signed((8'hb5)))));
                    end
                end
              else
                begin
                  for (forvar6221 = (1'h0); (forvar6221 < (2'h3)); forvar6221 = (forvar6221 + (1'h1)))
                    begin
                      reg6222 <= {$signed((reg6086[(3'h4):(2'h3)] ?
                              $unsigned(forvar6131) : reg6083))};
                      reg6223 <= ((forvar6123 && {reg6159}) <<< ($unsigned(reg6216[(1'h0):(1'h0)]) ?
                          (+$signed(forvar6120)) : $signed((forvar6209 >= forvar6209))));
                    end
                end
              for (forvar6232 = (1'h0); (forvar6232 < (2'h2)); forvar6232 = (forvar6232 + (1'h1)))
                begin
                  reg6233 <= forvar6049;
                  for (forvar6234 = (1'h0); (forvar6234 < (2'h2)); forvar6234 = (forvar6234 + (1'h1)))
                    begin
                      reg6235 <= (reg6153[(2'h3):(2'h2)] ~^ (((reg6082 ?
                              reg6190 : reg6052) ?
                          forvar6219[(2'h2):(1'h0)] : $unsigned(forvar6209)) >> reg6204[(1'h1):(1'h0)]));
                      reg6236 <= ((~^(reg6201[(1'h0):(1'h0)] | $unsigned((8'hb4)))) ^ $signed(reg6076[(3'h7):(3'h5)]));
                      reg6237 <= $signed($unsigned(forvar6111[(1'h0):(1'h0)]));
                      reg6238 <= forvar6121[(3'h7):(3'h7)];
                    end
                  if ((^~$unsigned($signed(wire5506))))
                    begin
                      reg6239 <= ($unsigned((^{reg6086})) ?
                          (^(~^$unsigned(reg6116))) : reg6174[(1'h1):(1'h0)]);
                      reg6240 <= (!reg6216);
                      reg6241 <= ((+$unsigned($unsigned(reg6238))) <= forvar6100[(4'h8):(3'h5)]);
                    end
                  else
                    begin
                      reg6239 <= {((reg6151[(3'h5):(1'h1)] ?
                                  (reg6113 ?
                                      reg6227 : reg6096) : {forvar6110}) ?
                              $signed($signed(reg6038)) : $unsigned((^~reg6121)))};
                      reg6240 <= reg6053;
                      reg6241 <= $signed(forvar6123[(2'h3):(1'h1)]);
                      reg6242 <= forvar6018[(4'hf):(3'h5)];
                    end
                end
              if (forvar6106)
                begin
                  reg6243 <= forvar6164;
                  for (forvar6244 = (1'h0); (forvar6244 < (2'h2)); forvar6244 = (forvar6244 + (1'h1)))
                    begin
                      reg6245 <= reg6111[(2'h2):(2'h2)];
                      reg6246 <= $signed({($unsigned(reg6077) ^ $signed(reg6237))});
                      reg6247 <= {$signed((~&(~^forvar6221)))};
                      reg6248 <= reg6148;
                    end
                  if ((~({reg6225[(3'h6):(3'h4)]} ?
                      reg6032 : ({reg6133} ~^ (reg6241 < forvar6045)))))
                    begin
                      reg6249 <= (&$signed($signed(forvar6026)));
                      reg6250 <= $signed({((|(8'ha5)) ?
                              reg6168[(3'h5):(3'h4)] : reg6187)});
                      reg6251 <= reg6168[(2'h2):(1'h1)];
                      reg6252 <= $unsigned(({(reg6173 > reg6051)} < (^(~|reg6090))));
                    end
                  else
                    begin
                      reg6249 <= (8'had);
                      reg6250 <= (($signed(reg6199[(1'h1):(1'h1)]) - (^(&forvar6131))) ?
                          (forvar6110[(4'h8):(4'h8)] >= $signed((+reg6229))) : (((!reg6038) & (wire5510 ?
                              forvar6210 : forvar6135)) <= ($unsigned(reg6174) ?
                              forvar6191 : $signed(forvar6018))));
                    end
                  for (forvar6253 = (1'h0); (forvar6253 < (1'h0)); forvar6253 = (forvar6253 + (1'h1)))
                    begin
                      reg6254 <= reg6211;
                      reg6255 <= {($unsigned((reg6147 ? reg6105 : reg6223)) ?
                              reg6213[(4'hd):(2'h3)] : $unsigned(forvar6186))};
                      reg6256 <= $unsigned($unsigned({$signed(reg6154)}));
                    end
                end
              else
                begin
                  for (forvar6243 = (1'h0); (forvar6243 < (1'h1)); forvar6243 = (forvar6243 + (1'h1)))
                    begin
                      reg6244 <= $unsigned({forvar6078});
                      reg6245 <= ((^reg6105) >> ($signed($unsigned(reg6254)) + $signed($signed(forvar6179))));
                    end
                end
              if ($signed($signed(((reg6170 ?
                  reg6140 : reg6248) ^~ $unsigned(forvar6136)))))
                begin
                  for (forvar6257 = (1'h0); (forvar6257 < (2'h3)); forvar6257 = (forvar6257 + (1'h1)))
                    begin
                      reg6258 <= ((~&(~|(reg6091 ? reg6111 : reg6225))) ?
                          ((((8'hb5) != reg6024) << reg6176) * $unsigned(reg6168)) : (^~(reg6114 ?
                              forvar6111[(2'h3):(2'h2)] : (reg6142 ?
                                  reg6040 : reg6084))));
                      reg6259 <= reg6113[(1'h1):(1'h1)];
                    end
                end
              else
                begin
                  reg6257 <= $signed((~|($signed(reg6153) ~^ $unsigned(wire6218))));
                  if ($unsigned((forvar6212 >> reg6046[(3'h7):(3'h5)])))
                    begin
                      reg6258 <= wire6016[(3'h5):(2'h2)];
                    end
                  else
                    begin
                      reg6258 <= $unsigned((reg6252 <<< (reg6206 ?
                          $unsigned(reg6141) : (reg6199 >> forvar6149))));
                      reg6259 <= $signed((8'ha3));
                      reg6260 <= (reg6082 ?
                          (~$unsigned(forvar6097)) : ((^~$signed(reg6063)) ?
                              (~|forvar6018[(4'hf):(4'hb)]) : ((reg6068 ?
                                  reg6148 : reg6140) + (!reg6190))));
                    end
                  if (reg6147)
                    begin
                      reg6261 <= forvar6081[(1'h0):(1'h0)];
                      reg6262 <= {reg6132[(1'h0):(1'h0)]};
                      reg6263 <= reg6167;
                      reg6264 <= reg6062[(3'h7):(3'h4)];
                    end
                  else
                    begin
                      reg6261 <= $signed(reg6136[(2'h3):(2'h2)]);
                      reg6262 <= reg6131[(3'h4):(3'h4)];
                      reg6263 <= $signed((reg6099[(3'h6):(3'h4)] != (~&reg6063[(5'h10):(4'hc)])));
                    end
                  if (($signed($unsigned(reg6197[(4'h9):(4'h8)])) ~^ ((^$unsigned((8'hb9))) | reg6162[(2'h2):(2'h2)])))
                    begin
                      reg6265 <= $signed($unsigned($signed({reg6181})));
                      reg6266 <= reg6145[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg6265 <= (~(-$unsigned((reg6107 - reg6225))));
                      reg6266 <= ($unsigned(((~reg6135) ?
                              {(8'hb7)} : reg6058)) ?
                          forvar6178 : (&(8'ha8)));
                      reg6267 <= (reg6187[(3'h4):(1'h0)] < ($unsigned((reg6037 >= reg6140)) <<< $unsigned(((8'haa) ?
                          reg6142 : reg6243))));
                      reg6268 <= (-$unsigned(($unsigned(reg6109) ?
                          $unsigned((8'hab)) : (reg6184 > reg6254))));
                    end
                end
            end
          for (forvar6269 = (1'h0); (forvar6269 < (2'h3)); forvar6269 = (forvar6269 + (1'h1)))
            begin
              if ((wire5510[(1'h0):(1'h0)] << forvar6195))
                begin
                  for (forvar6270 = (1'h0); (forvar6270 < (1'h0)); forvar6270 = (forvar6270 + (1'h1)))
                    begin
                      reg6271 <= $signed(forvar6061[(4'hb):(3'h6)]);
                      reg6272 <= (|(((8'haa) | $unsigned(reg6080)) == reg6247[(3'h6):(2'h3)]));
                    end
                  if ($unsigned((~^(~^{reg6050}))))
                    begin
                      reg6273 <= reg6102;
                    end
                  else
                    begin
                      reg6273 <= {(forvar6050[(4'hb):(3'h6)] ?
                              $unsigned($signed(reg6126)) : reg6199[(1'h0):(1'h0)])};
                      reg6274 <= $signed(reg6141[(2'h2):(1'h1)]);
                      reg6275 <= forvar6159[(2'h3):(1'h0)];
                      reg6276 <= (8'h9d);
                    end
                  for (forvar6277 = (1'h0); (forvar6277 < (1'h1)); forvar6277 = (forvar6277 + (1'h1)))
                    begin
                      reg6278 <= (~^$signed($signed(reg6144)));
                      reg6279 <= {$unsigned((reg6200[(3'h4):(3'h4)] < {reg6163}))};
                      reg6280 <= $signed($signed({reg6213[(4'ha):(4'ha)]}));
                      reg6281 <= ({reg6248} ?
                          $signed((forvar6164 ^~ forvar6139[(4'h8):(4'h8)])) : (~^reg6273));
                    end
                end
              else
                begin
                  for (forvar6270 = (1'h0); (forvar6270 < (1'h0)); forvar6270 = (forvar6270 + (1'h1)))
                    begin
                      reg6271 <= reg6225[(3'h7):(3'h4)];
                    end
                end
              for (forvar6282 = (1'h0); (forvar6282 < (1'h1)); forvar6282 = (forvar6282 + (1'h1)))
                begin
                  for (forvar6283 = (1'h0); (forvar6283 < (2'h3)); forvar6283 = (forvar6283 + (1'h1)))
                    begin
                      reg6284 <= (reg6144[(1'h0):(1'h0)] > reg6062);
                      reg6285 <= (reg6154 ?
                          (&($unsigned(reg6261) & (reg6140 ?
                              reg6044 : reg6080))) : reg6203);
                    end
                  for (forvar6286 = (1'h0); (forvar6286 < (1'h0)); forvar6286 = (forvar6286 + (1'h1)))
                    begin
                      reg6287 <= reg6231[(4'h8):(2'h2)];
                    end
                end
              for (forvar6288 = (1'h0); (forvar6288 < (2'h3)); forvar6288 = (forvar6288 + (1'h1)))
                begin
                  if ($unsigned((((reg6034 ?
                      forvar6283 : reg6226) && (~&reg6241)) - (~|reg6050[(3'h6):(2'h2)]))))
                    begin
                      reg6289 <= (~^(reg6136 && reg6100));
                    end
                  else
                    begin
                      reg6289 <= (~&(!$unsigned(((8'ha6) ?
                          (8'had) : forvar6243))));
                      reg6290 <= $signed((~|reg6265[(2'h2):(2'h2)]));
                      reg6291 <= (+{{$unsigned((8'had))}});
                      reg6292 <= $unsigned($unsigned(reg6093[(3'h4):(1'h1)]));
                    end
                end
              for (forvar6293 = (1'h0); (forvar6293 < (2'h2)); forvar6293 = (forvar6293 + (1'h1)))
                begin
                  reg6294 <= reg6175[(2'h2):(1'h1)];
                end
            end
        end
      for (forvar6295 = (1'h0); (forvar6295 < (2'h2)); forvar6295 = (forvar6295 + (1'h1)))
        begin
          for (forvar6296 = (1'h0); (forvar6296 < (1'h1)); forvar6296 = (forvar6296 + (1'h1)))
            begin
              for (forvar6297 = (1'h0); (forvar6297 < (2'h3)); forvar6297 = (forvar6297 + (1'h1)))
                begin
                  for (forvar6298 = (1'h0); (forvar6298 < (1'h1)); forvar6298 = (forvar6298 + (1'h1)))
                    begin
                      reg6299 <= $signed((^~reg6187));
                      reg6300 <= (8'ha1);
                      reg6301 <= $unsigned(reg6191[(2'h2):(1'h0)]);
                    end
                end
            end
          for (forvar6302 = (1'h0); (forvar6302 < (2'h2)); forvar6302 = (forvar6302 + (1'h1)))
            begin
              for (forvar6303 = (1'h0); (forvar6303 < (2'h3)); forvar6303 = (forvar6303 + (1'h1)))
                begin
                  reg6304 <= (8'hb1);
                end
              reg6305 <= $unsigned(($unsigned((forvar6209 ~^ reg6163)) ?
                  $signed($unsigned(reg6205)) : reg6077));
              for (forvar6306 = (1'h0); (forvar6306 < (1'h0)); forvar6306 = (forvar6306 + (1'h1)))
                begin
                  for (forvar6307 = (1'h0); (forvar6307 < (2'h3)); forvar6307 = (forvar6307 + (1'h1)))
                    begin
                      reg6308 <= $signed((~$signed(((8'hb2) ?
                          (8'hb1) : forvar6060))));
                      reg6309 <= (((~(forvar6277 <= reg6111)) ?
                          ((8'hac) ?
                              reg6154 : (reg6115 ?
                                  (8'h9d) : forvar6165)) : ($unsigned((8'ha0)) ?
                              forvar6220 : (forvar6036 > forvar6283))) != $signed($signed({(8'ha7)})));
                      reg6310 <= reg6222[(4'h9):(3'h6)];
                      reg6311 <= ((reg6222[(4'ha):(3'h6)] * $unsigned((reg6216 >= reg6117))) && $signed((forvar6298[(1'h0):(1'h0)] ?
                          ((8'ha3) ? reg6074 : reg6145) : (reg6153 ?
                              forvar6097 : forvar6055))));
                    end
                end
              if ((8'hb5))
                begin
                  for (forvar6312 = (1'h0); (forvar6312 < (2'h3)); forvar6312 = (forvar6312 + (1'h1)))
                    begin
                      reg6313 <= (forvar6178 * ((reg6291[(4'ha):(4'h8)] < (reg6163 ?
                              forvar6178 : reg6085)) ?
                          ((reg6187 ? reg6043 : forvar6178) ?
                              (+reg6241) : reg6163) : $unsigned($unsigned(reg6053))));
                      reg6314 <= $signed($signed((!(forvar6221 ?
                          reg6272 : forvar6021))));
                      reg6315 <= (-reg6261);
                      reg6316 <= ($unsigned($unsigned((reg6118 ?
                          forvar6170 : forvar6122))) & ($signed((forvar6097 ?
                              reg6040 : forvar6137)) ?
                          (reg6284[(2'h3):(1'h1)] < (&(8'hb8))) : ($unsigned((8'hb6)) ?
                              (~^forvar6302) : $signed(reg6027))));
                    end
                  for (forvar6317 = (1'h0); (forvar6317 < (1'h0)); forvar6317 = (forvar6317 + (1'h1)))
                    begin
                      reg6318 <= {{(8'h9f)}};
                    end
                  for (forvar6319 = (1'h0); (forvar6319 < (2'h2)); forvar6319 = (forvar6319 + (1'h1)))
                    begin
                      reg6320 <= ({$signed((+(8'hb6)))} ?
                          $unsigned($unsigned((reg6098 ?
                              (8'hba) : forvar6228))) : reg6230[(4'ha):(2'h2)]);
                      reg6321 <= {(reg6116[(4'ha):(4'h9)] & reg6175)};
                    end
                  for (forvar6322 = (1'h0); (forvar6322 < (2'h2)); forvar6322 = (forvar6322 + (1'h1)))
                    begin
                      reg6323 <= $unsigned({($unsigned(reg6153) || reg6148)});
                    end
                end
              else
                begin
                  reg6312 <= (($signed(reg6237) ?
                          $signed({reg6144}) : (8'hba)) ?
                      reg6162[(4'ha):(2'h2)] : ((&reg6321[(3'h4):(1'h0)]) & forvar6293[(2'h3):(2'h3)]));
                  if (({reg6110[(3'h7):(3'h7)]} ?
                      (~forvar6166) : $signed((~^{forvar6293}))))
                    begin
                      reg6313 <= (reg6148[(3'h4):(2'h2)] ?
                          $unsigned((reg6247 << reg6315)) : reg6239[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg6313 <= ({$unsigned((forvar6044 > reg6195))} << (~|(!$signed(forvar6104))));
                      reg6314 <= $signed((reg6174[(2'h2):(1'h1)] ?
                          {(8'hb8)} : reg6084[(4'hb):(1'h1)]));
                      reg6315 <= forvar6135;
                    end
                  for (forvar6316 = (1'h0); (forvar6316 < (2'h3)); forvar6316 = (forvar6316 + (1'h1)))
                    begin
                      reg6317 <= $unsigned((((+reg6164) ^ {forvar6191}) ?
                          $signed((forvar6050 >= reg6138)) : reg6034[(4'h8):(3'h4)]));
                    end
                end
            end
          for (forvar6324 = (1'h0); (forvar6324 < (2'h2)); forvar6324 = (forvar6324 + (1'h1)))
            begin
              for (forvar6325 = (1'h0); (forvar6325 < (1'h0)); forvar6325 = (forvar6325 + (1'h1)))
                begin
                  reg6326 <= ((8'had) ?
                      (($signed(reg6261) ~^ $unsigned(reg6049)) && reg6242[(2'h3):(2'h2)]) : ($unsigned((reg6064 >> forvar6079)) ?
                          reg6259 : (~$unsigned(forvar6270))));
                  for (forvar6327 = (1'h0); (forvar6327 < (2'h2)); forvar6327 = (forvar6327 + (1'h1)))
                    begin
                      reg6328 <= reg6285[(1'h1):(1'h1)];
                      reg6329 <= (reg6237 ?
                          (8'hb6) : {$unsigned(forvar6208[(3'h7):(1'h0)])});
                      reg6330 <= (!((~|reg6129[(3'h7):(1'h1)]) ?
                          ($signed(reg6184) > forvar6116[(4'h8):(2'h3)]) : (8'ha4)));
                      reg6331 <= reg6062[(2'h3):(1'h1)];
                    end
                end
              for (forvar6332 = (1'h0); (forvar6332 < (2'h3)); forvar6332 = (forvar6332 + (1'h1)))
                begin
                  reg6333 <= $signed((reg6032[(1'h1):(1'h0)] ?
                      {reg6310[(4'hc):(3'h5)]} : ($unsigned(forvar6117) ?
                          (reg6090 <<< (8'hba)) : (^reg6215))));
                end
            end
        end
      reg6334 <= $signed($signed($signed($unsigned(reg6130))));
    end
  always
    @(posedge clk) begin
      for (forvar6335 = (1'h0); (forvar6335 < (2'h2)); forvar6335 = (forvar6335 + (1'h1)))
        begin
          for (forvar6336 = (1'h0); (forvar6336 < (1'h1)); forvar6336 = (forvar6336 + (1'h1)))
            begin
              if (forvar6234[(2'h3):(2'h2)])
                begin
                  if (wire6218)
                    begin
                      reg6337 <= forvar6253[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg6337 <= (-($signed(forvar6324) > {$signed(reg6150)}));
                      reg6338 <= $unsigned(($signed((~(8'ha0))) ?
                          $signed($signed(reg6323)) : ($signed(forvar6021) > (8'hb6))));
                    end
                  reg6339 <= $signed((^forvar6104[(1'h1):(1'h1)]));
                end
              else
                begin
                  if ((($unsigned($signed(reg6261)) * reg6167) - (forvar6117 <= reg6027[(4'h9):(4'h9)])))
                    begin
                      reg6337 <= reg6137;
                      reg6338 <= reg6213[(4'hb):(4'hb)];
                    end
                  else
                    begin
                      reg6337 <= (8'hb4);
                      reg6338 <= ($unsigned($unsigned((forvar6298 < forvar6159))) <= reg6110);
                    end
                  for (forvar6339 = (1'h0); (forvar6339 < (1'h1)); forvar6339 = (forvar6339 + (1'h1)))
                    begin
                      reg6340 <= reg6323[(4'ha):(1'h1)];
                      reg6341 <= {(((~|forvar6120) * reg6323) << (~|(~|reg6255)))};
                      reg6342 <= $signed($signed((~|$signed(reg6136))));
                    end
                  if ($signed(reg6168[(1'h0):(1'h0)]))
                    begin
                      reg6343 <= reg6317[(4'he):(1'h0)];
                      reg6344 <= forvar6135;
                      reg6345 <= (((reg6123 ?
                              reg6243[(3'h4):(2'h2)] : reg6255[(2'h3):(1'h1)]) >>> ((^reg6203) | $unsigned(reg6107))) ?
                          (8'haa) : forvar6171);
                      reg6346 <= {{$signed((forvar6277 ?
                                  (8'hb0) : forvar6195))}};
                    end
                  else
                    begin
                      reg6343 <= $unsigned((&(^((8'h9e) ?
                          forvar6322 : reg6057))));
                      reg6344 <= $unsigned((({reg6093} ?
                              (~&(8'hb9)) : reg6314) ?
                          ((reg6265 >>> reg6136) ?
                              $signed(reg6069) : $signed(reg6279)) : $unsigned({forvar6159})));
                      reg6345 <= {(((&(8'hb1)) | reg6106) >>> $unsigned(reg6203))};
                      reg6346 <= ((^~(^~reg6243[(2'h3):(1'h0)])) * ($unsigned((forvar6228 ?
                              reg6109 : forvar6129)) ?
                          $signed(reg6059[(3'h5):(2'h3)]) : (8'hac)));
                    end
                  for (forvar6347 = (1'h0); (forvar6347 < (1'h1)); forvar6347 = (forvar6347 + (1'h1)))
                    begin
                      reg6348 <= reg6341[(1'h1):(1'h1)];
                    end
                end
              if ($unsigned($signed($unsigned($unsigned(reg6158)))))
                begin
                  for (forvar6349 = (1'h0); (forvar6349 < (1'h0)); forvar6349 = (forvar6349 + (1'h1)))
                    begin
                      reg6350 <= $signed($unsigned(($unsigned(forvar6307) ?
                          reg6123[(4'hd):(3'h6)] : {(8'ha2)})));
                      reg6351 <= (8'ha4);
                    end
                  for (forvar6352 = (1'h0); (forvar6352 < (1'h1)); forvar6352 = (forvar6352 + (1'h1)))
                    begin
                      reg6353 <= forvar6302;
                      reg6354 <= {reg6250};
                      reg6355 <= reg6108[(2'h3):(1'h0)];
                      reg6356 <= reg6077[(1'h1):(1'h1)];
                    end
                  for (forvar6357 = (1'h0); (forvar6357 < (1'h1)); forvar6357 = (forvar6357 + (1'h1)))
                    begin
                      reg6358 <= $unsigned(((&(forvar6293 ^~ reg6229)) ?
                          ((reg6034 < reg6225) ?
                              $signed((8'ha9)) : {(8'ha5)}) : reg6121));
                      reg6359 <= ($unsigned((&(8'hae))) ?
                          $unsigned(reg6137[(4'hb):(1'h0)]) : $unsigned(forvar6195[(4'hd):(3'h4)]));
                    end
                  reg6360 <= (($signed((forvar6117 * (8'hb0))) ~^ (!forvar6081)) >= forvar6202[(3'h7):(3'h5)]);
                end
              else
                begin
                  for (forvar6349 = (1'h0); (forvar6349 < (2'h3)); forvar6349 = (forvar6349 + (1'h1)))
                    begin
                      reg6350 <= forvar6322;
                      reg6351 <= ({$unsigned((reg6190 ?
                              (8'ha1) : (8'hae)))} >>> (!$signed(reg6321[(3'h4):(3'h4)])));
                      reg6352 <= {reg6185};
                      reg6353 <= (8'hba);
                    end
                end
              if (((~|reg6271) ? reg6110 : (|reg6266)))
                begin
                  for (forvar6361 = (1'h0); (forvar6361 < (2'h3)); forvar6361 = (forvar6361 + (1'h1)))
                    begin
                      reg6362 <= $signed(((&(~&(8'h9c))) ?
                          {reg6037[(1'h0):(1'h0)]} : reg6334));
                      reg6363 <= (~^reg6200[(4'hd):(4'hb)]);
                      reg6364 <= reg6030;
                      reg6365 <= (|(8'h9e));
                    end
                  for (forvar6366 = (1'h0); (forvar6366 < (1'h1)); forvar6366 = (forvar6366 + (1'h1)))
                    begin
                      reg6367 <= (reg6120 ? reg6185 : reg6284);
                      reg6368 <= forvar6296;
                      reg6369 <= $signed((-((8'ha6) ?
                          (~|reg6180) : $signed(reg6147))));
                      reg6370 <= reg6137[(4'hc):(3'h7)];
                    end
                  for (forvar6371 = (1'h0); (forvar6371 < (2'h2)); forvar6371 = (forvar6371 + (1'h1)))
                    begin
                      reg6372 <= ($unsigned(((reg6315 ? reg6308 : reg6117) ?
                          $signed(reg6150) : {reg6247})) <<< (reg6049 ?
                          $unsigned($signed(reg6163)) : $signed($unsigned(reg6071))));
                    end
                end
              else
                begin
                  reg6361 <= (8'h9f);
                end
            end
        end
      for (forvar6373 = (1'h0); (forvar6373 < (2'h2)); forvar6373 = (forvar6373 + (1'h1)))
        begin
          if ($unsigned((!$signed((reg6206 << forvar6373)))))
            begin
              for (forvar6374 = (1'h0); (forvar6374 < (1'h1)); forvar6374 = (forvar6374 + (1'h1)))
                begin
                  if ($signed(($unsigned($unsigned(reg6372)) || reg6305[(3'h5):(2'h2)])))
                    begin
                      reg6375 <= (reg6316 ?
                          (-$signed(reg6203[(1'h0):(1'h0)])) : $signed(reg6131[(2'h3):(2'h3)]));
                      reg6376 <= $signed(reg6150[(2'h2):(1'h0)]);
                      reg6377 <= (($unsigned(reg6273[(2'h3):(1'h0)]) <= (reg6274[(1'h1):(1'h0)] | ((8'hb4) ?
                              reg6229 : (8'haa)))) ?
                          $signed(((reg6163 ? (8'ha6) : (8'ha8)) ?
                              {forvar6100} : (reg6051 ?
                                  forvar6044 : (8'haf)))) : {$unsigned($signed(forvar6212))});
                    end
                  else
                    begin
                      reg6375 <= forvar6104;
                      reg6376 <= $unsigned(reg6377);
                      reg6377 <= {reg6125};
                      reg6378 <= $unsigned($signed(reg6190));
                    end
                  for (forvar6379 = (1'h0); (forvar6379 < (2'h3)); forvar6379 = (forvar6379 + (1'h1)))
                    begin
                      reg6380 <= forvar6122[(1'h1):(1'h1)];
                    end
                  for (forvar6381 = (1'h0); (forvar6381 < (1'h0)); forvar6381 = (forvar6381 + (1'h1)))
                    begin
                      reg6382 <= $signed(forvar6036);
                      reg6383 <= $signed(((reg6343[(3'h4):(3'h4)] ?
                          (forvar6091 ?
                              forvar6149 : reg6358) : forvar6129[(1'h1):(1'h0)]) != $signed((reg6364 ~^ reg6320))));
                      reg6384 <= (reg6076 ?
                          (forvar6306[(3'h7):(3'h5)] ?
                              (~(|reg6320)) : (-(reg6128 > reg6154))) : (8'haa));
                      reg6385 <= (~^(|reg6376[(1'h0):(1'h0)]));
                    end
                end
              if (((~&$unsigned((reg6305 ?
                  forvar6282 : (8'ha0)))) << $signed(reg6024)))
                begin
                  reg6386 <= {reg6361};
                  for (forvar6387 = (1'h0); (forvar6387 < (2'h2)); forvar6387 = (forvar6387 + (1'h1)))
                    begin
                      reg6388 <= (~^reg6231[(2'h3):(1'h1)]);
                      reg6389 <= (($unsigned(reg6205) ^~ (8'hba)) ?
                          $unsigned((forvar6288 ?
                              reg6237 : $unsigned(reg6151))) : $signed($unsigned($signed(reg6300))));
                      reg6390 <= $unsigned(reg6038);
                      reg6391 <= forvar6050[(4'hb):(4'ha)];
                    end
                  for (forvar6392 = (1'h0); (forvar6392 < (2'h2)); forvar6392 = (forvar6392 + (1'h1)))
                    begin
                      reg6393 <= reg6370;
                      reg6394 <= forvar6312[(4'hb):(4'hb)];
                    end
                  reg6395 <= reg6128;
                end
              else
                begin
                  if ({reg6041})
                    begin
                      reg6386 <= (!(forvar6293 ?
                          {$signed(reg6090)} : {{forvar6145}}));
                      reg6387 <= forvar6243;
                      reg6388 <= (|{forvar6371});
                    end
                  else
                    begin
                      reg6386 <= $signed(($unsigned(forvar6129[(1'h0):(1'h0)]) ?
                          $signed((~&reg6104)) : forvar6099[(4'h9):(3'h4)]));
                    end
                  if ((~^(((reg6144 ? reg6098 : reg6356) ?
                      $signed(reg6391) : reg6044[(1'h0):(1'h0)]) || forvar6097)))
                    begin
                      reg6389 <= (reg6329 ?
                          (~&($signed(forvar6349) & (|reg6343))) : ((reg6314 != $unsigned(reg6360)) ?
                              (forvar6195 != $signed(reg6239)) : reg6330[(1'h0):(1'h0)]));
                      reg6390 <= $signed(reg6064);
                      reg6391 <= (((^~$signed((8'haa))) << ((forvar6179 ?
                                  (8'ha3) : reg6224) ?
                              forvar6020 : $signed(reg6100))) ?
                          ($signed((forvar6137 >= reg6111)) || ((^reg6051) ^~ (reg6040 - reg6323))) : $signed(((reg6331 >= forvar6232) ?
                              $signed(wire5509) : {reg6268})));
                      reg6392 <= $unsigned(reg6246);
                    end
                  else
                    begin
                      reg6389 <= (|(($unsigned(forvar6123) ?
                              {reg6080} : (forvar6336 ^ reg6233)) ?
                          $signed((reg6383 ?
                              reg6383 : reg6031)) : $unsigned(((8'ha6) - forvar6161))));
                    end
                  if ($signed(reg6271))
                    begin
                      reg6393 <= reg6091[(4'hf):(4'hc)];
                      reg6394 <= (~^(^~reg6162));
                      reg6395 <= $unsigned($signed((forvar6049 > $unsigned(reg6194))));
                      reg6396 <= ((+$unsigned((reg6265 | reg6041))) < forvar6339);
                    end
                  else
                    begin
                      reg6393 <= $unsigned(reg6028);
                      reg6394 <= (($signed((reg6384 ?
                              forvar6361 : (8'hb5))) >> ($unsigned(reg6313) ?
                              reg6194[(4'ha):(4'h9)] : $unsigned(reg6034))) ?
                          ((8'hac) >> (reg6114[(4'hc):(3'h7)] << (reg6276 < (8'hb6)))) : {($signed(reg6310) != (-(8'ha0)))});
                    end
                end
            end
          else
            begin
              for (forvar6374 = (1'h0); (forvar6374 < (1'h1)); forvar6374 = (forvar6374 + (1'h1)))
                begin
                  for (forvar6375 = (1'h0); (forvar6375 < (1'h1)); forvar6375 = (forvar6375 + (1'h1)))
                    begin
                      reg6376 <= (~|((!forvar6257) | forvar6322[(3'h4):(3'h4)]));
                    end
                  for (forvar6377 = (1'h0); (forvar6377 < (1'h1)); forvar6377 = (forvar6377 + (1'h1)))
                    begin
                      reg6378 <= forvar6366;
                      reg6379 <= forvar6221[(2'h3):(2'h3)];
                      reg6380 <= (&reg6350);
                      reg6381 <= (forvar6155 ~^ $signed(({forvar6253} ?
                          $unsigned((8'hae)) : (reg6230 ? reg6205 : reg6313))));
                    end
                  if (({$unsigned((+(8'h9f)))} ?
                      $signed($unsigned($signed(reg6173))) : forvar6149))
                    begin
                      reg6382 <= (reg6276[(1'h1):(1'h1)] ?
                          (forvar6306 ?
                              (8'ha8) : ((reg6059 ? (8'ha1) : (8'h9f)) ?
                                  ((8'hac) & forvar6179) : (8'hb4))) : forvar6339[(4'hb):(3'h7)]);
                    end
                  else
                    begin
                      reg6382 <= ($unsigned(($unsigned(reg6169) ?
                              $signed(reg6105) : $signed(wire5506))) ?
                          (~$unsigned($signed((8'hb0)))) : $unsigned($unsigned($unsigned(reg6226))));
                      reg6383 <= $unsigned($unsigned(((~^forvar6126) || (forvar6243 ?
                          forvar6116 : (8'ha6)))));
                    end
                end
              for (forvar6384 = (1'h0); (forvar6384 < (1'h0)); forvar6384 = (forvar6384 + (1'h1)))
                begin
                  if ((-$signed((^$unsigned(wire5507)))))
                    begin
                      reg6385 <= reg6291[(3'h6):(3'h4)];
                      reg6386 <= forvar6379[(1'h1):(1'h1)];
                      reg6387 <= ((((^~reg6392) & $unsigned(reg6086)) ?
                              reg6355 : $signed(reg6370[(3'h5):(2'h3)])) ?
                          $unsigned({reg6356[(1'h1):(1'h0)]}) : reg6287[(1'h1):(1'h0)]);
                    end
                  else
                    begin
                      reg6385 <= $unsigned($unsigned(forvar6208[(1'h0):(1'h0)]));
                    end
                  if ($unsigned((-forvar6303)))
                    begin
                      reg6388 <= $signed($unsigned($signed(reg6180)));
                    end
                  else
                    begin
                      reg6388 <= (|reg6098[(4'hb):(3'h5)]);
                      reg6389 <= $signed($unsigned($signed((^forvar6381))));
                      reg6390 <= ((reg6367[(1'h0):(1'h0)] | reg6321) ?
                          ((((8'hb3) >> forvar6384) * reg6385[(2'h3):(2'h2)]) <<< forvar6145[(3'h4):(3'h4)]) : forvar6055);
                      reg6391 <= $unsigned({$signed(reg6080[(4'hc):(4'h8)])});
                    end
                  reg6392 <= (forvar6212 ?
                      reg6160[(1'h1):(1'h1)] : $signed({$signed(forvar6178)}));
                end
              for (forvar6393 = (1'h0); (forvar6393 < (2'h2)); forvar6393 = (forvar6393 + (1'h1)))
                begin
                  for (forvar6394 = (1'h0); (forvar6394 < (1'h0)); forvar6394 = (forvar6394 + (1'h1)))
                    begin
                      reg6395 <= reg6309[(1'h1):(1'h1)];
                    end
                  if (((^(reg6165[(2'h2):(1'h1)] - (|forvar6149))) - $unsigned({$unsigned(reg6130)})))
                    begin
                      reg6396 <= reg6353;
                    end
                  else
                    begin
                      reg6396 <= (|$signed((+$signed(reg6352))));
                      reg6397 <= {($unsigned((reg6258 < forvar6139)) ?
                              ($signed(reg6290) ?
                                  ((8'ha3) & reg6077) : reg6204[(1'h0):(1'h0)]) : $unsigned((forvar6297 ?
                                  reg6273 : reg6064)))};
                    end
                  for (forvar6398 = (1'h0); (forvar6398 < (2'h2)); forvar6398 = (forvar6398 + (1'h1)))
                    begin
                      reg6399 <= ((~^reg6238[(2'h2):(1'h1)]) >> reg6362);
                      reg6400 <= ($signed({reg6195[(3'h5):(2'h3)]}) >= $signed(($signed(reg6299) - ((8'haf) ^~ reg6187))));
                      reg6401 <= $unsigned($signed((&(+forvar6179))));
                      reg6402 <= ($signed((reg6281 ?
                              reg6090 : $unsigned(reg6117))) ?
                          $unsigned($unsigned({reg6089})) : ($signed((~forvar6065)) && $signed((reg6292 ?
                              forvar6065 : (8'ha5)))));
                    end
                  reg6403 <= reg6256;
                end
            end
          reg6404 <= (~|reg6059[(4'h8):(1'h0)]);
          for (forvar6405 = (1'h0); (forvar6405 < (1'h0)); forvar6405 = (forvar6405 + (1'h1)))
            begin
              if ((reg6241 ? (+($signed(reg6301) * reg6138)) : forvar6220))
                begin
                  for (forvar6406 = (1'h0); (forvar6406 < (2'h3)); forvar6406 = (forvar6406 + (1'h1)))
                    begin
                      reg6407 <= (reg6188[(2'h2):(2'h2)] ?
                          ((~&(forvar6269 != reg6370)) ?
                              reg6352[(1'h1):(1'h1)] : $unsigned($signed(reg6023))) : reg6217);
                      reg6408 <= (8'hab);
                    end
                end
              else
                begin
                  reg6406 <= ($signed($unsigned($unsigned(forvar6319))) ?
                      (8'hb2) : reg6351[(4'hf):(4'he)]);
                  for (forvar6407 = (1'h0); (forvar6407 < (2'h3)); forvar6407 = (forvar6407 + (1'h1)))
                    begin
                      reg6408 <= $unsigned({{(8'haf)}});
                      reg6409 <= (~^forvar6398);
                      reg6410 <= $unsigned(($unsigned($unsigned(reg6195)) >= ((reg6022 ?
                              reg6052 : reg6350) ?
                          ((8'hb7) ? forvar6306 : forvar6398) : (forvar6019 ?
                              reg6257 : wire5508))));
                    end
                  for (forvar6411 = (1'h0); (forvar6411 < (2'h2)); forvar6411 = (forvar6411 + (1'h1)))
                    begin
                      reg6412 <= {{($signed(reg6103) ~^ (reg6135 * reg6215))}};
                      reg6413 <= forvar6018;
                      reg6414 <= $signed(({(forvar6019 ?
                              reg6128 : reg6280)} || (-(!reg6104))));
                    end
                  reg6415 <= (forvar6078 ?
                      ($unsigned($signed((8'hb2))) ?
                          reg6243[(3'h6):(1'h0)] : (^reg6067)) : $signed({$unsigned(reg6236)}));
                end
              reg6416 <= forvar6094;
              for (forvar6417 = (1'h0); (forvar6417 < (2'h3)); forvar6417 = (forvar6417 + (1'h1)))
                begin
                  if (reg6268[(4'hd):(2'h2)])
                    begin
                      reg6418 <= forvar6210;
                    end
                  else
                    begin
                      reg6418 <= $signed({$signed(reg6364)});
                      reg6419 <= forvar6335[(2'h2):(2'h2)];
                      reg6420 <= $unsigned($signed(((reg6409 ?
                              reg6215 : reg6176) ?
                          (reg6206 ? reg6261 : reg6243) : $unsigned(reg6199))));
                      reg6421 <= reg6163;
                    end
                  if (({($unsigned(reg6144) >>> (~forvar6136))} ?
                      reg6321[(1'h1):(1'h0)] : (reg6122[(1'h1):(1'h1)] < (~&$signed(reg6257)))))
                    begin
                      reg6422 <= ((^((forvar6406 <<< reg6193) ?
                          (^reg6168) : $unsigned(forvar6392))) < reg6275);
                      reg6423 <= (((|forvar6282[(3'h5):(3'h4)]) ?
                          reg6114[(4'h9):(2'h3)] : ((8'hab) ?
                              (~^reg6124) : reg6330[(4'h8):(1'h0)])) != (8'hae));
                      reg6424 <= {$unsigned($signed(reg6276[(3'h6):(1'h0)]))};
                      reg6425 <= ((!((-reg6139) ?
                          $signed(reg6287) : ((8'hb5) << reg6414))) == (!{(8'h9d)}));
                    end
                  else
                    begin
                      reg6422 <= reg6350[(1'h1):(1'h1)];
                    end
                  for (forvar6426 = (1'h0); (forvar6426 < (2'h2)); forvar6426 = (forvar6426 + (1'h1)))
                    begin
                      reg6427 <= ({(~^$unsigned((8'ha7)))} * ((~forvar6049[(2'h2):(1'h1)]) ?
                          reg6244 : reg6248));
                      reg6428 <= {reg6384[(3'h6):(3'h5)]};
                      reg6429 <= $unsigned((8'hb6));
                    end
                end
            end
          for (forvar6430 = (1'h0); (forvar6430 < (2'h3)); forvar6430 = (forvar6430 + (1'h1)))
            begin
              for (forvar6431 = (1'h0); (forvar6431 < (1'h0)); forvar6431 = (forvar6431 + (1'h1)))
                begin
                  for (forvar6432 = (1'h0); (forvar6432 < (2'h3)); forvar6432 = (forvar6432 + (1'h1)))
                    begin
                      reg6433 <= forvar6312;
                      reg6434 <= ($unsigned($signed((+reg6427))) ?
                          (!(reg6368 ~^ {(8'ha5)})) : $signed(reg6304));
                    end
                  for (forvar6435 = (1'h0); (forvar6435 < (2'h2)); forvar6435 = (forvar6435 + (1'h1)))
                    begin
                      reg6436 <= forvar6155;
                    end
                  if ((reg6172[(4'h9):(4'h9)] ^ (+(reg6164 ?
                      reg6175 : forvar6099))))
                    begin
                      reg6437 <= $unsigned(($signed((reg6199 ?
                          reg6090 : (8'h9c))) || reg6147[(1'h1):(1'h1)]));
                      reg6438 <= (~^({$unsigned(reg6114)} ?
                          (-(^~reg6024)) : $signed(reg6123)));
                      reg6439 <= reg6135[(4'h8):(3'h7)];
                      reg6440 <= reg6314;
                    end
                  else
                    begin
                      reg6437 <= (($unsigned($signed(forvar6050)) <<< (^$unsigned(reg6091))) ?
                          (+$signed(reg6350)) : forvar6195);
                    end
                end
            end
        end
      reg6441 <= (forvar6244 ~^ $signed((|$signed(reg6369))));
      reg6442 <= reg6170;
    end
  assign wire6443 = reg6284[(2'h2):(2'h2)];
  assign wire6444 = $signed(reg6416[(2'h2):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar6445 = (1'h0); (forvar6445 < (2'h2)); forvar6445 = (forvar6445 + (1'h1)))
        begin
          for (forvar6446 = (1'h0); (forvar6446 < (2'h3)); forvar6446 = (forvar6446 + (1'h1)))
            begin
              for (forvar6447 = (1'h0); (forvar6447 < (1'h0)); forvar6447 = (forvar6447 + (1'h1)))
                begin
                  if ($signed({(~|forvar6405)}))
                    begin
                      reg6448 <= forvar6081[(1'h1):(1'h1)];
                      reg6449 <= {(!reg6331)};
                      reg6450 <= reg6238;
                      reg6451 <= (reg6442 <<< $unsigned(($unsigned(forvar6381) & $unsigned(forvar6302))));
                    end
                  else
                    begin
                      reg6448 <= (!{(&{reg6309})});
                      reg6449 <= forvar6347[(2'h2):(1'h1)];
                      reg6450 <= reg6276[(2'h3):(2'h2)];
                    end
                end
              for (forvar6452 = (1'h0); (forvar6452 < (2'h2)); forvar6452 = (forvar6452 + (1'h1)))
                begin
                  for (forvar6453 = (1'h0); (forvar6453 < (1'h0)); forvar6453 = (forvar6453 + (1'h1)))
                    begin
                      reg6454 <= (+reg6204[(3'h5):(2'h2)]);
                      reg6455 <= ($unsigned(((reg6339 ? (8'haa) : (8'hb1)) ?
                          forvar6104 : (reg6314 ?
                              reg6436 : wire6218))) < $signed((forvar6297 == reg6086[(3'h5):(1'h1)])));
                      reg6456 <= $unsigned((^forvar6430[(1'h1):(1'h0)]));
                    end
                  if (reg6229[(4'ha):(2'h2)])
                    begin
                      reg6457 <= (|$unsigned({$signed(reg6126)}));
                    end
                  else
                    begin
                      reg6457 <= reg6265[(2'h2):(1'h1)];
                      reg6458 <= (-{(|reg6231)});
                      reg6459 <= {((8'hba) && reg6183)};
                      reg6460 <= forvar6139[(2'h3):(1'h0)];
                    end
                end
            end
          reg6461 <= (((forvar6319[(2'h2):(2'h2)] ~^ (reg6216 ?
              forvar6319 : forvar6347)) * $signed({reg6157})) > reg6111);
          reg6462 <= $signed((reg6121[(4'hb):(4'h8)] ?
              $signed((reg6292 << reg6429)) : (forvar6210 < (forvar6379 ?
                  reg6182 : reg6278))));
        end
      for (forvar6463 = (1'h0); (forvar6463 < (2'h3)); forvar6463 = (forvar6463 + (1'h1)))
        begin
          for (forvar6464 = (1'h0); (forvar6464 < (2'h2)); forvar6464 = (forvar6464 + (1'h1)))
            begin
              if ((reg6182[(2'h2):(2'h2)] != (reg6383[(3'h5):(2'h3)] >> $signed($signed(reg6049)))))
                begin
                  if (($signed(((&(8'h9f)) | $signed(reg6059))) >= $unsigned((~&reg6262[(1'h0):(1'h0)]))))
                    begin
                      reg6465 <= ((($unsigned(forvar6411) ?
                                  (reg6341 ?
                                      reg6164 : reg6449) : $signed(reg6163)) ?
                              $signed(forvar6232) : $signed((8'hb0))) ?
                          (8'hb5) : forvar6111[(3'h5):(1'h1)]);
                      reg6466 <= {(reg6191 ? (8'hb3) : (+reg6068))};
                    end
                  else
                    begin
                      reg6465 <= forvar6131;
                      reg6466 <= (8'hb3);
                      reg6467 <= $signed(($signed((^~(8'h9c))) || reg6034));
                      reg6468 <= ($unsigned((reg6185[(3'h6):(1'h1)] >> reg6051[(3'h7):(1'h1)])) ?
                          forvar6387[(1'h1):(1'h1)] : $signed((+reg6356)));
                    end
                  for (forvar6469 = (1'h0); (forvar6469 < (2'h3)); forvar6469 = (forvar6469 + (1'h1)))
                    begin
                      reg6470 <= (~reg6124);
                      reg6471 <= (reg6176[(3'h4):(1'h0)] != reg6259[(3'h6):(3'h4)]);
                      reg6472 <= {$signed(($unsigned((8'hb5)) ?
                              $signed((8'hac)) : ((8'ha2) <<< wire5506)))};
                      reg6473 <= forvar6435;
                    end
                  if (($unsigned((&(forvar6210 ~^ forvar6212))) ?
                      reg6410 : {(|(^~reg6229))}))
                    begin
                      reg6474 <= $unsigned((((reg6043 | forvar6131) ?
                          reg6409[(2'h2):(1'h1)] : $unsigned(forvar6161)) || $signed((~reg6291))));
                      reg6475 <= reg6346;
                    end
                  else
                    begin
                      reg6474 <= reg6451[(2'h2):(1'h1)];
                      reg6475 <= reg6365[(2'h3):(1'h0)];
                      reg6476 <= (((~&forvar6283) >= ((forvar6122 & reg6400) && $signed(reg6034))) - reg6233);
                    end
                  for (forvar6477 = (1'h0); (forvar6477 < (2'h2)); forvar6477 = (forvar6477 + (1'h1)))
                    begin
                      reg6478 <= reg6261[(1'h1):(1'h1)];
                      reg6479 <= $signed($signed((^$signed(reg6139))));
                      reg6480 <= forvar6435;
                      reg6481 <= $signed($unsigned($unsigned((!reg6415))));
                    end
                end
              else
                begin
                  for (forvar6465 = (1'h0); (forvar6465 < (1'h0)); forvar6465 = (forvar6465 + (1'h1)))
                    begin
                      reg6466 <= $unsigned((8'hba));
                      reg6467 <= forvar6060;
                      reg6468 <= reg6072;
                      reg6469 <= reg6381;
                    end
                  for (forvar6470 = (1'h0); (forvar6470 < (1'h1)); forvar6470 = (forvar6470 + (1'h1)))
                    begin
                      reg6471 <= (^~($unsigned($unsigned(reg6034)) ?
                          $unsigned({reg6157}) : {(wire5507 > reg6043)}));
                      reg6472 <= ($signed(forvar6286[(3'h6):(1'h0)]) >>> reg6383[(3'h7):(2'h2)]);
                      reg6473 <= reg6203;
                    end
                end
            end
          for (forvar6482 = (1'h0); (forvar6482 < (1'h0)); forvar6482 = (forvar6482 + (1'h1)))
            begin
              for (forvar6483 = (1'h0); (forvar6483 < (2'h2)); forvar6483 = (forvar6483 + (1'h1)))
                begin
                  for (forvar6484 = (1'h0); (forvar6484 < (2'h3)); forvar6484 = (forvar6484 + (1'h1)))
                    begin
                      reg6485 <= (~&(&((|reg6147) ?
                          (forvar6407 ? reg6321 : wire6443) : (!reg6140))));
                      reg6486 <= (^~reg6457);
                    end
                end
            end
          for (forvar6487 = (1'h0); (forvar6487 < (2'h2)); forvar6487 = (forvar6487 + (1'h1)))
            begin
              for (forvar6488 = (1'h0); (forvar6488 < (1'h1)); forvar6488 = (forvar6488 + (1'h1)))
                begin
                  reg6489 <= forvar6470[(3'h7):(3'h4)];
                end
              reg6490 <= reg6113;
              for (forvar6491 = (1'h0); (forvar6491 < (2'h2)); forvar6491 = (forvar6491 + (1'h1)))
                begin
                  for (forvar6492 = (1'h0); (forvar6492 < (1'h0)); forvar6492 = (forvar6492 + (1'h1)))
                    begin
                      reg6493 <= ((8'ha3) <<< {$signed((reg6121 ?
                              reg6378 : reg6408))});
                      reg6494 <= reg6051[(4'h9):(4'h9)];
                    end
                end
            end
        end
      reg6495 <= (($signed(forvar6349) ?
              (!(forvar6136 ? reg6494 : reg6252)) : (+(reg6333 ?
                  reg6350 : reg6416))) ?
          (~&($unsigned(reg6454) ?
              (reg6171 & reg6313) : reg6069)) : (+{reg6476}));
      for (forvar6496 = (1'h0); (forvar6496 < (1'h0)); forvar6496 = (forvar6496 + (1'h1)))
        begin
          reg6497 <= forvar6488;
          for (forvar6498 = (1'h0); (forvar6498 < (1'h1)); forvar6498 = (forvar6498 + (1'h1)))
            begin
              reg6499 <= $signed((~reg6419[(2'h3):(1'h1)]));
              if (((~&({reg6039} ?
                      (reg6257 ? reg6172 : reg6107) : $unsigned(forvar6091))) ?
                  reg6395 : {forvar6195[(4'hc):(3'h5)]}))
                begin
                  if (reg6148[(2'h3):(1'h1)])
                    begin
                      reg6500 <= $unsigned((((reg6151 ? reg6314 : reg6394) ?
                          (reg6173 < reg6131) : reg6124) != {{reg6471}}));
                      reg6501 <= (forvar6375[(4'hc):(2'h2)] ?
                          (^$signed(forvar6496[(2'h2):(2'h2)])) : {$unsigned($signed(forvar6316))});
                    end
                  else
                    begin
                      reg6500 <= (^reg6370[(4'ha):(3'h4)]);
                    end
                end
              else
                begin
                  reg6500 <= (reg6486 & forvar6297[(1'h1):(1'h0)]);
                end
              for (forvar6502 = (1'h0); (forvar6502 < (2'h2)); forvar6502 = (forvar6502 + (1'h1)))
                begin
                  if (reg6024[(1'h1):(1'h0)])
                    begin
                      reg6503 <= $unsigned($unsigned($unsigned($unsigned(forvar6122))));
                      reg6504 <= reg6350;
                      reg6505 <= reg6387[(1'h0):(1'h0)];
                      reg6506 <= (reg6438 ?
                          $unsigned(((8'hac) ?
                              reg6414 : forvar6127)) : (reg6130 ?
                              (reg6252 != {forvar6198}) : reg6312[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg6503 <= (forvar6303 ?
                          (reg6300[(3'h6):(1'h0)] ?
                              $signed($unsigned(reg6308)) : $signed({reg6140})) : $signed((8'h9e)));
                      reg6504 <= $unsigned((((forvar6349 ?
                          reg6385 : reg6352) >> (-reg6069)) < forvar6094));
                    end
                  for (forvar6507 = (1'h0); (forvar6507 < (2'h3)); forvar6507 = (forvar6507 + (1'h1)))
                    begin
                      reg6508 <= $unsigned(reg6462);
                      reg6509 <= (((reg6160[(3'h4):(2'h3)] | (reg6190 ?
                                  (8'ha0) : reg6438)) ?
                              ((8'ha1) ?
                                  forvar6352[(3'h6):(1'h1)] : (reg6388 * reg6441)) : ($signed((8'hb7)) ?
                                  reg6042[(1'h0):(1'h0)] : $unsigned(forvar6484))) ?
                          reg6037[(3'h6):(1'h1)] : $unsigned(reg6131));
                      reg6510 <= {$unsigned({reg6377[(3'h6):(2'h2)]})};
                      reg6511 <= (((~|(reg6080 - reg6200)) ?
                          reg6504 : ((8'hb0) ?
                              reg6125 : $unsigned(reg6196))) >= reg6326[(2'h3):(1'h0)]);
                    end
                end
              if (reg6489)
                begin
                  for (forvar6512 = (1'h0); (forvar6512 < (1'h1)); forvar6512 = (forvar6512 + (1'h1)))
                    begin
                      reg6513 <= ({$unsigned(reg6194)} * (-((~|reg6129) ?
                          reg6390 : $signed(reg6058))));
                    end
                  for (forvar6514 = (1'h0); (forvar6514 < (2'h3)); forvar6514 = (forvar6514 + (1'h1)))
                    begin
                      reg6515 <= ((reg6138[(5'h10):(4'ha)] ?
                          $unsigned($signed(reg6363)) : (8'ha9)) != reg6132[(1'h0):(1'h0)]);
                    end
                  if (((wire5507 <= reg6064) ?
                      ((8'ha3) ?
                          $signed((~reg6233)) : $unsigned(reg6260)) : (!($unsigned(reg6046) ?
                          ((8'ha7) ?
                              reg6051 : wire6443) : (forvar6134 - reg6147)))))
                    begin
                      reg6516 <= $signed((forvar6392[(3'h6):(3'h4)] * (~|forvar6219[(3'h6):(2'h3)])));
                    end
                  else
                    begin
                      reg6516 <= ((reg6247 ^ $signed((~^wire6016))) <= (~(~|forvar6198[(1'h1):(1'h1)])));
                    end
                  if ({$signed(forvar6019)})
                    begin
                      reg6517 <= $unsigned(reg6085);
                      reg6518 <= ((((reg6216 <= reg6503) ?
                              reg6244[(2'h3):(2'h3)] : (~|reg6333)) ?
                          (reg6285 <= ((8'hb1) & reg6312)) : (reg6064[(4'ha):(4'ha)] ?
                              reg6074[(3'h7):(3'h7)] : reg6291[(1'h1):(1'h1)])) ^~ {(~(forvar6295 ?
                              forvar6379 : reg6101))});
                    end
                  else
                    begin
                      reg6517 <= forvar6136;
                      reg6518 <= ((({reg6025} != (reg6321 ?
                          (8'hba) : reg6224)) || ($unsigned(reg6267) ^ (^reg6377))) - reg6114);
                    end
                end
              else
                begin
                  reg6512 <= ((8'ha0) - (!(~&forvar6482)));
                  for (forvar6513 = (1'h0); (forvar6513 < (2'h2)); forvar6513 = (forvar6513 + (1'h1)))
                    begin
                      reg6514 <= {reg6418};
                      reg6515 <= forvar6026;
                      reg6516 <= {(!(^~(reg6394 < reg6146)))};
                    end
                  for (forvar6517 = (1'h0); (forvar6517 < (2'h2)); forvar6517 = (forvar6517 + (1'h1)))
                    begin
                      reg6518 <= {((!$signed(reg6205)) ?
                              forvar6325 : (-wire5508))};
                    end
                end
            end
          for (forvar6519 = (1'h0); (forvar6519 < (2'h2)); forvar6519 = (forvar6519 + (1'h1)))
            begin
              if ((|$unsigned(forvar6426[(1'h0):(1'h0)])))
                begin
                  reg6520 <= ($unsigned({reg6396}) ?
                      $unsigned(((~^reg6513) + (~|reg6351))) : (!((^reg6504) ?
                          forvar6465[(4'h8):(2'h2)] : {reg6352})));
                  for (forvar6521 = (1'h0); (forvar6521 < (2'h2)); forvar6521 = (forvar6521 + (1'h1)))
                    begin
                      reg6522 <= (~&(8'ha8));
                      reg6523 <= ((^~forvar6178[(2'h2):(2'h2)]) ?
                          $unsigned(($unsigned(reg6050) ?
                              (wire5510 ?
                                  forvar6519 : (8'hb7)) : ((8'ha8) > reg6263))) : ($unsigned(((8'h9e) ~^ forvar6164)) ?
                              $signed((reg6272 ?
                                  forvar6286 : reg6516)) : reg6077));
                      reg6524 <= (8'hb5);
                    end
                  for (forvar6525 = (1'h0); (forvar6525 < (1'h1)); forvar6525 = (forvar6525 + (1'h1)))
                    begin
                      reg6526 <= {forvar6366[(2'h2):(1'h0)]};
                      reg6527 <= $signed(((|(reg6481 && reg6523)) - ($unsigned(forvar6379) ^~ $unsigned(reg6171))));
                    end
                end
              else
                begin
                  reg6520 <= ($unsigned(forvar6220) ?
                      ($unsigned(((8'hac) ?
                          wire6016 : forvar6145)) - (((8'ha3) * forvar6379) ?
                          (forvar6257 * forvar6293) : reg6369)) : $signed($unsigned($signed((8'h9e)))));
                  if (($signed((~|(^reg6311))) ?
                      (forvar6122[(1'h1):(1'h1)] ?
                          forvar6131 : $unsigned(((8'hb2) || reg6455))) : $unsigned({$signed(forvar6452)})))
                    begin
                      reg6521 <= $signed(reg6361);
                    end
                  else
                    begin
                      reg6521 <= (wire5507 < ((8'ha9) ?
                          reg6125[(4'h8):(1'h1)] : ($unsigned(forvar6100) ?
                              (reg6388 && forvar6406) : ((8'ha8) >= reg6222))));
                    end
                  for (forvar6522 = (1'h0); (forvar6522 < (1'h0)); forvar6522 = (forvar6522 + (1'h1)))
                    begin
                      reg6523 <= $signed((8'hae));
                    end
                  if ((reg6337 ? (reg6470 >>> reg6246) : (8'hb0)))
                    begin
                      reg6524 <= (({$unsigned(forvar6322)} ?
                              {(reg6450 == forvar6208)} : $signed(reg6113[(3'h4):(3'h4)])) ?
                          forvar6522[(3'h6):(3'h6)] : reg6378);
                      reg6525 <= ($unsigned(reg6189) ?
                          (^($unsigned(reg6138) ?
                              $signed(reg6153) : (^reg6205))) : (~(|{reg6181})));
                      reg6526 <= $unsigned(($signed((reg6279 ?
                              forvar6121 : reg6039)) ?
                          (~^$unsigned(reg6362)) : ((reg6093 ^~ reg6390) >= forvar6453[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg6524 <= {$signed({$unsigned(reg6068)})};
                      reg6525 <= $signed((8'hac));
                      reg6526 <= (~|$unsigned(($unsigned(reg6255) >= reg6047)));
                      reg6527 <= (+$unsigned({(&(8'hb3))}));
                    end
                end
              for (forvar6528 = (1'h0); (forvar6528 < (1'h0)); forvar6528 = (forvar6528 + (1'h1)))
                begin
                  for (forvar6529 = (1'h0); (forvar6529 < (2'h2)); forvar6529 = (forvar6529 + (1'h1)))
                    begin
                      reg6530 <= $signed((!forvar6394));
                      reg6531 <= $unsigned(reg6278[(1'h1):(1'h0)]);
                      reg6532 <= ((forvar6371[(3'h5):(3'h4)] >> (+(forvar6517 ?
                          reg6490 : (8'ha9)))) << reg6239);
                      reg6533 <= (~{{(forvar6384 ? forvar6381 : reg6217)}});
                    end
                  for (forvar6534 = (1'h0); (forvar6534 < (1'h0)); forvar6534 = (forvar6534 + (1'h1)))
                    begin
                      reg6535 <= $signed($unsigned($signed((forvar6482 <<< forvar6431))));
                      reg6536 <= forvar6079[(3'h4):(3'h4)];
                      reg6537 <= reg6106;
                      reg6538 <= $unsigned(($signed((-forvar6035)) > reg6080));
                    end
                  reg6539 <= $unsigned(reg6515[(2'h3):(1'h1)]);
                  for (forvar6540 = (1'h0); (forvar6540 < (2'h3)); forvar6540 = (forvar6540 + (1'h1)))
                    begin
                      reg6541 <= forvar6302;
                      reg6542 <= (reg6536 + (~(^~$unsigned(reg6192))));
                      reg6543 <= $unsigned(($unsigned(reg6418) & $unsigned((reg6200 ?
                          reg6201 : reg6504))));
                    end
                end
              reg6544 <= $signed($unsigned($unsigned(reg6469[(1'h0):(1'h0)])));
            end
        end
    end
  assign wire6545 = forvar6498;
  always
    @(posedge clk) begin
      if ((~&reg6383))
        begin
          if (reg6076)
            begin
              for (forvar6546 = (1'h0); (forvar6546 < (1'h1)); forvar6546 = (forvar6546 + (1'h1)))
                begin
                  reg6547 <= reg6247;
                  reg6548 <= (reg6285[(1'h0):(1'h0)] - reg6350[(1'h0):(1'h0)]);
                end
              for (forvar6549 = (1'h0); (forvar6549 < (2'h2)); forvar6549 = (forvar6549 + (1'h1)))
                begin
                  if (reg6370[(2'h3):(2'h2)])
                    begin
                      reg6550 <= reg6068[(4'he):(4'hb)];
                      reg6551 <= $signed($signed((^(reg6505 ?
                          reg6115 : forvar6431))));
                    end
                  else
                    begin
                      reg6550 <= reg6465[(2'h3):(2'h2)];
                    end
                  if ($signed($unsigned($signed((-forvar6165)))))
                    begin
                      reg6552 <= ($unsigned(((reg6317 > reg6505) ?
                              reg6365 : (~^(8'hb6)))) ?
                          ((reg6254 ^ reg6230[(1'h0):(1'h0)]) >= (-forvar6079)) : forvar6521);
                    end
                  else
                    begin
                      reg6552 <= $unsigned(reg6326[(1'h0):(1'h0)]);
                      reg6553 <= $signed((8'hb2));
                    end
                  for (forvar6554 = (1'h0); (forvar6554 < (1'h0)); forvar6554 = (forvar6554 + (1'h1)))
                    begin
                      reg6555 <= ({$signed($signed(reg6434))} ?
                          $unsigned(forvar6166[(1'h0):(1'h0)]) : reg6125[(3'h4):(3'h4)]);
                      reg6556 <= $signed(reg6206);
                    end
                end
              for (forvar6557 = (1'h0); (forvar6557 < (2'h3)); forvar6557 = (forvar6557 + (1'h1)))
                begin
                  reg6558 <= $unsigned($signed(reg6231));
                  for (forvar6559 = (1'h0); (forvar6559 < (1'h0)); forvar6559 = (forvar6559 + (1'h1)))
                    begin
                      reg6560 <= ($unsigned(((~(8'ha6)) && {forvar6288})) ?
                          (8'ha4) : (reg6244[(4'hf):(2'h2)] ~^ $unsigned(reg6214)));
                      reg6561 <= (forvar6507 ?
                          forvar6177 : reg6181[(1'h0):(1'h0)]);
                      reg6562 <= $signed($signed(forvar6129[(2'h2):(2'h2)]));
                      reg6563 <= (~^(~|(8'ha6)));
                    end
                  for (forvar6564 = (1'h0); (forvar6564 < (1'h1)); forvar6564 = (forvar6564 + (1'h1)))
                    begin
                      reg6565 <= (((((8'hae) * (8'haf)) && $unsigned(reg6424)) ?
                              (-(~|wire5508)) : (reg6121[(4'h8):(3'h7)] ?
                                  (forvar6507 & reg6152) : (~&reg6053))) ?
                          (^reg6532[(1'h0):(1'h0)]) : (((8'ha9) ?
                              (reg6057 <= reg6064) : reg6388) <<< {reg6408[(2'h3):(2'h3)]}));
                    end
                  if (($unsigned(((wire5509 > reg6389) * $unsigned(reg6166))) == ($signed((+forvar6357)) ?
                      {(reg6342 ? reg6495 : (8'hb9))} : ((reg6539 ?
                          forvar6171 : (8'ha6)) != $unsigned(wire6545)))))
                    begin
                      reg6566 <= (-(&reg6226));
                      reg6567 <= $signed($signed((^reg6098[(3'h5):(1'h0)])));
                      reg6568 <= (-(+((forvar6228 ? reg6504 : (8'ha5)) ?
                          $unsigned(reg6486) : forvar6371[(3'h4):(3'h4)])));
                      reg6569 <= reg6193;
                    end
                  else
                    begin
                      reg6566 <= ((~{forvar6392}) <<< forvar6528[(3'h7):(1'h1)]);
                      reg6567 <= (forvar6445 ?
                          reg6375 : ($unsigned($signed((8'ha9))) ?
                              (8'ha0) : (!(reg6313 & forvar6522))));
                      reg6568 <= $signed(reg6556[(2'h3):(1'h1)]);
                    end
                end
            end
          else
            begin
              if ((8'hb1))
                begin
                  for (forvar6546 = (1'h0); (forvar6546 < (1'h1)); forvar6546 = (forvar6546 + (1'h1)))
                    begin
                      reg6547 <= $signed(({(+reg6407)} ^ (reg6203 ^~ (reg6460 | reg6082))));
                    end
                  for (forvar6548 = (1'h0); (forvar6548 < (2'h2)); forvar6548 = (forvar6548 + (1'h1)))
                    begin
                      reg6549 <= (((8'hb8) && forvar6061) ?
                          {reg6384[(4'ha):(4'h8)]} : forvar6470[(2'h3):(1'h1)]);
                    end
                  reg6550 <= ((8'ha0) ?
                      ({reg6505[(2'h2):(1'h0)]} ?
                          $unsigned((reg6166 ^ reg6292)) : reg6309[(1'h1):(1'h0)]) : reg6230);
                  if (forvar6352)
                    begin
                      reg6551 <= ($signed($signed((reg6368 | (8'ha1)))) ?
                          (~&(forvar6325[(4'hd):(3'h4)] ?
                              $signed(forvar6018) : $signed(forvar6312))) : forvar6228[(2'h3):(1'h0)]);
                      reg6552 <= $signed($unsigned($unsigned((&reg6109))));
                    end
                  else
                    begin
                      reg6551 <= reg6025;
                      reg6552 <= reg6337;
                      reg6553 <= $signed($unsigned((+(forvar6060 ^~ reg6369))));
                      reg6554 <= ((~forvar6477[(4'h8):(1'h0)]) << {(~$unsigned(reg6318))});
                    end
                end
              else
                begin
                  for (forvar6546 = (1'h0); (forvar6546 < (2'h2)); forvar6546 = (forvar6546 + (1'h1)))
                    begin
                      reg6547 <= reg6504;
                    end
                  for (forvar6548 = (1'h0); (forvar6548 < (1'h0)); forvar6548 = (forvar6548 + (1'h1)))
                    begin
                      reg6549 <= (wire5508 ?
                          ($unsigned(reg6389) ?
                              ($unsigned(reg6486) ?
                                  $unsigned(forvar6525) : $signed(reg6512)) : $signed($signed(reg6171))) : $unsigned(reg6169[(3'h5):(3'h5)]));
                      reg6550 <= ((({(8'ha9)} < (~|reg6289)) ~^ (|reg6517[(3'h5):(1'h0)])) >>> $signed(($signed(reg6530) ?
                          $signed(reg6275) : (reg6456 >= reg6138))));
                      reg6551 <= ($unsigned($signed($signed((8'hba)))) ?
                          ((~^$signed(forvar6170)) + $signed(((8'ha2) ?
                              (8'ha9) : reg6390))) : reg6394);
                    end
                end
              for (forvar6555 = (1'h0); (forvar6555 < (2'h2)); forvar6555 = (forvar6555 + (1'h1)))
                begin
                  if ((forvar6253[(4'hb):(3'h4)] ?
                      ((~|$unsigned(reg6457)) ?
                          $unsigned({forvar6491}) : reg6140[(3'h4):(2'h2)]) : $signed(($signed(reg6050) + $signed(forvar6339)))))
                    begin
                      reg6556 <= {(({forvar6555} ?
                                  reg6089 : ((8'ha8) ? reg6345 : (8'ha6))) ?
                              $signed($signed(forvar6228)) : (reg6556[(3'h4):(2'h3)] == {forvar6519}))};
                      reg6557 <= reg6260[(3'h7):(3'h4)];
                      reg6558 <= ((forvar6104[(3'h7):(3'h7)] ?
                          $unsigned((reg6281 >>> reg6258)) : (8'h9e)) >> $unsigned($signed((forvar6407 ?
                          reg6476 : forvar6430))));
                      reg6559 <= reg6049[(2'h2):(1'h1)];
                    end
                  else
                    begin
                      reg6556 <= (+forvar6020);
                      reg6557 <= forvar6221;
                      reg6558 <= forvar6210[(4'hd):(4'hb)];
                    end
                  reg6560 <= $signed((-forvar6078[(4'h9):(4'h9)]));
                  if (($unsigned((-(reg6116 ? reg6257 : reg6191))) ?
                      $unsigned(((reg6196 ?
                          forvar6234 : reg6493) >= (^(8'ha4)))) : ($signed($unsigned(forvar6453)) >> ($unsigned(reg6118) ?
                          (reg6425 ?
                              forvar6244 : forvar6519) : (&forvar6220)))))
                    begin
                      reg6561 <= {((!(reg6150 ? reg6031 : forvar6446)) ?
                              ($unsigned(reg6080) + forvar6317) : ((reg6495 > forvar6055) << (^~reg6272)))};
                    end
                  else
                    begin
                      reg6561 <= ((reg6338 >>> {$signed(reg6271)}) ?
                          $signed((forvar6498 > (reg6072 ~^ reg6162))) : $unsigned(((reg6226 ?
                              forvar6035 : reg6108) << ((8'ha9) ?
                              reg6523 : reg6356))));
                    end
                end
              if (forvar6221)
                begin
                  for (forvar6562 = (1'h0); (forvar6562 < (2'h2)); forvar6562 = (forvar6562 + (1'h1)))
                    begin
                      reg6563 <= $unsigned(((&wire6218[(4'hb):(3'h4)]) ?
                          reg6114 : $unsigned(forvar6430[(3'h4):(2'h3)])));
                      reg6564 <= (reg6448 ?
                          (+((^~reg6427) >>> $unsigned(reg6022))) : ((forvar6094[(3'h6):(1'h0)] > {reg6341}) ^~ $signed($signed((8'ha4)))));
                    end
                  if (forvar6099)
                    begin
                      reg6565 <= ((~&((reg6516 ^~ reg6121) ?
                          $signed(forvar6411) : (^~forvar6210))) - forvar6470[(4'hd):(4'hd)]);
                      reg6566 <= $unsigned(forvar6065);
                      reg6567 <= $unsigned(reg6197);
                      reg6568 <= (($unsigned($unsigned((8'hb8))) >>> reg6263) ?
                          wire5509 : $unsigned($unsigned((reg6419 ?
                              forvar6257 : forvar6127))));
                    end
                  else
                    begin
                      reg6565 <= $unsigned((forvar6445 ?
                          (reg6132[(2'h2):(1'h0)] <= (reg6425 ?
                              reg6125 : reg6415)) : (reg6095[(3'h6):(1'h1)] << {forvar6375})));
                      reg6566 <= (~|forvar6121);
                      reg6567 <= ((~$unsigned(reg6117)) ?
                          ($signed({reg6123}) >>> forvar6137[(3'h5):(1'h1)]) : reg6102);
                      reg6568 <= ($signed(reg6224) ?
                          (-$unsigned((reg6360 ?
                              reg6433 : reg6173))) : (+$unsigned(((8'ha5) ?
                              reg6472 : reg6311))));
                    end
                  if ((reg6158 > (((8'hb1) + $signed((8'ha1))) ?
                      reg6504[(4'ha):(3'h7)] : $unsigned((reg6407 != forvar6502)))))
                    begin
                      reg6569 <= forvar6317[(2'h2):(2'h2)];
                      reg6570 <= (~&$unsigned((^(|reg6175))));
                    end
                  else
                    begin
                      reg6569 <= (((~^$unsigned(reg6340)) == $signed({wire5509})) ?
                          {(~&reg6254[(1'h0):(1'h0)])} : reg6174);
                      reg6570 <= (~&((8'hb4) >= ($signed(forvar6088) ?
                          reg6301 : (reg6205 > reg6389))));
                    end
                end
              else
                begin
                  if (($unsigned($unsigned((+reg6262))) ?
                      $signed({$signed(reg6533)}) : {$unsigned((8'hb7))}))
                    begin
                      reg6562 <= reg6116[(4'h9):(3'h7)];
                      reg6563 <= $unsigned($unsigned((|forvar6557[(2'h2):(1'h0)])));
                      reg6564 <= ((!{(reg6199 ? reg6037 : reg6116)}) ?
                          forvar6312 : $signed(((^~reg6249) ?
                              $signed(reg6356) : (reg6369 ^~ (8'ha4)))));
                    end
                  else
                    begin
                      reg6562 <= $signed((~|reg6092));
                    end
                  reg6565 <= $unsigned(reg6326);
                  if ($unsigned(reg6091))
                    begin
                      reg6566 <= forvar6407;
                    end
                  else
                    begin
                      reg6566 <= reg6458;
                    end
                  reg6567 <= {(((forvar6371 ?
                          reg6068 : reg6501) | reg6524[(4'hd):(3'h6)]) <<< ((reg6118 | wire5508) >= $signed(reg6025)))};
                end
              if ({{(forvar6347[(2'h2):(2'h2)] << (~|reg6133))}})
                begin
                  for (forvar6571 = (1'h0); (forvar6571 < (1'h0)); forvar6571 = (forvar6571 + (1'h1)))
                    begin
                      reg6572 <= ((^(reg6194[(1'h1):(1'h0)] & reg6466[(3'h6):(2'h3)])) ?
                          (!((|forvar6555) ^ reg6413)) : (reg6068 ?
                              ((reg6518 || reg6358) && (reg6316 * (8'hab))) : reg6256));
                    end
                end
              else
                begin
                  if ((~&(reg6192 ?
                      ($signed(reg6264) ?
                          (reg6047 <<< reg6409) : $unsigned(reg6305)) : ((~&reg6263) < (forvar6384 ?
                          reg6252 : forvar6149)))))
                    begin
                      reg6571 <= ($unsigned(forvar6178) == reg6567);
                      reg6572 <= ($signed(forvar6327[(1'h0):(1'h0)]) ?
                          {(^~{reg6308})} : $unsigned(forvar6134));
                    end
                  else
                    begin
                      reg6571 <= ((reg6309[(1'h1):(1'h1)] ^~ forvar6021[(3'h5):(3'h5)]) ?
                          reg6064[(3'h7):(1'h0)] : (~$signed({reg6339})));
                      reg6572 <= $signed((~reg6506[(3'h4):(1'h0)]));
                      reg6573 <= reg6337;
                    end
                end
            end
        end
      else
        begin
          reg6546 <= reg6470;
        end
      for (forvar6574 = (1'h0); (forvar6574 < (1'h1)); forvar6574 = (forvar6574 + (1'h1)))
        begin
          reg6575 <= $unsigned(((((8'hae) != reg6290) ?
              $unsigned(forvar6374) : reg6418) + reg6419));
          for (forvar6576 = (1'h0); (forvar6576 < (1'h0)); forvar6576 = (forvar6576 + (1'h1)))
            begin
              reg6577 <= (&$signed($signed((+reg6301))));
              reg6578 <= reg6557;
              for (forvar6579 = (1'h0); (forvar6579 < (1'h1)); forvar6579 = (forvar6579 + (1'h1)))
                begin
                  if ((({$signed(reg6339)} == $signed($unsigned(reg6392))) ?
                      ((|reg6310[(4'hb):(4'h8)]) ^ (!$signed(reg6047))) : ((8'hb8) ?
                          forvar6398[(1'h1):(1'h1)] : (~|(forvar6159 ?
                              reg6514 : (8'ha8))))))
                    begin
                      reg6580 <= $signed((&((~&reg6340) <<< $signed(reg6450))));
                    end
                  else
                    begin
                      reg6580 <= (+($unsigned((reg6144 ?
                              forvar6021 : reg6091)) ?
                          ($signed(forvar6548) ^~ $unsigned((8'hae))) : ($signed(reg6469) <= {reg6214})));
                      reg6581 <= reg6056[(2'h3):(1'h1)];
                      reg6582 <= (~^reg6415[(3'h6):(3'h6)]);
                    end
                  for (forvar6583 = (1'h0); (forvar6583 < (2'h3)); forvar6583 = (forvar6583 + (1'h1)))
                    begin
                      reg6584 <= $signed($signed(($unsigned(forvar6202) | {reg6207})));
                      reg6585 <= $signed((reg6582[(3'h5):(1'h1)] ?
                          (forvar6159[(4'h9):(1'h0)] && reg6392[(1'h1):(1'h1)]) : forvar6296[(2'h2):(1'h1)]));
                    end
                  for (forvar6586 = (1'h0); (forvar6586 < (1'h1)); forvar6586 = (forvar6586 + (1'h1)))
                    begin
                      reg6587 <= (($unsigned(reg6425) | reg6159[(4'hd):(3'h7)]) < ((8'ha4) >= (reg6490[(1'h0):(1'h0)] ?
                          forvar6484[(3'h5):(1'h1)] : (reg6305 ?
                              reg6341 : reg6172))));
                    end
                  for (forvar6588 = (1'h0); (forvar6588 < (2'h2)); forvar6588 = (forvar6588 + (1'h1)))
                    begin
                      reg6589 <= (~|($signed((^reg6023)) << reg6326[(2'h2):(1'h0)]));
                      reg6590 <= (((^~{forvar6253}) ^ {$unsigned((8'haf))}) ?
                          (+$signed(forvar6091[(3'h6):(1'h0)])) : ({reg6145[(3'h7):(1'h1)]} ?
                              $signed((reg6542 != forvar6528)) : reg6343));
                    end
                end
              for (forvar6591 = (1'h0); (forvar6591 < (2'h2)); forvar6591 = (forvar6591 + (1'h1)))
                begin
                  for (forvar6592 = (1'h0); (forvar6592 < (1'h1)); forvar6592 = (forvar6592 + (1'h1)))
                    begin
                      reg6593 <= ({((forvar6283 ?
                              reg6578 : forvar6209) || reg6578)} * reg6557);
                      reg6594 <= $signed(((-(|(8'hac))) - $signed(reg6107[(1'h0):(1'h0)])));
                    end
                end
            end
          if (reg6497[(4'hc):(4'h9)])
            begin
              if ((reg6098[(4'h9):(1'h1)] < (8'h9e)))
                begin
                  for (forvar6595 = (1'h0); (forvar6595 < (2'h2)); forvar6595 = (forvar6595 + (1'h1)))
                    begin
                      reg6596 <= (&$unsigned(reg6316[(3'h7):(3'h6)]));
                      reg6597 <= (^(8'hae));
                      reg6598 <= (+$signed($signed(reg6501)));
                      reg6599 <= $unsigned($unsigned(forvar6502));
                    end
                end
              else
                begin
                  for (forvar6595 = (1'h0); (forvar6595 < (2'h2)); forvar6595 = (forvar6595 + (1'h1)))
                    begin
                      reg6596 <= forvar6332;
                      reg6597 <= (reg6364 ? reg6091 : wire5509);
                    end
                  if (((((8'ha6) ^ $signed(reg6278)) + ($signed(forvar6135) > $signed((8'h9d)))) ^~ ((8'ha0) >> (~^(reg6133 ?
                      reg6490 : forvar6282)))))
                    begin
                      reg6598 <= ($signed((~$signed(forvar6491))) >= ((~&(8'ha9)) ?
                          $signed(reg6341[(4'hb):(4'h9)]) : (|reg6341[(3'h6):(3'h4)])));
                      reg6599 <= (~|$unsigned($unsigned(reg6386[(2'h2):(1'h0)])));
                      reg6600 <= (forvar6302[(1'h0):(1'h0)] - {reg6455});
                      reg6601 <= reg6313;
                    end
                  else
                    begin
                      reg6598 <= (forvar6517[(1'h1):(1'h1)] >= reg6568);
                      reg6599 <= reg6119[(1'h0):(1'h0)];
                      reg6600 <= (reg6557 ?
                          {$signed((!forvar6073))} : (((~^reg6527) <<< $unsigned((8'hb2))) || $unsigned($unsigned(forvar6373))));
                      reg6601 <= {(8'ha8)};
                    end
                  for (forvar6602 = (1'h0); (forvar6602 < (2'h2)); forvar6602 = (forvar6602 + (1'h1)))
                    begin
                      reg6603 <= (~reg6181);
                    end
                  reg6604 <= {(((reg6543 & reg6131) ?
                              $unsigned(reg6080) : (reg6549 ?
                                  (8'had) : reg6560)) ?
                          forvar6212[(3'h6):(3'h6)] : $signed($signed(forvar6554)))};
                end
            end
          else
            begin
              for (forvar6595 = (1'h0); (forvar6595 < (2'h3)); forvar6595 = (forvar6595 + (1'h1)))
                begin
                  if (((+{(reg6133 ? reg6249 : reg6196)}) ?
                      {forvar6394[(4'he):(4'h9)]} : $unsigned({$signed(forvar6498)})))
                    begin
                      reg6596 <= ($unsigned(forvar6417[(4'hd):(3'h7)]) ?
                          (8'ha5) : ((~^(forvar6335 >>> forvar6270)) ?
                              (~&(reg6440 ?
                                  forvar6528 : reg6130)) : (!((8'hb3) ?
                                  reg6252 : reg6235))));
                    end
                  else
                    begin
                      reg6596 <= (reg6486 + $unsigned(reg6051[(4'h9):(3'h7)]));
                    end
                  for (forvar6597 = (1'h0); (forvar6597 < (2'h3)); forvar6597 = (forvar6597 + (1'h1)))
                    begin
                      reg6598 <= reg6238[(4'h8):(1'h1)];
                      reg6599 <= {reg6521[(4'he):(4'hc)]};
                    end
                  reg6600 <= $unsigned($signed($signed(reg6451)));
                end
              for (forvar6601 = (1'h0); (forvar6601 < (2'h3)); forvar6601 = (forvar6601 + (1'h1)))
                begin
                  reg6602 <= (forvar6453 ?
                      $signed(((forvar6549 ? (8'hb6) : (8'hb7)) ?
                          (+forvar6020) : forvar6191[(2'h3):(1'h1)])) : (((reg6213 ?
                              reg6121 : reg6500) && (reg6594 & (8'hb8))) ?
                          $signed(((8'hab) <<< forvar6357)) : reg6527[(2'h2):(1'h0)]));
                  for (forvar6603 = (1'h0); (forvar6603 < (2'h2)); forvar6603 = (forvar6603 + (1'h1)))
                    begin
                      reg6604 <= (8'hab);
                      reg6605 <= (|forvar6035);
                    end
                end
              for (forvar6606 = (1'h0); (forvar6606 < (2'h2)); forvar6606 = (forvar6606 + (1'h1)))
                begin
                  reg6607 <= reg6173[(1'h0):(1'h0)];
                end
              if ({$unsigned((8'hb1))})
                begin
                  reg6608 <= ($signed($unsigned($signed((8'ha8)))) ?
                      $signed(($signed(reg6400) ?
                          (8'hb5) : reg6271[(3'h6):(2'h2)])) : (&((forvar6178 ?
                              reg6429 : reg6581) ?
                          reg6279 : $unsigned(forvar6482))));
                  if ($signed((~^$signed(reg6578[(2'h2):(1'h0)]))))
                    begin
                      reg6609 <= (^~forvar6576[(1'h0):(1'h0)]);
                      reg6610 <= reg6533[(4'hc):(4'hb)];
                      reg6611 <= ($signed(((reg6400 <= (8'ha6)) && (reg6056 ?
                              reg6116 : reg6299))) ?
                          ($unsigned((reg6062 ?
                              reg6243 : reg6501)) >>> ({reg6508} ?
                              reg6401 : reg6326[(1'h1):(1'h1)])) : {$signed(reg6424)});
                      reg6612 <= (^reg6224);
                    end
                  else
                    begin
                      reg6609 <= (reg6594[(4'hb):(2'h2)] >> reg6439);
                      reg6610 <= {(^~reg6381)};
                    end
                  if ($unsigned(reg6121))
                    begin
                      reg6613 <= (|($signed($unsigned((8'ha2))) ?
                          {(~reg6346)} : reg6152[(4'ha):(2'h3)]));
                      reg6614 <= reg6278[(3'h4):(2'h2)];
                      reg6615 <= reg6594;
                    end
                  else
                    begin
                      reg6613 <= (8'h9c);
                    end
                end
              else
                begin
                  if (reg6329)
                    begin
                      reg6608 <= forvar6111[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg6608 <= reg6597;
                    end
                  for (forvar6609 = (1'h0); (forvar6609 < (1'h1)); forvar6609 = (forvar6609 + (1'h1)))
                    begin
                      reg6610 <= forvar6099;
                    end
                  reg6611 <= ((!((forvar6170 ?
                          (8'h9d) : reg6589) <= (reg6533 - (8'ha6)))) ?
                      reg6145 : $unsigned(reg6142[(4'hb):(4'ha)]));
                  reg6612 <= reg6611[(4'h8):(3'h5)];
                end
            end
        end
    end
  assign wire6616 = {$signed(((-reg6197) ? reg6461 : (~forvar6564)))};
  assign wire6617 = reg6509;
  assign wire6618 = (reg6365 ?
                        reg6505[(4'hf):(2'h2)] : $signed((+$unsigned(forvar6549))));
  always
    @(posedge clk) begin
      for (forvar6619 = (1'h0); (forvar6619 < (2'h2)); forvar6619 = (forvar6619 + (1'h1)))
        begin
          if (forvar6135[(2'h2):(1'h1)])
            begin
              for (forvar6620 = (1'h0); (forvar6620 < (2'h2)); forvar6620 = (forvar6620 + (1'h1)))
                begin
                  reg6621 <= {(reg6355 <= ({reg6394} ?
                          $unsigned((8'hb7)) : reg6114))};
                  if ((~&$signed(forvar6298[(1'h0):(1'h0)])))
                    begin
                      reg6622 <= reg6289;
                      reg6623 <= reg6556;
                    end
                  else
                    begin
                      reg6622 <= reg6459;
                      reg6623 <= ((+$unsigned($signed(reg6422))) ?
                          (^~$signed(reg6140)) : ($unsigned((~reg6370)) ?
                              $signed($unsigned(forvar6373)) : reg6159[(4'hc):(4'hc)]));
                      reg6624 <= $unsigned({reg6193[(1'h0):(1'h0)]});
                      reg6625 <= forvar6528[(1'h1):(1'h0)];
                    end
                  if (forvar6521[(3'h5):(3'h4)])
                    begin
                      reg6626 <= (^$signed((!(reg6448 ? (8'h9f) : reg6240))));
                      reg6627 <= ((reg6051[(4'ha):(3'h4)] <<< ($signed(reg6391) ?
                          $unsigned(forvar6081) : forvar6583)) * $unsigned(reg6581[(3'h5):(2'h3)]));
                      reg6628 <= (((&(reg6130 << reg6122)) ?
                          {$unsigned(reg6164)} : forvar6303) > (-$signed((&reg6258))));
                    end
                  else
                    begin
                      reg6626 <= reg6074;
                    end
                end
              if (reg6066)
                begin
                  if (reg6382[(4'he):(4'h9)])
                    begin
                      reg6629 <= reg6331;
                      reg6630 <= (forvar6049[(1'h0):(1'h0)] != reg6145);
                    end
                  else
                    begin
                      reg6629 <= (reg6478 >> $unsigned(reg6195[(3'h4):(2'h2)]));
                    end
                end
              else
                begin
                  for (forvar6629 = (1'h0); (forvar6629 < (2'h2)); forvar6629 = (forvar6629 + (1'h1)))
                    begin
                      reg6630 <= reg6101[(1'h0):(1'h0)];
                      reg6631 <= $signed(reg6041);
                      reg6632 <= forvar6554[(2'h3):(2'h3)];
                      reg6633 <= forvar6295[(1'h0):(1'h0)];
                    end
                  if ((&($unsigned((~forvar6549)) || reg6109)))
                    begin
                      reg6634 <= {$signed(reg6138[(4'hf):(3'h4)])};
                      reg6635 <= reg6360[(4'hc):(4'hb)];
                    end
                  else
                    begin
                      reg6634 <= (forvar6060[(2'h3):(1'h0)] & ($signed((+forvar6270)) ?
                          ((reg6318 ?
                              reg6279 : reg6564) ~^ reg6138[(3'h6):(1'h0)]) : (-$signed(reg6601))));
                      reg6635 <= $unsigned(((^~(+reg6098)) ?
                          {$signed(forvar6178)} : forvar6525[(4'h8):(3'h5)]));
                      reg6636 <= (&reg6167);
                      reg6637 <= reg6559;
                    end
                end
              reg6638 <= ({((reg6513 || (8'hb4)) ?
                          (reg6533 ?
                              reg6486 : reg6257) : ((8'haa) << forvar6564))} ?
                  ((8'hae) ?
                      $unsigned({wire6616}) : $unsigned(forvar6104[(4'hc):(2'h2)])) : reg6216[(2'h2):(2'h2)]);
              if (reg6229)
                begin
                  if ($unsigned((-reg6290[(2'h2):(1'h1)])))
                    begin
                      reg6639 <= reg6465;
                      reg6640 <= $signed(forvar6099);
                    end
                  else
                    begin
                      reg6639 <= reg6033;
                    end
                  for (forvar6641 = (1'h0); (forvar6641 < (2'h3)); forvar6641 = (forvar6641 + (1'h1)))
                    begin
                      reg6642 <= $unsigned(({(&reg6236)} ?
                          {reg6161} : (~|$signed(reg6382))));
                      reg6643 <= (reg6428[(2'h3):(1'h0)] ?
                          ($signed(reg6416) ~^ reg6460) : (reg6513[(3'h4):(2'h3)] ?
                              reg6326 : (reg6419 == forvar6149[(1'h1):(1'h0)])));
                      reg6644 <= (~&{$signed((~&reg6578))});
                    end
                  for (forvar6645 = (1'h0); (forvar6645 < (1'h1)); forvar6645 = (forvar6645 + (1'h1)))
                    begin
                      reg6646 <= {$signed(reg6243[(2'h2):(1'h1)])};
                    end
                  if ((reg6305[(2'h3):(2'h2)] ?
                      reg6524[(2'h3):(2'h2)] : $signed(((~|reg6392) ?
                          $unsigned(reg6475) : (reg6367 ? reg6494 : reg6083)))))
                    begin
                      reg6647 <= $unsigned($unsigned(reg6230[(3'h5):(2'h2)]));
                      reg6648 <= ($signed((^~((8'hab) ?
                          forvar6574 : forvar6534))) >= {(&{reg6121})});
                    end
                  else
                    begin
                      reg6647 <= ($unsigned($unsigned(((8'h9d) ?
                          reg6161 : reg6370))) - $unsigned($signed((reg6165 != reg6213))));
                      reg6648 <= (reg6107[(2'h3):(1'h0)] & (8'hab));
                    end
                end
              else
                begin
                  if (reg6420)
                    begin
                      reg6639 <= $unsigned(reg6612[(4'hd):(3'h5)]);
                      reg6640 <= (~{reg6226[(2'h3):(2'h2)]});
                      reg6641 <= {$signed({(reg6206 ? reg6025 : forvar6571)})};
                      reg6642 <= $unsigned($unsigned((reg6172 ^ (reg6341 | forvar6469))));
                    end
                  else
                    begin
                      reg6639 <= (^~($unsigned((~&(8'hb4))) || $unsigned(reg6356)));
                      reg6640 <= reg6224[(1'h1):(1'h0)];
                    end
                  if (reg6314)
                    begin
                      reg6643 <= reg6173[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg6643 <= (&$unsigned($unsigned((&reg6267))));
                    end
                  for (forvar6644 = (1'h0); (forvar6644 < (2'h3)); forvar6644 = (forvar6644 + (1'h1)))
                    begin
                      reg6645 <= reg6203[(1'h1):(1'h1)];
                    end
                  for (forvar6646 = (1'h0); (forvar6646 < (2'h2)); forvar6646 = (forvar6646 + (1'h1)))
                    begin
                      reg6647 <= $signed(forvar6106[(3'h4):(2'h2)]);
                    end
                end
            end
          else
            begin
              for (forvar6620 = (1'h0); (forvar6620 < (2'h3)); forvar6620 = (forvar6620 + (1'h1)))
                begin
                  for (forvar6621 = (1'h0); (forvar6621 < (2'h3)); forvar6621 = (forvar6621 + (1'h1)))
                    begin
                      reg6622 <= reg6563[(2'h3):(2'h3)];
                    end
                end
              for (forvar6623 = (1'h0); (forvar6623 < (1'h0)); forvar6623 = (forvar6623 + (1'h1)))
                begin
                  for (forvar6624 = (1'h0); (forvar6624 < (1'h1)); forvar6624 = (forvar6624 + (1'h1)))
                    begin
                      reg6625 <= $unsigned(reg6372);
                      reg6626 <= {reg6267[(2'h3):(1'h1)]};
                    end
                  if (reg6527)
                    begin
                      reg6627 <= (((reg6550 ?
                              $unsigned(reg6042) : (|reg6569)) | (reg6181[(2'h2):(2'h2)] ~^ reg6475[(4'h8):(3'h4)])) ?
                          (($unsigned((8'ha6)) ?
                              {reg6047} : $signed(reg6154)) * (8'ha8)) : (reg6437[(3'h4):(1'h1)] ?
                              (reg6467 ?
                                  ((8'ha2) >> reg6566) : $unsigned((8'hb4))) : (|(forvar6319 > reg6420))));
                      reg6628 <= reg6171;
                      reg6629 <= $signed($unsigned((~&{forvar6097})));
                      reg6630 <= $unsigned(reg6468[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg6627 <= (forvar6131[(2'h3):(2'h2)] ?
                          (forvar6574[(4'ha):(3'h6)] << (+((8'hac) ?
                              reg6563 : reg6313))) : ((^~(reg6207 > (8'h9e))) ?
                              ((reg6266 + (8'hab)) ?
                                  (reg6058 || reg6215) : {reg6459}) : ((forvar6221 ?
                                  reg6025 : reg6603) == $unsigned(reg6450))));
                    end
                  if ((~&((|reg6040) ? reg6111[(3'h4):(3'h4)] : reg6543)))
                    begin
                      reg6631 <= $unsigned($signed(forvar6212[(3'h4):(1'h0)]));
                      reg6632 <= (^forvar6406);
                      reg6633 <= (8'ha6);
                      reg6634 <= (($signed((~&reg6334)) ?
                              $signed($signed(reg6462)) : $unsigned((reg6395 ?
                                  reg6062 : (8'h9c)))) ?
                          {forvar6394} : reg6044[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg6631 <= ($signed(reg6344[(1'h1):(1'h1)]) > $signed((~|(+reg6113))));
                      reg6632 <= reg6637;
                      reg6633 <= ($signed(((~reg6538) ?
                          (reg6413 ?
                              reg6261 : forvar6277) : reg6450[(4'h8):(1'h0)])) - $unsigned(((reg6330 >= reg6195) & (forvar6469 << forvar6606))));
                    end
                end
              reg6635 <= reg6526[(4'h9):(1'h1)];
              for (forvar6636 = (1'h0); (forvar6636 < (2'h2)); forvar6636 = (forvar6636 + (1'h1)))
                begin
                  for (forvar6637 = (1'h0); (forvar6637 < (1'h0)); forvar6637 = (forvar6637 + (1'h1)))
                    begin
                      reg6638 <= (|$signed($signed({(8'hb1)})));
                    end
                  for (forvar6639 = (1'h0); (forvar6639 < (1'h0)); forvar6639 = (forvar6639 + (1'h1)))
                    begin
                      reg6640 <= $signed($signed((8'hac)));
                      reg6641 <= (reg6634 ?
                          $signed((forvar6165 ?
                              $signed((8'ha5)) : reg6548)) : ($signed(((8'hb5) ?
                              wire6618 : (8'h9e))) <= reg6154[(3'h7):(3'h4)]));
                      reg6642 <= $signed({$unsigned((~reg6625))});
                    end
                  if (reg6128)
                    begin
                      reg6643 <= ((((forvar6387 + forvar6546) ?
                                  {reg6287} : $signed(forvar6120)) ?
                              reg6370[(1'h1):(1'h1)] : {$unsigned(forvar6469)}) ?
                          reg6450[(2'h3):(2'h2)] : ($signed({forvar6121}) == $signed((|(8'ha7)))));
                      reg6644 <= reg6557[(3'h7):(2'h2)];
                      reg6645 <= reg6473[(4'ha):(1'h0)];
                    end
                  else
                    begin
                      reg6643 <= $signed((-reg6558[(3'h5):(1'h0)]));
                      reg6644 <= (~&$signed($signed($signed(reg6320))));
                      reg6645 <= forvar6521[(3'h5):(3'h5)];
                      reg6646 <= $signed($unsigned($signed($unsigned(reg6321))));
                    end
                end
            end
          if ((-reg6419[(1'h1):(1'h1)]))
            begin
              reg6649 <= (&($signed(forvar6018) >> {{forvar6483}}));
            end
          else
            begin
              for (forvar6649 = (1'h0); (forvar6649 < (1'h0)); forvar6649 = (forvar6649 + (1'h1)))
                begin
                  reg6650 <= $unsigned((reg6245 ?
                      $unsigned((forvar6296 ? reg6265 : reg6582)) : reg6530));
                end
              if (forvar6549)
                begin
                  if ((^~(reg6548[(2'h2):(1'h0)] ?
                      {(~|reg6098)} : {(forvar6375 ? reg6245 : reg6290)})))
                    begin
                      reg6651 <= (|(reg6638[(2'h3):(2'h2)] >> (^~forvar6121)));
                      reg6652 <= $unsigned($unsigned((+{reg6419})));
                      reg6653 <= (reg6566 >= reg6098);
                      reg6654 <= reg6448[(2'h3):(1'h0)];
                    end
                  else
                    begin
                      reg6651 <= $unsigned(((^~$signed((8'hb2))) <= reg6358));
                      reg6652 <= reg6213[(4'hd):(2'h2)];
                      reg6653 <= reg6274;
                    end
                end
              else
                begin
                  if ((~&reg6217[(2'h3):(2'h2)]))
                    begin
                      reg6651 <= reg6033[(3'h5):(3'h4)];
                      reg6652 <= (({$signed(reg6623)} - $unsigned((forvar6592 ?
                          forvar6488 : reg6196))) >> {(~(forvar6629 ^ reg6063))});
                    end
                  else
                    begin
                      reg6651 <= (wire6218 ?
                          (+forvar6143[(1'h0):(1'h0)]) : (|reg6066[(4'hc):(2'h2)]));
                      reg6652 <= {reg6596};
                      reg6653 <= (|((((8'hb9) ? reg6148 : forvar6591) ?
                          {forvar6637} : reg6654[(1'h0):(1'h0)]) * (&forvar6317)));
                      reg6654 <= (((forvar6134[(1'h0):(1'h0)] <= $unsigned(reg6536)) >> $signed($unsigned(reg6070))) >>> (+((reg6511 + (8'haf)) | forvar6116)));
                    end
                  if (reg6047[(2'h2):(1'h1)])
                    begin
                      reg6655 <= $unsigned(reg6459);
                    end
                  else
                    begin
                      reg6655 <= reg6422;
                      reg6656 <= $unsigned((8'h9e));
                      reg6657 <= reg6351;
                    end
                  for (forvar6658 = (1'h0); (forvar6658 < (2'h2)); forvar6658 = (forvar6658 + (1'h1)))
                    begin
                      reg6659 <= $signed($unsigned((reg6581[(4'hd):(1'h1)] ?
                          (forvar6295 ?
                              reg6564 : reg6048) : $signed(reg6080))));
                      reg6660 <= ($signed((^~(~|reg6594))) ?
                          $unsigned((^~reg6538)) : ((reg6383[(3'h6):(2'h3)] ?
                              forvar6317[(2'h2):(2'h2)] : (reg6554 ?
                                  reg6422 : (8'hac))) * reg6068));
                    end
                end
              for (forvar6661 = (1'h0); (forvar6661 < (2'h3)); forvar6661 = (forvar6661 + (1'h1)))
                begin
                  if ({(~&forvar6282)})
                    begin
                      reg6662 <= (^~(8'h9c));
                      reg6663 <= ($unsigned(reg6624) >> $unsigned((reg6659 ?
                          {forvar6298} : (reg6192 ~^ reg6527))));
                      reg6664 <= (($unsigned((!reg6563)) ?
                          reg6395 : (&$unsigned(reg6631))) << (^forvar6637[(3'h5):(1'h1)]));
                    end
                  else
                    begin
                      reg6662 <= reg6317[(1'h0):(1'h0)];
                    end
                  if ($unsigned(($unsigned((forvar6097 | forvar6574)) ?
                      reg6195 : forvar6588[(1'h0):(1'h0)])))
                    begin
                      reg6665 <= reg6471[(4'h8):(3'h5)];
                      reg6666 <= ($unsigned(($signed(reg6415) ?
                              reg6649 : reg6602)) ?
                          reg6530 : {reg6382});
                      reg6667 <= $signed((+($unsigned(forvar6295) ?
                          (~|reg6364) : (reg6313 ? reg6333 : reg6072))));
                    end
                  else
                    begin
                      reg6665 <= (forvar6512[(2'h2):(2'h2)] + forvar6116[(3'h7):(3'h6)]);
                      reg6666 <= reg6291;
                      reg6667 <= reg6301[(1'h1):(1'h0)];
                      reg6668 <= reg6379;
                    end
                  for (forvar6669 = (1'h0); (forvar6669 < (1'h0)); forvar6669 = (forvar6669 + (1'h1)))
                    begin
                      reg6670 <= {reg6152[(4'h9):(4'h9)]};
                    end
                  if ($unsigned(reg6440))
                    begin
                      reg6671 <= $signed($unsigned(reg6425[(4'hf):(2'h3)]));
                      reg6672 <= ($signed(((reg6187 ? reg6183 : reg6388) ?
                              reg6467 : (^~forvar6588))) ?
                          (8'hb2) : $unsigned(({forvar6639} ?
                              reg6285 : {reg6600})));
                    end
                  else
                    begin
                      reg6671 <= ({$signed(reg6511[(3'h5):(2'h2)])} - forvar6078[(3'h4):(2'h3)]);
                      reg6672 <= (((|(forvar6435 == reg6114)) ?
                              reg6116[(4'ha):(3'h5)] : ((8'hac) ~^ ((8'h9d) >> forvar6477))) ?
                          reg6539 : reg6428);
                      reg6673 <= $signed((&$signed(reg6440[(3'h4):(2'h3)])));
                      reg6674 <= (~&reg6304);
                    end
                end
              for (forvar6675 = (1'h0); (forvar6675 < (1'h0)); forvar6675 = (forvar6675 + (1'h1)))
                begin
                  for (forvar6676 = (1'h0); (forvar6676 < (1'h0)); forvar6676 = (forvar6676 + (1'h1)))
                    begin
                      reg6677 <= $signed($unsigned(forvar6564));
                    end
                  reg6678 <= $signed(reg6066);
                  reg6679 <= forvar6186;
                end
            end
          for (forvar6680 = (1'h0); (forvar6680 < (2'h3)); forvar6680 = (forvar6680 + (1'h1)))
            begin
              for (forvar6681 = (1'h0); (forvar6681 < (2'h3)); forvar6681 = (forvar6681 + (1'h1)))
                begin
                  for (forvar6682 = (1'h0); (forvar6682 < (1'h0)); forvar6682 = (forvar6682 + (1'h1)))
                    begin
                      reg6683 <= (|forvar6116[(3'h7):(3'h6)]);
                      reg6684 <= forvar6574;
                    end
                  for (forvar6685 = (1'h0); (forvar6685 < (1'h1)); forvar6685 = (forvar6685 + (1'h1)))
                    begin
                      reg6686 <= ((reg6292[(2'h2):(1'h0)] | $unsigned(reg6100[(3'h5):(2'h2)])) ?
                          (8'hab) : $signed(({forvar6179} ?
                              forvar6327[(1'h1):(1'h0)] : $signed((8'hab)))));
                    end
                  for (forvar6687 = (1'h0); (forvar6687 < (2'h3)); forvar6687 = (forvar6687 + (1'h1)))
                    begin
                      reg6688 <= (forvar6026 ? (8'h9f) : wire6616);
                      reg6689 <= ((($signed(reg6160) != $signed(reg6074)) ?
                          ({reg6480} ?
                              reg6075[(4'ha):(4'ha)] : (reg6275 > reg6117)) : forvar6548) == (~(&(reg6185 ?
                          (8'ha6) : reg6259))));
                      reg6690 <= (^~(~&(&reg6609[(4'h8):(3'h6)])));
                    end
                end
              if ((({forvar6512} ?
                  (8'hb1) : ($unsigned(forvar6049) ?
                      $signed(reg6456) : (forvar6357 ?
                          reg6637 : reg6471))) >= reg6110))
                begin
                  for (forvar6691 = (1'h0); (forvar6691 < (2'h3)); forvar6691 = (forvar6691 + (1'h1)))
                    begin
                      reg6692 <= $unsigned((($signed(reg6543) - $signed((8'h9f))) >> (&(reg6124 * reg6098))));
                      reg6693 <= {((^~forvar6361[(4'h9):(2'h3)]) < $unsigned($unsigned(forvar6244)))};
                      reg6694 <= (((8'hb8) ?
                              reg6376 : (reg6104[(4'h9):(3'h7)] ?
                                  forvar6195[(3'h4):(2'h2)] : (reg6239 ~^ (8'ha0)))) ?
                          forvar6540 : ((-(reg6456 && reg6039)) != $unsigned($signed(forvar6685))));
                    end
                  if ($signed(reg6380))
                    begin
                      reg6695 <= $unsigned($unsigned({((8'ha4) ^ (8'ha5))}));
                      reg6696 <= $signed($signed($signed($signed(forvar6303))));
                      reg6697 <= $unsigned({forvar6394[(4'hb):(4'h8)]});
                      reg6698 <= (~^(!$unsigned(reg6279[(3'h6):(3'h4)])));
                    end
                  else
                    begin
                      reg6695 <= ({(forvar6680 <<< reg6427[(4'h9):(3'h4)])} ^ $unsigned((reg6359[(3'h4):(2'h3)] < {reg6137})));
                    end
                end
              else
                begin
                  for (forvar6691 = (1'h0); (forvar6691 < (1'h1)); forvar6691 = (forvar6691 + (1'h1)))
                    begin
                      reg6692 <= (&{reg6605[(3'h4):(2'h2)]});
                      reg6693 <= (($signed(forvar6269[(3'h6):(1'h0)]) ?
                              {(8'hae)} : (~&forvar6161[(2'h2):(2'h2)])) ?
                          $unsigned(($signed(reg6522) ?
                              reg6168 : (forvar6483 ?
                                  reg6376 : reg6136))) : $signed($unsigned($signed((8'ha3)))));
                    end
                  if (wire6444)
                    begin
                      reg6694 <= (reg6458[(1'h0):(1'h0)] ?
                          (^~((|forvar6347) ?
                              $unsigned(reg6634) : forvar6482)) : (((reg6100 >> reg6241) > (reg6128 ?
                                  reg6165 : forvar6105)) ?
                              ($unsigned((8'h9d)) ?
                                  (reg6684 ?
                                      reg6659 : (8'hb2)) : $signed(forvar6221)) : (~^{reg6455})));
                      reg6695 <= {forvar6597[(1'h1):(1'h0)]};
                      reg6696 <= (reg6651 - (($unsigned((8'hb0)) ?
                              (&reg6197) : ((8'hb6) ~^ forvar6168)) ?
                          (reg6197[(3'h7):(2'h3)] ?
                              (forvar6073 || reg6203) : (~^reg6093)) : reg6194));
                    end
                  else
                    begin
                      reg6694 <= (+($unsigned((reg6421 ?
                              forvar6134 : forvar6253)) ?
                          reg6276[(1'h0):(1'h0)] : (8'ha3)));
                      reg6695 <= reg6578[(2'h3):(1'h1)];
                      reg6696 <= reg6152;
                    end
                  for (forvar6697 = (1'h0); (forvar6697 < (2'h3)); forvar6697 = (forvar6697 + (1'h1)))
                    begin
                      reg6698 <= (((~|(forvar6055 >>> reg6638)) ?
                              ($unsigned(reg6241) ?
                                  $unsigned(reg6052) : {(8'ha5)}) : {(forvar6562 & (8'ha9))}) ?
                          {$unsigned((reg6323 > reg6321))} : $unsigned($unsigned((forvar6658 ?
                              reg6683 : reg6589))));
                      reg6699 <= {$signed({reg6185[(3'h7):(3'h5)]})};
                      reg6700 <= ($unsigned($signed(((8'ha8) ?
                              reg6337 : reg6551))) ?
                          $signed(((reg6401 ?
                              reg6028 : reg6613) * ((8'hb7) >>> reg6022))) : reg6247);
                    end
                end
              for (forvar6701 = (1'h0); (forvar6701 < (2'h2)); forvar6701 = (forvar6701 + (1'h1)))
                begin
                  if ($signed($signed(reg6439[(4'h9):(3'h6)])))
                    begin
                      reg6702 <= {(~$unsigned((reg6427 * forvar6529)))};
                      reg6703 <= forvar6477[(3'h5):(3'h5)];
                      reg6704 <= {$signed($unsigned($unsigned(reg6038)))};
                    end
                  else
                    begin
                      reg6702 <= ($signed((((8'hb5) + reg6043) ^ (reg6462 & forvar6549))) - $signed({(reg6197 >= (8'ha8))}));
                      reg6703 <= (8'h9c);
                    end
                  reg6705 <= $unsigned($unsigned(forvar6073[(4'h8):(1'h1)]));
                  for (forvar6706 = (1'h0); (forvar6706 < (1'h0)); forvar6706 = (forvar6706 + (1'h1)))
                    begin
                      reg6707 <= {(+reg6420[(3'h5):(2'h3)])};
                      reg6708 <= (reg6139[(4'hf):(3'h4)] ?
                          forvar6379[(2'h3):(2'h2)] : ((8'hb5) - {reg6355[(2'h3):(1'h0)]}));
                      reg6709 <= $unsigned(((~&$unsigned(reg6651)) | ((&(8'ha5)) ?
                          (forvar6357 ? reg6543 : reg6612) : (forvar6170 ?
                              reg6427 : reg6115))));
                      reg6710 <= reg6514[(1'h1):(1'h1)];
                    end
                  reg6711 <= {$signed(reg6140)};
                end
              for (forvar6712 = (1'h0); (forvar6712 < (1'h1)); forvar6712 = (forvar6712 + (1'h1)))
                begin
                  if (forvar6646)
                    begin
                      reg6713 <= ({{(reg6111 ?
                                  reg6360 : forvar6603)}} < reg6672);
                    end
                  else
                    begin
                      reg6713 <= forvar6469[(4'h9):(1'h0)];
                      reg6714 <= forvar6522[(2'h2):(2'h2)];
                      reg6715 <= reg6361;
                    end
                  for (forvar6716 = (1'h0); (forvar6716 < (2'h2)); forvar6716 = (forvar6716 + (1'h1)))
                    begin
                      reg6717 <= $unsigned(reg6355[(1'h1):(1'h1)]);
                      reg6718 <= (reg6276 >> $unsigned(((reg6615 <<< forvar6540) ?
                          (^reg6318) : $signed(forvar6195))));
                      reg6719 <= (^$signed((&(-reg6272))));
                      reg6720 <= {forvar6100[(2'h3):(1'h1)]};
                    end
                  reg6721 <= (($unsigned((reg6064 >>> reg6628)) ?
                          $signed((reg6437 ?
                              reg6461 : reg6503)) : (&$unsigned(reg6501))) ?
                      (^(reg6493[(2'h3):(1'h1)] ?
                          {reg6170} : {reg6188})) : $unsigned(reg6427[(2'h2):(2'h2)]));
                end
            end
          for (forvar6722 = (1'h0); (forvar6722 < (2'h2)); forvar6722 = (forvar6722 + (1'h1)))
            begin
              if ((reg6609[(3'h4):(3'h4)] ?
                  reg6532[(1'h0):(1'h0)] : (forvar6018 <= ({reg6457} && $unsigned(reg6050)))))
                begin
                  for (forvar6723 = (1'h0); (forvar6723 < (1'h0)); forvar6723 = (forvar6723 + (1'h1)))
                    begin
                      reg6724 <= ((8'h9f) ?
                          (~|forvar6060[(2'h3):(1'h0)]) : (8'ha5));
                    end
                  if ((~^({(forvar6644 || (8'hb8))} >= reg6596[(3'h6):(2'h2)])))
                    begin
                      reg6725 <= $unsigned(reg6105);
                    end
                  else
                    begin
                      reg6725 <= (+({(^~(8'hb2))} ?
                          ($unsigned(reg6455) ?
                              $signed(reg6703) : reg6438) : (-reg6664[(4'h8):(2'h2)])));
                      reg6726 <= reg6140[(2'h2):(1'h0)];
                    end
                  if ($signed($signed(({reg6714} >> $signed(forvar6601)))))
                    begin
                      reg6727 <= reg6114;
                      reg6728 <= reg6284;
                      reg6729 <= (!reg6527[(3'h4):(2'h3)]);
                      reg6730 <= reg6043[(4'h8):(4'h8)];
                    end
                  else
                    begin
                      reg6727 <= (($signed(reg6572[(3'h6):(2'h3)]) >= ((|forvar6198) ?
                              $signed((8'ha3)) : (^~reg6478))) ?
                          (+reg6027[(3'h5):(1'h0)]) : $unsigned(($signed(reg6520) ?
                              reg6111[(1'h1):(1'h1)] : $signed(forvar6116))));
                    end
                end
              else
                begin
                  for (forvar6723 = (1'h0); (forvar6723 < (1'h1)); forvar6723 = (forvar6723 + (1'h1)))
                    begin
                      reg6724 <= ((reg6355 > reg6623) == (-{(reg6096 ~^ (8'hb7))}));
                      reg6725 <= (~($signed((reg6603 ?
                          forvar6177 : (8'ha4))) > ((8'ha1) ?
                          (reg6237 | (8'hb1)) : (~reg6679))));
                    end
                  for (forvar6726 = (1'h0); (forvar6726 < (2'h3)); forvar6726 = (forvar6726 + (1'h1)))
                    begin
                      reg6727 <= (|forvar6446);
                      reg6728 <= $unsigned($signed((~(forvar6549 < reg6348))));
                      reg6729 <= reg6486[(3'h5):(3'h5)];
                    end
                end
            end
        end
      if (forvar6514)
        begin
          for (forvar6731 = (1'h0); (forvar6731 < (1'h0)); forvar6731 = (forvar6731 + (1'h1)))
            begin
              reg6732 <= {(-reg6252)};
              reg6733 <= {$unsigned((|{reg6315}))};
              if ($signed(reg6438))
                begin
                  for (forvar6734 = (1'h0); (forvar6734 < (1'h1)); forvar6734 = (forvar6734 + (1'h1)))
                    begin
                      reg6735 <= ({forvar6149} || (~&(^~(^(8'ha6)))));
                      reg6736 <= $unsigned(($unsigned($unsigned(forvar6131)) ?
                          $signed($unsigned((8'ha9))) : (reg6555 ?
                              ((8'haf) || wire6545) : (reg6497 & reg6547))));
                      reg6737 <= ($unsigned(reg6328[(1'h1):(1'h0)]) & reg6451[(2'h2):(1'h0)]);
                      reg6738 <= reg6708[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar6734 = (1'h0); (forvar6734 < (1'h0)); forvar6734 = (forvar6734 + (1'h1)))
                    begin
                      reg6735 <= reg6259[(2'h3):(2'h3)];
                      reg6736 <= ({($signed(reg6418) - ((8'hb2) <= reg6047))} << ($signed(((8'ha4) & wire6218)) ?
                          reg6707[(4'h8):(4'h8)] : (^(+forvar6595))));
                    end
                end
            end
          for (forvar6739 = (1'h0); (forvar6739 < (1'h0)); forvar6739 = (forvar6739 + (1'h1)))
            begin
              for (forvar6740 = (1'h0); (forvar6740 < (1'h0)); forvar6740 = (forvar6740 + (1'h1)))
                begin
                  if ($unsigned((reg6351[(1'h0):(1'h0)] ^~ reg6028[(3'h6):(3'h5)])))
                    begin
                      reg6741 <= $signed(reg6285[(4'h9):(1'h1)]);
                      reg6742 <= ($unsigned(forvar6682[(4'ha):(3'h6)]) ?
                          reg6104 : reg6257);
                      reg6743 <= reg6113[(2'h2):(2'h2)];
                      reg6744 <= $signed($signed((reg6063 ~^ (+reg6275))));
                    end
                  else
                    begin
                      reg6741 <= $signed($signed(forvar6555));
                      reg6742 <= (8'h9e);
                      reg6743 <= (|$unsigned((^~(~&(8'hb5)))));
                      reg6744 <= ($unsigned(($unsigned(reg6472) ?
                          forvar6283 : ((8'ha4) <<< forvar6548))) ^ ((!reg6238) ?
                          $unsigned({wire6616}) : forvar6592[(1'h1):(1'h1)]));
                    end
                end
              if (({((~|(8'ha1)) ? reg6575 : $signed(reg6329))} ?
                  forvar6579[(2'h3):(2'h3)] : ((reg6246 || {reg6513}) ?
                      $signed(reg6508) : reg6589[(1'h0):(1'h0)])))
                begin
                  reg6745 <= $signed(($unsigned(reg6710) ?
                      {reg6174} : (forvar6177[(3'h7):(3'h4)] <<< reg6503[(4'hc):(4'ha)])));
                  for (forvar6746 = (1'h0); (forvar6746 < (2'h3)); forvar6746 = (forvar6746 + (1'h1)))
                    begin
                      reg6747 <= ({$unsigned({forvar6044})} ?
                          (|$unsigned(reg6076[(3'h7):(3'h5)])) : reg6196);
                      reg6748 <= $signed(((((8'hb5) ?
                              forvar6297 : forvar6706) || (reg6635 ^ reg6181)) ?
                          $unsigned($signed(forvar6491)) : reg6182));
                      reg6749 <= $signed((8'ha2));
                    end
                  for (forvar6750 = (1'h0); (forvar6750 < (2'h3)); forvar6750 = (forvar6750 + (1'h1)))
                    begin
                      reg6751 <= ($signed((8'hac)) ~^ $signed($unsigned((reg6449 ?
                          (8'hba) : forvar6209))));
                      reg6752 <= (reg6032[(4'hb):(2'h3)] ?
                          forvar6393[(3'h4):(2'h3)] : (+forvar6145));
                      reg6753 <= reg6694[(4'hf):(4'hd)];
                    end
                end
              else
                begin
                  for (forvar6745 = (1'h0); (forvar6745 < (1'h0)); forvar6745 = (forvar6745 + (1'h1)))
                    begin
                      reg6746 <= $unsigned(((|forvar6221) << reg6441[(4'he):(4'hd)]));
                    end
                  if (reg6368[(1'h0):(1'h0)])
                    begin
                      reg6747 <= forvar6557;
                      reg6748 <= $signed(((~^$unsigned(reg6695)) ?
                          $unsigned((~^reg6103)) : (((8'hb5) ?
                              forvar6295 : reg6251) <= $signed(reg6729))));
                      reg6749 <= reg6530[(1'h1):(1'h0)];
                      reg6750 <= {($unsigned((reg6138 >>> (8'h9f))) <<< ((^forvar6691) ?
                              reg6535 : {(8'had)}))};
                    end
                  else
                    begin
                      reg6747 <= $signed({reg6604});
                      reg6748 <= reg6526[(2'h2):(2'h2)];
                    end
                end
            end
          reg6754 <= reg6454;
          if (reg6104)
            begin
              if (forvar6166[(1'h1):(1'h1)])
                begin
                  if ($unsigned($signed((~&(reg6028 ? reg6039 : forvar6706)))))
                    begin
                      reg6755 <= {forvar6312};
                      reg6756 <= (^($unsigned(forvar6325[(4'h9):(2'h3)]) <= reg6243));
                    end
                  else
                    begin
                      reg6755 <= (8'ha8);
                      reg6756 <= (|(reg6428[(2'h3):(1'h1)] ~^ (8'hac)));
                      reg6757 <= ($unsigned($unsigned($signed(reg6109))) == forvar6131);
                      reg6758 <= (-(|$unsigned((reg6509 << reg6535))));
                    end
                end
              else
                begin
                  for (forvar6755 = (1'h0); (forvar6755 < (1'h1)); forvar6755 = (forvar6755 + (1'h1)))
                    begin
                      reg6756 <= reg6624;
                      reg6757 <= $signed((forvar6591[(3'h6):(3'h5)] ?
                          forvar6430[(2'h3):(2'h2)] : ({(8'h9d)} ?
                              reg6527[(2'h2):(1'h0)] : forvar6097[(3'h5):(3'h4)])));
                    end
                end
            end
          else
            begin
              for (forvar6755 = (1'h0); (forvar6755 < (1'h0)); forvar6755 = (forvar6755 + (1'h1)))
                begin
                  for (forvar6756 = (1'h0); (forvar6756 < (2'h2)); forvar6756 = (forvar6756 + (1'h1)))
                    begin
                      reg6757 <= reg6064;
                      reg6758 <= $unsigned($unsigned((~|$unsigned(reg6428))));
                      reg6759 <= reg6522;
                      reg6760 <= (^~($unsigned(forvar6045[(2'h2):(2'h2)]) || reg6074));
                    end
                  reg6761 <= reg6084[(5'h10):(3'h7)];
                  for (forvar6762 = (1'h0); (forvar6762 < (1'h0)); forvar6762 = (forvar6762 + (1'h1)))
                    begin
                      reg6763 <= reg6605;
                    end
                end
              for (forvar6764 = (1'h0); (forvar6764 < (2'h2)); forvar6764 = (forvar6764 + (1'h1)))
                begin
                  if ((8'hb9))
                    begin
                      reg6765 <= {({{reg6571}} ?
                              $signed($signed((8'hac))) : {((8'ha1) >>> (8'hb9))})};
                    end
                  else
                    begin
                      reg6765 <= (~&(reg6027 ~^ $unsigned($unsigned((8'ha6)))));
                      reg6766 <= forvar6398;
                      reg6767 <= reg6101;
                      reg6768 <= ((($signed(reg6454) >> forvar6139[(4'h8):(2'h3)]) ^ (reg6656[(4'hc):(4'hb)] ?
                              reg6499[(4'h9):(1'h1)] : {forvar6018})) ?
                          reg6345 : ((reg6226[(2'h3):(2'h3)] ?
                                  $unsigned(forvar6609) : reg6467) ?
                              $signed($signed(reg6695)) : reg6535));
                    end
                  for (forvar6769 = (1'h0); (forvar6769 < (1'h0)); forvar6769 = (forvar6769 + (1'h1)))
                    begin
                      reg6770 <= forvar6131;
                      reg6771 <= $signed($unsigned((reg6093 >= reg6100[(3'h4):(3'h4)])));
                    end
                end
            end
        end
      else
        begin
          for (forvar6731 = (1'h0); (forvar6731 < (2'h2)); forvar6731 = (forvar6731 + (1'h1)))
            begin
              for (forvar6732 = (1'h0); (forvar6732 < (2'h3)); forvar6732 = (forvar6732 + (1'h1)))
                begin
                  for (forvar6733 = (1'h0); (forvar6733 < (2'h3)); forvar6733 = (forvar6733 + (1'h1)))
                    begin
                      reg6734 <= $unsigned(forvar6079[(3'h4):(2'h2)]);
                      reg6735 <= reg6390[(2'h2):(1'h0)];
                      reg6736 <= $signed(({$signed(forvar6097)} ~^ reg6289));
                      reg6737 <= {$unsigned((forvar6557 & (forvar6756 && forvar6055)))};
                    end
                  reg6738 <= reg6138[(4'h9):(1'h1)];
                  reg6739 <= (8'hae);
                  if ($unsigned($unsigned((~&reg6575))))
                    begin
                      reg6740 <= (~|forvar6629);
                      reg6741 <= forvar6253[(3'h7):(3'h5)];
                      reg6742 <= reg6441[(4'h8):(4'h8)];
                      reg6743 <= {(~&reg6649)};
                    end
                  else
                    begin
                      reg6740 <= ({(~(reg6158 << reg6268))} - (reg6168[(1'h0):(1'h0)] && $unsigned((reg6033 ?
                          (8'h9f) : reg6381))));
                      reg6741 <= ($signed((~(reg6505 ~^ reg6621))) ?
                          reg6172 : forvar6134);
                      reg6742 <= ((reg6648 || $signed($signed(reg6749))) ?
                          (reg6563 ?
                              $signed((8'hba)) : ((reg6759 > forvar6514) ?
                                  {reg6771} : (&reg6175))) : (($unsigned(forvar6465) ?
                                  reg6092[(1'h1):(1'h0)] : $signed(reg6470)) ?
                              {reg6711[(1'h1):(1'h0)]} : $signed(reg6379[(3'h5):(2'h2)])));
                    end
                end
            end
          if (reg6046)
            begin
              reg6744 <= $unsigned($unsigned((^~reg6761[(4'hd):(4'hd)])));
              for (forvar6745 = (1'h0); (forvar6745 < (1'h1)); forvar6745 = (forvar6745 + (1'h1)))
                begin
                  for (forvar6746 = (1'h0); (forvar6746 < (1'h0)); forvar6746 = (forvar6746 + (1'h1)))
                    begin
                      reg6747 <= $signed($unsigned({$signed(forvar6470)}));
                    end
                  if ($signed((~^reg6397)))
                    begin
                      reg6748 <= $unsigned($unsigned((reg6033[(1'h1):(1'h0)] & reg6656[(1'h1):(1'h1)])));
                      reg6749 <= (($unsigned(((8'hb2) ?
                          reg6632 : reg6514)) & reg6171) >= ($unsigned((^reg6736)) ^~ $unsigned(forvar6020[(1'h1):(1'h1)])));
                    end
                  else
                    begin
                      reg6748 <= reg6451[(3'h5):(3'h4)];
                      reg6749 <= reg6289[(1'h0):(1'h0)];
                      reg6750 <= ($unsigned($unsigned(reg6304)) ?
                          $unsigned(reg6692[(2'h3):(2'h2)]) : $signed(((~forvar6111) ?
                              (forvar6649 ~^ forvar6232) : $signed((8'hb1)))));
                      reg6751 <= ($unsigned({(forvar6637 ?
                                  forvar6621 : reg6187)}) ?
                          reg6654[(2'h3):(1'h1)] : forvar6212[(1'h1):(1'h1)]);
                    end
                  for (forvar6752 = (1'h0); (forvar6752 < (1'h0)); forvar6752 = (forvar6752 + (1'h1)))
                    begin
                      reg6753 <= reg6333;
                      reg6754 <= $unsigned(reg6742);
                    end
                  for (forvar6755 = (1'h0); (forvar6755 < (2'h2)); forvar6755 = (forvar6755 + (1'h1)))
                    begin
                      reg6756 <= {(((forvar6732 ?
                              forvar6120 : forvar6110) >>> $signed(forvar6303)) == (reg6407 < ((8'hac) * reg6696)))};
                      reg6757 <= $unsigned(reg6110);
                    end
                end
            end
          else
            begin
              for (forvar6744 = (1'h0); (forvar6744 < (1'h1)); forvar6744 = (forvar6744 + (1'h1)))
                begin
                  if (({reg6320[(3'h5):(1'h1)]} >>> $unsigned(reg6034)))
                    begin
                      reg6745 <= $unsigned($unsigned($unsigned($signed(forvar6209))));
                      reg6746 <= reg6199[(3'h4):(1'h0)];
                      reg6747 <= (forvar6658[(2'h3):(2'h2)] ?
                          (!forvar6283) : $unsigned((^(reg6730 ?
                              (8'hae) : reg6200))));
                      reg6748 <= (8'hb9);
                    end
                  else
                    begin
                      reg6745 <= $signed((~&$unsigned(((8'hb6) ^~ reg6476))));
                      reg6746 <= $unsigned(reg6628[(3'h7):(3'h4)]);
                      reg6747 <= (wire6218[(4'hb):(3'h7)] ?
                          reg6102 : (($unsigned(reg6667) < (reg6263 & (8'hb7))) || reg6289));
                      reg6748 <= (reg6613 ?
                          $signed(reg6377) : forvar6081[(2'h2):(1'h1)]);
                    end
                  for (forvar6749 = (1'h0); (forvar6749 < (1'h1)); forvar6749 = (forvar6749 + (1'h1)))
                    begin
                      reg6750 <= forvar6347[(2'h2):(2'h2)];
                      reg6751 <= ((^~(reg6717 ?
                          $unsigned(forvar6639) : (forvar6745 ?
                              reg6551 : reg6580))) + {reg6183});
                      reg6752 <= (-(-reg6338));
                    end
                end
              if ((&$unsigned(($signed(reg6304) >= reg6334[(2'h2):(1'h0)]))))
                begin
                  if (((({(8'hab)} + forvar6055) || (8'ha3)) ?
                      $unsigned($signed(reg6759[(2'h2):(1'h1)])) : reg6667))
                    begin
                      reg6753 <= ($unsigned((reg6720 ?
                          (8'haf) : $signed(reg6614))) & forvar6592);
                      reg6754 <= {reg6041[(2'h3):(2'h3)]};
                      reg6755 <= $unsigned(reg6710);
                      reg6756 <= reg6739[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg6753 <= ($unsigned((forvar6726 ?
                          (reg6457 ?
                              forvar6512 : forvar6286) : {forvar6624})) > $unsigned((~|$signed(reg6136))));
                    end
                end
              else
                begin
                  for (forvar6753 = (1'h0); (forvar6753 < (2'h2)); forvar6753 = (forvar6753 + (1'h1)))
                    begin
                      reg6754 <= ((|reg6321[(1'h1):(1'h0)]) == {$signed((reg6086 == reg6466))});
                      reg6755 <= {$signed((reg6523 ?
                              $unsigned(forvar6332) : forvar6198[(2'h2):(1'h1)]))};
                      reg6756 <= reg6490[(1'h1):(1'h0)];
                    end
                end
            end
          reg6758 <= $signed((forvar6221[(3'h4):(3'h4)] ?
              $signed(reg6605[(4'h8):(1'h0)]) : forvar6393[(4'h8):(1'h1)]));
          for (forvar6759 = (1'h0); (forvar6759 < (2'h2)); forvar6759 = (forvar6759 + (1'h1)))
            begin
              for (forvar6760 = (1'h0); (forvar6760 < (2'h3)); forvar6760 = (forvar6760 + (1'h1)))
                begin
                  reg6761 <= ((^$signed(reg6243)) * reg6705);
                end
              reg6762 <= (reg6531 == ((|((8'hb4) ?
                  (8'hb8) : reg6348)) == ($unsigned(reg6474) ?
                  (~&forvar6463) : (reg6635 | (8'had)))));
              if ((|$signed({(^forvar6623)})))
                begin
                  if ($signed((8'h9c)))
                    begin
                      reg6763 <= {((reg6383 <<< (~reg6762)) ?
                              ((reg6649 >> reg6345) ^~ (forvar6571 == reg6734)) : {reg6535})};
                      reg6764 <= ((8'hb5) >= $unsigned((^reg6710)));
                      reg6765 <= $signed($signed(($signed(reg6714) ?
                          reg6505 : (reg6600 ? (8'ha0) : reg6539))));
                    end
                  else
                    begin
                      reg6763 <= reg6755[(4'h8):(2'h2)];
                    end
                  if ($unsigned((~|$signed(reg6205))))
                    begin
                      reg6766 <= reg6160[(2'h3):(2'h3)];
                      reg6767 <= {(~&$signed($signed(forvar6557)))};
                      reg6768 <= reg6278[(4'ha):(3'h7)];
                      reg6769 <= {forvar6534};
                    end
                  else
                    begin
                      reg6766 <= reg6077[(1'h0):(1'h0)];
                      reg6767 <= (($signed((reg6107 ~^ reg6266)) < {reg6741[(3'h4):(1'h1)]}) != reg6248[(3'h6):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar6763 = (1'h0); (forvar6763 < (2'h2)); forvar6763 = (forvar6763 + (1'h1)))
                    begin
                      reg6764 <= reg6112[(2'h2):(1'h0)];
                      reg6765 <= ($signed((reg6719[(1'h1):(1'h1)] ?
                          (-reg6761) : (forvar6649 ?
                              (8'hb6) : reg6597))) + $signed(forvar6431[(1'h0):(1'h0)]));
                    end
                  reg6766 <= (((^(reg6124 < reg6461)) ?
                      $signed(reg6093) : {(reg6523 >= reg6162)}) + (~^reg6683[(2'h2):(1'h0)]));
                end
              reg6770 <= $unsigned($signed(($signed((8'hb3)) <<< (reg6196 * reg6679))));
            end
        end
      for (forvar6772 = (1'h0); (forvar6772 < (2'h2)); forvar6772 = (forvar6772 + (1'h1)))
        begin
          if (reg6086[(3'h7):(3'h6)])
            begin
              if (reg6127)
                begin
                  reg6773 <= reg6380;
                  if ($unsigned((&$unsigned({reg6047}))))
                    begin
                      reg6774 <= reg6404[(2'h3):(1'h1)];
                      reg6775 <= forvar6583;
                      reg6776 <= reg6407[(3'h7):(2'h3)];
                      reg6777 <= forvar6209;
                    end
                  else
                    begin
                      reg6774 <= reg6408;
                      reg6775 <= $signed((~^$signed($unsigned((8'h9d)))));
                    end
                  if ((!(+forvar6492)))
                    begin
                      reg6778 <= (|reg6108);
                    end
                  else
                    begin
                      reg6778 <= $unsigned({(~&reg6663[(3'h7):(1'h1)])});
                      reg6779 <= $unsigned((($signed(reg6274) ?
                              (!reg6330) : forvar6164[(1'h0):(1'h0)]) ?
                          ((8'ha1) >>> (reg6769 && forvar6243)) : {forvar6452}));
                      reg6780 <= (((~&(~&reg6071)) ?
                          $signed((reg6110 ?
                              forvar6676 : (8'hac))) : $signed($unsigned(reg6067))) <= ($signed(reg6566) ?
                          $unsigned($unsigned(reg6419)) : reg6449));
                      reg6781 <= ((reg6663[(4'h9):(3'h5)] << (~(~|reg6255))) >= $signed({$unsigned(reg6109)}));
                    end
                  if ((reg6392 || $unsigned(reg6358[(1'h1):(1'h0)])))
                    begin
                      reg6782 <= (reg6640[(4'ha):(4'ha)] ?
                          forvar6649 : ($signed(reg6255[(2'h3):(1'h1)]) ^~ reg6358));
                    end
                  else
                    begin
                      reg6782 <= (|reg6747[(3'h6):(2'h3)]);
                    end
                end
              else
                begin
                  if ($unsigned(reg6514))
                    begin
                      reg6773 <= $unsigned($unsigned(reg6575[(3'h5):(1'h0)]));
                    end
                  else
                    begin
                      reg6773 <= $signed($signed(forvar6646[(3'h6):(3'h6)]));
                    end
                  for (forvar6774 = (1'h0); (forvar6774 < (2'h2)); forvar6774 = (forvar6774 + (1'h1)))
                    begin
                      reg6775 <= ((($unsigned(reg6150) | {reg6369}) > ($signed(reg6754) >= (reg6136 >> reg6732))) > $signed(($signed(forvar6020) ?
                          forvar6171[(1'h0):(1'h0)] : (~^reg6299))));
                      reg6776 <= reg6392[(2'h2):(2'h2)];
                      reg6777 <= $unsigned($signed((+(reg6082 >> reg6704))));
                      reg6778 <= $unsigned((((reg6382 ?
                          (8'h9f) : reg6402) - (~^(8'ha8))) - $unsigned((reg6181 & forvar6483))));
                    end
                  for (forvar6779 = (1'h0); (forvar6779 < (2'h3)); forvar6779 = (forvar6779 + (1'h1)))
                    begin
                      reg6780 <= ({(reg6250 ?
                              $unsigned(reg6383) : forvar6178)} || reg6753);
                      reg6781 <= reg6034;
                      reg6782 <= ((((reg6551 ~^ forvar6774) ?
                          $unsigned(forvar6609) : {reg6532}) && reg6642) >= ($unsigned($unsigned((8'ha0))) ?
                          reg6205 : ((reg6580 * reg6188) ?
                              (8'ha3) : $signed(forvar6772))));
                    end
                  for (forvar6783 = (1'h0); (forvar6783 < (2'h3)); forvar6783 = (forvar6783 + (1'h1)))
                    begin
                      reg6784 <= forvar6392;
                      reg6785 <= (^$signed((^~(reg6338 ?
                          forvar6641 : forvar6624))));
                      reg6786 <= {$unsigned(($unsigned(reg6048) ?
                              forvar6452[(3'h4):(1'h1)] : (reg6767 ?
                                  forvar6559 : reg6572)))};
                      reg6787 <= (~^forvar6394[(4'hd):(3'h4)]);
                    end
                end
              if (($unsigned(($signed(reg6604) ?
                  (~|reg6137) : (forvar6469 >> (8'hb9)))) >>> forvar6769))
                begin
                  reg6788 <= (8'ha7);
                  if (reg6285[(4'hb):(4'h9)])
                    begin
                      reg6789 <= {reg6326};
                      reg6790 <= $unsigned(reg6108);
                    end
                  else
                    begin
                      reg6789 <= reg6170[(3'h4):(2'h3)];
                      reg6790 <= $signed((+forvar6579[(2'h2):(2'h2)]));
                      reg6791 <= (^~{$unsigned((forvar6750 != forvar6073))});
                    end
                  reg6792 <= $unsigned($signed(reg6111));
                end
              else
                begin
                  if ((^(forvar6371 ? (8'hb0) : reg6185[(4'ha):(4'h8)])))
                    begin
                      reg6788 <= ((forvar6680 & (forvar6392[(1'h1):(1'h0)] ?
                              {reg6539} : $unsigned((8'hb4)))) ?
                          reg6536 : reg6738);
                    end
                  else
                    begin
                      reg6788 <= reg6294;
                      reg6789 <= $unsigned($unsigned(({forvar6491} >= reg6101[(2'h2):(1'h1)])));
                      reg6790 <= ($unsigned(reg6193[(1'h0):(1'h0)]) ?
                          (-reg6170) : $unsigned(reg6378));
                      reg6791 <= {(wire5508 || reg6189)};
                    end
                  reg6792 <= ($unsigned($unsigned((~&reg6194))) ~^ $unsigned(forvar6377));
                  for (forvar6793 = (1'h0); (forvar6793 < (2'h2)); forvar6793 = (forvar6793 + (1'h1)))
                    begin
                      reg6794 <= ((((reg6342 ?
                              reg6152 : (8'hab)) ~^ (~|(8'hb3))) < (+{forvar6464})) ?
                          $unsigned(reg6053[(2'h3):(2'h2)]) : ($unsigned($unsigned(reg6289)) == reg6590[(3'h4):(2'h2)]));
                    end
                end
              for (forvar6795 = (1'h0); (forvar6795 < (2'h2)); forvar6795 = (forvar6795 + (1'h1)))
                begin
                  for (forvar6796 = (1'h0); (forvar6796 < (1'h1)); forvar6796 = (forvar6796 + (1'h1)))
                    begin
                      reg6797 <= (^$unsigned((((8'h9d) ? forvar6701 : (8'ha3)) ?
                          (reg6167 ? reg6287 : forvar6161) : (8'hb6))));
                      reg6798 <= ($unsigned(($unsigned(forvar6179) ?
                          (reg6467 != (8'ha8)) : $unsigned(reg6399))) < {$unsigned($signed(reg6757))});
                      reg6799 <= $signed((^($unsigned(reg6394) << (reg6693 ?
                          reg6778 : (8'ha9)))));
                      reg6800 <= reg6222[(1'h1):(1'h0)];
                    end
                  for (forvar6801 = (1'h0); (forvar6801 < (2'h3)); forvar6801 = (forvar6801 + (1'h1)))
                    begin
                      reg6802 <= ({(!$unsigned(forvar6498))} ?
                          (!((reg6623 ?
                              forvar6234 : forvar6496) | (|forvar6453))) : ({reg6571[(1'h1):(1'h1)]} ^~ $signed($unsigned(forvar6324))));
                    end
                  if ((^~($signed((~^reg6129)) >> reg6124[(1'h0):(1'h0)])))
                    begin
                      reg6803 <= {reg6425};
                    end
                  else
                    begin
                      reg6803 <= ((-reg6063[(4'ha):(4'h9)]) ?
                          $unsigned(forvar6332) : $unsigned((+{reg6117})));
                    end
                  if ({(&reg6125[(4'hd):(3'h4)])})
                    begin
                      reg6804 <= ((8'had) < ((~&$unsigned(reg6593)) ^ ((reg6361 ?
                          (8'ha1) : reg6240) ^~ {reg6533})));
                      reg6805 <= {$signed((reg6758 <<< (|reg6771)))};
                      reg6806 <= {(^~($unsigned(forvar6393) - {reg6429}))};
                    end
                  else
                    begin
                      reg6804 <= $unsigned({$signed($signed((8'h9f)))});
                      reg6805 <= {$unsigned(forvar6507)};
                      reg6806 <= (reg6129 ^~ ($signed(reg6242) ?
                          ({reg6321} ?
                              ((8'hb7) ?
                                  reg6119 : forvar6168) : $signed(forvar6756)) : ($signed(reg6517) ?
                              forvar6366 : {reg6560})));
                    end
                end
            end
          else
            begin
              if ({{$unsigned((reg6700 * reg6503))}})
                begin
                  reg6773 <= {$unsigned($signed(reg6638[(3'h5):(3'h5)]))};
                  if (((-reg6677[(2'h3):(2'h2)]) ~^ (($signed(reg6688) < (~^reg6633)) ?
                      reg6350 : (8'ha2))))
                    begin
                      reg6774 <= (($unsigned(reg6660[(4'hc):(4'h9)]) | ((forvar6687 ?
                              forvar6253 : (8'h9d)) + (-forvar6597))) ?
                          (|reg6135) : $unsigned($unsigned($unsigned(reg6791))));
                      reg6775 <= $signed(reg6422);
                      reg6776 <= $signed(reg6485);
                      reg6777 <= ($unsigned((reg6182[(2'h2):(1'h0)] ?
                          $unsigned(reg6109) : $signed(reg6505))) ^~ (reg6199 + {reg6513}));
                    end
                  else
                    begin
                      reg6774 <= reg6346;
                      reg6775 <= ((~(+$unsigned(reg6390))) == (8'hb4));
                      reg6776 <= $unsigned((+$unsigned(reg6760)));
                    end
                  if ((reg6587 ?
                      (!$signed((-reg6409))) : ($signed(((8'ha1) ?
                              reg6274 : reg6512)) ?
                          ($signed(reg6259) ?
                              (8'ha5) : $signed(reg6657)) : (&$signed(forvar6122)))))
                    begin
                      reg6778 <= (forvar6202[(3'h7):(1'h1)] ?
                          {((forvar6195 ?
                                  reg6259 : reg6600) > $signed(forvar6120))} : $unsigned($signed((^~reg6508))));
                      reg6779 <= (~|forvar6762[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg6778 <= reg6436[(4'ha):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar6773 = (1'h0); (forvar6773 < (1'h1)); forvar6773 = (forvar6773 + (1'h1)))
                    begin
                      reg6774 <= (!{forvar6078});
                    end
                  for (forvar6775 = (1'h0); (forvar6775 < (2'h3)); forvar6775 = (forvar6775 + (1'h1)))
                    begin
                      reg6776 <= reg6696[(1'h1):(1'h0)];
                      reg6777 <= {(reg6256[(4'he):(3'h6)] ?
                              $unsigned((wire6443 ?
                                  forvar6513 : reg6207)) : ((8'ha6) ?
                                  (+forvar6579) : (wire6218 ?
                                      forvar6111 : forvar6502)))};
                      reg6778 <= ($signed((reg6503[(3'h4):(1'h0)] < reg6022[(2'h2):(1'h1)])) ?
                          reg6254[(1'h1):(1'h0)] : {reg6375});
                    end
                  if ((reg6732 ?
                      reg6640 : ((reg6032[(4'h8):(2'h2)] ?
                          (forvar6312 + forvar6435) : $unsigned(reg6271)) * reg6080)))
                    begin
                      reg6779 <= {reg6359};
                    end
                  else
                    begin
                      reg6779 <= $unsigned(reg6797);
                      reg6780 <= ((&(8'haa)) ?
                          $signed(reg6717[(2'h3):(1'h1)]) : reg6203[(2'h2):(2'h2)]);
                      reg6781 <= $unsigned(((&$unsigned(reg6643)) ?
                          $unsigned(((8'hab) ?
                              (8'ha5) : (8'ha6))) : ($signed(reg6112) >= (8'h9f))));
                    end
                  if (forvar6522[(1'h1):(1'h1)])
                    begin
                      reg6782 <= reg6489;
                      reg6783 <= reg6070[(3'h7):(1'h1)];
                    end
                  else
                    begin
                      reg6782 <= reg6275[(1'h1):(1'h1)];
                      reg6783 <= (^$signed(reg6093[(3'h7):(1'h0)]));
                    end
                end
              for (forvar6784 = (1'h0); (forvar6784 < (1'h1)); forvar6784 = (forvar6784 + (1'h1)))
                begin
                  reg6785 <= $signed($signed($signed((~&reg6285))));
                end
              reg6786 <= (8'haa);
            end
          if ((~&{{$unsigned(reg6607)}}))
            begin
              for (forvar6807 = (1'h0); (forvar6807 < (1'h1)); forvar6807 = (forvar6807 + (1'h1)))
                begin
                  for (forvar6808 = (1'h0); (forvar6808 < (1'h0)); forvar6808 = (forvar6808 + (1'h1)))
                    begin
                      reg6809 <= reg6557[(2'h2):(2'h2)];
                    end
                  for (forvar6810 = (1'h0); (forvar6810 < (1'h1)); forvar6810 = (forvar6810 + (1'h1)))
                    begin
                      reg6811 <= {(8'ha3)};
                      reg6812 <= $unsigned(($signed($unsigned((8'haa))) ?
                          reg6656[(4'hb):(2'h3)] : $signed($unsigned((8'hba)))));
                    end
                  if ({forvar6411})
                    begin
                      reg6813 <= (reg6395[(3'h6):(3'h4)] ?
                          (^(-{forvar6387})) : (reg6101[(3'h6):(3'h4)] ?
                              {reg6174[(1'h0):(1'h0)]} : reg6354));
                      reg6814 <= (reg6501 ?
                          ((8'hb5) ?
                              $signed(forvar6317[(1'h0):(1'h0)]) : reg6505[(3'h6):(1'h0)]) : $unsigned({$unsigned(reg6259)}));
                    end
                  else
                    begin
                      reg6813 <= forvar6564[(3'h4):(1'h1)];
                      reg6814 <= (reg6572[(1'h0):(1'h0)] + reg6670);
                      reg6815 <= wire6617;
                    end
                  if (forvar6111[(3'h6):(2'h2)])
                    begin
                      reg6816 <= (^$unsigned(forvar6521));
                      reg6817 <= reg6600;
                    end
                  else
                    begin
                      reg6816 <= $unsigned((^$unsigned((reg6123 ?
                          (8'haf) : reg6449))));
                    end
                end
            end
          else
            begin
              for (forvar6807 = (1'h0); (forvar6807 < (1'h1)); forvar6807 = (forvar6807 + (1'h1)))
                begin
                  for (forvar6808 = (1'h0); (forvar6808 < (1'h0)); forvar6808 = (forvar6808 + (1'h1)))
                    begin
                      reg6809 <= ($signed(reg6113[(1'h0):(1'h0)]) + reg6514);
                    end
                  if (($signed($signed(reg6741[(1'h0):(1'h0)])) ?
                      (((!(8'ha7)) && (~^reg6148)) ?
                          reg6647[(4'hc):(4'h8)] : $signed((reg6040 > reg6697))) : $signed($signed((forvar6406 ?
                          forvar6405 : forvar6045)))))
                    begin
                      reg6810 <= forvar6592[(1'h0):(1'h0)];
                      reg6811 <= $signed(reg6064);
                      reg6812 <= {($unsigned({reg6740}) ^ ({reg6679} ?
                              (+(8'hb0)) : {(8'hb2)}))};
                    end
                  else
                    begin
                      reg6810 <= ({(forvar6307 ?
                              (reg6672 > (8'ha3)) : (+reg6031))} & reg6115[(2'h3):(1'h0)]);
                      reg6811 <= (~^reg6381[(3'h6):(2'h2)]);
                      reg6812 <= reg6355[(3'h7):(2'h2)];
                      reg6813 <= forvar6327[(2'h3):(1'h1)];
                    end
                  if ($unsigned($signed(forvar6680[(1'h1):(1'h1)])))
                    begin
                      reg6814 <= (reg6673 ?
                          reg6354[(2'h2):(1'h1)] : $unsigned(reg6117[(4'h9):(1'h1)]));
                      reg6815 <= $unsigned($signed(((reg6408 ?
                              reg6625 : (8'hae)) ?
                          reg6506[(3'h6):(3'h4)] : $signed(reg6333))));
                      reg6816 <= $signed($unsigned($signed($unsigned(reg6478))));
                      reg6817 <= (^~(|reg6403));
                    end
                  else
                    begin
                      reg6814 <= {$unsigned(reg6134[(3'h7):(3'h6)])};
                      reg6815 <= $unsigned((~|{forvar6595[(2'h2):(1'h0)]}));
                      reg6816 <= $signed((((8'h9d) ?
                              $unsigned(reg6780) : (^forvar6097)) ?
                          $unsigned((reg6272 ?
                              reg6647 : forvar6270)) : $signed((+reg6475))));
                      reg6817 <= ((&$signed((reg6128 ?
                          reg6473 : (8'hba)))) + reg6376[(3'h4):(3'h4)]);
                    end
                  reg6818 <= $signed((^~reg6125[(4'hc):(3'h5)]));
                end
              for (forvar6819 = (1'h0); (forvar6819 < (2'h2)); forvar6819 = (forvar6819 + (1'h1)))
                begin
                  reg6820 <= $unsigned(reg6151[(4'hd):(4'hc)]);
                  if ($unsigned($signed((8'hae))))
                    begin
                      reg6821 <= (&$signed($unsigned((8'hb3))));
                      reg6822 <= reg6821[(3'h4):(2'h3)];
                    end
                  else
                    begin
                      reg6821 <= reg6580;
                      reg6822 <= ($signed($unsigned($unsigned(forvar6411))) ^ $unsigned((reg6063[(4'hb):(3'h7)] ?
                          reg6547 : (forvar6644 <<< (8'hae)))));
                    end
                end
            end
          reg6823 <= (reg6091[(3'h7):(2'h2)] ^~ $signed((reg6117 ?
              (reg6565 ? forvar6645 : reg6551) : forvar6087)));
          for (forvar6824 = (1'h0); (forvar6824 < (1'h0)); forvar6824 = (forvar6824 + (1'h1)))
            begin
              for (forvar6825 = (1'h0); (forvar6825 < (2'h3)); forvar6825 = (forvar6825 + (1'h1)))
                begin
                  for (forvar6826 = (1'h0); (forvar6826 < (2'h2)); forvar6826 = (forvar6826 + (1'h1)))
                    begin
                      reg6827 <= reg6612;
                      reg6828 <= $signed(forvar6732[(2'h2):(1'h0)]);
                    end
                  for (forvar6829 = (1'h0); (forvar6829 < (1'h1)); forvar6829 = (forvar6829 + (1'h1)))
                    begin
                      reg6830 <= $signed(reg6473);
                      reg6831 <= {reg6059};
                    end
                  reg6832 <= $unsigned(reg6621);
                  for (forvar6833 = (1'h0); (forvar6833 < (2'h3)); forvar6833 = (forvar6833 + (1'h1)))
                    begin
                      reg6834 <= (((forvar6035 - (&forvar6269)) < reg6308) - (+$unsigned($unsigned(reg6784))));
                      reg6835 <= (&($unsigned((^~wire5506)) * $unsigned(reg6630[(1'h1):(1'h1)])));
                      reg6836 <= (reg6080[(4'h8):(3'h5)] ?
                          forvar6220[(4'he):(4'h8)] : (+$unsigned({forvar6744})));
                      reg6837 <= reg6294[(1'h0):(1'h0)];
                    end
                end
            end
        end
      for (forvar6838 = (1'h0); (forvar6838 < (1'h1)); forvar6838 = (forvar6838 + (1'h1)))
        begin
          for (forvar6839 = (1'h0); (forvar6839 < (1'h1)); forvar6839 = (forvar6839 + (1'h1)))
            begin
              for (forvar6840 = (1'h0); (forvar6840 < (2'h3)); forvar6840 = (forvar6840 + (1'h1)))
                begin
                  if (reg6268[(4'ha):(3'h7)])
                    begin
                      reg6841 <= (~^($signed(reg6385[(2'h2):(1'h0)]) ?
                          $unsigned(reg6369) : (^~$unsigned(forvar6452))));
                      reg6842 <= reg6631;
                      reg6843 <= ($unsigned((~(forvar6629 >= reg6381))) ?
                          {(~&((8'h9c) ? reg6525 : forvar6088))} : ((!(reg6130 ?
                                  forvar6134 : (8'ha6))) ?
                              wire6443[(3'h6):(3'h4)] : reg6173[(4'hc):(3'h5)]));
                      reg6844 <= (!$signed($unsigned({reg6689})));
                    end
                  else
                    begin
                      reg6841 <= (!reg6605);
                      reg6842 <= forvar6335[(1'h0):(1'h0)];
                      reg6843 <= $signed({$unsigned((forvar6464 == reg6378))});
                      reg6844 <= ({$unsigned((reg6262 & (8'hb5)))} ^ (((forvar6562 ~^ forvar6209) ?
                          {forvar6825} : reg6399[(1'h1):(1'h0)]) | ($unsigned(forvar6745) ?
                          $unsigned(reg6356) : (reg6315 ?
                              reg6433 : forvar6808))));
                    end
                  for (forvar6845 = (1'h0); (forvar6845 < (1'h0)); forvar6845 = (forvar6845 + (1'h1)))
                    begin
                      reg6846 <= $unsigned($unsigned($signed((forvar6352 ?
                          reg6656 : (8'ha3)))));
                      reg6847 <= $unsigned(((reg6533 ^ $unsigned((8'h9e))) >> reg6717[(3'h5):(3'h5)]));
                    end
                  reg6848 <= (+{forvar6164});
                end
            end
          for (forvar6849 = (1'h0); (forvar6849 < (2'h3)); forvar6849 = (forvar6849 + (1'h1)))
            begin
              for (forvar6850 = (1'h0); (forvar6850 < (2'h2)); forvar6850 = (forvar6850 + (1'h1)))
                begin
                  for (forvar6851 = (1'h0); (forvar6851 < (1'h1)); forvar6851 = (forvar6851 + (1'h1)))
                    begin
                      reg6852 <= $signed((8'ha2));
                    end
                  for (forvar6853 = (1'h0); (forvar6853 < (1'h0)); forvar6853 = (forvar6853 + (1'h1)))
                    begin
                      reg6854 <= $signed(reg6564);
                      reg6855 <= forvar6453[(3'h5):(1'h1)];
                      reg6856 <= reg6468;
                    end
                  if (($unsigned(reg6466[(1'h1):(1'h1)]) ?
                      reg6512 : forvar6772))
                    begin
                      reg6857 <= $signed(($unsigned(forvar6808[(1'h0):(1'h0)]) ?
                          ((forvar6094 ? reg6313 : reg6638) ?
                              (reg6601 * reg6756) : (8'h9c)) : (reg6650 ?
                              $signed(reg6251) : (8'ha8))));
                    end
                  else
                    begin
                      reg6857 <= $unsigned((((^reg6755) > forvar6680) > ($signed(reg6396) ?
                          ((8'ha3) ? reg6527 : reg6747) : ((8'hba) ?
                              reg6098 : reg6448))));
                      reg6858 <= (~|(+$signed(reg6321[(2'h2):(1'h0)])));
                      reg6859 <= $unsigned($unsigned($signed(reg6170[(3'h4):(2'h2)])));
                      reg6860 <= $unsigned($signed(((reg6032 * reg6666) + (reg6510 | forvar6637))));
                    end
                end
            end
        end
    end
  assign wire6861 = $unsigned(reg6406[(1'h0):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module5511
#( parameter param6015 = ((-(((8'hba) | (8'ha6)) < (~(8'ha3)))) ? (&({(8'had)} >= (~|(8'ha2)))) : (~^(((8'ha8) ? (8'hae) : (8'haa)) ? ((8'hb5) ? (8'hb0) : (8'haf)) : (|(8'ha7))))) )
(y, clk, wire5515, wire5514, wire5513, wire5512);
  output wire [(32'h151c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire5515;
  input wire signed [(3'h5):(1'h0)] wire5514;
  input wire signed [(4'h8):(1'h0)] wire5513;
  input wire signed [(3'h6):(1'h0)] wire5512;
  reg [(5'h10):(1'h0)] reg6014 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6013 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6002 = (1'h0);
  reg [(4'he):(1'h0)] reg6012 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar6011 = (1'h0);
  reg [(4'h8):(1'h0)] reg6010 = (1'h0);
  reg [(2'h2):(1'h0)] reg6009 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg6008 = (1'h0);
  reg [(4'hd):(1'h0)] reg6007 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg6006 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg6005 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6004 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg6003 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6002 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6001 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar6000 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5999 = (1'h0);
  reg [(4'hd):(1'h0)] reg5998 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5997 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5996 = (1'h0);
  reg [(4'he):(1'h0)] forvar5995 = (1'h0);
  reg [(5'h10):(1'h0)] reg5994 = (1'h0);
  reg [(4'hb):(1'h0)] reg5993 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5992 = (1'h0);
  reg [(3'h4):(1'h0)] reg5991 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5990 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5989 = (1'h0);
  reg [(4'h9):(1'h0)] reg5989 = (1'h0);
  reg [(4'ha):(1'h0)] reg5988 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5987 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5986 = (1'h0);
  reg [(4'hb):(1'h0)] reg5985 = (1'h0);
  reg [(4'hd):(1'h0)] reg5984 = (1'h0);
  reg [(4'ha):(1'h0)] reg5983 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5982 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5981 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5980 = (1'h0);
  reg [(4'hd):(1'h0)] reg5979 = (1'h0);
  reg [(3'h5):(1'h0)] reg5978 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5977 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5976 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5975 = (1'h0);
  reg [(4'hc):(1'h0)] reg5974 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5973 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5972 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5971 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5970 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5969 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5968 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5967 = (1'h0);
  reg [(4'h8):(1'h0)] reg5966 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5965 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar5964 = (1'h0);
  reg [(4'h8):(1'h0)] reg5963 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5962 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5961 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5960 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5959 = (1'h0);
  reg [(4'h9):(1'h0)] reg5958 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5957 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5956 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5955 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5954 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5953 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5952 = (1'h0);
  reg [(3'h7):(1'h0)] reg5951 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5950 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5949 = (1'h0);
  reg [(4'hf):(1'h0)] reg5948 = (1'h0);
  reg [(3'h7):(1'h0)] reg5947 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5946 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5945 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5944 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5943 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5942 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5941 = (1'h0);
  reg [(3'h5):(1'h0)] reg5940 = (1'h0);
  reg [(4'hc):(1'h0)] reg5939 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5938 = (1'h0);
  reg [(3'h6):(1'h0)] reg5937 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5936 = (1'h0);
  reg [(3'h5):(1'h0)] reg5935 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5934 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5933 = (1'h0);
  reg [(3'h7):(1'h0)] reg5932 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5931 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5930 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5929 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5928 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5927 = (1'h0);
  reg [(4'h9):(1'h0)] reg5926 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5919 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5918 = (1'h0);
  reg [(4'hd):(1'h0)] reg5925 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5924 = (1'h0);
  reg [(3'h6):(1'h0)] reg5923 = (1'h0);
  reg [(3'h6):(1'h0)] reg5922 = (1'h0);
  reg [(4'he):(1'h0)] reg5921 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5920 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5919 = (1'h0);
  reg [(4'hb):(1'h0)] reg5918 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5917 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5916 = (1'h0);
  reg [(4'h9):(1'h0)] reg5915 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5914 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5913 = (1'h0);
  reg [(3'h4):(1'h0)] reg5912 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5911 = (1'h0);
  reg [(5'h10):(1'h0)] reg5910 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5909 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5908 = (1'h0);
  reg [(4'hc):(1'h0)] reg5907 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5906 = (1'h0);
  reg [(4'ha):(1'h0)] reg5905 = (1'h0);
  reg [(3'h7):(1'h0)] reg5904 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5903 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5902 = (1'h0);
  reg [(5'h10):(1'h0)] reg5901 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5900 = (1'h0);
  reg [(4'hf):(1'h0)] reg5899 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5898 = (1'h0);
  reg [(3'h7):(1'h0)] reg5897 = (1'h0);
  reg [(3'h5):(1'h0)] reg5896 = (1'h0);
  reg [(4'ha):(1'h0)] reg5895 = (1'h0);
  reg [(2'h3):(1'h0)] reg5894 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5893 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5892 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5891 = (1'h0);
  reg [(4'he):(1'h0)] forvar5890 = (1'h0);
  reg [(5'h10):(1'h0)] reg5889 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5888 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5887 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5886 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5885 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5884 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5883 = (1'h0);
  reg [(4'hd):(1'h0)] reg5882 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5881 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5880 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5879 = (1'h0);
  reg [(4'ha):(1'h0)] reg5878 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5875 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5870 = (1'h0);
  reg [(4'h8):(1'h0)] reg5877 = (1'h0);
  reg [(3'h7):(1'h0)] reg5876 = (1'h0);
  reg [(4'he):(1'h0)] reg5875 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5874 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5873 = (1'h0);
  reg [(4'hd):(1'h0)] reg5872 = (1'h0);
  reg [(4'hf):(1'h0)] reg5871 = (1'h0);
  reg [(4'hf):(1'h0)] reg5870 = (1'h0);
  reg [(4'hc):(1'h0)] reg5869 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5868 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5867 = (1'h0);
  wire [(3'h5):(1'h0)] wire5866;
  wire signed [(3'h5):(1'h0)] wire5865;
  wire [(4'h8):(1'h0)] wire5864;
  wire signed [(2'h2):(1'h0)] wire5863;
  reg signed [(5'h10):(1'h0)] reg5832 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5830 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5828 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5827 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5819 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5818 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5862 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5848 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5847 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5846 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5843 = (1'h0);
  reg [(2'h2):(1'h0)] reg5840 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5839 = (1'h0);
  reg [(4'hb):(1'h0)] reg5861 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5860 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5859 = (1'h0);
  reg [(2'h2):(1'h0)] reg5858 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5857 = (1'h0);
  reg [(4'ha):(1'h0)] reg5856 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5855 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5854 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5853 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5852 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5851 = (1'h0);
  reg [(3'h5):(1'h0)] reg5850 = (1'h0);
  reg [(4'h8):(1'h0)] reg5849 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5848 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5847 = (1'h0);
  reg [(5'h10):(1'h0)] reg5846 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5845 = (1'h0);
  reg [(3'h5):(1'h0)] reg5844 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5843 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5842 = (1'h0);
  reg [(4'h8):(1'h0)] reg5841 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5840 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5839 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5838 = (1'h0);
  reg [(4'ha):(1'h0)] reg5837 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5836 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5820 = (1'h0);
  reg [(3'h6):(1'h0)] reg5826 = (1'h0);
  reg [(4'hb):(1'h0)] reg5823 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5829 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5835 = (1'h0);
  reg [(5'h10):(1'h0)] reg5834 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5833 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5832 = (1'h0);
  reg [(4'hf):(1'h0)] reg5831 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5830 = (1'h0);
  reg [(4'h9):(1'h0)] reg5829 = (1'h0);
  reg [(3'h7):(1'h0)] reg5828 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5827 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5826 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5817 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5825 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5824 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5823 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5822 = (1'h0);
  reg [(3'h5):(1'h0)] reg5821 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5820 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5819 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5818 = (1'h0);
  reg [(4'hb):(1'h0)] reg5817 = (1'h0);
  reg [(5'h10):(1'h0)] reg5816 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5815 = (1'h0);
  reg [(3'h7):(1'h0)] reg5814 = (1'h0);
  reg [(4'hf):(1'h0)] reg5813 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5812 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5811 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5810 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5809 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5808 = (1'h0);
  reg [(4'h8):(1'h0)] reg5807 = (1'h0);
  reg [(4'hd):(1'h0)] reg5806 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5805 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5804 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5803 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5802 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5801 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5800 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5799 = (1'h0);
  reg [(4'he):(1'h0)] reg5798 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5797 = (1'h0);
  reg [(2'h2):(1'h0)] reg5796 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5795 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5794 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5793 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5792 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5791 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5790 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5789 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5788 = (1'h0);
  reg [(4'hf):(1'h0)] reg5787 = (1'h0);
  reg [(4'h9):(1'h0)] reg5786 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5785 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5784 = (1'h0);
  reg [(4'ha):(1'h0)] reg5783 = (1'h0);
  reg [(2'h2):(1'h0)] reg5782 = (1'h0);
  reg [(2'h3):(1'h0)] reg5781 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5780 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5779 = (1'h0);
  reg [(4'h9):(1'h0)] reg5778 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5777 = (1'h0);
  reg [(3'h5):(1'h0)] reg5776 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5775 = (1'h0);
  reg [(4'hc):(1'h0)] reg5774 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5773 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5772 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5771 = (1'h0);
  reg [(3'h6):(1'h0)] reg5770 = (1'h0);
  reg [(4'ha):(1'h0)] reg5769 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5768 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5767 = (1'h0);
  reg [(3'h5):(1'h0)] reg5766 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5765 = (1'h0);
  reg [(3'h7):(1'h0)] reg5764 = (1'h0);
  reg [(4'he):(1'h0)] forvar5763 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5762 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5761 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5741 = (1'h0);
  reg [(4'hc):(1'h0)] reg5746 = (1'h0);
  reg [(3'h7):(1'h0)] reg5739 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5725 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5721 = (1'h0);
  reg [(4'he):(1'h0)] reg5730 = (1'h0);
  reg [(4'ha):(1'h0)] reg5738 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5734 = (1'h0);
  reg [(4'h9):(1'h0)] reg5733 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5726 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5720 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5718 = (1'h0);
  reg [(4'h8):(1'h0)] reg5716 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5760 = (1'h0);
  reg [(4'hc):(1'h0)] reg5759 = (1'h0);
  reg [(3'h7):(1'h0)] reg5758 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5757 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5756 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5752 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5751 = (1'h0);
  reg [(3'h6):(1'h0)] reg5756 = (1'h0);
  reg [(4'he):(1'h0)] reg5755 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5754 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5753 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5752 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5751 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5750 = (1'h0);
  reg [(4'hb):(1'h0)] reg5749 = (1'h0);
  reg [(4'hc):(1'h0)] reg5748 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5747 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5746 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5745 = (1'h0);
  reg [(2'h2):(1'h0)] reg5744 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5743 = (1'h0);
  reg [(4'hd):(1'h0)] reg5742 = (1'h0);
  reg [(4'h8):(1'h0)] reg5741 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5740 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5739 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5738 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5737 = (1'h0);
  reg [(4'hb):(1'h0)] reg5736 = (1'h0);
  reg [(4'hb):(1'h0)] reg5735 = (1'h0);
  reg [(3'h6):(1'h0)] reg5734 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5733 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5732 = (1'h0);
  reg [(4'ha):(1'h0)] reg5731 = (1'h0);
  reg [(3'h6):(1'h0)] forvar5730 = (1'h0);
  reg [(5'h10):(1'h0)] reg5729 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5728 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5727 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5726 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5725 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5724 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5723 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5722 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5721 = (1'h0);
  reg [(4'hb):(1'h0)] reg5720 = (1'h0);
  reg [(4'hf):(1'h0)] reg5719 = (1'h0);
  reg [(5'h10):(1'h0)] reg5718 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5717 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5717 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5716 = (1'h0);
  reg [(4'h8):(1'h0)] reg5715 = (1'h0);
  reg [(4'h8):(1'h0)] reg5714 = (1'h0);
  reg [(4'h8):(1'h0)] reg5713 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5712 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5709 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5703 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5700 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5695 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5687 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5683 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5679 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5670 = (1'h0);
  reg [(3'h5):(1'h0)] forvar5669 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5668 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5658 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5655 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5650 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5646 = (1'h0);
  reg [(2'h2):(1'h0)] reg5652 = (1'h0);
  reg [(3'h4):(1'h0)] reg5647 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5645 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5711 = (1'h0);
  reg [(4'h8):(1'h0)] reg5699 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5694 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5710 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5709 = (1'h0);
  reg [(2'h2):(1'h0)] reg5708 = (1'h0);
  reg [(3'h4):(1'h0)] reg5707 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5706 = (1'h0);
  reg [(2'h3):(1'h0)] reg5705 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5704 = (1'h0);
  reg [(4'h9):(1'h0)] reg5703 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5702 = (1'h0);
  reg [(4'hb):(1'h0)] reg5701 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5700 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar5699 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5698 = (1'h0);
  reg [(4'hf):(1'h0)] reg5697 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5696 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5695 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5694 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5693 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5692 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5691 = (1'h0);
  reg [(4'he):(1'h0)] reg5690 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5686 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5684 = (1'h0);
  reg [(4'hb):(1'h0)] forvar5681 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5680 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5677 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5675 = (1'h0);
  reg [(4'h8):(1'h0)] forvar5673 = (1'h0);
  reg [(4'hb):(1'h0)] reg5671 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5689 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5688 = (1'h0);
  reg [(4'hf):(1'h0)] reg5687 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5686 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5685 = (1'h0);
  reg [(5'h10):(1'h0)] reg5684 = (1'h0);
  reg [(3'h5):(1'h0)] reg5683 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5682 = (1'h0);
  reg [(4'hd):(1'h0)] reg5681 = (1'h0);
  reg [(4'hf):(1'h0)] reg5680 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5679 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5678 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5677 = (1'h0);
  reg [(3'h5):(1'h0)] reg5676 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5675 = (1'h0);
  reg [(2'h3):(1'h0)] reg5674 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5673 = (1'h0);
  reg [(4'h9):(1'h0)] reg5672 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5671 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar5670 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5663 = (1'h0);
  reg [(4'h9):(1'h0)] reg5662 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5669 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar5668 = (1'h0);
  reg [(4'he):(1'h0)] reg5667 = (1'h0);
  reg [(3'h6):(1'h0)] reg5666 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5665 = (1'h0);
  reg [(3'h4):(1'h0)] reg5664 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5663 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar5662 = (1'h0);
  reg [(4'he):(1'h0)] reg5661 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5660 = (1'h0);
  reg [(3'h5):(1'h0)] reg5659 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5658 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5657 = (1'h0);
  reg [(3'h4):(1'h0)] reg5656 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5655 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5654 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5653 = (1'h0);
  reg [(4'he):(1'h0)] forvar5652 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5651 = (1'h0);
  reg [(4'h9):(1'h0)] reg5650 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5649 = (1'h0);
  reg [(4'hf):(1'h0)] reg5648 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5647 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5646 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5645 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg5644 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire5643;
  wire signed [(4'h9):(1'h0)] wire5642;
  wire [(4'he):(1'h0)] wire5641;
  reg [(3'h7):(1'h0)] reg5640 = (1'h0);
  reg [(2'h2):(1'h0)] reg5639 = (1'h0);
  reg [(4'hc):(1'h0)] reg5638 = (1'h0);
  reg [(4'hf):(1'h0)] reg5637 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5636 = (1'h0);
  reg [(3'h4):(1'h0)] reg5635 = (1'h0);
  reg [(4'hd):(1'h0)] reg5634 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5633 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5632 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5631 = (1'h0);
  reg [(5'h10):(1'h0)] reg5630 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5629 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5628 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5627 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5626 = (1'h0);
  reg [(4'hd):(1'h0)] reg5625 = (1'h0);
  reg [(3'h7):(1'h0)] reg5624 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5623 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5622 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5621 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5620 = (1'h0);
  reg [(3'h7):(1'h0)] reg5619 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5618 = (1'h0);
  reg [(4'h8):(1'h0)] reg5617 = (1'h0);
  reg [(5'h10):(1'h0)] reg5616 = (1'h0);
  reg [(4'ha):(1'h0)] reg5615 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5614 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5613 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5612 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5611 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5610 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5609 = (1'h0);
  reg [(2'h2):(1'h0)] reg5608 = (1'h0);
  reg [(4'ha):(1'h0)] reg5607 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5606 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5605 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5604 = (1'h0);
  reg [(4'ha):(1'h0)] reg5603 = (1'h0);
  reg [(5'h10):(1'h0)] reg5602 = (1'h0);
  reg [(4'ha):(1'h0)] forvar5601 = (1'h0);
  reg [(4'h8):(1'h0)] reg5600 = (1'h0);
  reg [(4'h8):(1'h0)] reg5599 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5596 = (1'h0);
  reg [(4'hd):(1'h0)] reg5594 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5593 = (1'h0);
  reg [(2'h3):(1'h0)] reg5590 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5589 = (1'h0);
  reg [(4'hb):(1'h0)] reg5598 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg5597 = (1'h0);
  reg [(4'he):(1'h0)] reg5596 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg5595 = (1'h0);
  reg [(4'hc):(1'h0)] forvar5594 = (1'h0);
  reg [(4'hb):(1'h0)] reg5593 = (1'h0);
  reg [(4'hc):(1'h0)] reg5592 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5591 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar5590 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5589 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5588 = (1'h0);
  reg [(4'h9):(1'h0)] forvar5587 = (1'h0);
  reg [(4'hb):(1'h0)] reg5586 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5585 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5584 = (1'h0);
  reg [(4'h8):(1'h0)] reg5583 = (1'h0);
  reg [(4'ha):(1'h0)] reg5582 = (1'h0);
  reg [(2'h3):(1'h0)] reg5580 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5578 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg5581 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5580 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5579 = (1'h0);
  reg [(3'h4):(1'h0)] reg5578 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5577 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5576 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5575 = (1'h0);
  reg [(4'h9):(1'h0)] reg5574 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5573 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5572 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5571 = (1'h0);
  reg [(2'h3):(1'h0)] reg5570 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar5569 = (1'h0);
  reg [(4'hf):(1'h0)] reg5568 = (1'h0);
  reg [(4'hd):(1'h0)] reg5567 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5566 = (1'h0);
  reg [(3'h5):(1'h0)] reg5565 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar5564 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5563 = (1'h0);
  reg [(3'h7):(1'h0)] reg5562 = (1'h0);
  reg [(4'hc):(1'h0)] reg5561 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5560 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5558 = (1'h0);
  reg [(4'hc):(1'h0)] reg5555 = (1'h0);
  reg [(4'hd):(1'h0)] forvar5552 = (1'h0);
  reg [(2'h2):(1'h0)] reg5559 = (1'h0);
  reg [(3'h7):(1'h0)] reg5558 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5557 = (1'h0);
  reg [(5'h10):(1'h0)] reg5556 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar5555 = (1'h0);
  reg [(3'h7):(1'h0)] reg5554 = (1'h0);
  reg [(4'h9):(1'h0)] reg5553 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5552 = (1'h0);
  reg [(2'h2):(1'h0)] reg5551 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar5549 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5547 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5546 = (1'h0);
  reg [(4'he):(1'h0)] forvar5540 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar5529 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5527 = (1'h0);
  reg [(3'h4):(1'h0)] forvar5526 = (1'h0);
  reg [(4'hf):(1'h0)] forvar5521 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5519 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5518 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar5537 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5538 = (1'h0);
  reg [(4'hb):(1'h0)] reg5536 = (1'h0);
  reg [(4'h9):(1'h0)] reg5550 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5549 = (1'h0);
  reg [(3'h4):(1'h0)] reg5548 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg5547 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5543 = (1'h0);
  reg [(3'h5):(1'h0)] reg5542 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg5546 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5545 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg5544 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5543 = (1'h0);
  reg [(2'h2):(1'h0)] forvar5542 = (1'h0);
  reg [(2'h3):(1'h0)] reg5541 = (1'h0);
  reg [(4'hf):(1'h0)] reg5540 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5539 = (1'h0);
  reg [(2'h2):(1'h0)] reg5538 = (1'h0);
  reg [(4'h9):(1'h0)] reg5537 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar5536 = (1'h0);
  reg [(2'h3):(1'h0)] reg5535 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5534 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg5533 = (1'h0);
  reg [(2'h3):(1'h0)] reg5532 = (1'h0);
  reg [(4'ha):(1'h0)] reg5531 = (1'h0);
  reg [(4'h8):(1'h0)] reg5530 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg5529 = (1'h0);
  reg [(3'h7):(1'h0)] reg5528 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar5527 = (1'h0);
  reg [(3'h7):(1'h0)] reg5526 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5525 = (1'h0);
  reg [(3'h5):(1'h0)] reg5524 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5523 = (1'h0);
  reg [(4'hc):(1'h0)] reg5522 = (1'h0);
  reg signed [(4'he):(1'h0)] reg5521 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg5520 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5519 = (1'h0);
  reg [(2'h3):(1'h0)] forvar5518 = (1'h0);
  reg [(5'h10):(1'h0)] forvar5517 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg5516 = (1'h0);
  assign y = {reg6014,
                 reg6013,
                 reg6002,
                 reg6012,
                 forvar6011,
                 reg6010,
                 reg6009,
                 reg6008,
                 reg6007,
                 reg6006,
                 reg6005,
                 reg6004,
                 reg6003,
                 forvar6002,
                 forvar6001,
                 forvar6000,
                 reg5999,
                 reg5998,
                 forvar5997,
                 reg5996,
                 forvar5995,
                 reg5994,
                 reg5993,
                 forvar5992,
                 reg5991,
                 reg5990,
                 forvar5989,
                 reg5989,
                 reg5988,
                 reg5987,
                 reg5986,
                 reg5985,
                 reg5984,
                 reg5983,
                 reg5982,
                 forvar5981,
                 forvar5980,
                 reg5979,
                 reg5978,
                 reg5977,
                 reg5976,
                 forvar5975,
                 reg5974,
                 reg5973,
                 reg5972,
                 forvar5971,
                 reg5970,
                 forvar5969,
                 forvar5968,
                 reg5967,
                 reg5966,
                 reg5965,
                 forvar5964,
                 reg5963,
                 reg5962,
                 forvar5961,
                 reg5960,
                 reg5959,
                 reg5958,
                 forvar5957,
                 reg5956,
                 reg5955,
                 reg5954,
                 reg5953,
                 forvar5952,
                 reg5951,
                 forvar5950,
                 reg5949,
                 reg5948,
                 reg5947,
                 forvar5946,
                 reg5945,
                 reg5944,
                 reg5943,
                 forvar5942,
                 reg5941,
                 reg5940,
                 reg5939,
                 forvar5938,
                 reg5937,
                 reg5936,
                 reg5935,
                 forvar5934,
                 reg5933,
                 reg5932,
                 reg5931,
                 reg5930,
                 forvar5929,
                 forvar5928,
                 forvar5927,
                 reg5926,
                 reg5919,
                 forvar5918,
                 reg5925,
                 forvar5924,
                 reg5923,
                 reg5922,
                 reg5921,
                 reg5920,
                 forvar5919,
                 reg5918,
                 reg5917,
                 forvar5916,
                 reg5915,
                 forvar5914,
                 reg5913,
                 reg5912,
                 reg5911,
                 reg5910,
                 forvar5909,
                 reg5908,
                 reg5907,
                 reg5906,
                 reg5905,
                 reg5904,
                 forvar5903,
                 forvar5902,
                 reg5901,
                 reg5900,
                 reg5899,
                 forvar5898,
                 reg5897,
                 reg5896,
                 reg5895,
                 reg5894,
                 reg5893,
                 forvar5892,
                 forvar5891,
                 forvar5890,
                 reg5889,
                 reg5888,
                 reg5887,
                 forvar5886,
                 reg5885,
                 reg5884,
                 reg5883,
                 reg5882,
                 forvar5881,
                 reg5880,
                 reg5879,
                 reg5878,
                 forvar5875,
                 forvar5870,
                 reg5877,
                 reg5876,
                 reg5875,
                 reg5874,
                 reg5873,
                 reg5872,
                 reg5871,
                 reg5870,
                 reg5869,
                 forvar5868,
                 forvar5867,
                 wire5866,
                 wire5865,
                 wire5864,
                 wire5863,
                 reg5832,
                 forvar5830,
                 forvar5828,
                 reg5827,
                 forvar5819,
                 forvar5818,
                 reg5862,
                 reg5848,
                 forvar5847,
                 forvar5846,
                 reg5843,
                 reg5840,
                 reg5839,
                 reg5861,
                 reg5860,
                 reg5859,
                 reg5858,
                 forvar5857,
                 reg5856,
                 reg5855,
                 forvar5854,
                 forvar5853,
                 reg5852,
                 reg5851,
                 reg5850,
                 reg5849,
                 forvar5848,
                 reg5847,
                 reg5846,
                 reg5845,
                 reg5844,
                 forvar5843,
                 reg5842,
                 reg5841,
                 forvar5840,
                 forvar5839,
                 reg5838,
                 reg5837,
                 forvar5836,
                 forvar5820,
                 reg5826,
                 reg5823,
                 forvar5829,
                 reg5835,
                 reg5834,
                 reg5833,
                 forvar5832,
                 reg5831,
                 reg5830,
                 reg5829,
                 reg5828,
                 forvar5827,
                 forvar5826,
                 forvar5817,
                 reg5825,
                 reg5824,
                 forvar5823,
                 reg5822,
                 reg5821,
                 reg5820,
                 reg5819,
                 reg5818,
                 reg5817,
                 reg5816,
                 reg5815,
                 reg5814,
                 reg5813,
                 reg5812,
                 reg5811,
                 reg5810,
                 reg5809,
                 reg5808,
                 reg5807,
                 reg5806,
                 forvar5805,
                 forvar5804,
                 reg5803,
                 reg5802,
                 forvar5801,
                 reg5800,
                 forvar5799,
                 reg5798,
                 reg5797,
                 reg5796,
                 reg5795,
                 reg5794,
                 reg5793,
                 reg5792,
                 forvar5791,
                 forvar5790,
                 forvar5789,
                 reg5788,
                 reg5787,
                 reg5786,
                 forvar5785,
                 reg5784,
                 reg5783,
                 reg5782,
                 reg5781,
                 forvar5780,
                 reg5779,
                 reg5778,
                 forvar5777,
                 reg5776,
                 reg5775,
                 reg5774,
                 forvar5773,
                 forvar5772,
                 forvar5771,
                 reg5770,
                 reg5769,
                 forvar5768,
                 reg5767,
                 reg5766,
                 reg5765,
                 reg5764,
                 forvar5763,
                 forvar5762,
                 forvar5761,
                 forvar5741,
                 reg5746,
                 reg5739,
                 reg5725,
                 forvar5721,
                 reg5730,
                 reg5738,
                 forvar5734,
                 reg5733,
                 forvar5726,
                 forvar5720,
                 forvar5718,
                 reg5716,
                 reg5760,
                 reg5759,
                 reg5758,
                 reg5757,
                 forvar5756,
                 reg5752,
                 forvar5751,
                 reg5756,
                 reg5755,
                 reg5754,
                 reg5753,
                 forvar5752,
                 reg5751,
                 reg5750,
                 reg5749,
                 reg5748,
                 reg5747,
                 forvar5746,
                 reg5745,
                 reg5744,
                 reg5743,
                 reg5742,
                 reg5741,
                 reg5740,
                 forvar5739,
                 forvar5738,
                 reg5737,
                 reg5736,
                 reg5735,
                 reg5734,
                 forvar5733,
                 reg5732,
                 reg5731,
                 forvar5730,
                 reg5729,
                 reg5728,
                 reg5727,
                 reg5726,
                 forvar5725,
                 reg5724,
                 reg5723,
                 reg5722,
                 reg5721,
                 reg5720,
                 reg5719,
                 reg5718,
                 forvar5717,
                 reg5717,
                 forvar5716,
                 reg5715,
                 reg5714,
                 reg5713,
                 reg5712,
                 forvar5709,
                 forvar5703,
                 forvar5700,
                 forvar5695,
                 forvar5687,
                 forvar5683,
                 forvar5679,
                 reg5670,
                 forvar5669,
                 reg5668,
                 forvar5658,
                 forvar5655,
                 forvar5650,
                 reg5646,
                 reg5652,
                 reg5647,
                 reg5645,
                 reg5711,
                 reg5699,
                 reg5694,
                 reg5710,
                 reg5709,
                 reg5708,
                 reg5707,
                 reg5706,
                 reg5705,
                 forvar5704,
                 reg5703,
                 reg5702,
                 reg5701,
                 reg5700,
                 forvar5699,
                 reg5698,
                 reg5697,
                 reg5696,
                 reg5695,
                 forvar5694,
                 reg5693,
                 forvar5692,
                 reg5691,
                 reg5690,
                 reg5686,
                 forvar5684,
                 forvar5681,
                 forvar5680,
                 forvar5677,
                 reg5675,
                 forvar5673,
                 reg5671,
                 reg5689,
                 reg5688,
                 reg5687,
                 forvar5686,
                 reg5685,
                 reg5684,
                 reg5683,
                 reg5682,
                 reg5681,
                 reg5680,
                 reg5679,
                 reg5678,
                 reg5677,
                 reg5676,
                 forvar5675,
                 reg5674,
                 reg5673,
                 reg5672,
                 forvar5671,
                 forvar5670,
                 forvar5663,
                 reg5662,
                 reg5669,
                 forvar5668,
                 reg5667,
                 reg5666,
                 forvar5665,
                 reg5664,
                 reg5663,
                 forvar5662,
                 reg5661,
                 reg5660,
                 reg5659,
                 reg5658,
                 forvar5657,
                 reg5656,
                 reg5655,
                 reg5654,
                 reg5653,
                 forvar5652,
                 reg5651,
                 reg5650,
                 reg5649,
                 reg5648,
                 forvar5647,
                 forvar5646,
                 forvar5645,
                 reg5644,
                 wire5643,
                 wire5642,
                 wire5641,
                 reg5640,
                 reg5639,
                 reg5638,
                 reg5637,
                 forvar5636,
                 reg5635,
                 reg5634,
                 reg5633,
                 reg5632,
                 forvar5631,
                 reg5630,
                 forvar5629,
                 forvar5628,
                 forvar5627,
                 reg5626,
                 reg5625,
                 reg5624,
                 reg5623,
                 reg5622,
                 reg5621,
                 forvar5620,
                 reg5619,
                 forvar5618,
                 reg5617,
                 reg5616,
                 reg5615,
                 reg5614,
                 forvar5613,
                 reg5612,
                 forvar5611,
                 forvar5610,
                 reg5609,
                 reg5608,
                 reg5607,
                 reg5606,
                 forvar5605,
                 reg5604,
                 reg5603,
                 reg5602,
                 forvar5601,
                 reg5600,
                 reg5599,
                 forvar5596,
                 reg5594,
                 forvar5593,
                 reg5590,
                 forvar5589,
                 reg5598,
                 reg5597,
                 reg5596,
                 reg5595,
                 forvar5594,
                 reg5593,
                 reg5592,
                 reg5591,
                 forvar5590,
                 reg5589,
                 forvar5588,
                 forvar5587,
                 reg5586,
                 reg5585,
                 reg5584,
                 reg5583,
                 reg5582,
                 reg5580,
                 forvar5578,
                 reg5581,
                 forvar5580,
                 reg5579,
                 reg5578,
                 reg5577,
                 reg5576,
                 forvar5575,
                 reg5574,
                 forvar5573,
                 reg5572,
                 reg5571,
                 reg5570,
                 forvar5569,
                 reg5568,
                 reg5567,
                 reg5566,
                 reg5565,
                 forvar5564,
                 reg5563,
                 reg5562,
                 reg5561,
                 reg5560,
                 forvar5558,
                 reg5555,
                 forvar5552,
                 reg5559,
                 reg5558,
                 reg5557,
                 reg5556,
                 forvar5555,
                 reg5554,
                 reg5553,
                 reg5552,
                 reg5551,
                 forvar5549,
                 forvar5547,
                 forvar5546,
                 forvar5540,
                 forvar5529,
                 reg5527,
                 forvar5526,
                 forvar5521,
                 reg5519,
                 reg5518,
                 forvar5537,
                 forvar5538,
                 reg5536,
                 reg5550,
                 reg5549,
                 reg5548,
                 reg5547,
                 forvar5543,
                 reg5542,
                 reg5546,
                 reg5545,
                 reg5544,
                 reg5543,
                 forvar5542,
                 reg5541,
                 reg5540,
                 reg5539,
                 reg5538,
                 reg5537,
                 forvar5536,
                 reg5535,
                 reg5534,
                 reg5533,
                 reg5532,
                 reg5531,
                 reg5530,
                 reg5529,
                 reg5528,
                 forvar5527,
                 reg5526,
                 reg5525,
                 reg5524,
                 reg5523,
                 reg5522,
                 reg5521,
                 reg5520,
                 forvar5519,
                 forvar5518,
                 forvar5517,
                 reg5516,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((^($unsigned((wire5514 ? (8'ha1) : wire5514)) ?
          $signed($unsigned(wire5513)) : ((wire5513 ? wire5513 : wire5515) ?
              $unsigned(wire5515) : (wire5513 ? wire5513 : wire5515)))))
        begin
          reg5516 <= ($unsigned($signed($unsigned(wire5514))) ?
              (8'h9d) : {((8'h9d) ? $signed((8'ha1)) : $signed(wire5513))});
          for (forvar5517 = (1'h0); (forvar5517 < (1'h1)); forvar5517 = (forvar5517 + (1'h1)))
            begin
              for (forvar5518 = (1'h0); (forvar5518 < (1'h0)); forvar5518 = (forvar5518 + (1'h1)))
                begin
                  for (forvar5519 = (1'h0); (forvar5519 < (2'h3)); forvar5519 = (forvar5519 + (1'h1)))
                    begin
                      reg5520 <= (!wire5512);
                      reg5521 <= wire5513[(4'h8):(2'h3)];
                      reg5522 <= wire5512[(1'h0):(1'h0)];
                    end
                end
              if ($signed((^$signed((wire5515 <= (8'ha9))))))
                begin
                  reg5523 <= ($unsigned((((8'ha6) ? reg5521 : forvar5518) ?
                          forvar5517[(2'h3):(1'h0)] : (-(8'ha4)))) ?
                      (8'hae) : $signed((wire5512 <= {(8'hb4)})));
                end
              else
                begin
                  if (wire5513[(2'h2):(2'h2)])
                    begin
                      reg5523 <= (^(wire5514 ?
                          {(forvar5518 ^ wire5512)} : (reg5520 & reg5522)));
                    end
                  else
                    begin
                      reg5523 <= (($signed((~^wire5513)) ?
                              wire5513 : (^wire5514)) ?
                          (^~$signed($signed(forvar5518))) : wire5514);
                      reg5524 <= ($signed($signed((wire5515 ?
                          (8'hba) : forvar5518))) << (((reg5521 ~^ reg5520) ~^ {reg5516}) ^ wire5513));
                      reg5525 <= (((^(reg5524 >= reg5516)) + (8'hab)) ?
                          $signed($unsigned((^~reg5523))) : (|(^reg5522)));
                    end
                  reg5526 <= $unsigned($unsigned($signed((!wire5513))));
                  for (forvar5527 = (1'h0); (forvar5527 < (1'h0)); forvar5527 = (forvar5527 + (1'h1)))
                    begin
                      reg5528 <= ((~(-(~&forvar5527))) == wire5515);
                    end
                  if ($unsigned(wire5514))
                    begin
                      reg5529 <= (((~|$signed(forvar5519)) ?
                              $unsigned((-(8'h9d))) : (reg5525 || (wire5513 | wire5515))) ?
                          ($signed((reg5526 ?
                              forvar5518 : wire5515)) < (~|(+wire5512))) : (8'ha2));
                      reg5530 <= ((|$unsigned($signed(reg5526))) ?
                          forvar5519[(2'h2):(1'h0)] : reg5524[(2'h2):(1'h1)]);
                      reg5531 <= (reg5520[(1'h0):(1'h0)] ?
                          (8'ha1) : ($unsigned(wire5512[(1'h0):(1'h0)]) ?
                              forvar5517 : (~&forvar5517[(2'h3):(2'h3)])));
                      reg5532 <= $unsigned((((reg5528 ? reg5516 : reg5526) ?
                          ((8'ha5) ?
                              reg5530 : reg5531) : wire5515[(3'h7):(3'h5)]) || reg5526));
                    end
                  else
                    begin
                      reg5529 <= ($signed((8'hb0)) != wire5514[(1'h1):(1'h0)]);
                      reg5530 <= ($signed($signed({wire5512})) ?
                          $unsigned($signed((^~reg5530))) : $signed(({reg5522} ~^ $signed(forvar5517))));
                      reg5531 <= (!wire5515);
                      reg5532 <= $signed($unsigned(($unsigned(reg5525) ^~ {wire5513})));
                    end
                end
              reg5533 <= ($signed(forvar5518[(1'h0):(1'h0)]) ^ reg5530[(1'h0):(1'h0)]);
              reg5534 <= ($signed($unsigned((8'h9d))) ?
                  (~&$unsigned((reg5531 ?
                      (8'hb0) : wire5514))) : {$signed($unsigned((8'ha9)))});
            end
          if ((~wire5514[(2'h2):(1'h1)]))
            begin
              reg5535 <= {forvar5517[(3'h5):(2'h3)]};
              for (forvar5536 = (1'h0); (forvar5536 < (1'h0)); forvar5536 = (forvar5536 + (1'h1)))
                begin
                  reg5537 <= ((($signed(reg5522) >= (reg5533 < reg5526)) << $signed(reg5532)) > ($signed((reg5520 ?
                          wire5513 : wire5515)) ?
                      {(^~reg5528)} : $signed($signed(reg5525))));
                  if ($unsigned($signed({{wire5513}})))
                    begin
                      reg5538 <= ($signed({(reg5516 ^~ reg5534)}) <<< $unsigned((8'hb0)));
                      reg5539 <= ((8'hb0) ?
                          $signed((reg5521 - reg5530[(1'h0):(1'h0)])) : $signed(((reg5537 ?
                                  reg5529 : (8'h9d)) ?
                              $unsigned(reg5521) : (~forvar5519))));
                      reg5540 <= ((8'hb1) ~^ wire5512);
                      reg5541 <= reg5529;
                    end
                  else
                    begin
                      reg5538 <= $signed($signed(($unsigned((8'ha0)) | reg5528)));
                      reg5539 <= {({((8'hb0) ? wire5515 : reg5537)} ?
                              ($signed((8'ha5)) << forvar5517) : $signed((|forvar5517)))};
                      reg5540 <= wire5512;
                    end
                end
              if ((((+(reg5522 ? reg5529 : wire5514)) ?
                      (|$unsigned((8'hb5))) : ((~&reg5533) ?
                          {reg5534} : reg5523[(1'h1):(1'h0)])) ?
                  (-((8'ha4) + reg5516)) : reg5522[(2'h3):(1'h1)]))
                begin
                  for (forvar5542 = (1'h0); (forvar5542 < (2'h2)); forvar5542 = (forvar5542 + (1'h1)))
                    begin
                      reg5543 <= wire5512;
                      reg5544 <= reg5540[(4'h9):(3'h7)];
                      reg5545 <= (8'ha8);
                      reg5546 <= reg5525[(4'hd):(1'h1)];
                    end
                end
              else
                begin
                  reg5542 <= reg5543;
                  for (forvar5543 = (1'h0); (forvar5543 < (2'h2)); forvar5543 = (forvar5543 + (1'h1)))
                    begin
                      reg5544 <= ((($signed(forvar5543) ?
                              {reg5539} : (reg5523 >= reg5544)) | $signed((^(8'hb4)))) ?
                          $signed({wire5515}) : {(reg5531[(3'h6):(3'h5)] ~^ (reg5545 ?
                                  reg5534 : (8'ha4)))});
                      reg5545 <= (&$signed(reg5525[(4'h9):(2'h3)]));
                      reg5546 <= ({wire5514} ~^ (&forvar5542[(1'h1):(1'h1)]));
                    end
                  reg5547 <= {(-$unsigned((forvar5536 | reg5521)))};
                  if (($unsigned($unsigned((reg5522 + reg5538))) - {(8'hb9)}))
                    begin
                      reg5548 <= ($signed(reg5546) ?
                          $unsigned($unsigned({wire5513})) : (reg5539 < (8'haf)));
                    end
                  else
                    begin
                      reg5548 <= (^(!forvar5517[(1'h1):(1'h0)]));
                      reg5549 <= (~&$signed(((reg5543 ? (8'ha9) : reg5516) ?
                          $signed(reg5537) : reg5548)));
                      reg5550 <= $signed(reg5544[(2'h3):(1'h0)]);
                    end
                end
            end
          else
            begin
              reg5535 <= ((-reg5537[(1'h1):(1'h1)]) == (&reg5545[(1'h1):(1'h1)]));
              reg5536 <= $unsigned(reg5547[(3'h4):(1'h0)]);
              if (reg5533)
                begin
                  reg5537 <= $signed(forvar5518);
                  for (forvar5538 = (1'h0); (forvar5538 < (2'h2)); forvar5538 = (forvar5538 + (1'h1)))
                    begin
                      reg5539 <= (($unsigned((|reg5520)) | {(reg5549 ?
                                  reg5524 : reg5533)}) ?
                          $signed((reg5523 & $signed(reg5548))) : (^$signed($unsigned(reg5542))));
                      reg5540 <= (~^(($signed((8'hb0)) ?
                              {reg5538} : forvar5536[(4'hc):(1'h1)]) ?
                          forvar5518 : $unsigned((|(8'hb7)))));
                    end
                end
              else
                begin
                  for (forvar5537 = (1'h0); (forvar5537 < (1'h0)); forvar5537 = (forvar5537 + (1'h1)))
                    begin
                      reg5538 <= $unsigned($unsigned(reg5548));
                      reg5539 <= $unsigned((({reg5538} ?
                              (reg5543 ?
                                  reg5523 : reg5531) : $signed(reg5546)) ?
                          ((~^forvar5519) ?
                              (^reg5532) : (reg5548 & (8'ha6))) : ($signed(forvar5538) >>> forvar5542[(1'h0):(1'h0)])));
                      reg5540 <= ((((8'h9f) > (forvar5517 ?
                              reg5523 : reg5532)) && $signed($unsigned((8'ha2)))) ?
                          (&$unsigned((wire5514 ^ reg5549))) : ($signed({reg5546}) & ($signed(reg5549) ?
                              (reg5548 ~^ wire5514) : $unsigned(reg5525))));
                      reg5541 <= wire5513[(3'h7):(2'h2)];
                    end
                  reg5542 <= (!$unsigned(($unsigned(forvar5518) ?
                      (forvar5536 || wire5514) : (forvar5538 <= reg5524))));
                  for (forvar5543 = (1'h0); (forvar5543 < (2'h2)); forvar5543 = (forvar5543 + (1'h1)))
                    begin
                      reg5544 <= $signed($unsigned(reg5528));
                      reg5545 <= (8'ha0);
                      reg5546 <= (~|{reg5520});
                      reg5547 <= $unsigned(((|reg5550) ?
                          {reg5520} : forvar5517[(3'h7):(1'h0)]));
                    end
                end
            end
        end
      else
        begin
          reg5516 <= (-$signed((~^reg5529)));
          for (forvar5517 = (1'h0); (forvar5517 < (2'h3)); forvar5517 = (forvar5517 + (1'h1)))
            begin
              if ($unsigned(reg5525))
                begin
                  if (((8'hb4) ?
                      $signed(forvar5542) : (forvar5519[(3'h5):(3'h5)] ?
                          $signed((8'haf)) : (|forvar5542))))
                    begin
                      reg5518 <= reg5520[(1'h1):(1'h0)];
                      reg5519 <= (forvar5518 > forvar5517[(4'he):(4'ha)]);
                    end
                  else
                    begin
                      reg5518 <= reg5539;
                      reg5519 <= (+reg5544[(1'h1):(1'h0)]);
                      reg5520 <= $signed(reg5521);
                    end
                  for (forvar5521 = (1'h0); (forvar5521 < (2'h3)); forvar5521 = (forvar5521 + (1'h1)))
                    begin
                      reg5522 <= ($unsigned(($signed(reg5524) - (&reg5536))) << forvar5538);
                      reg5523 <= {$unsigned(reg5529[(2'h2):(1'h0)])};
                      reg5524 <= ((^((reg5532 ?
                          reg5541 : (8'ha0)) ^~ (-reg5542))) - {$signed($signed(reg5549))});
                      reg5525 <= $unsigned({(+{reg5524})});
                    end
                  for (forvar5526 = (1'h0); (forvar5526 < (2'h3)); forvar5526 = (forvar5526 + (1'h1)))
                    begin
                      reg5527 <= (~{$unsigned((forvar5521 || reg5544))});
                      reg5528 <= reg5529;
                    end
                end
              else
                begin
                  reg5518 <= {reg5550};
                  for (forvar5519 = (1'h0); (forvar5519 < (1'h0)); forvar5519 = (forvar5519 + (1'h1)))
                    begin
                      reg5520 <= $signed(reg5521);
                      reg5521 <= $unsigned($signed((~^(reg5541 + (8'hac)))));
                      reg5522 <= wire5513;
                      reg5523 <= $unsigned(reg5523[(1'h1):(1'h0)]);
                    end
                end
              if ($unsigned((~&$unsigned(reg5543[(1'h1):(1'h0)]))))
                begin
                  for (forvar5529 = (1'h0); (forvar5529 < (2'h3)); forvar5529 = (forvar5529 + (1'h1)))
                    begin
                      reg5530 <= ($unsigned(({reg5546} != reg5550)) << forvar5536);
                      reg5531 <= reg5546;
                    end
                end
              else
                begin
                  if (reg5549)
                    begin
                      reg5529 <= ((^~($unsigned(reg5535) ?
                          {forvar5543} : (wire5515 ?
                              forvar5526 : reg5516))) * (reg5519[(3'h4):(2'h2)] ?
                          ($unsigned(wire5513) | $signed((8'hae))) : {$signed(reg5519)}));
                    end
                  else
                    begin
                      reg5529 <= $signed($signed((reg5541[(2'h3):(2'h2)] >> (forvar5537 ^~ reg5542))));
                      reg5530 <= (forvar5527 ?
                          $signed($unsigned($signed(reg5532))) : forvar5538);
                      reg5531 <= ((^($signed(reg5519) >> $unsigned((8'hac)))) != $unsigned((^~wire5512[(2'h2):(1'h1)])));
                      reg5532 <= forvar5538;
                    end
                  reg5533 <= (-$unsigned((8'hb5)));
                  if (($unsigned($signed(reg5549)) | (forvar5538[(4'h8):(3'h7)] ?
                      (reg5534 ?
                          $unsigned(reg5537) : (|(8'ha9))) : wire5514[(3'h5):(2'h2)])))
                    begin
                      reg5534 <= reg5540[(3'h5):(2'h3)];
                      reg5535 <= {{((reg5532 ? (8'hac) : reg5547) ?
                                  (8'hb5) : forvar5527)}};
                      reg5536 <= (8'ha6);
                    end
                  else
                    begin
                      reg5534 <= $unsigned($unsigned($signed({reg5537})));
                      reg5535 <= reg5530[(2'h2):(1'h0)];
                      reg5536 <= (8'h9e);
                      reg5537 <= reg5533[(2'h2):(1'h0)];
                    end
                  if ($unsigned($unsigned($unsigned($unsigned((8'ha6))))))
                    begin
                      reg5538 <= reg5519[(4'ha):(2'h3)];
                      reg5539 <= $unsigned((~(~$signed(forvar5517))));
                    end
                  else
                    begin
                      reg5538 <= $unsigned(reg5546[(4'hf):(4'h9)]);
                    end
                end
              for (forvar5540 = (1'h0); (forvar5540 < (1'h1)); forvar5540 = (forvar5540 + (1'h1)))
                begin
                  if ($signed($unsigned($unsigned((~forvar5538)))))
                    begin
                      reg5541 <= reg5528;
                      reg5542 <= $unsigned((reg5520[(4'hb):(4'h9)] * $signed((reg5522 ~^ reg5540))));
                      reg5543 <= (forvar5536 ~^ ($signed((reg5518 <<< forvar5537)) <<< reg5523[(4'ha):(4'h9)]));
                      reg5544 <= $unsigned((reg5549 && $unsigned($signed((8'ha1)))));
                    end
                  else
                    begin
                      reg5541 <= reg5544[(2'h3):(1'h1)];
                      reg5542 <= ($unsigned(forvar5542[(1'h0):(1'h0)]) ?
                          reg5516[(1'h1):(1'h0)] : (((wire5515 ?
                              forvar5518 : reg5539) != (reg5529 ?
                              forvar5538 : forvar5538)) <<< (~^wire5515)));
                      reg5543 <= (8'hba);
                      reg5544 <= $signed($signed($unsigned({wire5515})));
                    end
                  reg5545 <= (reg5523 > {((reg5538 ?
                          reg5541 : reg5538) >= $signed(forvar5527))});
                end
              for (forvar5546 = (1'h0); (forvar5546 < (2'h3)); forvar5546 = (forvar5546 + (1'h1)))
                begin
                  for (forvar5547 = (1'h0); (forvar5547 < (1'h1)); forvar5547 = (forvar5547 + (1'h1)))
                    begin
                      reg5548 <= reg5540[(4'h9):(2'h2)];
                    end
                end
            end
          if ({({((8'hb9) + forvar5529)} ?
                  $unsigned(((8'ha0) ? forvar5518 : reg5546)) : ({(8'ha3)} ?
                      (-(8'hb4)) : (^reg5541)))})
            begin
              for (forvar5549 = (1'h0); (forvar5549 < (1'h1)); forvar5549 = (forvar5549 + (1'h1)))
                begin
                  reg5550 <= forvar5527;
                  if ((&$signed((&forvar5540))))
                    begin
                      reg5551 <= wire5512[(3'h6):(2'h3)];
                      reg5552 <= $signed((8'h9d));
                      reg5553 <= (&forvar5517);
                      reg5554 <= forvar5526;
                    end
                  else
                    begin
                      reg5551 <= (8'ha0);
                      reg5552 <= forvar5526[(1'h0):(1'h0)];
                    end
                  for (forvar5555 = (1'h0); (forvar5555 < (1'h1)); forvar5555 = (forvar5555 + (1'h1)))
                    begin
                      reg5556 <= (^reg5523);
                      reg5557 <= ($unsigned(forvar5549) * reg5553);
                      reg5558 <= reg5549;
                    end
                end
              reg5559 <= (~&reg5521[(3'h6):(3'h5)]);
            end
          else
            begin
              if (reg5537[(1'h0):(1'h0)])
                begin
                  if (($signed($signed(reg5533[(3'h6):(3'h6)])) ?
                      reg5519 : forvar5546[(5'h10):(4'hf)]))
                    begin
                      reg5549 <= wire5515[(3'h4):(2'h2)];
                      reg5550 <= (~&$signed((8'ha4)));
                    end
                  else
                    begin
                      reg5549 <= $unsigned({{(reg5525 ^~ (8'hb6))}});
                      reg5550 <= {(^(((8'ha6) <= reg5559) ?
                              forvar5540 : (reg5544 < forvar5542)))};
                      reg5551 <= $unsigned(($signed((^(8'ha6))) ?
                          (reg5522 ?
                              (reg5528 ?
                                  reg5516 : forvar5521) : forvar5536[(4'hd):(4'ha)]) : reg5528));
                    end
                  for (forvar5552 = (1'h0); (forvar5552 < (2'h2)); forvar5552 = (forvar5552 + (1'h1)))
                    begin
                      reg5553 <= $unsigned(reg5549);
                      reg5554 <= forvar5546;
                      reg5555 <= ((~|{{reg5522}}) & {(8'ha7)});
                      reg5556 <= $signed(reg5555[(4'h9):(3'h5)]);
                    end
                end
              else
                begin
                  reg5549 <= $unsigned(($signed(((8'hb9) ?
                      reg5552 : reg5529)) >>> (8'hb7)));
                end
              reg5557 <= forvar5521[(3'h6):(2'h2)];
              if (reg5548[(1'h1):(1'h1)])
                begin
                  for (forvar5558 = (1'h0); (forvar5558 < (2'h3)); forvar5558 = (forvar5558 + (1'h1)))
                    begin
                      reg5559 <= {forvar5543[(1'h1):(1'h1)]};
                      reg5560 <= ((~&{((8'hae) << forvar5537)}) == reg5527[(4'he):(3'h7)]);
                    end
                  if ((wire5512 >= $unsigned((+reg5549))))
                    begin
                      reg5561 <= (~^$unsigned(reg5522[(4'hc):(3'h4)]));
                      reg5562 <= ($signed(reg5527[(4'ha):(1'h0)]) ?
                          reg5560[(1'h1):(1'h1)] : forvar5558);
                      reg5563 <= (8'ha4);
                    end
                  else
                    begin
                      reg5561 <= $unsigned(({((8'hb6) ?
                              reg5534 : reg5548)} ^ (8'hb9)));
                      reg5562 <= $unsigned(($signed($signed(reg5561)) || $unsigned(forvar5543[(2'h2):(2'h2)])));
                    end
                end
              else
                begin
                  if (((~|(((8'hb0) ? forvar5538 : forvar5540) ?
                      $signed(forvar5542) : $signed(reg5556))) * (((~(8'ha2)) ?
                      (reg5527 - reg5550) : wire5512) || {reg5559})))
                    begin
                      reg5558 <= $unsigned($signed(reg5527[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg5558 <= (!(8'ha5));
                      reg5559 <= reg5556[(3'h4):(1'h1)];
                    end
                end
              for (forvar5564 = (1'h0); (forvar5564 < (2'h3)); forvar5564 = (forvar5564 + (1'h1)))
                begin
                  reg5565 <= {$signed($unsigned((+reg5544)))};
                  if (reg5525[(4'h8):(4'h8)])
                    begin
                      reg5566 <= reg5540[(4'h9):(4'h8)];
                      reg5567 <= (-(+(~(reg5521 ? (8'haf) : reg5559))));
                      reg5568 <= ({((forvar5546 ?
                                  reg5548 : reg5535) - (reg5565 ?
                                  reg5535 : (8'hb9)))} ?
                          (~|((reg5541 ?
                              reg5536 : reg5562) && (~forvar5540))) : forvar5542[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg5566 <= $unsigned(forvar5527[(2'h3):(2'h2)]);
                      reg5567 <= reg5555;
                    end
                  for (forvar5569 = (1'h0); (forvar5569 < (2'h2)); forvar5569 = (forvar5569 + (1'h1)))
                    begin
                      reg5570 <= $signed(($signed(reg5537) ?
                          reg5533 : ((~^forvar5546) ?
                              $unsigned(reg5552) : (wire5515 <<< reg5561))));
                      reg5571 <= (&({(8'hb7)} ?
                          reg5568[(1'h1):(1'h0)] : $signed($unsigned(reg5567))));
                    end
                  reg5572 <= reg5527[(2'h3):(1'h0)];
                end
            end
          for (forvar5573 = (1'h0); (forvar5573 < (1'h0)); forvar5573 = (forvar5573 + (1'h1)))
            begin
              reg5574 <= ((reg5519 << $signed({reg5535})) ?
                  $unsigned($unsigned($signed(wire5512))) : ((~&(~|forvar5543)) ?
                      reg5550 : $signed((+forvar5537))));
              if (((~|(~^reg5530[(2'h3):(2'h3)])) ?
                  $unsigned($signed((~reg5534))) : ($unsigned((reg5567 ?
                      reg5558 : reg5562)) || $unsigned((~^(8'hac))))))
                begin
                  for (forvar5575 = (1'h0); (forvar5575 < (2'h2)); forvar5575 = (forvar5575 + (1'h1)))
                    begin
                      reg5576 <= (~&$signed((((8'h9d) << (8'hb8)) ^ (reg5557 >> reg5547))));
                      reg5577 <= (-{$signed(reg5536[(1'h0):(1'h0)])});
                      reg5578 <= ($signed(($signed(forvar5538) <<< (8'hab))) ?
                          (8'hb6) : reg5521);
                    end
                  reg5579 <= ((~((forvar5575 ?
                      reg5519 : reg5521) & reg5577[(2'h2):(1'h1)])) ^~ reg5554);
                  for (forvar5580 = (1'h0); (forvar5580 < (2'h2)); forvar5580 = (forvar5580 + (1'h1)))
                    begin
                      reg5581 <= (|reg5521);
                    end
                end
              else
                begin
                  for (forvar5575 = (1'h0); (forvar5575 < (2'h2)); forvar5575 = (forvar5575 + (1'h1)))
                    begin
                      reg5576 <= (reg5524[(3'h4):(2'h2)] <= $unsigned((8'h9d)));
                      reg5577 <= $unsigned(((+reg5531[(1'h1):(1'h0)]) ?
                          ($unsigned(reg5559) ?
                              $unsigned(reg5577) : (reg5538 ?
                                  reg5541 : forvar5555)) : $signed($unsigned(reg5528))));
                    end
                  for (forvar5578 = (1'h0); (forvar5578 < (1'h0)); forvar5578 = (forvar5578 + (1'h1)))
                    begin
                      reg5579 <= $unsigned((~|(reg5550 ?
                          (reg5537 <= reg5547) : (^~reg5566))));
                      reg5580 <= (({(reg5554 ? reg5539 : reg5565)} ?
                          $unsigned(reg5579) : ((&(8'hb2)) ?
                              reg5534 : (reg5571 ?
                                  (8'ha3) : (8'hb4)))) ^ $signed(($unsigned(forvar5546) ?
                          {reg5556} : $unsigned(forvar5543))));
                      reg5581 <= reg5576[(1'h1):(1'h1)];
                      reg5582 <= $signed(forvar5538);
                    end
                  if (forvar5552)
                    begin
                      reg5583 <= ((reg5548[(2'h2):(1'h0)] ?
                              $signed(reg5523) : {forvar5543[(2'h2):(1'h1)]}) ?
                          reg5578 : reg5562[(2'h3):(2'h3)]);
                      reg5584 <= $unsigned(($unsigned($unsigned(reg5576)) ?
                          reg5582 : $signed($signed(forvar5542))));
                      reg5585 <= $unsigned($unsigned($signed({reg5549})));
                    end
                  else
                    begin
                      reg5583 <= (~&$signed(((~reg5563) || (reg5553 ?
                          forvar5569 : reg5518))));
                      reg5584 <= (forvar5527[(2'h3):(2'h3)] ?
                          reg5538 : ((~&((8'had) ? forvar5569 : reg5532)) ?
                              $signed((reg5556 ?
                                  reg5535 : reg5535)) : reg5535));
                      reg5585 <= {(^$signed((+forvar5518)))};
                      reg5586 <= reg5540;
                    end
                end
            end
        end
      for (forvar5587 = (1'h0); (forvar5587 < (2'h3)); forvar5587 = (forvar5587 + (1'h1)))
        begin
          for (forvar5588 = (1'h0); (forvar5588 < (2'h3)); forvar5588 = (forvar5588 + (1'h1)))
            begin
              if ((~&$signed($signed(((8'ha7) < reg5522)))))
                begin
                  reg5589 <= $unsigned(forvar5555);
                  for (forvar5590 = (1'h0); (forvar5590 < (2'h2)); forvar5590 = (forvar5590 + (1'h1)))
                    begin
                      reg5591 <= reg5536;
                      reg5592 <= $signed(((|forvar5540) ~^ $unsigned(wire5512[(1'h0):(1'h0)])));
                      reg5593 <= $unsigned((~&{$signed(reg5554)}));
                    end
                  for (forvar5594 = (1'h0); (forvar5594 < (1'h0)); forvar5594 = (forvar5594 + (1'h1)))
                    begin
                      reg5595 <= (!wire5513[(3'h5):(3'h5)]);
                      reg5596 <= reg5547;
                      reg5597 <= ((~reg5570) >> ((8'ha0) >>> ($unsigned(forvar5542) || (&reg5543))));
                      reg5598 <= {(~&$unsigned(reg5593[(1'h1):(1'h1)]))};
                    end
                end
              else
                begin
                  for (forvar5589 = (1'h0); (forvar5589 < (2'h3)); forvar5589 = (forvar5589 + (1'h1)))
                    begin
                      reg5590 <= (($signed((-reg5539)) ^~ (^~$signed(reg5534))) ?
                          $unsigned((!(reg5528 <= forvar5543))) : $signed($signed({(8'ha7)})));
                      reg5591 <= $signed($unsigned((^(reg5537 * reg5557))));
                      reg5592 <= reg5578[(2'h3):(1'h0)];
                    end
                  for (forvar5593 = (1'h0); (forvar5593 < (1'h1)); forvar5593 = (forvar5593 + (1'h1)))
                    begin
                      reg5594 <= ({({reg5570} * (reg5545 < reg5555))} || {$signed(((8'hb2) ?
                              reg5519 : reg5550))});
                      reg5595 <= (($signed((reg5543 ^ reg5553)) ?
                          forvar5589 : $signed($signed((8'hb4)))) != (((reg5557 == reg5586) ?
                              (reg5535 > reg5541) : (-reg5558)) ?
                          reg5561 : $signed($unsigned(forvar5526))));
                    end
                  for (forvar5596 = (1'h0); (forvar5596 < (2'h2)); forvar5596 = (forvar5596 + (1'h1)))
                    begin
                      reg5597 <= ((reg5595 || ((^forvar5558) ?
                              {reg5548} : reg5539)) ?
                          (~&reg5524) : (forvar5521 ?
                              $signed(((8'hae) >>> reg5551)) : (forvar5527[(3'h4):(3'h4)] ?
                                  $signed(reg5594) : {reg5535})));
                      reg5598 <= (-((8'ha1) << (|(forvar5593 ?
                          forvar5589 : reg5537))));
                      reg5599 <= $signed({reg5519});
                      reg5600 <= (reg5536 ?
                          (~&reg5563) : (((reg5532 - (8'hb7)) ?
                                  $unsigned(reg5541) : $unsigned(reg5552)) ?
                              $unsigned($unsigned((8'ha9))) : ((forvar5593 << reg5520) ?
                                  forvar5526 : (reg5535 ?
                                      (8'hb4) : forvar5546))));
                    end
                  for (forvar5601 = (1'h0); (forvar5601 < (1'h0)); forvar5601 = (forvar5601 + (1'h1)))
                    begin
                      reg5602 <= (-forvar5526);
                      reg5603 <= (^~(($unsigned((8'h9d)) <<< {reg5562}) ?
                          ((~&reg5594) ?
                              $signed(reg5581) : reg5526) : {(reg5585 ?
                                  reg5516 : reg5531)}));
                      reg5604 <= forvar5546[(3'h5):(1'h0)];
                    end
                end
              for (forvar5605 = (1'h0); (forvar5605 < (1'h1)); forvar5605 = (forvar5605 + (1'h1)))
                begin
                  if ($signed($unsigned({((8'h9f) ? (8'ha0) : forvar5540)})))
                    begin
                      reg5606 <= {(~&(&(reg5555 ? reg5529 : reg5540)))};
                      reg5607 <= $signed(reg5557);
                      reg5608 <= $signed($unsigned(((reg5546 ?
                              forvar5578 : reg5591) ?
                          reg5560 : (reg5577 == reg5571))));
                    end
                  else
                    begin
                      reg5606 <= forvar5589[(1'h0):(1'h0)];
                      reg5607 <= {forvar5589};
                      reg5608 <= (~$unsigned({forvar5601[(2'h3):(2'h2)]}));
                      reg5609 <= forvar5540[(4'hd):(1'h1)];
                    end
                end
            end
          for (forvar5610 = (1'h0); (forvar5610 < (1'h1)); forvar5610 = (forvar5610 + (1'h1)))
            begin
              for (forvar5611 = (1'h0); (forvar5611 < (1'h0)); forvar5611 = (forvar5611 + (1'h1)))
                begin
                  reg5612 <= (^($unsigned(forvar5521[(4'hd):(3'h7)]) >>> $signed(reg5516)));
                  for (forvar5613 = (1'h0); (forvar5613 < (2'h3)); forvar5613 = (forvar5613 + (1'h1)))
                    begin
                      reg5614 <= reg5551;
                      reg5615 <= forvar5521[(1'h0):(1'h0)];
                      reg5616 <= $unsigned(wire5514[(3'h5):(3'h5)]);
                      reg5617 <= reg5582;
                    end
                  for (forvar5618 = (1'h0); (forvar5618 < (2'h3)); forvar5618 = (forvar5618 + (1'h1)))
                    begin
                      reg5619 <= (^(^$signed(forvar5537[(1'h0):(1'h0)])));
                    end
                end
              for (forvar5620 = (1'h0); (forvar5620 < (2'h3)); forvar5620 = (forvar5620 + (1'h1)))
                begin
                  if (((^~($signed((8'haa)) ?
                      (8'hb1) : (reg5537 & reg5549))) ^ reg5533))
                    begin
                      reg5621 <= forvar5521;
                      reg5622 <= forvar5580[(4'ha):(1'h1)];
                      reg5623 <= $unsigned(reg5580);
                    end
                  else
                    begin
                      reg5621 <= $unsigned((-((8'ha3) ?
                          {reg5537} : (~reg5530))));
                      reg5622 <= $signed($unsigned(forvar5519[(3'h6):(2'h2)]));
                    end
                  if ($unsigned(reg5555))
                    begin
                      reg5624 <= {$signed(((reg5558 ? reg5520 : reg5556) ?
                              (forvar5578 == reg5529) : $signed(reg5622)))};
                    end
                  else
                    begin
                      reg5624 <= ((^(&(~^forvar5518))) ?
                          $unsigned(($unsigned(reg5558) ?
                              ((8'hb5) ?
                                  reg5592 : reg5616) : (reg5593 >= reg5577))) : $signed((-(wire5513 ?
                              (8'ha5) : (8'hb1)))));
                      reg5625 <= $unsigned(reg5607);
                      reg5626 <= {$signed(($signed((8'ha9)) == $signed(reg5555)))};
                    end
                end
            end
          for (forvar5627 = (1'h0); (forvar5627 < (1'h1)); forvar5627 = (forvar5627 + (1'h1)))
            begin
              for (forvar5628 = (1'h0); (forvar5628 < (2'h2)); forvar5628 = (forvar5628 + (1'h1)))
                begin
                  for (forvar5629 = (1'h0); (forvar5629 < (2'h3)); forvar5629 = (forvar5629 + (1'h1)))
                    begin
                      reg5630 <= ((&reg5550) ?
                          {($signed(reg5580) | (~|reg5534))} : (^~$unsigned(reg5616[(1'h1):(1'h0)])));
                    end
                  for (forvar5631 = (1'h0); (forvar5631 < (2'h2)); forvar5631 = (forvar5631 + (1'h1)))
                    begin
                      reg5632 <= forvar5518[(1'h1):(1'h0)];
                      reg5633 <= $signed(($unsigned(reg5533) ?
                          (8'hb5) : reg5547));
                      reg5634 <= {((~&$unsigned(reg5516)) ?
                              forvar5555[(2'h2):(2'h2)] : $signed(reg5550))};
                    end
                  if ($unsigned(((|(reg5532 * reg5562)) ?
                      ($signed((8'hb9)) ?
                          forvar5631[(2'h3):(2'h2)] : $unsigned(reg5544)) : {{reg5539}})))
                    begin
                      reg5635 <= reg5568[(4'ha):(4'h9)];
                    end
                  else
                    begin
                      reg5635 <= (&((((8'hb5) ?
                          reg5545 : reg5609) - forvar5521[(4'hd):(2'h2)]) >>> ($signed(reg5579) >= $unsigned(forvar5589))));
                    end
                  for (forvar5636 = (1'h0); (forvar5636 < (1'h0)); forvar5636 = (forvar5636 + (1'h1)))
                    begin
                      reg5637 <= (+forvar5589[(2'h3):(1'h0)]);
                      reg5638 <= (!$signed((reg5553[(3'h6):(3'h4)] ?
                          forvar5549[(3'h4):(2'h3)] : $unsigned(reg5544))));
                      reg5639 <= $signed((reg5580 <<< reg5612[(4'hc):(3'h5)]));
                    end
                end
              reg5640 <= {(reg5632[(1'h0):(1'h0)] ?
                      {reg5572[(1'h0):(1'h0)]} : (8'haf))};
            end
        end
    end
  assign wire5641 = {((~^(+reg5630)) ?
                            reg5546[(2'h3):(1'h1)] : (reg5521 ?
                                (~reg5519) : $signed((8'hab))))};
  assign wire5642 = (reg5630[(5'h10):(1'h1)] ?
                        (&reg5635[(2'h3):(1'h1)]) : forvar5555[(1'h0):(1'h0)]);
  assign wire5643 = (&(~$unsigned($unsigned(reg5518))));
  always
    @(posedge clk) begin
      reg5644 <= forvar5573[(3'h5):(2'h3)];
      if ((+(($unsigned((8'ha3)) ~^ reg5556[(3'h7):(3'h5)]) ?
          (reg5540[(4'he):(3'h4)] ? $signed(reg5599) : reg5608) : {(reg5560 ?
                  reg5519 : (8'h9d))})))
        begin
          for (forvar5645 = (1'h0); (forvar5645 < (2'h3)); forvar5645 = (forvar5645 + (1'h1)))
            begin
              for (forvar5646 = (1'h0); (forvar5646 < (2'h2)); forvar5646 = (forvar5646 + (1'h1)))
                begin
                  for (forvar5647 = (1'h0); (forvar5647 < (2'h3)); forvar5647 = (forvar5647 + (1'h1)))
                    begin
                      reg5648 <= forvar5519[(3'h7):(3'h4)];
                      reg5649 <= reg5586;
                      reg5650 <= (reg5533 ? reg5648[(3'h7):(2'h2)] : reg5638);
                      reg5651 <= reg5566;
                    end
                  for (forvar5652 = (1'h0); (forvar5652 < (1'h0)); forvar5652 = (forvar5652 + (1'h1)))
                    begin
                      reg5653 <= $signed(forvar5620);
                      reg5654 <= $unsigned((&(reg5555[(2'h2):(1'h1)] ?
                          forvar5519[(3'h6):(2'h2)] : $signed(reg5614))));
                      reg5655 <= ($unsigned({forvar5611[(2'h2):(1'h1)]}) ?
                          (reg5560[(3'h5):(3'h4)] ?
                              reg5525 : reg5538[(2'h2):(2'h2)]) : ((reg5633 == ((8'ha1) ?
                              reg5558 : forvar5601)) && ($unsigned((8'hb7)) >>> (-(8'hb0)))));
                      reg5656 <= (~&$signed($signed(reg5563[(4'h9):(4'h9)])));
                    end
                  for (forvar5657 = (1'h0); (forvar5657 < (2'h3)); forvar5657 = (forvar5657 + (1'h1)))
                    begin
                      reg5658 <= reg5579[(4'hd):(3'h7)];
                      reg5659 <= $unsigned($signed(reg5557[(1'h1):(1'h1)]));
                      reg5660 <= (~|reg5651);
                    end
                end
              if (reg5560)
                begin
                  reg5661 <= $unsigned($unsigned({(reg5516 >>> reg5556)}));
                  for (forvar5662 = (1'h0); (forvar5662 < (1'h1)); forvar5662 = (forvar5662 + (1'h1)))
                    begin
                      reg5663 <= (reg5608[(2'h2):(1'h1)] >> $unsigned((((8'hb5) & reg5580) ?
                          (~^(8'ha1)) : (&reg5597))));
                      reg5664 <= {forvar5629[(4'ha):(2'h3)]};
                    end
                  for (forvar5665 = (1'h0); (forvar5665 < (1'h0)); forvar5665 = (forvar5665 + (1'h1)))
                    begin
                      reg5666 <= ((reg5574[(1'h0):(1'h0)] ~^ {reg5664}) >= ($signed(reg5606) <<< reg5612[(4'hc):(1'h1)]));
                      reg5667 <= $unsigned({($unsigned((8'ha6)) ?
                              (^~forvar5610) : $unsigned(reg5530))});
                    end
                  for (forvar5668 = (1'h0); (forvar5668 < (1'h1)); forvar5668 = (forvar5668 + (1'h1)))
                    begin
                      reg5669 <= reg5658;
                    end
                end
              else
                begin
                  if (reg5574)
                    begin
                      reg5661 <= ((reg5639 == reg5544[(1'h1):(1'h1)]) >>> $signed($signed($signed((8'hb2)))));
                      reg5662 <= ((|(~|$signed(reg5546))) >= (8'ha0));
                    end
                  else
                    begin
                      reg5661 <= reg5530[(3'h7):(2'h2)];
                      reg5662 <= reg5589;
                    end
                  for (forvar5663 = (1'h0); (forvar5663 < (2'h3)); forvar5663 = (forvar5663 + (1'h1)))
                    begin
                      reg5664 <= (|$unsigned(reg5639[(1'h1):(1'h1)]));
                    end
                end
            end
          if ($signed(reg5664))
            begin
              for (forvar5670 = (1'h0); (forvar5670 < (1'h0)); forvar5670 = (forvar5670 + (1'h1)))
                begin
                  for (forvar5671 = (1'h0); (forvar5671 < (1'h0)); forvar5671 = (forvar5671 + (1'h1)))
                    begin
                      reg5672 <= $signed(($signed($signed((8'hb9))) == (|$unsigned(forvar5657))));
                      reg5673 <= (reg5622 | ({$unsigned(reg5614)} ?
                          reg5630[(4'he):(2'h2)] : ((+reg5632) ?
                              (&(8'haf)) : (~^reg5653))));
                      reg5674 <= $signed({{(reg5669 << reg5519)}});
                    end
                end
              for (forvar5675 = (1'h0); (forvar5675 < (2'h3)); forvar5675 = (forvar5675 + (1'h1)))
                begin
                  reg5676 <= ((~^($unsigned(forvar5587) >= (reg5594 ?
                      reg5549 : forvar5588))) ^ $unsigned(reg5623[(4'hb):(4'h8)]));
                  if ((~|(forvar5542[(2'h2):(2'h2)] ?
                      (~&{reg5608}) : reg5656[(2'h3):(1'h1)])))
                    begin
                      reg5677 <= (($unsigned((~(8'h9e))) ?
                          reg5617 : forvar5611) <<< (~^{$unsigned(forvar5578)}));
                    end
                  else
                    begin
                      reg5677 <= (|(+forvar5538));
                    end
                end
              if ($unsigned(reg5650[(4'h8):(3'h5)]))
                begin
                  reg5678 <= forvar5671[(3'h5):(1'h1)];
                end
              else
                begin
                  if ($signed(reg5580[(1'h1):(1'h0)]))
                    begin
                      reg5678 <= $unsigned((~&(!$signed(forvar5587))));
                      reg5679 <= (reg5677 ~^ ((^~{forvar5662}) ?
                          $signed((~|(8'ha2))) : $signed((forvar5594 ?
                              reg5661 : forvar5596))));
                      reg5680 <= reg5600[(4'h8):(1'h0)];
                    end
                  else
                    begin
                      reg5678 <= {((+{reg5672}) | wire5512[(1'h1):(1'h0)])};
                      reg5679 <= reg5634[(3'h7):(1'h0)];
                      reg5680 <= forvar5610[(4'ha):(2'h2)];
                    end
                  reg5681 <= reg5559[(1'h1):(1'h1)];
                  if (forvar5546)
                    begin
                      reg5682 <= ((|((^reg5658) ?
                          $unsigned(reg5536) : (forvar5663 << forvar5636))) * reg5634[(1'h0):(1'h0)]);
                      reg5683 <= reg5533;
                      reg5684 <= reg5661[(3'h6):(3'h5)];
                      reg5685 <= (reg5522[(2'h3):(1'h1)] ?
                          (forvar5652[(4'he):(4'hc)] ?
                              reg5654[(4'h9):(1'h0)] : $unsigned(wire5642)) : (({reg5560} ?
                              (reg5648 ?
                                  (8'h9d) : reg5640) : $signed((8'hb1))) >>> $signed((reg5566 - reg5648))));
                    end
                  else
                    begin
                      reg5682 <= forvar5549;
                      reg5683 <= (reg5566 >= {forvar5663[(1'h0):(1'h0)]});
                      reg5684 <= (8'hb7);
                    end
                  for (forvar5686 = (1'h0); (forvar5686 < (1'h0)); forvar5686 = (forvar5686 + (1'h1)))
                    begin
                      reg5687 <= (8'h9c);
                      reg5688 <= (reg5617 | forvar5546[(1'h0):(1'h0)]);
                      reg5689 <= ({$signed(reg5609[(1'h1):(1'h1)])} ?
                          {forvar5573[(3'h4):(1'h1)]} : $unsigned((reg5661 ?
                              reg5583[(1'h1):(1'h1)] : (reg5558 ?
                                  (8'hb9) : reg5622))));
                    end
                end
            end
          else
            begin
              for (forvar5670 = (1'h0); (forvar5670 < (1'h1)); forvar5670 = (forvar5670 + (1'h1)))
                begin
                  if ($signed(($signed({wire5643}) ?
                      $signed((reg5604 ?
                          forvar5647 : (8'h9d))) : $unsigned($signed(reg5662)))))
                    begin
                      reg5671 <= (8'hab);
                      reg5672 <= $unsigned((reg5633[(4'hb):(3'h4)] ~^ reg5678));
                    end
                  else
                    begin
                      reg5671 <= ((|$signed({(8'hb4)})) ?
                          {(|$signed((8'hb2)))} : $unsigned($signed((!reg5677))));
                      reg5672 <= $signed($signed((+((8'ha9) << reg5609))));
                    end
                end
              if ((forvar5564 ? forvar5605[(2'h2):(2'h2)] : (-reg5664)))
                begin
                  for (forvar5673 = (1'h0); (forvar5673 < (1'h0)); forvar5673 = (forvar5673 + (1'h1)))
                    begin
                      reg5674 <= (forvar5590[(4'ha):(3'h6)] != wire5512);
                      reg5675 <= $signed(reg5571[(1'h1):(1'h1)]);
                      reg5676 <= reg5537;
                    end
                end
              else
                begin
                  if ($unsigned(forvar5517[(4'hf):(2'h2)]))
                    begin
                      reg5673 <= ($signed($unsigned(reg5598)) ?
                          reg5626[(3'h7):(1'h0)] : ((((8'hab) ?
                              reg5556 : reg5689) < (~|forvar5546)) >> (^~forvar5529[(3'h7):(1'h1)])));
                      reg5674 <= reg5576[(3'h4):(1'h0)];
                      reg5675 <= forvar5686;
                      reg5676 <= $signed($signed(reg5673[(2'h2):(1'h1)]));
                    end
                  else
                    begin
                      reg5673 <= $signed(((~^(reg5666 ?
                          forvar5588 : reg5617)) * $unsigned((~forvar5665))));
                      reg5674 <= (reg5602 ?
                          ($unsigned(reg5678) ^~ $unsigned($unsigned(reg5606))) : reg5525[(4'hb):(4'h8)]);
                      reg5675 <= ((~^reg5603) <= $unsigned(($unsigned((8'hb6)) ?
                          $signed(reg5606) : reg5582)));
                      reg5676 <= (^~reg5566[(3'h5):(1'h1)]);
                    end
                  for (forvar5677 = (1'h0); (forvar5677 < (1'h0)); forvar5677 = (forvar5677 + (1'h1)))
                    begin
                      reg5678 <= {forvar5527};
                      reg5679 <= forvar5668;
                    end
                end
              for (forvar5680 = (1'h0); (forvar5680 < (2'h2)); forvar5680 = (forvar5680 + (1'h1)))
                begin
                  for (forvar5681 = (1'h0); (forvar5681 < (2'h2)); forvar5681 = (forvar5681 + (1'h1)))
                    begin
                      reg5682 <= ({reg5614} ? $unsigned(forvar5543) : reg5669);
                      reg5683 <= forvar5573[(4'hd):(3'h4)];
                    end
                  for (forvar5684 = (1'h0); (forvar5684 < (2'h2)); forvar5684 = (forvar5684 + (1'h1)))
                    begin
                      reg5685 <= forvar5521[(3'h4):(3'h4)];
                      reg5686 <= ($unsigned($signed(reg5598)) | reg5623);
                      reg5687 <= forvar5580[(3'h4):(2'h2)];
                    end
                  if (($unsigned((!(~|reg5666))) ?
                      (|forvar5588) : $unsigned(((forvar5537 ?
                          (8'ha5) : reg5568) ^~ (~&reg5662)))))
                    begin
                      reg5688 <= ((~|(8'hb6)) <= reg5538);
                      reg5689 <= reg5654;
                      reg5690 <= reg5667[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg5688 <= reg5538;
                      reg5689 <= reg5572[(1'h0):(1'h0)];
                      reg5690 <= (~&$signed(forvar5610));
                      reg5691 <= ($signed($signed(reg5545[(1'h1):(1'h0)])) | reg5673[(1'h0):(1'h0)]);
                    end
                  for (forvar5692 = (1'h0); (forvar5692 < (2'h2)); forvar5692 = (forvar5692 + (1'h1)))
                    begin
                      reg5693 <= $signed(reg5673[(1'h1):(1'h1)]);
                    end
                end
            end
          if ({$signed({$unsigned(reg5591)})})
            begin
              for (forvar5694 = (1'h0); (forvar5694 < (2'h2)); forvar5694 = (forvar5694 + (1'h1)))
                begin
                  if (((reg5689[(1'h0):(1'h0)] << $signed(((8'hb6) ?
                      forvar5526 : reg5585))) != (-reg5671)))
                    begin
                      reg5695 <= $signed(reg5667[(3'h7):(3'h6)]);
                      reg5696 <= (reg5630[(5'h10):(4'h9)] ?
                          reg5520 : $signed(reg5584));
                      reg5697 <= {$unsigned((~(reg5520 > wire5514)))};
                      reg5698 <= ((reg5528[(3'h6):(3'h4)] <<< (^~(8'hb3))) ?
                          $signed(forvar5594) : {$signed(reg5632[(1'h1):(1'h0)])});
                    end
                  else
                    begin
                      reg5695 <= ((((reg5597 & reg5606) ^~ forvar5646) ^ $unsigned((+forvar5647))) ~^ (~&$unsigned((~^reg5559))));
                      reg5696 <= $signed((($signed((8'h9c)) | (reg5545 || forvar5611)) ?
                          (reg5675 ?
                              (forvar5529 >= forvar5646) : {(8'hb3)}) : {(8'hb9)}));
                      reg5697 <= (~&(forvar5573 ?
                          reg5625[(4'hd):(1'h0)] : ({(8'hae)} ~^ {forvar5681})));
                    end
                end
              for (forvar5699 = (1'h0); (forvar5699 < (1'h1)); forvar5699 = (forvar5699 + (1'h1)))
                begin
                  if (forvar5605)
                    begin
                      reg5700 <= $signed(reg5594);
                      reg5701 <= $signed(reg5570[(2'h3):(2'h3)]);
                      reg5702 <= $unsigned(reg5592);
                      reg5703 <= (forvar5549[(2'h3):(2'h3)] >= {wire5513});
                    end
                  else
                    begin
                      reg5700 <= ((8'hba) && reg5684);
                      reg5701 <= forvar5589[(2'h3):(1'h0)];
                      reg5702 <= (reg5574 ?
                          $unsigned({{forvar5663}}) : ($signed(((8'hb0) >> reg5640)) ?
                              forvar5662[(4'hd):(4'hb)] : (~|((8'hb6) ~^ reg5703))));
                    end
                  for (forvar5704 = (1'h0); (forvar5704 < (1'h0)); forvar5704 = (forvar5704 + (1'h1)))
                    begin
                      reg5705 <= (forvar5543 ?
                          $signed((~|$signed((8'hb1)))) : ($signed((reg5527 >>> reg5622)) - (+$signed(reg5527))));
                    end
                  reg5706 <= $signed(($unsigned((reg5523 ?
                      reg5536 : reg5538)) << $unsigned(forvar5620)));
                  if ({$signed({(8'ha3)})})
                    begin
                      reg5707 <= (reg5677 ?
                          $signed(($unsigned(reg5679) ?
                              reg5695[(5'h10):(2'h2)] : (+reg5686))) : reg5577[(1'h0):(1'h0)]);
                      reg5708 <= reg5696;
                    end
                  else
                    begin
                      reg5707 <= (((8'hb6) == reg5677) ?
                          $signed(reg5686) : ($unsigned({reg5559}) ?
                              ($unsigned(reg5566) && reg5597[(4'hd):(4'hb)]) : (forvar5540 <<< (reg5541 ?
                                  reg5682 : reg5612))));
                      reg5708 <= (~^reg5673);
                      reg5709 <= (forvar5611 + $unsigned(($unsigned(reg5538) ?
                          (8'hb5) : (~|wire5642))));
                      reg5710 <= reg5586;
                    end
                end
            end
          else
            begin
              if ((($unsigned(reg5558) >> reg5608[(1'h1):(1'h0)]) & ((reg5574[(3'h5):(2'h2)] ?
                      reg5644[(3'h4):(2'h2)] : reg5593) ?
                  ((!reg5516) && ((8'hb0) ? reg5560 : reg5536)) : (8'hb2))))
                begin
                  if ((((-reg5648) ?
                          $signed($signed(wire5512)) : $signed({forvar5536})) ?
                      ($signed($unsigned(reg5661)) || forvar5677[(2'h2):(2'h2)]) : (~^({reg5671} ?
                          reg5648 : $unsigned(reg5683)))))
                    begin
                      reg5694 <= reg5708;
                      reg5695 <= reg5530;
                      reg5696 <= (8'ha5);
                      reg5697 <= (^reg5706);
                    end
                  else
                    begin
                      reg5694 <= (((forvar5671 ? $signed(reg5679) : reg5624) ?
                              $unsigned((reg5559 < reg5581)) : $unsigned((|reg5682))) ?
                          reg5664[(3'h4):(2'h2)] : reg5615[(4'h8):(4'h8)]);
                      reg5695 <= forvar5629;
                      reg5696 <= ((((forvar5564 ? (8'hb6) : reg5542) ?
                                  (reg5696 ?
                                      reg5675 : reg5591) : (reg5640 - forvar5665)) ?
                              ((reg5675 * forvar5668) - $unsigned((8'ha3))) : (~^$unsigned(reg5706))) ?
                          (reg5608 < (^(wire5514 ?
                              reg5637 : forvar5589))) : (((reg5531 <= reg5623) ?
                              {reg5542} : ((8'ha1) ?
                                  (8'hb2) : reg5566)) << reg5583[(2'h2):(2'h2)]));
                    end
                  reg5698 <= ($signed(reg5550) | {$signed((^forvar5675))});
                  if ($unsigned($unsigned({(forvar5611 ? (8'hba) : reg5594)})))
                    begin
                      reg5699 <= ((reg5567 ^~ $signed($signed(reg5687))) ?
                          (((&reg5526) ?
                                  (forvar5519 * reg5579) : $unsigned(reg5659)) ?
                              (~^((8'h9c) ^ reg5661)) : forvar5587) : (8'haf));
                    end
                  else
                    begin
                      reg5699 <= forvar5527;
                      reg5700 <= reg5531;
                      reg5701 <= $signed($signed(reg5710));
                    end
                end
              else
                begin
                  if ($signed(((8'had) >= ((+reg5684) < reg5555[(4'ha):(3'h7)]))))
                    begin
                      reg5694 <= reg5708[(1'h1):(1'h0)];
                      reg5695 <= $unsigned(($signed($signed(reg5669)) < $unsigned((+forvar5645))));
                    end
                  else
                    begin
                      reg5694 <= ({((reg5684 ? forvar5521 : forvar5636) ?
                              reg5586[(3'h4):(3'h4)] : $unsigned(forvar5555))} || ($unsigned({forvar5613}) || ($signed(reg5619) ?
                          (|forvar5521) : reg5597)));
                      reg5695 <= (!{$unsigned($unsigned(reg5523))});
                      reg5696 <= (+$signed((|((8'ha6) != (8'ha6)))));
                    end
                end
              reg5702 <= reg5600;
            end
          reg5711 <= ($unsigned(reg5656[(1'h0):(1'h0)]) ^~ ((reg5524 * $unsigned(reg5549)) ?
              reg5545[(4'ha):(3'h4)] : (~|$signed((8'ha2)))));
        end
      else
        begin
          if ($unsigned(reg5625[(3'h4):(3'h4)]))
            begin
              reg5645 <= ($signed($signed((+reg5572))) < reg5516[(1'h1):(1'h1)]);
              for (forvar5646 = (1'h0); (forvar5646 < (2'h3)); forvar5646 = (forvar5646 + (1'h1)))
                begin
                  if (forvar5657[(4'h9):(4'h9)])
                    begin
                      reg5647 <= forvar5552[(1'h1):(1'h1)];
                      reg5648 <= ((8'had) ?
                          ($unsigned((~(8'h9c))) | ((~|(8'hae)) ?
                              ((8'haa) == reg5637) : (forvar5575 ?
                                  reg5649 : (8'h9e)))) : $signed(((reg5560 ?
                              reg5630 : forvar5549) + $unsigned(reg5695))));
                      reg5649 <= (reg5516 ?
                          (^~((reg5663 ? forvar5542 : forvar5587) ?
                              (reg5693 ^~ forvar5552) : reg5638)) : forvar5546[(4'hd):(4'h8)]);
                    end
                  else
                    begin
                      reg5647 <= (&(($signed(reg5612) <= forvar5628[(2'h3):(1'h0)]) >> $signed((reg5683 ?
                          reg5644 : reg5702))));
                    end
                  reg5650 <= reg5654[(4'h8):(2'h2)];
                  if (reg5562)
                    begin
                      reg5651 <= $signed(($signed({reg5521}) ?
                          ((~^reg5625) >>> reg5644) : ($unsigned(forvar5593) >> (!forvar5590))));
                      reg5652 <= {$unsigned(reg5695[(3'h5):(1'h1)])};
                      reg5653 <= $signed(reg5586);
                    end
                  else
                    begin
                      reg5651 <= (~reg5609);
                      reg5652 <= $unsigned(((forvar5647[(1'h0):(1'h0)] ?
                              (&(8'haf)) : ((8'haf) - reg5681)) ?
                          $unsigned($unsigned((8'h9c))) : (reg5675[(2'h2):(1'h0)] ?
                              $unsigned(reg5675) : $signed(reg5554))));
                      reg5653 <= {reg5532[(1'h1):(1'h1)]};
                    end
                end
              reg5654 <= $signed((reg5598 | $signed((!(8'hae)))));
            end
          else
            begin
              if ($unsigned(reg5574[(1'h0):(1'h0)]))
                begin
                  reg5645 <= (((-(~&forvar5575)) ?
                      ($signed((8'ha9)) - $signed(reg5561)) : reg5550) ~^ $unsigned(reg5554));
                  for (forvar5646 = (1'h0); (forvar5646 < (2'h3)); forvar5646 = (forvar5646 + (1'h1)))
                    begin
                      reg5647 <= ($unsigned(reg5648) ?
                          {reg5565} : $signed($unsigned(reg5559[(1'h0):(1'h0)])));
                      reg5648 <= reg5549[(1'h1):(1'h0)];
                      reg5649 <= $unsigned(((8'hac) == reg5691[(3'h4):(1'h1)]));
                    end
                end
              else
                begin
                  if (((~&$signed((&(8'ha5)))) ~^ $signed((((8'hb9) ?
                          reg5681 : forvar5618) ?
                      reg5660[(1'h1):(1'h0)] : reg5538[(2'h2):(2'h2)]))))
                    begin
                      reg5645 <= forvar5663[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg5645 <= (~&reg5675);
                      reg5646 <= forvar5549[(3'h7):(3'h6)];
                    end
                end
              for (forvar5650 = (1'h0); (forvar5650 < (2'h2)); forvar5650 = (forvar5650 + (1'h1)))
                begin
                  reg5651 <= reg5632[(1'h1):(1'h0)];
                  for (forvar5652 = (1'h0); (forvar5652 < (1'h0)); forvar5652 = (forvar5652 + (1'h1)))
                    begin
                      reg5653 <= reg5709[(2'h3):(1'h0)];
                      reg5654 <= $signed((^~({reg5518} ?
                          $signed((8'ha3)) : reg5664[(3'h4):(2'h2)])));
                    end
                  for (forvar5655 = (1'h0); (forvar5655 < (2'h2)); forvar5655 = (forvar5655 + (1'h1)))
                    begin
                      reg5656 <= reg5644;
                    end
                end
              for (forvar5657 = (1'h0); (forvar5657 < (1'h1)); forvar5657 = (forvar5657 + (1'h1)))
                begin
                  for (forvar5658 = (1'h0); (forvar5658 < (2'h2)); forvar5658 = (forvar5658 + (1'h1)))
                    begin
                      reg5659 <= $unsigned($unsigned(forvar5646[(3'h7):(2'h3)]));
                      reg5660 <= reg5577[(4'hb):(4'h8)];
                      reg5661 <= ($signed((-(~&forvar5580))) * $signed((^$unsigned(reg5659))));
                    end
                  for (forvar5662 = (1'h0); (forvar5662 < (2'h2)); forvar5662 = (forvar5662 + (1'h1)))
                    begin
                      reg5663 <= reg5677[(3'h7):(3'h4)];
                      reg5664 <= (~^((reg5581[(3'h6):(1'h0)] != reg5532) | ((^forvar5588) ?
                          (reg5597 ? reg5664 : reg5553) : $unsigned(reg5586))));
                    end
                end
            end
          for (forvar5665 = (1'h0); (forvar5665 < (2'h3)); forvar5665 = (forvar5665 + (1'h1)))
            begin
              if ($unsigned(reg5550))
                begin
                  if ((reg5526 ?
                      (~($unsigned(reg5615) ?
                          $unsigned((8'hae)) : $unsigned(reg5584))) : (~$signed((reg5603 >>> reg5599)))))
                    begin
                      reg5666 <= $signed((((reg5540 + (8'ha3)) <= reg5626[(3'h7):(2'h3)]) ?
                          reg5691 : ($signed((8'hb5)) & (reg5534 <= reg5580))));
                      reg5667 <= reg5684;
                    end
                  else
                    begin
                      reg5666 <= reg5527[(4'ha):(2'h2)];
                      reg5667 <= reg5669;
                      reg5668 <= $unsigned(($signed((reg5684 ?
                          reg5518 : reg5675)) < ((wire5641 ~^ (8'ha4)) == {reg5578})));
                    end
                  reg5669 <= $signed(wire5642);
                  for (forvar5670 = (1'h0); (forvar5670 < (1'h1)); forvar5670 = (forvar5670 + (1'h1)))
                    begin
                      reg5671 <= {reg5664[(1'h1):(1'h0)]};
                      reg5672 <= {((reg5644 ^~ reg5678) <<< (reg5531[(3'h5):(3'h4)] ?
                              (|reg5684) : $signed(forvar5671)))};
                      reg5673 <= ((8'hae) ?
                          reg5684 : {$unsigned((reg5666 * reg5571))});
                      reg5674 <= (forvar5650[(2'h2):(2'h2)] && ((^((8'hb4) ?
                              reg5681 : reg5635)) ?
                          $unsigned((^~forvar5605)) : ((forvar5613 == reg5626) ?
                              (|reg5702) : (reg5708 ? reg5541 : forvar5657))));
                    end
                  if ($unsigned(($signed($unsigned(reg5519)) | (&{reg5534}))))
                    begin
                      reg5675 <= $signed($signed(($signed(reg5658) ?
                          reg5677 : (reg5586 >= reg5538))));
                      reg5676 <= reg5554[(3'h6):(3'h6)];
                      reg5677 <= $unsigned(({(reg5652 && forvar5629)} > (!$signed(forvar5564))));
                      reg5678 <= reg5687;
                    end
                  else
                    begin
                      reg5675 <= (reg5526 ?
                          reg5710 : $signed((reg5632[(1'h1):(1'h0)] <= $signed(reg5695))));
                      reg5676 <= (-(8'hb6));
                    end
                end
              else
                begin
                  reg5666 <= reg5669[(4'ha):(3'h7)];
                  if (($unsigned($signed($unsigned(reg5710))) ?
                      ((~|(^reg5551)) >= $signed({forvar5575})) : forvar5704))
                    begin
                      reg5667 <= (((8'hb0) >> $signed((|reg5598))) ^ forvar5569[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg5667 <= reg5619[(3'h5):(1'h1)];
                      reg5668 <= {(^$signed($signed(wire5515)))};
                    end
                  for (forvar5669 = (1'h0); (forvar5669 < (2'h2)); forvar5669 = (forvar5669 + (1'h1)))
                    begin
                      reg5670 <= (reg5545 ?
                          reg5556[(2'h3):(2'h2)] : (reg5680 < reg5640));
                    end
                  for (forvar5671 = (1'h0); (forvar5671 < (1'h0)); forvar5671 = (forvar5671 + (1'h1)))
                    begin
                      reg5672 <= $signed(($signed($unsigned(reg5621)) <= ((forvar5680 || reg5647) ?
                          reg5710 : (~|reg5525))));
                      reg5673 <= ((~&reg5677[(3'h6):(3'h4)]) ~^ reg5621[(2'h2):(1'h1)]);
                    end
                end
              for (forvar5679 = (1'h0); (forvar5679 < (2'h2)); forvar5679 = (forvar5679 + (1'h1)))
                begin
                  if ((^~(8'hb1)))
                    begin
                      reg5680 <= $signed((($signed(reg5530) | {reg5523}) << {$signed(forvar5610)}));
                      reg5681 <= $signed(reg5621[(3'h7):(3'h4)]);
                      reg5682 <= ((~$signed(reg5676)) > $signed(reg5658));
                    end
                  else
                    begin
                      reg5680 <= $unsigned($signed(forvar5575));
                      reg5681 <= (reg5662 && $unsigned(reg5676[(2'h2):(2'h2)]));
                    end
                  for (forvar5683 = (1'h0); (forvar5683 < (1'h1)); forvar5683 = (forvar5683 + (1'h1)))
                    begin
                      reg5684 <= $signed(((forvar5588 != (8'haa)) ?
                          ((reg5593 ?
                              reg5630 : reg5595) && (+reg5711)) : ($unsigned(forvar5519) ?
                              (8'hac) : (|(8'ha0)))));
                    end
                end
              reg5685 <= (reg5651 ?
                  (reg5697[(2'h2):(2'h2)] ^~ $unsigned(reg5586[(1'h1):(1'h1)])) : (8'hb7));
              for (forvar5686 = (1'h0); (forvar5686 < (1'h0)); forvar5686 = (forvar5686 + (1'h1)))
                begin
                  for (forvar5687 = (1'h0); (forvar5687 < (2'h2)); forvar5687 = (forvar5687 + (1'h1)))
                    begin
                      reg5688 <= reg5698[(1'h0):(1'h0)];
                      reg5689 <= (~|(($unsigned(reg5699) ?
                          forvar5646 : $unsigned(reg5597)) ^~ ($unsigned((8'hb3)) ?
                          reg5711 : $signed(forvar5542))));
                      reg5690 <= reg5669[(1'h1):(1'h0)];
                      reg5691 <= ((reg5702[(1'h1):(1'h1)] == reg5523[(3'h5):(1'h1)]) * reg5584);
                    end
                  for (forvar5692 = (1'h0); (forvar5692 < (2'h3)); forvar5692 = (forvar5692 + (1'h1)))
                    begin
                      reg5693 <= forvar5540[(1'h1):(1'h0)];
                    end
                end
            end
          for (forvar5694 = (1'h0); (forvar5694 < (1'h0)); forvar5694 = (forvar5694 + (1'h1)))
            begin
              for (forvar5695 = (1'h0); (forvar5695 < (2'h3)); forvar5695 = (forvar5695 + (1'h1)))
                begin
                  if (forvar5628[(2'h3):(1'h1)])
                    begin
                      reg5696 <= $unsigned((+({forvar5618} <= (forvar5596 < reg5662))));
                      reg5697 <= (&(+$unsigned($unsigned((8'ha2)))));
                    end
                  else
                    begin
                      reg5696 <= {(((wire5642 || reg5536) ?
                                  reg5644 : reg5702[(3'h6):(2'h2)]) ?
                              $unsigned($signed(forvar5669)) : forvar5662)};
                      reg5697 <= reg5606;
                      reg5698 <= ($signed(reg5568) ?
                          (reg5538 ?
                              ((forvar5590 >> reg5540) > $unsigned(forvar5663)) : $unsigned({reg5705})) : $signed(forvar5555));
                    end
                  reg5699 <= (reg5615[(2'h2):(1'h1)] ?
                      reg5669 : (reg5693[(2'h2):(1'h1)] + $unsigned((-(8'h9e)))));
                  for (forvar5700 = (1'h0); (forvar5700 < (1'h0)); forvar5700 = (forvar5700 + (1'h1)))
                    begin
                      reg5701 <= (($signed((reg5554 ? forvar5589 : reg5531)) ?
                              (8'h9c) : forvar5663) ?
                          (&(-(reg5536 != reg5667))) : forvar5564);
                      reg5702 <= reg5590[(1'h0):(1'h0)];
                    end
                end
              for (forvar5703 = (1'h0); (forvar5703 < (1'h0)); forvar5703 = (forvar5703 + (1'h1)))
                begin
                  for (forvar5704 = (1'h0); (forvar5704 < (1'h1)); forvar5704 = (forvar5704 + (1'h1)))
                    begin
                      reg5705 <= $signed($unsigned((~^reg5559)));
                      reg5706 <= reg5520[(3'h6):(3'h5)];
                      reg5707 <= (-$unsigned(reg5689));
                    end
                  reg5708 <= $unsigned((~^$unsigned(reg5678[(4'h8):(3'h7)])));
                  for (forvar5709 = (1'h0); (forvar5709 < (1'h0)); forvar5709 = (forvar5709 + (1'h1)))
                    begin
                      reg5710 <= (^~reg5711[(1'h1):(1'h0)]);
                      reg5711 <= reg5688[(1'h1):(1'h0)];
                      reg5712 <= $unsigned(((8'hb4) ?
                          reg5536[(4'h9):(1'h0)] : reg5656));
                    end
                  reg5713 <= (reg5553[(4'h9):(3'h6)] ?
                      $unsigned($signed((forvar5517 ?
                          (8'ha7) : forvar5610))) : $unsigned((^$signed(forvar5587))));
                end
              reg5714 <= $unsigned($signed($unsigned((&reg5552))));
            end
        end
      reg5715 <= $unsigned(reg5651[(4'hb):(4'h9)]);
      if ($unsigned({(-(+reg5600))}))
        begin
          for (forvar5716 = (1'h0); (forvar5716 < (1'h1)); forvar5716 = (forvar5716 + (1'h1)))
            begin
              if ((($signed({reg5685}) ?
                  ((reg5708 ? reg5615 : reg5652) ?
                      wire5643 : wire5513) : ((8'ha0) ?
                      forvar5629 : $signed(reg5590))) + $unsigned(reg5520)))
                begin
                  reg5717 <= $signed($unsigned($signed((forvar5543 ?
                      reg5703 : reg5572))));
                end
              else
                begin
                  for (forvar5717 = (1'h0); (forvar5717 < (1'h1)); forvar5717 = (forvar5717 + (1'h1)))
                    begin
                      reg5718 <= ({((8'hb9) ? (|reg5525) : forvar5587)} ?
                          (reg5537[(4'h9):(2'h3)] <<< reg5561) : $signed($unsigned((reg5612 & forvar5662))));
                      reg5719 <= (({$signed(reg5706)} ?
                              reg5557 : $unsigned(reg5651)) ?
                          (8'hb3) : reg5700);
                      reg5720 <= $unsigned((8'ha4));
                      reg5721 <= (+{{$signed(forvar5703)}});
                    end
                  if (({(|reg5584)} == ((^~(^reg5565)) & $signed(reg5520[(4'hc):(3'h7)]))))
                    begin
                      reg5722 <= (^~(~&reg5533));
                    end
                  else
                    begin
                      reg5722 <= $signed({forvar5646});
                      reg5723 <= reg5622;
                      reg5724 <= reg5570;
                    end
                  for (forvar5725 = (1'h0); (forvar5725 < (2'h3)); forvar5725 = (forvar5725 + (1'h1)))
                    begin
                      reg5726 <= (&(^~$signed((reg5649 ?
                          wire5513 : forvar5519))));
                    end
                end
              if ($unsigned({{$signed(forvar5636)}}))
                begin
                  reg5727 <= {$unsigned($unsigned($unsigned((8'h9f))))};
                end
              else
                begin
                  if ((!(($unsigned((8'h9f)) >>> forvar5529) == $unsigned(forvar5536[(3'h5):(2'h2)]))))
                    begin
                      reg5727 <= $unsigned((!$signed(reg5608)));
                      reg5728 <= (~&(((reg5715 <<< reg5596) < $signed(reg5690)) >>> $unsigned($unsigned(reg5713))));
                      reg5729 <= {reg5593[(3'h7):(3'h5)]};
                    end
                  else
                    begin
                      reg5727 <= $unsigned(forvar5538[(3'h5):(3'h4)]);
                    end
                  for (forvar5730 = (1'h0); (forvar5730 < (2'h3)); forvar5730 = (forvar5730 + (1'h1)))
                    begin
                      reg5731 <= reg5584;
                      reg5732 <= $unsigned($unsigned((8'ha4)));
                    end
                  for (forvar5733 = (1'h0); (forvar5733 < (1'h0)); forvar5733 = (forvar5733 + (1'h1)))
                    begin
                      reg5734 <= (8'ha5);
                      reg5735 <= reg5578;
                      reg5736 <= $unsigned($signed(reg5660[(4'hf):(4'h8)]));
                      reg5737 <= ($signed((reg5676 ?
                          {reg5713} : (&forvar5646))) != reg5633[(4'hb):(1'h1)]);
                    end
                end
            end
          for (forvar5738 = (1'h0); (forvar5738 < (2'h3)); forvar5738 = (forvar5738 + (1'h1)))
            begin
              for (forvar5739 = (1'h0); (forvar5739 < (1'h0)); forvar5739 = (forvar5739 + (1'h1)))
                begin
                  if (reg5580)
                    begin
                      reg5740 <= reg5653[(1'h0):(1'h0)];
                      reg5741 <= $signed($signed(reg5566[(1'h0):(1'h0)]));
                      reg5742 <= (^forvar5546[(4'he):(2'h3)]);
                      reg5743 <= $signed(reg5589);
                    end
                  else
                    begin
                      reg5740 <= reg5666;
                      reg5741 <= reg5525[(1'h1):(1'h0)];
                      reg5742 <= $signed($signed({(reg5674 <<< reg5679)}));
                    end
                  reg5744 <= {$unsigned(reg5552)};
                  reg5745 <= (forvar5611[(1'h1):(1'h0)] != (($signed((8'ha7)) - (reg5672 || reg5638)) ?
                      {((8'hb8) + reg5562)} : $signed($signed(forvar5683))));
                  for (forvar5746 = (1'h0); (forvar5746 < (1'h1)); forvar5746 = (forvar5746 + (1'h1)))
                    begin
                      reg5747 <= reg5633;
                    end
                end
              reg5748 <= $unsigned($unsigned($unsigned((reg5570 ?
                  reg5669 : forvar5699))));
              if ($signed($signed({$unsigned(reg5531)})))
                begin
                  if (reg5727)
                    begin
                      reg5749 <= forvar5687[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg5749 <= forvar5686;
                      reg5750 <= wire5514[(3'h4):(2'h3)];
                      reg5751 <= forvar5662;
                    end
                  for (forvar5752 = (1'h0); (forvar5752 < (2'h2)); forvar5752 = (forvar5752 + (1'h1)))
                    begin
                      reg5753 <= ((|({(8'hab)} ?
                          (-reg5559) : {reg5687})) < $unsigned($unsigned(forvar5628[(4'h9):(4'h8)])));
                      reg5754 <= (reg5558[(3'h6):(2'h3)] ?
                          (($signed(forvar5733) ?
                              (forvar5739 != reg5522) : reg5524[(2'h2):(1'h1)]) ^ ((~&reg5713) ?
                              (reg5578 ?
                                  reg5719 : forvar5547) : $signed(forvar5669))) : (forvar5694 ?
                              {(8'ha3)} : (&{forvar5529})));
                    end
                  reg5755 <= reg5706[(1'h0):(1'h0)];
                  reg5756 <= $signed(((~reg5736) && forvar5686[(1'h1):(1'h0)]));
                end
              else
                begin
                  if (reg5753)
                    begin
                      reg5749 <= reg5662;
                    end
                  else
                    begin
                      reg5749 <= $signed((~^({(8'h9f)} && (|(8'hb2)))));
                      reg5750 <= $unsigned($unsigned(reg5694[(1'h1):(1'h0)]));
                    end
                  for (forvar5751 = (1'h0); (forvar5751 < (2'h2)); forvar5751 = (forvar5751 + (1'h1)))
                    begin
                      reg5752 <= reg5685[(3'h4):(1'h0)];
                      reg5753 <= ((~$unsigned((8'hb2))) <= wire5512);
                      reg5754 <= $unsigned(({(^~reg5666)} ?
                          $unsigned({reg5714}) : {reg5597}));
                      reg5755 <= {(^~((-reg5593) ?
                              forvar5526 : forvar5703[(2'h2):(2'h2)]))};
                    end
                  for (forvar5756 = (1'h0); (forvar5756 < (2'h2)); forvar5756 = (forvar5756 + (1'h1)))
                    begin
                      reg5757 <= ($unsigned((reg5670 - {reg5592})) >>> $signed((~|(reg5682 ?
                          (8'ha9) : forvar5668))));
                      reg5758 <= forvar5578[(1'h0):(1'h0)];
                      reg5759 <= (^$unsigned(($signed((8'h9e)) ?
                          (reg5520 ? (8'ha4) : reg5527) : $signed(wire5512))));
                      reg5760 <= ($signed($signed($unsigned(forvar5519))) && (^{{(8'ha6)}}));
                    end
                end
            end
        end
      else
        begin
          reg5716 <= {$signed((forvar5546[(4'hc):(4'h9)] ? reg5671 : reg5754))};
          if ((~|(|((forvar5569 ? forvar5704 : forvar5558) | (~^reg5608)))))
            begin
              reg5717 <= reg5577[(4'hc):(3'h7)];
              for (forvar5718 = (1'h0); (forvar5718 < (1'h1)); forvar5718 = (forvar5718 + (1'h1)))
                begin
                  reg5719 <= reg5535;
                  for (forvar5720 = (1'h0); (forvar5720 < (1'h1)); forvar5720 = (forvar5720 + (1'h1)))
                    begin
                      reg5721 <= (~^$unsigned(forvar5588));
                      reg5722 <= ($signed(reg5699) < reg5709);
                      reg5723 <= (forvar5542[(1'h0):(1'h0)] <<< reg5654);
                      reg5724 <= (((forvar5517[(2'h3):(2'h2)] ?
                          $signed((8'hb3)) : $signed(reg5752)) ^ ((reg5740 <<< forvar5620) ?
                          (reg5674 ? forvar5580 : reg5556) : (reg5581 ?
                              reg5563 : reg5708))) - (($unsigned(reg5714) ?
                              ((8'hb4) + forvar5647) : $signed(reg5582)) ?
                          $signed($signed(reg5679)) : ((reg5670 ?
                              reg5744 : (8'hb6)) == forvar5752)));
                    end
                end
              for (forvar5725 = (1'h0); (forvar5725 < (2'h3)); forvar5725 = (forvar5725 + (1'h1)))
                begin
                  for (forvar5726 = (1'h0); (forvar5726 < (1'h0)); forvar5726 = (forvar5726 + (1'h1)))
                    begin
                      reg5727 <= (reg5592 ?
                          reg5551 : forvar5679[(4'hf):(4'hb)]);
                      reg5728 <= (!$signed((((8'ha9) == reg5721) | $unsigned(reg5742))));
                      reg5729 <= $signed(reg5530);
                    end
                  for (forvar5730 = (1'h0); (forvar5730 < (2'h2)); forvar5730 = (forvar5730 + (1'h1)))
                    begin
                      reg5731 <= wire5641;
                      reg5732 <= ({reg5606} * reg5719);
                      reg5733 <= reg5656;
                    end
                  for (forvar5734 = (1'h0); (forvar5734 < (1'h1)); forvar5734 = (forvar5734 + (1'h1)))
                    begin
                      reg5735 <= $unsigned(reg5603);
                      reg5736 <= reg5678;
                      reg5737 <= $signed(reg5622);
                      reg5738 <= (~&reg5626);
                    end
                  for (forvar5739 = (1'h0); (forvar5739 < (1'h1)); forvar5739 = (forvar5739 + (1'h1)))
                    begin
                      reg5740 <= forvar5652[(3'h5):(2'h2)];
                    end
                end
            end
          else
            begin
              if ((~|$signed({(^~(8'hb0))})))
                begin
                  if (($signed({reg5751[(3'h5):(2'h3)]}) & (forvar5549 > reg5579[(2'h3):(1'h0)])))
                    begin
                      reg5717 <= {$signed(forvar5538)};
                      reg5718 <= ($signed(reg5688[(2'h3):(1'h1)]) ?
                          (($unsigned(reg5675) ^~ $unsigned(reg5527)) ?
                              forvar5716[(3'h7):(1'h1)] : (-forvar5628)) : forvar5564);
                    end
                  else
                    begin
                      reg5717 <= reg5560;
                    end
                end
              else
                begin
                  for (forvar5717 = (1'h0); (forvar5717 < (1'h0)); forvar5717 = (forvar5717 + (1'h1)))
                    begin
                      reg5718 <= ($signed(forvar5537[(1'h1):(1'h1)]) ?
                          (({(8'ha1)} ? (!(8'ha5)) : $unsigned(reg5599)) ?
                              (8'hac) : forvar5699[(3'h7):(3'h6)]) : (&(reg5568[(3'h6):(2'h2)] ?
                              (wire5643 ? reg5734 : reg5744) : (|reg5584))));
                      reg5719 <= $signed(forvar5546);
                      reg5720 <= $unsigned((&$unsigned($unsigned(reg5541))));
                    end
                end
              if ($signed(reg5608[(2'h2):(1'h1)]))
                begin
                  if (((~|(|{reg5516})) ?
                      reg5707[(2'h2):(1'h0)] : $signed((~|forvar5627[(1'h0):(1'h0)]))))
                    begin
                      reg5721 <= $unsigned($unsigned($unsigned((reg5644 & forvar5558))));
                      reg5722 <= forvar5673;
                    end
                  else
                    begin
                      reg5721 <= reg5581[(4'h9):(1'h0)];
                      reg5722 <= $unsigned($signed((-((8'ha8) ?
                          forvar5650 : reg5578))));
                      reg5723 <= (^~$signed($unsigned(reg5691[(3'h4):(2'h3)])));
                      reg5724 <= (~|((wire5641 ?
                          $unsigned(reg5706) : ((8'h9f) + (8'ha4))) | $signed(reg5659)));
                    end
                  for (forvar5725 = (1'h0); (forvar5725 < (1'h1)); forvar5725 = (forvar5725 + (1'h1)))
                    begin
                      reg5726 <= (~^$unsigned((8'hb1)));
                      reg5727 <= reg5624;
                    end
                  if (reg5625[(2'h3):(1'h1)])
                    begin
                      reg5728 <= forvar5665[(1'h1):(1'h1)];
                      reg5729 <= ($unsigned((&$unsigned(reg5635))) ^ {{$unsigned(forvar5564)}});
                    end
                  else
                    begin
                      reg5728 <= (reg5623 - {(~|{reg5753})});
                    end
                  if ((-($unsigned((reg5519 ? forvar5605 : forvar5673)) ?
                      (~^(reg5599 == reg5531)) : ((~&reg5711) == $unsigned(reg5630)))))
                    begin
                      reg5730 <= (-$unsigned($unsigned(reg5699)));
                      reg5731 <= reg5683;
                    end
                  else
                    begin
                      reg5730 <= (^((8'hba) ^ ($signed(forvar5657) && $unsigned(reg5689))));
                      reg5731 <= $unsigned((($signed(wire5642) != (reg5614 ^ reg5756)) >= $signed(reg5709[(4'hf):(4'ha)])));
                      reg5732 <= (+(^~(reg5551 <<< reg5710[(2'h2):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar5721 = (1'h0); (forvar5721 < (1'h1)); forvar5721 = (forvar5721 + (1'h1)))
                    begin
                      reg5722 <= {$signed((~(forvar5549 && reg5676)))};
                    end
                  if ($unsigned((($signed(forvar5726) ?
                          ((8'hba) != forvar5668) : reg5723) ?
                      (~|(reg5710 ?
                          forvar5646 : reg5597)) : (+reg5685[(3'h6):(3'h4)]))))
                    begin
                      reg5723 <= (8'haf);
                      reg5724 <= ((^~$unsigned((reg5716 ? (8'hb2) : reg5600))) ?
                          $signed($unsigned(reg5721[(1'h0):(1'h0)])) : (^$unsigned(reg5567[(4'h9):(1'h0)])));
                      reg5725 <= $signed((reg5592 ?
                          ((~reg5666) ?
                              $unsigned(reg5670) : {reg5705}) : forvar5652[(3'h6):(2'h3)]));
                    end
                  else
                    begin
                      reg5723 <= reg5589[(3'h5):(2'h2)];
                      reg5724 <= (8'ha9);
                    end
                  if ((~{((reg5626 && (8'haa)) ?
                          {reg5710} : (forvar5519 ^~ forvar5596))}))
                    begin
                      reg5726 <= (reg5520[(3'h7):(3'h4)] ?
                          $signed(((~&reg5718) ?
                              $unsigned(forvar5730) : reg5687[(4'hc):(3'h6)])) : $unsigned($unsigned(((8'h9d) >= reg5592))));
                    end
                  else
                    begin
                      reg5726 <= {reg5681};
                      reg5727 <= ((-$signed(forvar5717)) ?
                          $unsigned({(forvar5695 ?
                                  reg5562 : forvar5673)}) : forvar5540);
                      reg5728 <= $signed({reg5649[(3'h5):(2'h2)]});
                    end
                  if (((reg5599 ?
                          (|(reg5669 ?
                              reg5532 : reg5721)) : $signed($unsigned(reg5523))) ?
                      forvar5681 : reg5551))
                    begin
                      reg5729 <= $signed($unsigned(forvar5718));
                      reg5730 <= (8'h9d);
                      reg5731 <= ({$unsigned((reg5757 ~^ reg5529))} <<< {(((8'h9d) ?
                              reg5718 : forvar5684) << $signed(forvar5725))});
                    end
                  else
                    begin
                      reg5729 <= (&(((^reg5622) ? reg5602 : forvar5721) ?
                          $unsigned(((8'h9f) << reg5743)) : $signed($unsigned(reg5634))));
                      reg5730 <= (wire5513 ?
                          $signed((|(reg5633 ? (8'had) : reg5616))) : (reg5659 ?
                              reg5725 : $signed($signed(reg5738))));
                      reg5731 <= {(+$signed((forvar5590 ? reg5677 : (8'ha0))))};
                      reg5732 <= (reg5742[(4'h8):(2'h3)] > ($signed(forvar5700) ?
                          (forvar5631 || $signed(reg5619)) : $signed(reg5659[(2'h2):(2'h2)])));
                    end
                end
              for (forvar5733 = (1'h0); (forvar5733 < (2'h3)); forvar5733 = (forvar5733 + (1'h1)))
                begin
                  for (forvar5734 = (1'h0); (forvar5734 < (1'h0)); forvar5734 = (forvar5734 + (1'h1)))
                    begin
                      reg5735 <= reg5701;
                      reg5736 <= wire5641[(3'h5):(2'h2)];
                    end
                  reg5737 <= (^~(8'hac));
                end
              if ((8'hb2))
                begin
                  if (forvar5695[(4'h9):(1'h0)])
                    begin
                      reg5738 <= (((!(~^(8'hb6))) >> reg5553[(1'h1):(1'h1)]) && {$signed((reg5745 ?
                              reg5589 : reg5689))});
                      reg5739 <= reg5625[(1'h1):(1'h0)];
                      reg5740 <= {$signed($unsigned({(8'hb6)}))};
                      reg5741 <= (({forvar5529[(4'h9):(3'h4)]} ?
                              ((-reg5638) ?
                                  {reg5732} : (+forvar5593)) : $signed((forvar5718 != reg5572))) ?
                          reg5598[(3'h5):(2'h2)] : reg5729[(4'h8):(4'h8)]);
                    end
                  else
                    begin
                      reg5738 <= (+$unsigned(((|reg5612) >> reg5712[(1'h1):(1'h0)])));
                    end
                  if ($signed($signed($signed({forvar5704}))))
                    begin
                      reg5742 <= (forvar5645 ?
                          forvar5725 : $signed(forvar5527));
                      reg5743 <= (reg5722 ?
                          reg5687 : $signed($unsigned(reg5733[(3'h5):(1'h1)])));
                    end
                  else
                    begin
                      reg5742 <= reg5740;
                      reg5743 <= reg5693[(3'h4):(1'h0)];
                      reg5744 <= $unsigned((reg5751[(2'h2):(1'h1)] | (-$signed((8'hab)))));
                      reg5745 <= reg5759;
                    end
                  reg5746 <= $signed(((forvar5631 ?
                      $unsigned(reg5640) : $unsigned((8'hb0))) != $unsigned((&(8'h9f)))));
                end
              else
                begin
                  for (forvar5738 = (1'h0); (forvar5738 < (1'h1)); forvar5738 = (forvar5738 + (1'h1)))
                    begin
                      reg5739 <= ((!$signed(forvar5593[(1'h1):(1'h1)])) ?
                          (forvar5645 && (reg5590 >= {wire5514})) : $signed(reg5721));
                    end
                  reg5740 <= (reg5550 ?
                      ((8'h9e) + ($signed(reg5586) <= (8'hb6))) : ((&{(8'hb9)}) ?
                          $unsigned((reg5681 ?
                              forvar5681 : reg5541)) : $unsigned($signed((8'ha9)))));
                  for (forvar5741 = (1'h0); (forvar5741 < (1'h1)); forvar5741 = (forvar5741 + (1'h1)))
                    begin
                      reg5742 <= {forvar5620[(3'h4):(3'h4)]};
                      reg5743 <= {$unsigned((8'hb9))};
                      reg5744 <= $signed(($signed(((8'hb5) && forvar5540)) ?
                          (~^{reg5701}) : $unsigned((reg5670 >> reg5699))));
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar5761 = (1'h0); (forvar5761 < (2'h2)); forvar5761 = (forvar5761 + (1'h1)))
        begin
          for (forvar5762 = (1'h0); (forvar5762 < (2'h2)); forvar5762 = (forvar5762 + (1'h1)))
            begin
              for (forvar5763 = (1'h0); (forvar5763 < (1'h0)); forvar5763 = (forvar5763 + (1'h1)))
                begin
                  if (reg5600)
                    begin
                      reg5764 <= {(~|(^~reg5530))};
                    end
                  else
                    begin
                      reg5764 <= $signed((|(((8'hb5) > forvar5738) << reg5689)));
                      reg5765 <= {reg5542[(1'h1):(1'h1)]};
                      reg5766 <= (-($unsigned((reg5608 ?
                              forvar5669 : reg5759)) ?
                          forvar5716[(1'h1):(1'h1)] : reg5609[(1'h0):(1'h0)]));
                      reg5767 <= ((8'ha7) != reg5531[(3'h5):(2'h2)]);
                    end
                  for (forvar5768 = (1'h0); (forvar5768 < (1'h1)); forvar5768 = (forvar5768 + (1'h1)))
                    begin
                      reg5769 <= (|(reg5645 ~^ ((reg5590 ^ reg5536) ?
                          $signed((8'h9c)) : $unsigned((8'hae)))));
                    end
                end
              reg5770 <= ((forvar5518 ?
                      (+$signed(forvar5646)) : $unsigned(reg5551)) ?
                  (!forvar5762) : (((8'hb9) <<< forvar5613[(2'h3):(1'h1)]) && (reg5557[(2'h2):(2'h2)] > forvar5655)));
            end
        end
      for (forvar5771 = (1'h0); (forvar5771 < (1'h0)); forvar5771 = (forvar5771 + (1'h1)))
        begin
          for (forvar5772 = (1'h0); (forvar5772 < (2'h2)); forvar5772 = (forvar5772 + (1'h1)))
            begin
              for (forvar5773 = (1'h0); (forvar5773 < (2'h2)); forvar5773 = (forvar5773 + (1'h1)))
                begin
                  if (({$signed(((8'h9c) ? forvar5636 : reg5568))} ?
                      $signed(forvar5529[(4'ha):(1'h1)]) : reg5718))
                    begin
                      reg5774 <= forvar5590;
                      reg5775 <= (((reg5674 << reg5521) || reg5524[(2'h3):(2'h3)]) ?
                          (-reg5599) : {({forvar5652} ?
                                  (reg5633 ?
                                      reg5520 : (8'haf)) : (&forvar5746))});
                      reg5776 <= $unsigned((|$unsigned(reg5741[(3'h5):(3'h5)])));
                    end
                  else
                    begin
                      reg5774 <= $signed($signed(((reg5755 < reg5714) ?
                          (8'hb5) : {reg5563})));
                      reg5775 <= ((|reg5712[(3'h6):(2'h3)]) ~^ $unsigned(reg5565));
                    end
                  for (forvar5777 = (1'h0); (forvar5777 < (1'h0)); forvar5777 = (forvar5777 + (1'h1)))
                    begin
                      reg5778 <= reg5680[(1'h1):(1'h1)];
                      reg5779 <= (~|$unsigned(($signed(reg5546) ^ reg5652)));
                    end
                  for (forvar5780 = (1'h0); (forvar5780 < (2'h3)); forvar5780 = (forvar5780 + (1'h1)))
                    begin
                      reg5781 <= reg5532;
                      reg5782 <= ($unsigned($unsigned($signed(forvar5613))) * ($signed((&reg5703)) ~^ reg5664[(3'h4):(1'h1)]));
                      reg5783 <= (reg5708[(2'h2):(2'h2)] ?
                          (reg5523 ?
                              $signed($signed(forvar5741)) : reg5606[(3'h4):(2'h3)]) : (((reg5720 >= reg5673) ?
                              $signed(reg5639) : $unsigned(forvar5771)) + reg5578));
                      reg5784 <= (reg5571[(4'h8):(4'h8)] - $signed($signed((reg5653 ?
                          forvar5780 : forvar5679))));
                    end
                  for (forvar5785 = (1'h0); (forvar5785 < (1'h0)); forvar5785 = (forvar5785 + (1'h1)))
                    begin
                      reg5786 <= (reg5760[(3'h6):(2'h2)] & reg5632[(1'h1):(1'h1)]);
                      reg5787 <= ({$unsigned((reg5639 >>> reg5578))} ?
                          (8'hab) : reg5774[(1'h1):(1'h0)]);
                    end
                end
            end
          reg5788 <= (8'haa);
          for (forvar5789 = (1'h0); (forvar5789 < (1'h1)); forvar5789 = (forvar5789 + (1'h1)))
            begin
              for (forvar5790 = (1'h0); (forvar5790 < (2'h3)); forvar5790 = (forvar5790 + (1'h1)))
                begin
                  for (forvar5791 = (1'h0); (forvar5791 < (2'h3)); forvar5791 = (forvar5791 + (1'h1)))
                    begin
                      reg5792 <= {(reg5745 <<< forvar5668)};
                      reg5793 <= reg5766[(2'h2):(2'h2)];
                      reg5794 <= (forvar5777 ~^ (forvar5699[(3'h7):(1'h1)] ?
                          reg5516 : (((8'hba) ? (8'hb9) : reg5774) ?
                              reg5616 : (reg5602 + (8'ha0)))));
                    end
                  if ($signed((reg5784 * $unsigned(forvar5726))))
                    begin
                      reg5795 <= (&(reg5526 ?
                          (reg5640[(1'h1):(1'h1)] ?
                              reg5555[(2'h2):(2'h2)] : reg5530) : $unsigned($signed(reg5634))));
                    end
                  else
                    begin
                      reg5795 <= (reg5567[(4'ha):(3'h5)] ?
                          $unsigned((((8'ha1) ^ reg5661) >> (~|reg5595))) : wire5641);
                      reg5796 <= ((8'hb0) + forvar5611);
                      reg5797 <= $unsigned(((reg5746[(1'h0):(1'h0)] + (reg5744 & reg5545)) ?
                          {$unsigned(forvar5741)} : reg5582[(4'h9):(3'h7)]));
                      reg5798 <= (~&$unsigned(reg5522));
                    end
                  for (forvar5799 = (1'h0); (forvar5799 < (2'h2)); forvar5799 = (forvar5799 + (1'h1)))
                    begin
                      reg5800 <= (reg5529[(2'h2):(2'h2)] * $unsigned(reg5535));
                    end
                  for (forvar5801 = (1'h0); (forvar5801 < (2'h3)); forvar5801 = (forvar5801 + (1'h1)))
                    begin
                      reg5802 <= $unsigned($unsigned(((+reg5672) ?
                          forvar5655 : $unsigned(forvar5763))));
                      reg5803 <= {((reg5651[(1'h1):(1'h1)] ?
                              $signed((8'ha9)) : reg5598) >>> ($signed(forvar5761) ?
                              reg5687 : (8'hac)))};
                    end
                end
              for (forvar5804 = (1'h0); (forvar5804 < (1'h1)); forvar5804 = (forvar5804 + (1'h1)))
                begin
                  for (forvar5805 = (1'h0); (forvar5805 < (1'h0)); forvar5805 = (forvar5805 + (1'h1)))
                    begin
                      reg5806 <= $signed($unsigned({reg5776[(1'h1):(1'h1)]}));
                    end
                  if (reg5724)
                    begin
                      reg5807 <= reg5767;
                      reg5808 <= $unsigned((forvar5647 ? reg5568 : reg5599));
                      reg5809 <= forvar5668;
                      reg5810 <= ((^{(^~reg5578)}) ?
                          (({forvar5575} ?
                                  (forvar5675 ?
                                      reg5607 : reg5524) : ((8'ha6) <= reg5547)) ?
                              ({forvar5752} ?
                                  (wire5514 * reg5764) : (~forvar5537)) : ((~&forvar5805) >>> wire5515)) : ({{(8'ha0)}} ?
                              reg5568 : ((forvar5589 ? (8'hb6) : reg5593) ?
                                  (~&forvar5790) : {forvar5772})));
                    end
                  else
                    begin
                      reg5807 <= (^~reg5615);
                      reg5808 <= $signed(($signed({forvar5620}) ?
                          ($signed(reg5730) ^~ forvar5587[(3'h7):(1'h0)]) : {(reg5727 != forvar5799)}));
                      reg5809 <= $signed(($signed((reg5770 | reg5557)) && reg5732));
                    end
                end
              if (reg5671)
                begin
                  reg5811 <= (^~reg5676[(1'h1):(1'h0)]);
                  if ($unsigned(reg5539[(3'h4):(2'h2)]))
                    begin
                      reg5812 <= reg5532[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg5812 <= reg5572[(1'h0):(1'h0)];
                    end
                  if (reg5758[(3'h4):(2'h3)])
                    begin
                      reg5813 <= $unsigned(reg5774);
                      reg5814 <= (reg5658[(2'h3):(2'h2)] ?
                          reg5646[(3'h6):(3'h5)] : $signed((reg5732[(4'he):(4'h8)] ?
                              (reg5706 ? reg5689 : reg5604) : reg5809)));
                      reg5815 <= reg5746[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg5813 <= reg5604;
                    end
                end
              else
                begin
                  if ((^~(((~|reg5709) ?
                      $unsigned(reg5662) : (!forvar5547)) != (~&(forvar5610 ?
                      reg5614 : reg5586)))))
                    begin
                      reg5811 <= {reg5637};
                      reg5812 <= (($signed($unsigned(reg5765)) * ($unsigned(reg5796) - (|(8'hb3)))) & (reg5738 ?
                          reg5652 : forvar5657));
                    end
                  else
                    begin
                      reg5811 <= reg5707;
                    end
                end
            end
          reg5816 <= reg5794[(2'h2):(2'h2)];
        end
      if (($signed(reg5732) ? reg5648[(4'he):(1'h0)] : forvar5575))
        begin
          if ((reg5634 ?
              reg5545 : $unsigned(($unsigned(forvar5761) && {reg5659}))))
            begin
              if (($signed($signed((reg5671 ?
                  reg5534 : forvar5655))) <= (((-forvar5558) <<< ((8'haf) ?
                  reg5650 : reg5655)) || (reg5625 ?
                  $signed(forvar5709) : (reg5716 >> reg5565)))))
                begin
                  if ($signed(reg5784[(2'h3):(1'h1)]))
                    begin
                      reg5817 <= (~|forvar5680[(1'h1):(1'h0)]);
                      reg5818 <= $signed(forvar5620[(2'h2):(1'h0)]);
                      reg5819 <= $unsigned({($unsigned(forvar5751) << forvar5683[(4'h8):(4'h8)])});
                    end
                  else
                    begin
                      reg5817 <= (((^~(&reg5775)) < reg5609) & (((reg5676 ?
                              reg5529 : reg5579) ?
                          $signed((8'hae)) : $signed(reg5539)) <<< (wire5513 >>> {(8'hb3)})));
                      reg5818 <= $unsigned((({reg5576} >= (reg5700 || forvar5673)) | $unsigned($signed(reg5521))));
                      reg5819 <= $signed({{$unsigned(forvar5670)}});
                      reg5820 <= $unsigned(reg5705);
                    end
                  reg5821 <= {((+(reg5591 ?
                          (8'ha8) : reg5714)) >> (~^(wire5513 ?
                          reg5728 : reg5798)))};
                  reg5822 <= $unsigned(forvar5610[(2'h3):(1'h0)]);
                  for (forvar5823 = (1'h0); (forvar5823 < (2'h2)); forvar5823 = (forvar5823 + (1'h1)))
                    begin
                      reg5824 <= (reg5687[(3'h5):(2'h2)] ?
                          (^((reg5590 ?
                              forvar5605 : forvar5594) || (-forvar5593))) : ((((8'ha9) <= forvar5537) ^ (wire5641 > reg5607)) | (forvar5773 ?
                              (-(8'h9e)) : (&forvar5675))));
                      reg5825 <= ({$unsigned((reg5651 ? reg5696 : reg5687))} ?
                          $unsigned($signed((reg5746 ^ forvar5718))) : $unsigned((^forvar5543[(2'h3):(1'h1)])));
                    end
                end
              else
                begin
                  for (forvar5817 = (1'h0); (forvar5817 < (2'h3)); forvar5817 = (forvar5817 + (1'h1)))
                    begin
                      reg5818 <= reg5738[(4'ha):(1'h1)];
                    end
                end
              for (forvar5826 = (1'h0); (forvar5826 < (2'h2)); forvar5826 = (forvar5826 + (1'h1)))
                begin
                  for (forvar5827 = (1'h0); (forvar5827 < (1'h0)); forvar5827 = (forvar5827 + (1'h1)))
                    begin
                      reg5828 <= $signed($unsigned(reg5607[(4'h9):(2'h2)]));
                    end
                end
              if ((($unsigned((8'hb6)) ?
                  (&reg5547[(3'h5):(3'h4)]) : $signed(forvar5587[(1'h0):(1'h0)])) ^ reg5814))
                begin
                  if (((((^forvar5680) ?
                          (reg5537 >>> reg5652) : $signed(reg5639)) ?
                      ((~|reg5800) ?
                          $unsigned(reg5532) : (~^forvar5518)) : ((reg5798 ?
                          reg5645 : (8'ha6)) ^ reg5807)) < reg5563[(4'hb):(3'h5)]))
                    begin
                      reg5829 <= (+reg5599[(2'h3):(1'h0)]);
                    end
                  else
                    begin
                      reg5829 <= (forvar5763 ?
                          ((8'ha7) ?
                              reg5541 : forvar5700[(1'h1):(1'h0)]) : $unsigned($unsigned((~&forvar5791))));
                      reg5830 <= (|(+(8'haa)));
                      reg5831 <= (forvar5655 > reg5820[(4'h9):(2'h2)]);
                    end
                  for (forvar5832 = (1'h0); (forvar5832 < (1'h0)); forvar5832 = (forvar5832 + (1'h1)))
                    begin
                      reg5833 <= ((~&reg5541) <<< $signed(((+reg5558) ?
                          (forvar5680 ? reg5708 : reg5765) : (reg5523 ?
                              reg5737 : reg5750))));
                      reg5834 <= $signed(reg5729[(3'h6):(3'h5)]);
                      reg5835 <= $unsigned(reg5670[(4'h9):(4'h8)]);
                    end
                end
              else
                begin
                  for (forvar5829 = (1'h0); (forvar5829 < (2'h2)); forvar5829 = (forvar5829 + (1'h1)))
                    begin
                      reg5830 <= (((+(forvar5746 ?
                          reg5528 : forvar5601)) - (forvar5721 ?
                          reg5516 : reg5678[(1'h0):(1'h0)])) >>> forvar5771[(1'h0):(1'h0)]);
                      reg5831 <= (8'ha3);
                    end
                end
            end
          else
            begin
              if ($unsigned(reg5591[(1'h0):(1'h0)]))
                begin
                  if ($signed($signed(($unsigned(forvar5578) < (forvar5665 ?
                      reg5678 : reg5624)))))
                    begin
                      reg5817 <= (^~$unsigned((~^(forvar5673 == reg5626))));
                      reg5818 <= ($signed(reg5614[(2'h3):(1'h1)]) != $unsigned(reg5677));
                      reg5819 <= forvar5671[(4'h8):(1'h0)];
                    end
                  else
                    begin
                      reg5817 <= $signed(((8'hb9) ?
                          reg5803 : ({forvar5538} << reg5685)));
                      reg5818 <= (^~(((reg5623 ?
                          reg5784 : (8'ha3)) >>> (forvar5675 ?
                          reg5720 : reg5552)) >> (-reg5798[(4'he):(3'h6)])));
                      reg5819 <= ((!$unsigned((reg5695 ?
                              forvar5601 : (8'hb1)))) ?
                          forvar5580 : ((reg5679 <= forvar5618) || forvar5620));
                      reg5820 <= {((^~(&reg5690)) && (reg5630[(4'h8):(3'h4)] >= (reg5534 ?
                              reg5720 : reg5828)))};
                    end
                  if (reg5675[(1'h0):(1'h0)])
                    begin
                      reg5821 <= reg5635;
                      reg5822 <= ($signed((forvar5756 < (forvar5519 >= (8'hb7)))) || {(8'hb9)});
                    end
                  else
                    begin
                      reg5821 <= forvar5601[(4'h8):(2'h3)];
                      reg5822 <= {$unsigned(((reg5539 ?
                              reg5821 : reg5765) | reg5566))};
                      reg5823 <= (forvar5611 ?
                          (~^reg5711[(3'h4):(1'h0)]) : forvar5658[(2'h2):(1'h0)]);
                      reg5824 <= reg5678[(3'h4):(1'h1)];
                    end
                  reg5825 <= $unsigned(((^~forvar5564[(1'h1):(1'h1)]) >> reg5728));
                  reg5826 <= reg5651;
                end
              else
                begin
                  reg5817 <= ((~&(reg5548[(2'h3):(2'h3)] ?
                          (&reg5697) : reg5630)) ?
                      (^~$unsigned((reg5678 ?
                          forvar5529 : reg5824))) : (reg5680[(4'hd):(2'h2)] ?
                          reg5654[(2'h3):(1'h0)] : {((8'hac) ?
                                  reg5597 : reg5616)}));
                  if (forvar5543[(2'h2):(1'h0)])
                    begin
                      reg5818 <= reg5622[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg5818 <= ($unsigned((|(|reg5658))) < ((forvar5756 ?
                              $signed(forvar5549) : reg5797) ?
                          ((forvar5527 ~^ reg5732) != $signed(reg5679)) : $unsigned($unsigned(forvar5652))));
                      reg5819 <= $signed(((~(reg5599 + reg5681)) | $signed((forvar5692 ?
                          reg5833 : forvar5658))));
                    end
                  for (forvar5820 = (1'h0); (forvar5820 < (2'h2)); forvar5820 = (forvar5820 + (1'h1)))
                    begin
                      reg5821 <= reg5593;
                      reg5822 <= $unsigned((~^reg5731));
                      reg5823 <= {($signed(reg5663[(3'h6):(2'h2)]) ^ $signed({reg5547}))};
                    end
                end
            end
          for (forvar5836 = (1'h0); (forvar5836 < (2'h2)); forvar5836 = (forvar5836 + (1'h1)))
            begin
              reg5837 <= reg5796;
            end
          if (({$unsigned(reg5647)} ? reg5524 : $signed((^~$signed(reg5516)))))
            begin
              reg5838 <= $unsigned(({$signed(forvar5699)} != forvar5700[(2'h2):(1'h0)]));
              for (forvar5839 = (1'h0); (forvar5839 < (2'h3)); forvar5839 = (forvar5839 + (1'h1)))
                begin
                  for (forvar5840 = (1'h0); (forvar5840 < (1'h0)); forvar5840 = (forvar5840 + (1'h1)))
                    begin
                      reg5841 <= (reg5570[(1'h0):(1'h0)] ?
                          $unsigned($unsigned({forvar5629})) : reg5626);
                      reg5842 <= ((|reg5776[(1'h0):(1'h0)]) ?
                          ((~(8'ha7)) & (^forvar5540)) : (reg5654[(4'hb):(3'h7)] * ($unsigned(forvar5733) + reg5753[(2'h2):(1'h0)])));
                    end
                  for (forvar5843 = (1'h0); (forvar5843 < (2'h3)); forvar5843 = (forvar5843 + (1'h1)))
                    begin
                      reg5844 <= $signed($unsigned(reg5556[(4'hd):(2'h3)]));
                      reg5845 <= $signed((^(reg5736[(3'h4):(2'h3)] ?
                          (reg5758 ? reg5560 : forvar5684) : forvar5547)));
                      reg5846 <= $unsigned($unsigned((+(^~forvar5629))));
                    end
                  reg5847 <= $unsigned(reg5819[(4'hd):(2'h3)]);
                  for (forvar5848 = (1'h0); (forvar5848 < (1'h0)); forvar5848 = (forvar5848 + (1'h1)))
                    begin
                      reg5849 <= $unsigned((~|reg5824[(3'h4):(1'h0)]));
                      reg5850 <= {forvar5662};
                      reg5851 <= (($unsigned((~&reg5621)) ^~ {(reg5536 >= forvar5610)}) ?
                          ($unsigned($unsigned(reg5609)) * ($unsigned((8'hac)) ?
                              $signed(reg5784) : reg5526[(3'h7):(3'h7)])) : reg5754[(1'h0):(1'h0)]);
                    end
                end
              reg5852 <= $signed($signed($signed(forvar5763[(2'h2):(1'h0)])));
              for (forvar5853 = (1'h0); (forvar5853 < (1'h0)); forvar5853 = (forvar5853 + (1'h1)))
                begin
                  for (forvar5854 = (1'h0); (forvar5854 < (2'h2)); forvar5854 = (forvar5854 + (1'h1)))
                    begin
                      reg5855 <= reg5699;
                      reg5856 <= (^{((~^forvar5738) ?
                              $signed(reg5540) : (^reg5726))});
                    end
                  for (forvar5857 = (1'h0); (forvar5857 < (1'h1)); forvar5857 = (forvar5857 + (1'h1)))
                    begin
                      reg5858 <= $signed(forvar5801[(2'h3):(1'h0)]);
                      reg5859 <= (-$signed(forvar5687));
                      reg5860 <= reg5751[(2'h2):(2'h2)];
                      reg5861 <= (|reg5576);
                    end
                end
            end
          else
            begin
              reg5838 <= (reg5604 ? (8'h9c) : $unsigned(reg5675));
              if ((~&((+(^~reg5524)) < $signed(reg5684[(1'h1):(1'h0)]))))
                begin
                  if ((^(-(8'haa))))
                    begin
                      reg5839 <= reg5796;
                      reg5840 <= ($signed({$signed(reg5649)}) < forvar5789);
                      reg5841 <= ($unsigned(reg5861) ?
                          reg5706 : (-reg5520[(4'hc):(4'ha)]));
                    end
                  else
                    begin
                      reg5839 <= (reg5577[(4'hd):(1'h0)] || $signed($signed((~reg5781))));
                      reg5840 <= ($signed(forvar5590) > (reg5673[(1'h1):(1'h1)] ?
                          reg5835 : ({reg5600} ?
                              (forvar5658 >> (8'hb7)) : reg5788[(4'h9):(2'h2)])));
                    end
                  if ($signed({((wire5515 ?
                          reg5582 : reg5753) || $signed(reg5758))}))
                    begin
                      reg5842 <= {$unsigned(($signed(reg5745) ?
                              (|reg5737) : $unsigned(wire5512)))};
                      reg5843 <= {reg5518[(3'h4):(2'h3)]};
                      reg5844 <= $signed($signed(reg5577));
                      reg5845 <= {reg5678[(2'h2):(1'h1)]};
                    end
                  else
                    begin
                      reg5842 <= (!reg5590[(1'h1):(1'h1)]);
                      reg5843 <= (reg5660 ?
                          $signed(reg5592[(3'h4):(1'h1)]) : reg5557);
                      reg5844 <= reg5834[(5'h10):(4'he)];
                    end
                end
              else
                begin
                  for (forvar5839 = (1'h0); (forvar5839 < (2'h2)); forvar5839 = (forvar5839 + (1'h1)))
                    begin
                      reg5840 <= forvar5683;
                      reg5841 <= $signed($unsigned({reg5607[(4'h9):(2'h2)]}));
                      reg5842 <= ((reg5597 <<< reg5716[(4'h8):(3'h4)]) == reg5714);
                    end
                  reg5843 <= $unsigned($signed($unsigned(reg5807[(3'h4):(3'h4)])));
                end
              for (forvar5846 = (1'h0); (forvar5846 < (1'h0)); forvar5846 = (forvar5846 + (1'h1)))
                begin
                  for (forvar5847 = (1'h0); (forvar5847 < (1'h0)); forvar5847 = (forvar5847 + (1'h1)))
                    begin
                      reg5848 <= ((~&(8'haf)) && (+forvar5827));
                    end
                end
            end
          reg5862 <= {(reg5570 ~^ (&$signed(reg5612)))};
        end
      else
        begin
          for (forvar5817 = (1'h0); (forvar5817 < (1'h1)); forvar5817 = (forvar5817 + (1'h1)))
            begin
              for (forvar5818 = (1'h0); (forvar5818 < (1'h0)); forvar5818 = (forvar5818 + (1'h1)))
                begin
                  for (forvar5819 = (1'h0); (forvar5819 < (2'h2)); forvar5819 = (forvar5819 + (1'h1)))
                    begin
                      reg5820 <= forvar5817;
                    end
                  if ((-(^~{(^reg5522)})))
                    begin
                      reg5821 <= forvar5684[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg5821 <= forvar5575[(3'h5):(1'h1)];
                      reg5822 <= (((&$unsigned((8'hb4))) ?
                              reg5614[(3'h6):(3'h4)] : (8'hb1)) ?
                          ($unsigned(forvar5687) ^ {$unsigned(forvar5777)}) : (^$unsigned(reg5852[(3'h5):(3'h4)])));
                      reg5823 <= (forvar5789[(1'h0):(1'h0)] == $signed({forvar5677}));
                    end
                  if ($unsigned({(!$unsigned(forvar5780))}))
                    begin
                      reg5824 <= $unsigned(({forvar5658[(2'h2):(2'h2)]} ^ $signed($signed((8'ha1)))));
                      reg5825 <= (reg5648 >= (^~(reg5798 > $signed(reg5537))));
                    end
                  else
                    begin
                      reg5824 <= $signed(reg5598[(2'h3):(2'h3)]);
                      reg5825 <= (((8'hb4) == reg5548[(1'h0):(1'h0)]) || reg5559[(1'h1):(1'h0)]);
                      reg5826 <= (((~&$unsigned((8'ha6))) ?
                          $unsigned(reg5675) : (reg5850[(2'h3):(1'h0)] >>> (reg5567 ^~ reg5737))) ^ reg5532[(2'h3):(1'h1)]);
                      reg5827 <= (((((8'ha7) ? (8'hb5) : forvar5739) ?
                          forvar5773 : (8'ha5)) >>> forvar5529) == {(reg5722[(2'h2):(1'h1)] ?
                              reg5700 : (reg5754 + reg5579))});
                    end
                end
              for (forvar5828 = (1'h0); (forvar5828 < (2'h2)); forvar5828 = (forvar5828 + (1'h1)))
                begin
                  reg5829 <= $unsigned(reg5749[(2'h3):(1'h1)]);
                  for (forvar5830 = (1'h0); (forvar5830 < (2'h2)); forvar5830 = (forvar5830 + (1'h1)))
                    begin
                      reg5831 <= forvar5790;
                    end
                  reg5832 <= reg5565[(2'h3):(2'h3)];
                end
            end
          reg5833 <= $signed($signed(((forvar5791 ?
              (8'ha4) : reg5823) != $unsigned(reg5725))));
        end
    end
  assign wire5863 = $unsigned((~$signed((reg5720 != forvar5670))));
  assign wire5864 = (+(!(!$unsigned((8'ha2)))));
  assign wire5865 = ((|((|forvar5538) && reg5732[(4'hc):(2'h2)])) ?
                        reg5670 : {$signed((reg5645 < reg5745))});
  assign wire5866 = reg5570;
  always
    @(posedge clk) begin
      for (forvar5867 = (1'h0); (forvar5867 < (2'h2)); forvar5867 = (forvar5867 + (1'h1)))
        begin
          if (reg5679[(4'he):(4'he)])
            begin
              for (forvar5868 = (1'h0); (forvar5868 < (2'h2)); forvar5868 = (forvar5868 + (1'h1)))
                begin
                  reg5869 <= $signed((reg5746 ?
                      ((-reg5527) ~^ forvar5549[(2'h3):(1'h0)]) : reg5713[(3'h4):(1'h0)]));
                  if ((^($signed((reg5671 ?
                      reg5851 : reg5720)) - (reg5827[(3'h4):(1'h1)] ^ (!reg5651)))))
                    begin
                      reg5870 <= {((8'hb2) ?
                              (forvar5679 == forvar5772[(1'h0):(1'h0)]) : forvar5588)};
                      reg5871 <= (-$unsigned($unsigned(reg5570)));
                    end
                  else
                    begin
                      reg5870 <= (|forvar5790[(3'h6):(2'h3)]);
                      reg5871 <= forvar5540[(4'h8):(2'h3)];
                    end
                  if (((reg5524[(1'h0):(1'h0)] ?
                      reg5847[(2'h3):(2'h3)] : $signed((wire5515 > reg5816))) == ($unsigned((!reg5719)) ?
                      reg5802[(3'h7):(1'h0)] : (~&(8'h9d)))))
                    begin
                      reg5872 <= forvar5542;
                      reg5873 <= (~^(~reg5531));
                      reg5874 <= ((((reg5674 * reg5812) ?
                              reg5681[(1'h1):(1'h0)] : (reg5723 ?
                                  reg5647 : reg5572)) ?
                          ((+reg5753) ?
                              (-reg5743) : $unsigned(reg5703)) : (~$unsigned(reg5784))) ^ {reg5715[(1'h0):(1'h0)]});
                    end
                  else
                    begin
                      reg5872 <= reg5606[(4'ha):(4'h9)];
                      reg5873 <= forvar5529;
                      reg5874 <= ($signed((+forvar5636)) >> forvar5540[(2'h3):(2'h3)]);
                      reg5875 <= {((((8'hb2) ?
                                  reg5539 : forvar5738) >= reg5654[(3'h6):(1'h1)]) ?
                              {(forvar5594 <<< reg5640)} : (8'hb3))};
                    end
                  if ($unsigned($unsigned(reg5608[(1'h0):(1'h0)])))
                    begin
                      reg5876 <= $signed((!(|$unsigned(forvar5716))));
                      reg5877 <= (~&({(forvar5832 * forvar5610)} ^~ $signed(reg5738)));
                    end
                  else
                    begin
                      reg5876 <= $signed($unsigned((^~reg5536)));
                    end
                end
            end
          else
            begin
              for (forvar5868 = (1'h0); (forvar5868 < (1'h0)); forvar5868 = (forvar5868 + (1'h1)))
                begin
                  reg5869 <= (forvar5840[(3'h7):(2'h2)] < ((|reg5520) ?
                      reg5648 : forvar5658));
                  for (forvar5870 = (1'h0); (forvar5870 < (2'h2)); forvar5870 = (forvar5870 + (1'h1)))
                    begin
                      reg5871 <= (^~((~{(8'ha4)}) && reg5876));
                      reg5872 <= $unsigned(($unsigned(reg5528[(3'h4):(2'h3)]) >= reg5810[(1'h1):(1'h0)]));
                      reg5873 <= ($unsigned($signed((~&reg5729))) ?
                          (~|($signed(reg5589) - (reg5812 ^ reg5676))) : ($unsigned((forvar5555 >>> reg5644)) ?
                              (reg5776[(3'h5):(3'h4)] ?
                                  (reg5630 | reg5810) : $signed(reg5576)) : $unsigned($unsigned(reg5574))));
                    end
                  reg5874 <= {reg5597};
                  for (forvar5875 = (1'h0); (forvar5875 < (2'h2)); forvar5875 = (forvar5875 + (1'h1)))
                    begin
                      reg5876 <= reg5541;
                      reg5877 <= ({((reg5675 | forvar5538) ?
                                  (~&reg5551) : $unsigned(reg5524))} ?
                          $unsigned(($unsigned((8'h9f)) ?
                              $unsigned(wire5865) : $unsigned(forvar5848))) : $unsigned((&forvar5627)));
                      reg5878 <= (&$unsigned($signed(forvar5671)));
                      reg5879 <= (8'hb2);
                    end
                end
              if ((~^reg5810))
                begin
                  reg5880 <= ({reg5576} ?
                      ($unsigned($unsigned(reg5602)) ?
                          reg5878 : {(|forvar5829)}) : $signed(reg5858));
                  for (forvar5881 = (1'h0); (forvar5881 < (2'h2)); forvar5881 = (forvar5881 + (1'h1)))
                    begin
                      reg5882 <= reg5559;
                    end
                end
              else
                begin
                  if ((((~&(reg5562 ? (8'hb0) : reg5741)) ?
                      (^(~forvar5791)) : {(reg5698 <= reg5553)}) <<< $signed((&$signed(reg5824)))))
                    begin
                      reg5880 <= (^$unsigned((!$signed(reg5872))));
                    end
                  else
                    begin
                      reg5880 <= $signed(reg5808);
                    end
                  for (forvar5881 = (1'h0); (forvar5881 < (2'h3)); forvar5881 = (forvar5881 + (1'h1)))
                    begin
                      reg5882 <= forvar5671[(3'h5):(2'h2)];
                      reg5883 <= (reg5850[(3'h4):(2'h3)] ^~ $signed((forvar5613[(3'h6):(1'h1)] ?
                          (forvar5881 >= forvar5668) : forvar5756[(4'hb):(4'h9)])));
                      reg5884 <= (+reg5734);
                      reg5885 <= forvar5542;
                    end
                  for (forvar5886 = (1'h0); (forvar5886 < (2'h3)); forvar5886 = (forvar5886 + (1'h1)))
                    begin
                      reg5887 <= $unsigned((8'ha7));
                      reg5888 <= reg5633[(3'h7):(1'h1)];
                      reg5889 <= $unsigned((((wire5515 <= (8'hac)) ?
                          (8'hba) : (reg5870 ?
                              (8'hb7) : reg5806)) >> {$unsigned((8'ha7))}));
                    end
                end
            end
        end
      for (forvar5890 = (1'h0); (forvar5890 < (2'h2)); forvar5890 = (forvar5890 + (1'h1)))
        begin
          for (forvar5891 = (1'h0); (forvar5891 < (2'h2)); forvar5891 = (forvar5891 + (1'h1)))
            begin
              if ($signed($signed(reg5732)))
                begin
                  for (forvar5892 = (1'h0); (forvar5892 < (1'h1)); forvar5892 = (forvar5892 + (1'h1)))
                    begin
                      reg5893 <= {($unsigned(reg5840) > $signed({forvar5542}))};
                      reg5894 <= reg5760[(2'h3):(2'h2)];
                      reg5895 <= ({((reg5594 ?
                                  reg5812 : reg5802) >= (^~forvar5662))} ?
                          (forvar5647[(5'h10):(1'h1)] && ($unsigned(reg5552) ?
                              (!reg5845) : (&forvar5771))) : (8'hb1));
                    end
                end
              else
                begin
                  for (forvar5892 = (1'h0); (forvar5892 < (1'h0)); forvar5892 = (forvar5892 + (1'h1)))
                    begin
                      reg5893 <= reg5729;
                      reg5894 <= reg5536[(1'h1):(1'h0)];
                    end
                  if ({reg5615[(3'h6):(3'h5)]})
                    begin
                      reg5895 <= (+reg5583);
                      reg5896 <= reg5831;
                      reg5897 <= $signed(reg5602[(4'ha):(4'h8)]);
                    end
                  else
                    begin
                      reg5895 <= ((-(reg5590 ?
                          reg5630 : (!reg5544))) * {{(reg5765 > reg5558)}});
                    end
                  for (forvar5898 = (1'h0); (forvar5898 < (1'h1)); forvar5898 = (forvar5898 + (1'h1)))
                    begin
                      reg5899 <= (reg5661 != ($signed(((8'h9e) ~^ forvar5898)) ?
                          reg5874[(1'h1):(1'h1)] : (8'hb8)));
                      reg5900 <= wire5865;
                      reg5901 <= $signed($unsigned((forvar5699 >> {(8'h9d)})));
                    end
                end
              for (forvar5902 = (1'h0); (forvar5902 < (2'h2)); forvar5902 = (forvar5902 + (1'h1)))
                begin
                  for (forvar5903 = (1'h0); (forvar5903 < (2'h2)); forvar5903 = (forvar5903 + (1'h1)))
                    begin
                      reg5904 <= reg5565[(2'h2):(2'h2)];
                      reg5905 <= (($signed(forvar5790) < ((+reg5747) ?
                          forvar5627 : (&(8'ha5)))) <= reg5626);
                      reg5906 <= ((|$unsigned($unsigned(forvar5657))) <<< reg5756[(3'h5):(1'h1)]);
                      reg5907 <= (~^(((~|reg5784) ?
                          {reg5806} : reg5576[(2'h3):(1'h0)]) + reg5706));
                    end
                  reg5908 <= reg5893;
                  for (forvar5909 = (1'h0); (forvar5909 < (2'h2)); forvar5909 = (forvar5909 + (1'h1)))
                    begin
                      reg5910 <= forvar5663[(1'h0):(1'h0)];
                      reg5911 <= {((&$unsigned(reg5737)) ?
                              $unsigned(((8'haa) ^~ reg5726)) : $unsigned((forvar5768 == reg5633)))};
                      reg5912 <= ($signed(reg5766) ?
                          reg5521[(4'h9):(4'h8)] : reg5678[(4'h9):(1'h1)]);
                      reg5913 <= forvar5558;
                    end
                  for (forvar5914 = (1'h0); (forvar5914 < (2'h3)); forvar5914 = (forvar5914 + (1'h1)))
                    begin
                      reg5915 <= ({($unsigned(reg5840) || (reg5796 <= reg5689))} ?
                          (&(-((8'hac) ?
                              reg5696 : reg5764))) : ($signed({(8'ha0)}) & {reg5781[(2'h2):(1'h0)]}));
                    end
                end
              if (reg5719)
                begin
                  for (forvar5916 = (1'h0); (forvar5916 < (1'h0)); forvar5916 = (forvar5916 + (1'h1)))
                    begin
                      reg5917 <= (reg5803 <<< (+(8'h9c)));
                      reg5918 <= (((~&(8'hb4)) ?
                          $signed((reg5676 && reg5647)) : ((^reg5598) ?
                              $unsigned(forvar5662) : reg5615)) > (forvar5785[(3'h4):(1'h0)] ?
                          reg5653 : ((reg5806 ?
                              forvar5629 : reg5694) == reg5820[(3'h4):(2'h2)])));
                    end
                  for (forvar5919 = (1'h0); (forvar5919 < (1'h0)); forvar5919 = (forvar5919 + (1'h1)))
                    begin
                      reg5920 <= (($unsigned((reg5848 ?
                          (8'hb2) : reg5574)) & (reg5792 ^~ (reg5717 != forvar5890))) ~^ $signed((~(forvar5594 ~^ forvar5699))));
                      reg5921 <= (($signed((forvar5588 >>> reg5527)) ?
                              $signed((forvar5677 == reg5888)) : $unsigned((~|reg5578))) ?
                          {wire5512} : forvar5687);
                      reg5922 <= ((~|reg5671[(4'ha):(2'h2)]) - (+reg5677[(1'h1):(1'h1)]));
                    end
                  reg5923 <= $unsigned($unsigned($signed((~|reg5562))));
                  for (forvar5924 = (1'h0); (forvar5924 < (1'h0)); forvar5924 = (forvar5924 + (1'h1)))
                    begin
                      reg5925 <= forvar5881[(3'h5):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar5916 = (1'h0); (forvar5916 < (1'h0)); forvar5916 = (forvar5916 + (1'h1)))
                    begin
                      reg5917 <= $unsigned((reg5555 < reg5579));
                    end
                  for (forvar5918 = (1'h0); (forvar5918 < (1'h1)); forvar5918 = (forvar5918 + (1'h1)))
                    begin
                      reg5919 <= forvar5854[(3'h4):(2'h3)];
                      reg5920 <= $unsigned($signed(reg5748[(3'h6):(3'h4)]));
                      reg5921 <= (^~((reg5837 >> (+(8'hac))) > ((reg5540 ?
                              reg5755 : reg5521) ?
                          (reg5586 ? reg5837 : reg5879) : (~&(8'hba)))));
                    end
                end
              reg5926 <= $signed(wire5866[(3'h5):(2'h2)]);
            end
          for (forvar5927 = (1'h0); (forvar5927 < (2'h3)); forvar5927 = (forvar5927 + (1'h1)))
            begin
              for (forvar5928 = (1'h0); (forvar5928 < (1'h1)); forvar5928 = (forvar5928 + (1'h1)))
                begin
                  for (forvar5929 = (1'h0); (forvar5929 < (2'h2)); forvar5929 = (forvar5929 + (1'h1)))
                    begin
                      reg5930 <= reg5537;
                      reg5931 <= ($unsigned((!(8'hb9))) < forvar5527);
                    end
                  if (reg5807)
                    begin
                      reg5932 <= forvar5739;
                    end
                  else
                    begin
                      reg5932 <= forvar5546;
                      reg5933 <= reg5820[(3'h6):(2'h2)];
                    end
                  for (forvar5934 = (1'h0); (forvar5934 < (2'h2)); forvar5934 = (forvar5934 + (1'h1)))
                    begin
                      reg5935 <= $signed((((~|reg5584) ? {reg5555} : reg5739) ?
                          ($unsigned(reg5841) | reg5660[(1'h1):(1'h0)]) : forvar5725));
                      reg5936 <= (reg5519 ^ $signed($signed((reg5694 <= forvar5819))));
                    end
                  reg5937 <= (forvar5791[(1'h0):(1'h0)] <<< $unsigned($signed($signed(reg5525))));
                end
              if (((!($signed(reg5654) ~^ reg5686)) ^ ((reg5679[(4'h8):(4'h8)] ~^ reg5921) || $unsigned(forvar5868[(4'hb):(4'h9)]))))
                begin
                  for (forvar5938 = (1'h0); (forvar5938 < (2'h3)); forvar5938 = (forvar5938 + (1'h1)))
                    begin
                      reg5939 <= $unsigned(reg5765[(3'h4):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar5938 = (1'h0); (forvar5938 < (1'h1)); forvar5938 = (forvar5938 + (1'h1)))
                    begin
                      reg5939 <= $unsigned((~^{$unsigned((8'hb0))}));
                      reg5940 <= wire5513;
                      reg5941 <= reg5539;
                    end
                  for (forvar5942 = (1'h0); (forvar5942 < (2'h3)); forvar5942 = (forvar5942 + (1'h1)))
                    begin
                      reg5943 <= (forvar5636[(1'h0):(1'h0)] >>> reg5873);
                      reg5944 <= $unsigned($signed($unsigned(reg5581[(3'h6):(3'h6)])));
                      reg5945 <= $unsigned($unsigned($unsigned((reg5581 ?
                          reg5882 : forvar5695))));
                    end
                  for (forvar5946 = (1'h0); (forvar5946 < (1'h1)); forvar5946 = (forvar5946 + (1'h1)))
                    begin
                      reg5947 <= (reg5549 ?
                          (((!reg5850) && {reg5684}) == reg5767[(3'h4):(2'h2)]) : {$signed(((8'ha1) <<< forvar5519))});
                      reg5948 <= ((^~$signed((8'had))) ?
                          reg5779 : $unsigned(((reg5540 ?
                              reg5819 : forvar5771) * (forvar5846 ?
                              reg5583 : reg5745))));
                      reg5949 <= ((~^(forvar5564[(2'h2):(1'h1)] && reg5703[(3'h5):(1'h1)])) ?
                          $signed(((forvar5683 ? forvar5549 : reg5912) ?
                              reg5603[(4'ha):(4'ha)] : reg5675)) : $unsigned((!(reg5616 | reg5677))));
                    end
                  for (forvar5950 = (1'h0); (forvar5950 < (2'h2)); forvar5950 = (forvar5950 + (1'h1)))
                    begin
                      reg5951 <= ((wire5515[(1'h0):(1'h0)] ?
                          (reg5738 ?
                              reg5930[(4'hf):(4'ha)] : (^~forvar5558)) : reg5746) && reg5654);
                    end
                end
              for (forvar5952 = (1'h0); (forvar5952 < (2'h3)); forvar5952 = (forvar5952 + (1'h1)))
                begin
                  if (((($unsigned(forvar5771) ?
                      $unsigned(wire5641) : $unsigned(forvar5650)) >>> {$signed(reg5856)}) >= (8'h9e)))
                    begin
                      reg5953 <= (reg5722 ?
                          reg5516 : (reg5538[(2'h2):(1'h1)] ?
                              (~(~|forvar5647)) : ((reg5802 ?
                                      reg5560 : reg5720) ?
                                  $unsigned((8'hb0)) : (+forvar5699))));
                    end
                  else
                    begin
                      reg5953 <= ($signed(($unsigned(reg5590) ~^ (&reg5612))) != $signed(($signed(reg5861) ?
                          ((8'ha3) == reg5741) : (reg5522 >= reg5844))));
                    end
                  if ($signed($signed((^~((8'ha7) ? forvar5817 : forvar5804)))))
                    begin
                      reg5954 <= reg5698[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg5954 <= $unsigned((((forvar5909 ? reg5516 : reg5591) ?
                          (~&reg5878) : (forvar5655 > reg5648)) || reg5882));
                      reg5955 <= forvar5589[(2'h3):(2'h2)];
                      reg5956 <= $signed(reg5541[(1'h0):(1'h0)]);
                    end
                end
            end
          for (forvar5957 = (1'h0); (forvar5957 < (1'h0)); forvar5957 = (forvar5957 + (1'h1)))
            begin
              if ((((~&(~&reg5931)) ?
                  ($signed(reg5543) ^~ {reg5637}) : reg5662) <<< (~^$unsigned(((8'ha4) ?
                  reg5534 : (8'hb4))))))
                begin
                  if ($signed(((~|(^forvar5547)) + ((forvar5739 ?
                      reg5551 : reg5633) | reg5861[(3'h6):(3'h6)]))))
                    begin
                      reg5958 <= $unsigned((reg5832[(4'hb):(1'h1)] & reg5555));
                      reg5959 <= reg5889;
                    end
                  else
                    begin
                      reg5958 <= $signed(wire5864);
                      reg5959 <= (8'ha5);
                      reg5960 <= ((reg5945[(4'ha):(3'h4)] ?
                          forvar5768[(3'h6):(3'h6)] : (8'h9f)) >>> reg5846);
                    end
                  for (forvar5961 = (1'h0); (forvar5961 < (1'h0)); forvar5961 = (forvar5961 + (1'h1)))
                    begin
                      reg5962 <= (!reg5956[(4'hc):(3'h4)]);
                      reg5963 <= forvar5675[(2'h2):(1'h1)];
                    end
                  for (forvar5964 = (1'h0); (forvar5964 < (1'h1)); forvar5964 = (forvar5964 + (1'h1)))
                    begin
                      reg5965 <= {{forvar5618[(3'h7):(3'h7)]}};
                      reg5966 <= $signed(reg5941);
                      reg5967 <= reg5540[(4'hc):(3'h4)];
                    end
                end
              else
                begin
                  reg5958 <= reg5562;
                  reg5959 <= ((-reg5614[(2'h3):(1'h1)]) ?
                      $signed($unsigned(((8'ha8) * forvar5870))) : (|(forvar5957 ?
                          $signed(forvar5832) : reg5682[(2'h2):(2'h2)])));
                end
              for (forvar5968 = (1'h0); (forvar5968 < (2'h3)); forvar5968 = (forvar5968 + (1'h1)))
                begin
                  for (forvar5969 = (1'h0); (forvar5969 < (2'h2)); forvar5969 = (forvar5969 + (1'h1)))
                    begin
                      reg5970 <= forvar5924[(1'h1):(1'h1)];
                    end
                  for (forvar5971 = (1'h0); (forvar5971 < (1'h1)); forvar5971 = (forvar5971 + (1'h1)))
                    begin
                      reg5972 <= $unsigned((($signed(forvar5611) ?
                          (reg5809 ? reg5843 : reg5633) : (wire5866 ?
                              (8'hac) : reg5875)) & (~^(reg5555 ?
                          reg5615 : forvar5646))));
                      reg5973 <= (&reg5749);
                      reg5974 <= $unsigned(reg5845[(3'h5):(3'h4)]);
                    end
                  for (forvar5975 = (1'h0); (forvar5975 < (1'h0)); forvar5975 = (forvar5975 + (1'h1)))
                    begin
                      reg5976 <= forvar5909;
                      reg5977 <= reg5630[(3'h4):(2'h3)];
                      reg5978 <= reg5705;
                    end
                  reg5979 <= (&$signed($unsigned((8'hb6))));
                end
              for (forvar5980 = (1'h0); (forvar5980 < (1'h0)); forvar5980 = (forvar5980 + (1'h1)))
                begin
                  for (forvar5981 = (1'h0); (forvar5981 < (1'h1)); forvar5981 = (forvar5981 + (1'h1)))
                    begin
                      reg5982 <= reg5787[(4'ha):(4'h9)];
                      reg5983 <= (~{(8'ha3)});
                      reg5984 <= {reg5596};
                    end
                  reg5985 <= $unsigned((reg5705[(1'h1):(1'h1)] ?
                      ((forvar5964 ?
                          reg5956 : forvar5898) * reg5960[(3'h7):(1'h0)]) : {$unsigned(forvar5892)}));
                  if ((+(((|reg5672) ?
                      (forvar5680 ?
                          reg5797 : reg5710) : reg5687) | (|(^(8'h9f))))))
                    begin
                      reg5986 <= (~^reg5519[(2'h3):(2'h3)]);
                      reg5987 <= (8'hb1);
                      reg5988 <= (forvar5751[(1'h0):(1'h0)] != $signed($unsigned(reg5630)));
                    end
                  else
                    begin
                      reg5986 <= $signed((reg5656[(1'h1):(1'h0)] << ((^reg5917) - $unsigned(reg5745))));
                      reg5987 <= ({forvar5870[(3'h4):(1'h0)]} ?
                          $signed(reg5630) : $signed(((-reg5676) != $unsigned(forvar5975))));
                      reg5988 <= (((^(forvar5717 ? reg5793 : reg5676)) ?
                          ({reg5676} | $signed(forvar5886)) : {(^reg5524)}) - (~^(~$signed(reg5782))));
                    end
                end
              if (reg5935)
                begin
                  reg5989 <= ((($signed(forvar5517) ?
                      forvar5646[(4'hb):(1'h1)] : (8'h9e)) ^ reg5747) < $signed(reg5874[(3'h7):(2'h3)]));
                end
              else
                begin
                  for (forvar5989 = (1'h0); (forvar5989 < (2'h2)); forvar5989 = (forvar5989 + (1'h1)))
                    begin
                      reg5990 <= $unsigned((forvar5927[(1'h1):(1'h0)] >> (8'hba)));
                      reg5991 <= $unsigned(reg5825[(4'ha):(3'h4)]);
                    end
                  for (forvar5992 = (1'h0); (forvar5992 < (2'h3)); forvar5992 = (forvar5992 + (1'h1)))
                    begin
                      reg5993 <= $signed($unsigned($unsigned($signed(reg5932))));
                      reg5994 <= reg5526[(2'h2):(1'h1)];
                    end
                end
            end
          for (forvar5995 = (1'h0); (forvar5995 < (2'h2)); forvar5995 = (forvar5995 + (1'h1)))
            begin
              reg5996 <= reg5523;
              for (forvar5997 = (1'h0); (forvar5997 < (1'h1)); forvar5997 = (forvar5997 + (1'h1)))
                begin
                  reg5998 <= (8'hb8);
                end
              reg5999 <= $unsigned($unsigned($signed(forvar5677[(3'h7):(1'h1)])));
            end
        end
      for (forvar6000 = (1'h0); (forvar6000 < (2'h2)); forvar6000 = (forvar6000 + (1'h1)))
        begin
          for (forvar6001 = (1'h0); (forvar6001 < (2'h3)); forvar6001 = (forvar6001 + (1'h1)))
            begin
              if (reg5677)
                begin
                  for (forvar6002 = (1'h0); (forvar6002 < (1'h0)); forvar6002 = (forvar6002 + (1'h1)))
                    begin
                      reg6003 <= ($signed($unsigned($unsigned((8'ha0)))) * (~(forvar5518 + (forvar5820 << reg5734))));
                      reg6004 <= reg5598;
                      reg6005 <= ((-((reg5988 ?
                          forvar5929 : forvar5823) <= (forvar5590 ?
                          (8'ha2) : forvar5854))) > (forvar5848 ?
                          $signed((+reg5686)) : reg5796[(1'h1):(1'h1)]));
                    end
                  if (($unsigned((forvar5751 ~^ reg5544)) ?
                      (~&(8'hb9)) : (-$signed($signed((8'ha0))))))
                    begin
                      reg6006 <= (reg5729[(4'h8):(4'h8)] ^~ (reg5549[(3'h7):(1'h0)] ?
                          (~&$signed((8'hb0))) : reg5694));
                    end
                  else
                    begin
                      reg6006 <= $unsigned(($signed({reg5885}) ?
                          forvar5679 : $signed((~&reg5724))));
                      reg6007 <= $signed((($unsigned(wire5864) ~^ reg5812) ?
                          ($signed(reg5901) | forvar6001) : {$unsigned(reg5566)}));
                      reg6008 <= $signed((((^~forvar5679) | (&(8'had))) && reg5897[(1'h0):(1'h0)]));
                    end
                  if (((($signed(forvar5752) ? $signed(forvar5721) : (8'hb9)) ?
                          ((reg5529 ?
                              forvar5971 : reg5669) != (forvar5552 ^ reg5559)) : reg5684) ?
                      reg5583 : (~^(^$signed(reg5662)))))
                    begin
                      reg6009 <= forvar6001[(2'h2):(1'h0)];
                      reg6010 <= (~|$unsigned({(^reg5977)}));
                    end
                  else
                    begin
                      reg6009 <= $unsigned($unsigned($signed((reg5654 ^ reg5721))));
                      reg6010 <= reg5883[(3'h4):(3'h4)];
                    end
                  for (forvar6011 = (1'h0); (forvar6011 < (2'h2)); forvar6011 = (forvar6011 + (1'h1)))
                    begin
                      reg6012 <= reg5572[(3'h4):(1'h0)];
                    end
                end
              else
                begin
                  reg6002 <= reg5675;
                  if ($unsigned($unsigned($signed({reg5912}))))
                    begin
                      reg6003 <= reg5962;
                      reg6004 <= (($signed((reg5614 ? reg5676 : reg5527)) ?
                          $unsigned($unsigned(reg5829)) : ((8'hab) != $unsigned(forvar6001))) >> ($signed((reg5949 * forvar5843)) == (^((8'h9e) || reg5547))));
                    end
                  else
                    begin
                      reg6003 <= (&(($signed(forvar5843) ?
                              (-reg5539) : (~&reg5758)) ?
                          $unsigned($signed(reg5831)) : forvar5898[(3'h4):(2'h2)]));
                      reg6004 <= ((((8'ha6) ?
                              reg5920 : $unsigned(reg5750)) | $unsigned($signed(reg5693))) ?
                          (~^(^(reg5841 ?
                              reg5682 : forvar5848))) : $signed({$signed(reg5778)}));
                      reg6005 <= reg5551;
                      reg6006 <= (8'had);
                    end
                  reg6007 <= $unsigned(reg5798[(4'hc):(4'hc)]);
                end
              reg6013 <= $unsigned(reg5876[(3'h7):(2'h2)]);
            end
          reg6014 <= $signed(($unsigned((^~reg5825)) ?
              ($signed(forvar5700) + (!forvar5762)) : $signed($unsigned(reg5783))));
        end
    end
endmodule