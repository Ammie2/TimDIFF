module inverter (
    input in,
    output out
);
    assign out = ~in;
endmodule