(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h1335):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hf):(1'h0)] wire4;
  input wire [(4'hd):(1'h0)] wire3;
  input wire [(4'hf):(1'h0)] wire2;
  input wire [(4'h8):(1'h0)] wire1;
  input wire signed [(4'hb):(1'h0)] wire0;
  reg signed [(3'h6):(1'h0)] reg1902 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1901 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1900 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1899 = (1'h0);
  reg [(3'h6):(1'h0)] reg1898 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1897 = (1'h0);
  reg [(2'h3):(1'h0)] reg1896 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1895 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1894 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1893 = (1'h0);
  reg [(3'h5):(1'h0)] reg1892 = (1'h0);
  reg [(4'hb):(1'h0)] reg1891 = (1'h0);
  reg [(3'h6):(1'h0)] reg1890 = (1'h0);
  reg [(3'h6):(1'h0)] reg1889 = (1'h0);
  reg [(4'h9):(1'h0)] reg1888 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1887 = (1'h0);
  reg [(3'h4):(1'h0)] reg1886 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1885 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1884 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1883 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1882 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1881 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1880 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1879 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1878 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1843 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1841 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1839 = (1'h0);
  reg [(3'h7):(1'h0)] reg1877 = (1'h0);
  reg [(4'hb):(1'h0)] reg1876 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1875 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1874 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1873 = (1'h0);
  reg [(4'h9):(1'h0)] reg1872 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1871 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1870 = (1'h0);
  reg [(3'h7):(1'h0)] reg1869 = (1'h0);
  reg [(4'ha):(1'h0)] reg1868 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1867 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1866 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1865 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1864 = (1'h0);
  reg [(4'hb):(1'h0)] reg1863 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1862 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1861 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1860 = (1'h0);
  reg [(4'he):(1'h0)] forvar1859 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1858 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1857 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1856 = (1'h0);
  reg [(2'h2):(1'h0)] reg1855 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1852 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1850 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1854 = (1'h0);
  reg [(4'hf):(1'h0)] reg1853 = (1'h0);
  reg [(4'h8):(1'h0)] reg1852 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1851 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1850 = (1'h0);
  reg [(2'h3):(1'h0)] reg1849 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1848 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1847 = (1'h0);
  reg [(4'hb):(1'h0)] reg1846 = (1'h0);
  reg [(4'he):(1'h0)] reg1845 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1844 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1843 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1842 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1841 = (1'h0);
  reg [(4'he):(1'h0)] reg1840 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1839 = (1'h0);
  reg [(4'hb):(1'h0)] reg1838 = (1'h0);
  reg [(2'h2):(1'h0)] reg1837 = (1'h0);
  reg [(4'ha):(1'h0)] reg1836 = (1'h0);
  reg [(4'hf):(1'h0)] reg1835 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1834 = (1'h0);
  reg [(2'h2):(1'h0)] reg1833 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1832 = (1'h0);
  reg [(2'h3):(1'h0)] reg1831 = (1'h0);
  reg [(4'hc):(1'h0)] reg1830 = (1'h0);
  reg [(4'he):(1'h0)] reg1829 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1828 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1827 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1826 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1825 = (1'h0);
  reg [(4'hb):(1'h0)] reg1824 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1823 = (1'h0);
  reg [(3'h6):(1'h0)] reg1822 = (1'h0);
  reg [(3'h7):(1'h0)] reg1821 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1820 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1819 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1818 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1817 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1816 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1815 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1814 = (1'h0);
  reg [(4'h8):(1'h0)] reg1813 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1812 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1811 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1810 = (1'h0);
  wire [(4'hf):(1'h0)] wire1809;
  wire [(3'h5):(1'h0)] wire1808;
  wire signed [(3'h6):(1'h0)] wire1807;
  reg signed [(4'hc):(1'h0)] forvar1782 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1787 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1785 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1770 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1769 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1768 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1766 = (1'h0);
  reg [(3'h4):(1'h0)] reg1765 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1762 = (1'h0);
  reg [(4'h9):(1'h0)] reg1760 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1806 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1805 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1804 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1803 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1802 = (1'h0);
  reg [(2'h2):(1'h0)] reg1801 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1800 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1799 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1798 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1797 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1791 = (1'h0);
  reg [(4'hc):(1'h0)] reg1796 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1795 = (1'h0);
  reg [(4'h8):(1'h0)] reg1794 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1793 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1792 = (1'h0);
  reg [(5'h10):(1'h0)] reg1791 = (1'h0);
  reg [(4'hb):(1'h0)] reg1790 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1783 = (1'h0);
  reg [(3'h4):(1'h0)] reg1789 = (1'h0);
  reg [(4'hf):(1'h0)] reg1788 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1787 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1786 = (1'h0);
  reg [(4'hc):(1'h0)] reg1785 = (1'h0);
  reg [(3'h7):(1'h0)] reg1784 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1783 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1782 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1776 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1781 = (1'h0);
  reg [(2'h2):(1'h0)] reg1780 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1779 = (1'h0);
  reg [(3'h5):(1'h0)] reg1778 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1775 = (1'h0);
  reg [(2'h2):(1'h0)] reg1774 = (1'h0);
  reg [(2'h2):(1'h0)] reg1777 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1776 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1775 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1774 = (1'h0);
  reg [(5'h10):(1'h0)] reg1773 = (1'h0);
  reg [(4'ha):(1'h0)] reg1772 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1771 = (1'h0);
  reg [(4'h9):(1'h0)] reg1770 = (1'h0);
  reg [(4'ha):(1'h0)] reg1769 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1768 = (1'h0);
  reg [(4'hb):(1'h0)] reg1767 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1766 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1765 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1761 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1764 = (1'h0);
  reg [(3'h7):(1'h0)] reg1763 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1762 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1761 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1760 = (1'h0);
  reg [(4'h9):(1'h0)] reg1752 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1749 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1748 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1739 = (1'h0);
  reg [(4'he):(1'h0)] reg1736 = (1'h0);
  reg [(3'h7):(1'h0)] reg1759 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1758 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1757 = (1'h0);
  reg [(4'h9):(1'h0)] reg1756 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1755 = (1'h0);
  reg [(4'hd):(1'h0)] reg1754 = (1'h0);
  reg [(2'h2):(1'h0)] reg1753 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1752 = (1'h0);
  reg [(4'h8):(1'h0)] reg1751 = (1'h0);
  reg [(4'hb):(1'h0)] reg1750 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1749 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1744 = (1'h0);
  reg [(4'hb):(1'h0)] reg1748 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1747 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1746 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1745 = (1'h0);
  reg [(5'h10):(1'h0)] reg1744 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1743 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1742 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1741 = (1'h0);
  reg [(4'hc):(1'h0)] reg1740 = (1'h0);
  reg [(3'h7):(1'h0)] reg1739 = (1'h0);
  reg [(4'h9):(1'h0)] reg1738 = (1'h0);
  reg [(4'hf):(1'h0)] reg1737 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1736 = (1'h0);
  reg [(2'h2):(1'h0)] reg1735 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1734 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1733 = (1'h0);
  reg [(4'he):(1'h0)] reg1732 = (1'h0);
  reg [(4'hb):(1'h0)] reg1731 = (1'h0);
  reg [(4'ha):(1'h0)] reg1730 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1729 = (1'h0);
  reg [(3'h4):(1'h0)] reg1728 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1727 = (1'h0);
  reg [(3'h6):(1'h0)] reg1726 = (1'h0);
  reg [(3'h6):(1'h0)] reg1725 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1724 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1723 = (1'h0);
  reg [(3'h6):(1'h0)] reg1722 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1721 = (1'h0);
  reg [(4'he):(1'h0)] reg1720 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1719 = (1'h0);
  reg [(4'hb):(1'h0)] reg1718 = (1'h0);
  reg [(4'hf):(1'h0)] reg1717 = (1'h0);
  reg [(4'hd):(1'h0)] reg1716 = (1'h0);
  reg [(3'h5):(1'h0)] reg1715 = (1'h0);
  reg [(4'hb):(1'h0)] reg1714 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1713 = (1'h0);
  reg [(4'he):(1'h0)] forvar1712 = (1'h0);
  reg [(2'h3):(1'h0)] reg1711 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1710 = (1'h0);
  reg [(4'h8):(1'h0)] reg1709 = (1'h0);
  reg [(3'h7):(1'h0)] reg1708 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1705 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1704 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1707 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1706 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1705 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1704 = (1'h0);
  reg [(4'h8):(1'h0)] reg1703 = (1'h0);
  reg [(4'hc):(1'h0)] reg1702 = (1'h0);
  reg [(4'he):(1'h0)] reg1701 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1700 = (1'h0);
  reg [(4'hc):(1'h0)] reg1699 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1698 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1697 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1696 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1695 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1694 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1693 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1692 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1685 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1683 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1682 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1691 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1690 = (1'h0);
  reg [(3'h6):(1'h0)] reg1689 = (1'h0);
  reg [(4'hc):(1'h0)] reg1688 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1687 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1686 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1685 = (1'h0);
  reg [(4'h8):(1'h0)] reg1684 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1683 = (1'h0);
  reg [(2'h3):(1'h0)] reg1682 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1681 = (1'h0);
  reg [(4'h9):(1'h0)] reg1680 = (1'h0);
  reg [(4'hc):(1'h0)] reg1679 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1676 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1671 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1669 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1668 = (1'h0);
  reg [(4'h8):(1'h0)] reg1667 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1664 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1666 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1660 = (1'h0);
  reg [(4'he):(1'h0)] reg1678 = (1'h0);
  reg [(3'h6):(1'h0)] reg1677 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1676 = (1'h0);
  reg [(4'hf):(1'h0)] reg1675 = (1'h0);
  reg [(4'h9):(1'h0)] reg1674 = (1'h0);
  reg [(4'h9):(1'h0)] reg1673 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1672 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1671 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1670 = (1'h0);
  reg [(4'hd):(1'h0)] reg1669 = (1'h0);
  reg [(4'h8):(1'h0)] reg1668 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1667 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1666 = (1'h0);
  reg [(2'h3):(1'h0)] reg1665 = (1'h0);
  reg [(2'h3):(1'h0)] reg1664 = (1'h0);
  reg [(4'ha):(1'h0)] reg1663 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1662 = (1'h0);
  reg [(3'h6):(1'h0)] reg1661 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1660 = (1'h0);
  reg [(4'hc):(1'h0)] reg1659 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1657 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1655 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1653 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1651 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1646 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1642 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1641 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1639 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1636 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1633 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1658 = (1'h0);
  reg [(2'h2):(1'h0)] reg1657 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1656 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1655 = (1'h0);
  reg [(4'h8):(1'h0)] reg1654 = (1'h0);
  reg [(4'hc):(1'h0)] reg1653 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1652 = (1'h0);
  reg [(4'hb):(1'h0)] reg1651 = (1'h0);
  reg [(3'h7):(1'h0)] reg1650 = (1'h0);
  reg [(3'h4):(1'h0)] reg1649 = (1'h0);
  reg [(5'h10):(1'h0)] reg1648 = (1'h0);
  reg [(4'hb):(1'h0)] reg1647 = (1'h0);
  reg [(2'h3):(1'h0)] reg1646 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1645 = (1'h0);
  reg [(4'he):(1'h0)] reg1644 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1643 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1642 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1641 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1640 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1639 = (1'h0);
  reg [(4'hc):(1'h0)] reg1638 = (1'h0);
  reg [(3'h7):(1'h0)] reg1637 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1636 = (1'h0);
  reg [(3'h7):(1'h0)] reg1635 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1634 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1633 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1632 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1631 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1630 = (1'h0);
  reg [(3'h4):(1'h0)] reg1627 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1626 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1625 = (1'h0);
  reg [(2'h2):(1'h0)] reg1624 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1623 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1631 = (1'h0);
  reg [(4'h9):(1'h0)] reg1630 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1629 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1628 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1627 = (1'h0);
  reg [(3'h5):(1'h0)] reg1626 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1625 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1624 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1623 = (1'h0);
  reg [(4'h9):(1'h0)] reg1622 = (1'h0);
  reg [(2'h3):(1'h0)] reg1621 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1620 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1619 = (1'h0);
  wire [(4'ha):(1'h0)] wire1618;
  reg [(4'hb):(1'h0)] reg1617 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1616 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1615 = (1'h0);
  reg [(4'hb):(1'h0)] reg1614 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1613 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1612 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1611 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1610 = (1'h0);
  reg [(3'h7):(1'h0)] reg1609 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1608 = (1'h0);
  reg [(4'he):(1'h0)] reg1607 = (1'h0);
  reg [(4'hb):(1'h0)] reg1606 = (1'h0);
  reg [(2'h2):(1'h0)] reg1605 = (1'h0);
  reg [(4'he):(1'h0)] reg1604 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1603 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1602 = (1'h0);
  reg [(4'hc):(1'h0)] reg1601 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1600 = (1'h0);
  reg [(4'hc):(1'h0)] reg1599 = (1'h0);
  reg [(4'he):(1'h0)] forvar1598 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1597 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1596 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1595 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1594 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1592 = (1'h0);
  reg [(2'h2):(1'h0)] reg1593 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1592 = (1'h0);
  reg [(3'h6):(1'h0)] reg1591 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1590 = (1'h0);
  reg [(4'hb):(1'h0)] reg1589 = (1'h0);
  reg [(5'h10):(1'h0)] reg1588 = (1'h0);
  reg [(3'h6):(1'h0)] reg1587 = (1'h0);
  reg [(4'h8):(1'h0)] reg1586 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1585 = (1'h0);
  reg [(4'he):(1'h0)] reg1584 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1583 = (1'h0);
  reg [(3'h4):(1'h0)] reg1567 = (1'h0);
  reg [(4'hd):(1'h0)] reg1582 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1581 = (1'h0);
  reg [(4'hf):(1'h0)] reg1580 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1577 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1572 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1560 = (1'h0);
  reg [(4'hf):(1'h0)] reg1558 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1571 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1579 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1578 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1577 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1576 = (1'h0);
  reg [(4'hc):(1'h0)] reg1575 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1574 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1573 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1572 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1571 = (1'h0);
  reg [(4'he):(1'h0)] reg1570 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1569 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1568 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1567 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1566 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1565 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1564 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1563 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1562 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1561 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1560 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1559 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1558 = (1'h0);
  reg [(4'he):(1'h0)] reg1557 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1556 = (1'h0);
  reg [(4'h8):(1'h0)] reg1555 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1554 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1550 = (1'h0);
  reg [(4'ha):(1'h0)] reg1548 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1546 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1545 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1543 = (1'h0);
  reg [(4'h9):(1'h0)] reg1541 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1540 = (1'h0);
  reg [(4'hd):(1'h0)] reg1538 = (1'h0);
  reg [(4'ha):(1'h0)] reg1553 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1552 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1551 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1550 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1549 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1548 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1547 = (1'h0);
  reg [(3'h4):(1'h0)] reg1546 = (1'h0);
  reg [(4'hb):(1'h0)] reg1545 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1544 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1543 = (1'h0);
  reg [(4'he):(1'h0)] reg1542 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1541 = (1'h0);
  reg [(4'hf):(1'h0)] reg1540 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1539 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1538 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1537 = (1'h0);
  reg [(4'hf):(1'h0)] reg1536 = (1'h0);
  reg [(2'h3):(1'h0)] reg1535 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1534 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1533 = (1'h0);
  reg [(4'hd):(1'h0)] reg1532 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1531 = (1'h0);
  reg [(4'hc):(1'h0)] reg1531 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1530 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1529 = (1'h0);
  reg [(4'hb):(1'h0)] reg1528 = (1'h0);
  reg [(4'hf):(1'h0)] reg1527 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1526 = (1'h0);
  reg [(4'ha):(1'h0)] reg1525 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1524 = (1'h0);
  reg [(4'he):(1'h0)] reg1523 = (1'h0);
  reg [(4'ha):(1'h0)] reg1522 = (1'h0);
  reg [(3'h5):(1'h0)] reg1521 = (1'h0);
  reg [(4'hb):(1'h0)] reg1520 = (1'h0);
  reg [(4'hc):(1'h0)] reg1519 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1518 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1517 = (1'h0);
  reg [(3'h4):(1'h0)] reg1516 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1515 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1514 = (1'h0);
  reg [(4'hb):(1'h0)] reg1513 = (1'h0);
  reg [(3'h7):(1'h0)] reg1512 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1511 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1510 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1509 = (1'h0);
  reg [(4'hb):(1'h0)] reg1508 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1507 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1506 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1505 = (1'h0);
  reg [(4'ha):(1'h0)] reg1504 = (1'h0);
  reg [(4'hb):(1'h0)] reg1503 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1502 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1501 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1499 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1495 = (1'h0);
  reg [(4'h9):(1'h0)] reg1494 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1485 = (1'h0);
  reg [(2'h2):(1'h0)] reg1502 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1501 = (1'h0);
  reg [(3'h4):(1'h0)] reg1500 = (1'h0);
  reg [(4'hc):(1'h0)] reg1499 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1490 = (1'h0);
  reg [(2'h2):(1'h0)] reg1486 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1498 = (1'h0);
  reg [(2'h2):(1'h0)] reg1497 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1496 = (1'h0);
  reg [(2'h3):(1'h0)] reg1495 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1494 = (1'h0);
  reg [(3'h4):(1'h0)] reg1493 = (1'h0);
  reg [(3'h6):(1'h0)] reg1492 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1491 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1490 = (1'h0);
  reg [(4'he):(1'h0)] reg1489 = (1'h0);
  reg [(4'hb):(1'h0)] reg1488 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1487 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1486 = (1'h0);
  reg [(4'hc):(1'h0)] reg1485 = (1'h0);
  reg [(4'he):(1'h0)] reg1484 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1483 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1482 = (1'h0);
  reg [(4'hf):(1'h0)] reg1481 = (1'h0);
  reg [(4'hf):(1'h0)] reg1480 = (1'h0);
  reg [(4'hb):(1'h0)] reg1479 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1478 = (1'h0);
  reg [(2'h3):(1'h0)] reg1477 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1476 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1472 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1470 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1467 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1475 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1474 = (1'h0);
  reg [(4'h8):(1'h0)] reg1473 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1472 = (1'h0);
  reg [(2'h2):(1'h0)] reg1471 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1470 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1469 = (1'h0);
  reg [(4'hd):(1'h0)] reg1468 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1467 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1466 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1465 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1464 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1461 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1456 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1459 = (1'h0);
  reg [(2'h3):(1'h0)] reg1463 = (1'h0);
  reg [(4'hf):(1'h0)] reg1462 = (1'h0);
  reg [(4'hc):(1'h0)] reg1461 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1460 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1459 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1455 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1458 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1457 = (1'h0);
  reg [(2'h3):(1'h0)] reg1456 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1455 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1454 = (1'h0);
  wire [(4'ha):(1'h0)] wire1453;
  wire [(4'hc):(1'h0)] wire1295;
  wire signed [(4'hf):(1'h0)] wire6;
  wire [(5'h10):(1'h0)] wire5;
  wire signed [(5'h10):(1'h0)] wire1451;
  assign y = {reg1902,
                 forvar1901,
                 reg1900,
                 forvar1899,
                 reg1898,
                 reg1897,
                 reg1896,
                 forvar1895,
                 forvar1894,
                 reg1893,
                 reg1892,
                 reg1891,
                 reg1890,
                 reg1889,
                 reg1888,
                 reg1887,
                 reg1886,
                 forvar1885,
                 forvar1884,
                 forvar1883,
                 reg1882,
                 reg1881,
                 forvar1880,
                 forvar1879,
                 forvar1878,
                 forvar1843,
                 reg1841,
                 reg1839,
                 reg1877,
                 reg1876,
                 forvar1875,
                 reg1874,
                 forvar1873,
                 reg1872,
                 reg1871,
                 forvar1870,
                 reg1869,
                 reg1868,
                 reg1867,
                 reg1866,
                 reg1865,
                 forvar1864,
                 reg1863,
                 reg1862,
                 reg1861,
                 forvar1860,
                 forvar1859,
                 reg1858,
                 forvar1857,
                 reg1856,
                 reg1855,
                 forvar1852,
                 reg1850,
                 reg1854,
                 reg1853,
                 reg1852,
                 reg1851,
                 forvar1850,
                 reg1849,
                 reg1848,
                 reg1847,
                 reg1846,
                 reg1845,
                 reg1844,
                 reg1843,
                 reg1842,
                 forvar1841,
                 reg1840,
                 forvar1839,
                 reg1838,
                 reg1837,
                 reg1836,
                 reg1835,
                 reg1834,
                 reg1833,
                 forvar1832,
                 reg1831,
                 reg1830,
                 reg1829,
                 forvar1828,
                 forvar1827,
                 reg1826,
                 reg1825,
                 reg1824,
                 reg1823,
                 reg1822,
                 reg1821,
                 reg1820,
                 forvar1819,
                 reg1818,
                 reg1817,
                 reg1816,
                 reg1815,
                 reg1814,
                 reg1813,
                 forvar1812,
                 forvar1811,
                 forvar1810,
                 wire1809,
                 wire1808,
                 wire1807,
                 forvar1782,
                 reg1787,
                 forvar1785,
                 forvar1770,
                 forvar1769,
                 reg1768,
                 forvar1766,
                 reg1765,
                 forvar1762,
                 reg1760,
                 reg1806,
                 reg1805,
                 reg1804,
                 reg1803,
                 reg1802,
                 reg1801,
                 reg1800,
                 reg1799,
                 forvar1798,
                 forvar1797,
                 forvar1791,
                 reg1796,
                 reg1795,
                 reg1794,
                 reg1793,
                 reg1792,
                 reg1791,
                 reg1790,
                 forvar1783,
                 reg1789,
                 reg1788,
                 forvar1787,
                 reg1786,
                 reg1785,
                 reg1784,
                 reg1783,
                 reg1782,
                 forvar1776,
                 reg1781,
                 reg1780,
                 reg1779,
                 reg1778,
                 reg1775,
                 reg1774,
                 reg1777,
                 reg1776,
                 forvar1775,
                 forvar1774,
                 reg1773,
                 reg1772,
                 reg1771,
                 reg1770,
                 reg1769,
                 forvar1768,
                 reg1767,
                 reg1766,
                 forvar1765,
                 forvar1761,
                 reg1764,
                 reg1763,
                 reg1762,
                 reg1761,
                 forvar1760,
                 reg1752,
                 forvar1749,
                 forvar1748,
                 forvar1739,
                 reg1736,
                 reg1759,
                 forvar1758,
                 forvar1757,
                 reg1756,
                 forvar1755,
                 reg1754,
                 reg1753,
                 forvar1752,
                 reg1751,
                 reg1750,
                 reg1749,
                 forvar1744,
                 reg1748,
                 reg1747,
                 reg1746,
                 reg1745,
                 reg1744,
                 reg1743,
                 reg1742,
                 reg1741,
                 reg1740,
                 reg1739,
                 reg1738,
                 reg1737,
                 forvar1736,
                 reg1735,
                 forvar1734,
                 reg1733,
                 reg1732,
                 reg1731,
                 reg1730,
                 reg1729,
                 reg1728,
                 forvar1727,
                 reg1726,
                 reg1725,
                 reg1724,
                 reg1723,
                 reg1722,
                 forvar1721,
                 reg1720,
                 reg1719,
                 reg1718,
                 reg1717,
                 reg1716,
                 reg1715,
                 reg1714,
                 forvar1713,
                 forvar1712,
                 reg1711,
                 reg1710,
                 reg1709,
                 reg1708,
                 forvar1705,
                 reg1704,
                 reg1707,
                 reg1706,
                 reg1705,
                 forvar1704,
                 reg1703,
                 reg1702,
                 reg1701,
                 reg1700,
                 reg1699,
                 reg1698,
                 reg1697,
                 reg1696,
                 forvar1695,
                 forvar1694,
                 forvar1693,
                 reg1692,
                 forvar1685,
                 reg1683,
                 forvar1682,
                 reg1691,
                 reg1690,
                 reg1689,
                 reg1688,
                 reg1687,
                 reg1686,
                 reg1685,
                 reg1684,
                 forvar1683,
                 reg1682,
                 forvar1681,
                 reg1680,
                 reg1679,
                 forvar1676,
                 reg1671,
                 forvar1669,
                 forvar1668,
                 reg1667,
                 forvar1664,
                 reg1666,
                 forvar1660,
                 reg1678,
                 reg1677,
                 reg1676,
                 reg1675,
                 reg1674,
                 reg1673,
                 reg1672,
                 forvar1671,
                 reg1670,
                 reg1669,
                 reg1668,
                 forvar1667,
                 forvar1666,
                 reg1665,
                 reg1664,
                 reg1663,
                 forvar1662,
                 reg1661,
                 reg1660,
                 reg1659,
                 forvar1657,
                 reg1655,
                 forvar1653,
                 forvar1651,
                 forvar1646,
                 reg1642,
                 reg1641,
                 forvar1639,
                 reg1636,
                 reg1633,
                 forvar1629,
                 reg1658,
                 reg1657,
                 reg1656,
                 forvar1655,
                 reg1654,
                 reg1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 reg1647,
                 reg1646,
                 reg1645,
                 reg1644,
                 reg1643,
                 forvar1642,
                 forvar1641,
                 reg1640,
                 reg1639,
                 reg1638,
                 reg1637,
                 forvar1636,
                 reg1635,
                 reg1634,
                 forvar1633,
                 reg1632,
                 forvar1631,
                 forvar1630,
                 reg1627,
                 forvar1626,
                 reg1625,
                 reg1624,
                 forvar1623,
                 reg1631,
                 reg1630,
                 reg1629,
                 reg1628,
                 forvar1627,
                 reg1626,
                 forvar1625,
                 forvar1624,
                 reg1623,
                 reg1622,
                 reg1621,
                 reg1620,
                 forvar1619,
                 wire1618,
                 reg1617,
                 forvar1616,
                 reg1615,
                 reg1614,
                 forvar1613,
                 forvar1612,
                 reg1611,
                 reg1610,
                 reg1609,
                 forvar1608,
                 reg1607,
                 reg1606,
                 reg1605,
                 reg1604,
                 forvar1603,
                 reg1602,
                 reg1601,
                 forvar1600,
                 reg1599,
                 forvar1598,
                 forvar1597,
                 reg1596,
                 reg1595,
                 reg1594,
                 forvar1592,
                 reg1593,
                 reg1592,
                 reg1591,
                 forvar1590,
                 reg1589,
                 reg1588,
                 reg1587,
                 reg1586,
                 forvar1585,
                 reg1584,
                 forvar1583,
                 reg1567,
                 reg1582,
                 reg1581,
                 reg1580,
                 reg1577,
                 forvar1572,
                 forvar1560,
                 reg1558,
                 reg1571,
                 reg1579,
                 reg1578,
                 forvar1577,
                 reg1576,
                 reg1575,
                 reg1574,
                 reg1573,
                 reg1572,
                 forvar1571,
                 reg1570,
                 reg1569,
                 reg1568,
                 forvar1567,
                 reg1566,
                 reg1565,
                 reg1564,
                 reg1563,
                 reg1562,
                 reg1561,
                 reg1560,
                 forvar1559,
                 forvar1558,
                 reg1557,
                 reg1556,
                 reg1555,
                 forvar1554,
                 reg1550,
                 reg1548,
                 forvar1546,
                 forvar1545,
                 forvar1543,
                 reg1541,
                 forvar1540,
                 reg1538,
                 reg1553,
                 reg1552,
                 reg1551,
                 forvar1550,
                 reg1549,
                 forvar1548,
                 reg1547,
                 reg1546,
                 reg1545,
                 reg1544,
                 reg1543,
                 reg1542,
                 forvar1541,
                 reg1540,
                 reg1539,
                 forvar1538,
                 reg1537,
                 reg1536,
                 reg1535,
                 forvar1534,
                 forvar1533,
                 reg1532,
                 forvar1531,
                 reg1531,
                 reg1530,
                 forvar1529,
                 reg1528,
                 reg1527,
                 reg1526,
                 reg1525,
                 forvar1524,
                 reg1523,
                 reg1522,
                 reg1521,
                 reg1520,
                 reg1519,
                 forvar1518,
                 reg1517,
                 reg1516,
                 reg1515,
                 forvar1514,
                 reg1513,
                 reg1512,
                 reg1511,
                 forvar1510,
                 reg1509,
                 reg1508,
                 reg1507,
                 forvar1506,
                 reg1505,
                 reg1504,
                 reg1503,
                 forvar1502,
                 forvar1501,
                 forvar1499,
                 forvar1495,
                 reg1494,
                 forvar1485,
                 reg1502,
                 reg1501,
                 reg1500,
                 reg1499,
                 forvar1490,
                 reg1486,
                 reg1498,
                 reg1497,
                 reg1496,
                 reg1495,
                 forvar1494,
                 reg1493,
                 reg1492,
                 reg1491,
                 reg1490,
                 reg1489,
                 reg1488,
                 reg1487,
                 forvar1486,
                 reg1485,
                 reg1484,
                 forvar1483,
                 forvar1482,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1478,
                 reg1477,
                 forvar1476,
                 forvar1472,
                 reg1470,
                 forvar1467,
                 reg1475,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1471,
                 forvar1470,
                 reg1469,
                 reg1468,
                 reg1467,
                 reg1466,
                 reg1465,
                 reg1464,
                 forvar1461,
                 forvar1456,
                 reg1459,
                 reg1463,
                 reg1462,
                 reg1461,
                 reg1460,
                 forvar1459,
                 reg1455,
                 reg1458,
                 reg1457,
                 reg1456,
                 forvar1455,
                 forvar1454,
                 wire1453,
                 wire1295,
                 wire6,
                 wire5,
                 wire1451,
                 (1'h0)};
  assign wire5 = (wire2 || ($signed((wire0 <<< wire1)) ?
                     $signed(wire4) : $unsigned((~^wire1))));
  assign wire6 = wire1[(3'h4):(1'h1)];
  module7 modinst1296 (wire1295, clk, wire3, wire2, wire6, wire0, wire4);
  module1297 modinst1452 (.wire1299(wire1295), .wire1300(wire5), .wire1302(wire1), .clk(clk), .wire1301(wire6), .wire1298(wire4), .y(wire1451));
  assign wire1453 = ({{((8'hac) & wire5)}} == wire1451[(3'h7):(3'h6)]);
  always
    @(posedge clk) begin
      for (forvar1454 = (1'h0); (forvar1454 < (1'h0)); forvar1454 = (forvar1454 + (1'h1)))
        begin
          if (($signed($signed((~^wire3))) ?
              (8'hb0) : $unsigned($signed((~&wire1)))))
            begin
              if (((((wire6 ?
                  forvar1454 : wire1) | wire0) & wire1451[(3'h5):(1'h0)]) << wire3))
                begin
                  for (forvar1455 = (1'h0); (forvar1455 < (1'h0)); forvar1455 = (forvar1455 + (1'h1)))
                    begin
                      reg1456 <= wire3;
                      reg1457 <= ($signed(({forvar1454} & wire5)) ?
                          $unsigned(wire6[(4'ha):(3'h7)]) : (wire6 ?
                              {(~^reg1456)} : $unsigned({reg1456})));
                      reg1458 <= $unsigned({wire1[(1'h0):(1'h0)]});
                    end
                end
              else
                begin
                  if ((wire0[(1'h1):(1'h0)] || $unsigned(wire2[(4'hd):(3'h5)])))
                    begin
                      reg1455 <= (~|($unsigned($unsigned(wire1451)) ?
                          (~wire1295[(2'h2):(1'h0)]) : $unsigned((forvar1454 ^~ wire6))));
                      reg1456 <= forvar1455[(3'h5):(2'h3)];
                    end
                  else
                    begin
                      reg1455 <= (8'hb1);
                      reg1456 <= wire4[(4'he):(2'h3)];
                    end
                  if ($signed(reg1458))
                    begin
                      reg1457 <= wire4[(4'h8):(3'h5)];
                      reg1458 <= wire5[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg1457 <= $signed(($signed($signed((8'ha7))) && $unsigned({wire1451})));
                    end
                  for (forvar1459 = (1'h0); (forvar1459 < (2'h2)); forvar1459 = (forvar1459 + (1'h1)))
                    begin
                      reg1460 <= $unsigned(({(^~reg1457)} >= {(wire0 ?
                              reg1456 : reg1457)}));
                      reg1461 <= ((~(((8'hb8) >> forvar1455) - (forvar1454 >= wire1453))) || (($signed(wire1) ^ (reg1457 ?
                          (8'ha6) : forvar1459)) && (|wire2)));
                      reg1462 <= wire3;
                      reg1463 <= (reg1460[(2'h3):(1'h1)] == ({wire1451[(4'hc):(4'h8)]} && (-{forvar1459})));
                    end
                end
            end
          else
            begin
              if (($unsigned($signed((~^wire1))) ^~ reg1462[(4'hc):(4'hb)]))
                begin
                  if (wire1451[(5'h10):(4'hb)])
                    begin
                      reg1455 <= reg1463[(1'h0):(1'h0)];
                      reg1456 <= $signed((+$unsigned(reg1455)));
                      reg1457 <= reg1460;
                    end
                  else
                    begin
                      reg1455 <= (~(8'hb4));
                      reg1456 <= forvar1455[(3'h4):(1'h0)];
                    end
                  if ((~^wire0))
                    begin
                      reg1458 <= reg1458[(3'h4):(3'h4)];
                      reg1459 <= reg1463[(1'h1):(1'h1)];
                      reg1460 <= wire3;
                    end
                  else
                    begin
                      reg1458 <= wire1;
                      reg1459 <= (($unsigned((wire5 << wire2)) ?
                          ($signed(reg1458) ?
                              $signed((8'hb0)) : (wire6 ?
                                  reg1463 : wire1)) : (reg1458 ?
                              ((8'hac) >= wire5) : wire4)) ^~ $signed((reg1456 ?
                          (-wire1295) : $unsigned(reg1455))));
                    end
                end
              else
                begin
                  reg1455 <= (^~wire4[(4'hf):(4'h9)]);
                  for (forvar1456 = (1'h0); (forvar1456 < (1'h1)); forvar1456 = (forvar1456 + (1'h1)))
                    begin
                      reg1457 <= (({(wire2 && (8'hae))} ?
                              wire1[(2'h2):(1'h1)] : ($unsigned((8'hb9)) ?
                                  (wire5 ? wire3 : wire1295) : (~&reg1458))) ?
                          ($unsigned($unsigned(reg1458)) ?
                              $signed($unsigned(forvar1459)) : (reg1463[(1'h1):(1'h0)] ?
                                  (!wire2) : (8'ha6))) : (+({reg1456} ?
                              (!wire1451) : {wire3})));
                      reg1458 <= wire6;
                      reg1459 <= {($signed($unsigned(wire3)) * wire4[(3'h7):(2'h3)])};
                      reg1460 <= ((^(reg1463 & wire1453[(4'h9):(2'h3)])) ?
                          (&reg1456) : (reg1456[(1'h0):(1'h0)] & reg1463));
                    end
                  for (forvar1461 = (1'h0); (forvar1461 < (2'h2)); forvar1461 = (forvar1461 + (1'h1)))
                    begin
                      reg1462 <= wire0;
                      reg1463 <= reg1462;
                      reg1464 <= $unsigned($unsigned($unsigned(reg1459)));
                      reg1465 <= forvar1455;
                    end
                end
              reg1466 <= ((~{{(8'hb4)}}) ?
                  (~^(reg1457[(1'h0):(1'h0)] == $signed((8'hb2)))) : {$unsigned((^~wire4))});
              if (wire3)
                begin
                  if ($signed((!reg1457[(1'h1):(1'h1)])))
                    begin
                      reg1467 <= $signed(({(forvar1455 <<< reg1465)} << ((wire2 | reg1459) ?
                          $unsigned((8'ha7)) : (~wire1453))));
                      reg1468 <= forvar1459[(1'h1):(1'h0)];
                      reg1469 <= {reg1460};
                    end
                  else
                    begin
                      reg1467 <= (~$signed({((8'hb6) < wire1295)}));
                      reg1468 <= (|wire1295[(1'h1):(1'h0)]);
                      reg1469 <= (^~(((reg1461 ?
                              wire1453 : wire1453) ^~ (reg1460 <<< reg1464)) ?
                          ($signed((8'ha7)) + (wire5 ?
                              wire1453 : reg1460)) : $unsigned({reg1457})));
                    end
                  for (forvar1470 = (1'h0); (forvar1470 < (1'h1)); forvar1470 = (forvar1470 + (1'h1)))
                    begin
                      reg1471 <= (((~|{forvar1470}) ?
                          ((reg1459 ?
                              (8'hac) : wire1451) <= forvar1470) : (~^(^(8'ha7)))) | $unsigned(((forvar1459 - reg1456) != (8'hb5))));
                      reg1472 <= reg1471[(1'h0):(1'h0)];
                      reg1473 <= (|$signed($unsigned((!(8'hba)))));
                      reg1474 <= (|(($signed(wire6) <= (reg1459 < reg1463)) ?
                          forvar1459 : {$signed(reg1473)}));
                    end
                  reg1475 <= $unsigned($unsigned($unsigned(reg1465[(2'h2):(2'h2)])));
                end
              else
                begin
                  for (forvar1467 = (1'h0); (forvar1467 < (2'h2)); forvar1467 = (forvar1467 + (1'h1)))
                    begin
                      reg1468 <= ((reg1457[(2'h2):(1'h0)] | ($unsigned((8'ha1)) == (~wire1451))) ?
                          $unsigned(((wire2 && reg1467) ?
                              $unsigned(forvar1459) : reg1473)) : $signed($unsigned((~|reg1471))));
                      reg1469 <= ({forvar1459[(4'ha):(3'h4)]} ~^ wire4);
                      reg1470 <= ({forvar1454} + $signed(forvar1461[(3'h6):(3'h4)]));
                      reg1471 <= reg1474[(1'h0):(1'h0)];
                    end
                  for (forvar1472 = (1'h0); (forvar1472 < (2'h3)); forvar1472 = (forvar1472 + (1'h1)))
                    begin
                      reg1473 <= (~($unsigned(reg1472) * (wire2[(3'h6):(1'h0)] ?
                          {(8'ha4)} : (forvar1470 ? reg1461 : (8'h9c)))));
                      reg1474 <= reg1461[(1'h1):(1'h1)];
                      reg1475 <= (~&$unsigned(wire6));
                    end
                  for (forvar1476 = (1'h0); (forvar1476 < (1'h0)); forvar1476 = (forvar1476 + (1'h1)))
                    begin
                      reg1477 <= forvar1467;
                      reg1478 <= $signed({reg1458});
                      reg1479 <= $signed({forvar1459});
                      reg1480 <= ($unsigned(((8'hb8) != (wire1451 ?
                              (8'ha7) : reg1455))) ?
                          $signed(((wire0 | wire2) || (reg1478 <<< (8'ha3)))) : {(^~{reg1468})});
                    end
                  reg1481 <= forvar1454;
                end
            end
        end
      for (forvar1482 = (1'h0); (forvar1482 < (1'h0)); forvar1482 = (forvar1482 + (1'h1)))
        begin
          for (forvar1483 = (1'h0); (forvar1483 < (2'h3)); forvar1483 = (forvar1483 + (1'h1)))
            begin
              reg1484 <= ($signed(reg1469) ?
                  forvar1470[(1'h1):(1'h0)] : reg1474[(1'h0):(1'h0)]);
            end
          if ((!((+(&forvar1454)) | (reg1468 ?
              $unsigned(forvar1472) : {reg1466}))))
            begin
              reg1485 <= $unsigned($signed(wire6[(4'hb):(1'h1)]));
              if ({((+$unsigned(reg1478)) ? (^wire2) : reg1472)})
                begin
                  for (forvar1486 = (1'h0); (forvar1486 < (2'h2)); forvar1486 = (forvar1486 + (1'h1)))
                    begin
                      reg1487 <= $signed((-($signed(reg1480) ?
                          $unsigned(forvar1476) : (forvar1456 <<< reg1469))));
                      reg1488 <= (^~(|$signed((reg1461 * reg1464))));
                      reg1489 <= forvar1483;
                    end
                  if ((reg1467 ^~ ($signed((reg1467 ?
                      reg1466 : reg1459)) ^ reg1484)))
                    begin
                      reg1490 <= reg1467;
                    end
                  else
                    begin
                      reg1490 <= (^wire1);
                      reg1491 <= (({(reg1484 ? forvar1454 : wire5)} ?
                          (!$signed(reg1460)) : reg1480[(1'h1):(1'h1)]) ^ $signed(($unsigned((8'hb1)) ?
                          $unsigned((8'haa)) : (forvar1482 * reg1465))));
                      reg1492 <= $signed(wire1295);
                      reg1493 <= $signed(($signed($signed(forvar1476)) ?
                          {(reg1457 ?
                                  reg1468 : reg1487)} : $unsigned($unsigned(forvar1486))));
                    end
                  for (forvar1494 = (1'h0); (forvar1494 < (1'h1)); forvar1494 = (forvar1494 + (1'h1)))
                    begin
                      reg1495 <= (($signed($signed(reg1468)) ^ forvar1456) ?
                          (reg1455 ?
                              (+(8'ha1)) : ($signed(reg1459) >= (!reg1458))) : $signed((wire6[(4'hf):(1'h1)] ~^ (reg1477 ?
                              wire2 : forvar1467))));
                      reg1496 <= (reg1493[(1'h0):(1'h0)] ?
                          wire2 : (~|forvar1486));
                      reg1497 <= $signed(($signed(((8'h9f) ?
                              reg1461 : reg1460)) ?
                          ($signed(reg1473) ?
                              $signed(wire3) : (wire1 == forvar1454)) : $unsigned((reg1461 ?
                              reg1467 : reg1474))));
                      reg1498 <= wire4;
                    end
                end
              else
                begin
                  if ((8'h9d))
                    begin
                      reg1486 <= (8'hb8);
                      reg1487 <= wire2;
                      reg1488 <= $signed((^$unsigned((reg1481 << reg1492))));
                      reg1489 <= $unsigned((8'hac));
                    end
                  else
                    begin
                      reg1486 <= ($unsigned(((8'had) ^ $signed(forvar1472))) ?
                          $signed(((reg1495 != wire5) ?
                              (forvar1482 ?
                                  wire5 : wire5) : reg1481)) : reg1471);
                      reg1487 <= $unsigned({$signed($signed((8'haa)))});
                      reg1488 <= $signed(reg1497[(1'h1):(1'h1)]);
                    end
                  for (forvar1490 = (1'h0); (forvar1490 < (1'h1)); forvar1490 = (forvar1490 + (1'h1)))
                    begin
                      reg1491 <= {reg1475};
                      reg1492 <= $unsigned($signed(($signed(reg1470) ?
                          (~&reg1463) : {forvar1486})));
                      reg1493 <= $signed(reg1475[(2'h2):(1'h0)]);
                    end
                  for (forvar1494 = (1'h0); (forvar1494 < (2'h2)); forvar1494 = (forvar1494 + (1'h1)))
                    begin
                      reg1495 <= ($signed(((reg1492 | (8'hb2)) ?
                              (8'h9e) : (~&reg1484))) ?
                          reg1470[(1'h1):(1'h0)] : ((^(reg1485 & reg1477)) ?
                              reg1460 : reg1459[(2'h2):(1'h0)]));
                      reg1496 <= (!reg1484);
                      reg1497 <= ($signed($signed((reg1461 && reg1465))) == $unsigned(((~^reg1477) ^~ wire5)));
                    end
                  if (reg1462[(2'h3):(2'h3)])
                    begin
                      reg1498 <= $signed($signed(((wire2 ? wire5 : wire1295) ?
                          $unsigned(forvar1455) : (reg1458 <= reg1490))));
                      reg1499 <= ($signed((reg1459 + reg1492)) ^ reg1486[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1498 <= (~{(&$unsigned(reg1474))});
                      reg1499 <= wire1;
                      reg1500 <= {(|reg1484[(1'h0):(1'h0)])};
                      reg1501 <= ($signed(($signed(forvar1494) ?
                              forvar1476[(2'h2):(1'h1)] : $unsigned(reg1455))) ?
                          $signed((+$unsigned(reg1488))) : reg1499[(3'h7):(3'h4)]);
                    end
                end
              reg1502 <= {($signed($unsigned(reg1479)) ?
                      forvar1455 : {$unsigned(reg1461)})};
            end
          else
            begin
              for (forvar1485 = (1'h0); (forvar1485 < (1'h1)); forvar1485 = (forvar1485 + (1'h1)))
                begin
                  for (forvar1486 = (1'h0); (forvar1486 < (1'h0)); forvar1486 = (forvar1486 + (1'h1)))
                    begin
                      reg1487 <= reg1486[(2'h2):(2'h2)];
                      reg1488 <= (reg1465 - forvar1483[(2'h2):(1'h0)]);
                      reg1489 <= ($signed({$unsigned(reg1486)}) < ($signed($signed(reg1500)) - ($signed((8'hac)) | $unsigned(reg1477))));
                      reg1490 <= (wire4 ?
                          ($unsigned((|reg1488)) >>> ((reg1459 ?
                                  reg1491 : reg1466) ?
                              (reg1473 && reg1502) : reg1464)) : (reg1470[(3'h5):(3'h4)] || (+reg1462)));
                    end
                  if ((&(reg1466 != $signed($signed(wire0)))))
                    begin
                      reg1491 <= ($unsigned((wire1453[(1'h0):(1'h0)] <<< (^~reg1466))) ?
                          forvar1470[(3'h4):(1'h0)] : reg1491[(3'h6):(3'h5)]);
                      reg1492 <= (($unsigned($signed(reg1481)) & reg1480[(3'h5):(1'h1)]) ?
                          (8'hb2) : (reg1469 ? wire6 : forvar1494));
                      reg1493 <= forvar1470;
                      reg1494 <= (reg1472 ?
                          $unsigned($unsigned($signed((8'hb9)))) : $unsigned((|wire3[(4'hb):(3'h5)])));
                    end
                  else
                    begin
                      reg1491 <= $unsigned(($unsigned($signed(wire1453)) ?
                          ((forvar1459 ~^ wire1451) ?
                              (forvar1485 >> (8'hb0)) : $unsigned(reg1480)) : reg1456));
                    end
                  for (forvar1495 = (1'h0); (forvar1495 < (1'h1)); forvar1495 = (forvar1495 + (1'h1)))
                    begin
                      reg1496 <= (~reg1457[(4'h8):(2'h2)]);
                      reg1497 <= (-($unsigned(reg1493) ?
                          ((reg1463 >>> forvar1455) & (reg1502 || (8'ha7))) : (&(reg1464 || forvar1483))));
                      reg1498 <= reg1498[(3'h5):(3'h4)];
                    end
                end
              if ($unsigned(reg1472[(3'h4):(3'h4)]))
                begin
                  for (forvar1499 = (1'h0); (forvar1499 < (1'h0)); forvar1499 = (forvar1499 + (1'h1)))
                    begin
                      reg1500 <= ($signed(forvar1490) ^ ({reg1462} && ((reg1495 ?
                              wire1295 : reg1471) ?
                          (~&forvar1455) : forvar1482[(4'h9):(3'h7)])));
                    end
                end
              else
                begin
                  reg1499 <= {reg1472[(4'h8):(2'h2)]};
                end
              for (forvar1501 = (1'h0); (forvar1501 < (1'h1)); forvar1501 = (forvar1501 + (1'h1)))
                begin
                  for (forvar1502 = (1'h0); (forvar1502 < (2'h2)); forvar1502 = (forvar1502 + (1'h1)))
                    begin
                      reg1503 <= $signed({(reg1491 - (reg1478 ?
                              (8'ha0) : forvar1476))});
                      reg1504 <= forvar1501[(1'h1):(1'h0)];
                      reg1505 <= forvar1495;
                    end
                  for (forvar1506 = (1'h0); (forvar1506 < (2'h2)); forvar1506 = (forvar1506 + (1'h1)))
                    begin
                      reg1507 <= reg1474[(1'h0):(1'h0)];
                      reg1508 <= $unsigned((~reg1477[(1'h0):(1'h0)]));
                      reg1509 <= $unsigned(reg1459[(1'h0):(1'h0)]);
                    end
                  for (forvar1510 = (1'h0); (forvar1510 < (1'h1)); forvar1510 = (forvar1510 + (1'h1)))
                    begin
                      reg1511 <= $unsigned((^~(+reg1467)));
                      reg1512 <= forvar1510[(4'h9):(2'h2)];
                      reg1513 <= $signed(((8'h9f) ?
                          (reg1455[(4'hc):(3'h6)] ?
                              $signed(reg1499) : reg1466[(2'h3):(2'h2)]) : $unsigned(reg1485[(2'h2):(2'h2)])));
                    end
                  for (forvar1514 = (1'h0); (forvar1514 < (1'h0)); forvar1514 = (forvar1514 + (1'h1)))
                    begin
                      reg1515 <= forvar1490;
                      reg1516 <= (|$signed((+reg1484[(4'hb):(1'h1)])));
                      reg1517 <= reg1457;
                    end
                end
              for (forvar1518 = (1'h0); (forvar1518 < (2'h3)); forvar1518 = (forvar1518 + (1'h1)))
                begin
                  if (($signed({$signed(reg1505)}) + $unsigned(($unsigned((8'ha8)) ?
                      (reg1504 ? wire1453 : wire2) : $unsigned((8'haf))))))
                    begin
                      reg1519 <= $unsigned(forvar1494);
                      reg1520 <= reg1494[(3'h6):(3'h4)];
                      reg1521 <= $signed($unsigned((~&(reg1519 || reg1497))));
                      reg1522 <= $unsigned($unsigned(({forvar1514} << (reg1466 ?
                          forvar1482 : (8'hb1)))));
                    end
                  else
                    begin
                      reg1519 <= (reg1484 ?
                          $unsigned($unsigned({reg1521})) : reg1507);
                    end
                  reg1523 <= (reg1517[(4'ha):(2'h3)] >> (^$unsigned($signed(reg1455))));
                  for (forvar1524 = (1'h0); (forvar1524 < (1'h1)); forvar1524 = (forvar1524 + (1'h1)))
                    begin
                      reg1525 <= (8'ha7);
                    end
                  reg1526 <= $signed(reg1495);
                end
            end
          reg1527 <= $unsigned({$signed((reg1519 ? forvar1518 : (8'hba)))});
          reg1528 <= $unsigned($unsigned(($signed(wire2) == reg1512)));
        end
      for (forvar1529 = (1'h0); (forvar1529 < (2'h3)); forvar1529 = (forvar1529 + (1'h1)))
        begin
          reg1530 <= (forvar1483[(1'h0):(1'h0)] ?
              reg1465[(3'h6):(3'h6)] : wire1451[(4'h9):(4'h9)]);
        end
      if ((|(|{(forvar1506 << reg1501)})))
        begin
          reg1531 <= (8'h9c);
        end
      else
        begin
          for (forvar1531 = (1'h0); (forvar1531 < (1'h0)); forvar1531 = (forvar1531 + (1'h1)))
            begin
              reg1532 <= reg1456[(2'h3):(2'h2)];
            end
          if ({forvar1486[(4'ha):(3'h5)]})
            begin
              for (forvar1533 = (1'h0); (forvar1533 < (1'h0)); forvar1533 = (forvar1533 + (1'h1)))
                begin
                  for (forvar1534 = (1'h0); (forvar1534 < (1'h0)); forvar1534 = (forvar1534 + (1'h1)))
                    begin
                      reg1535 <= reg1461;
                      reg1536 <= {reg1499};
                      reg1537 <= ($unsigned({(&forvar1495)}) ?
                          ($signed(wire3) - ((reg1521 >> forvar1534) + $unsigned(reg1502))) : $unsigned((^(reg1470 ?
                              reg1484 : reg1468))));
                    end
                  for (forvar1538 = (1'h0); (forvar1538 < (1'h0)); forvar1538 = (forvar1538 + (1'h1)))
                    begin
                      reg1539 <= (forvar1494[(3'h6):(3'h5)] ~^ $unsigned((reg1480 ?
                          $unsigned(forvar1472) : {wire6})));
                      reg1540 <= wire0;
                    end
                  for (forvar1541 = (1'h0); (forvar1541 < (1'h1)); forvar1541 = (forvar1541 + (1'h1)))
                    begin
                      reg1542 <= (!$unsigned((forvar1461[(3'h5):(2'h2)] >>> (forvar1495 <= reg1522))));
                      reg1543 <= $signed($unsigned(((+reg1460) == (!wire5))));
                      reg1544 <= (^~$signed($signed($signed(wire1))));
                    end
                  if ((forvar1506 ?
                      forvar1482[(2'h2):(1'h1)] : $unsigned({(!reg1458)})))
                    begin
                      reg1545 <= reg1459[(3'h6):(3'h5)];
                      reg1546 <= (forvar1455[(1'h1):(1'h1)] & ((|reg1495[(2'h3):(2'h3)]) != $signed((reg1473 ?
                          reg1505 : forvar1461))));
                      reg1547 <= reg1488;
                    end
                  else
                    begin
                      reg1545 <= (&(|(|forvar1467)));
                      reg1546 <= (~((reg1463[(2'h2):(1'h0)] ?
                          $signed((8'hb1)) : (|(8'h9c))) != (reg1474[(1'h0):(1'h0)] << reg1542[(3'h6):(1'h0)])));
                      reg1547 <= reg1521;
                    end
                end
              for (forvar1548 = (1'h0); (forvar1548 < (1'h0)); forvar1548 = (forvar1548 + (1'h1)))
                begin
                  reg1549 <= $unsigned((^~{reg1494}));
                  for (forvar1550 = (1'h0); (forvar1550 < (2'h3)); forvar1550 = (forvar1550 + (1'h1)))
                    begin
                      reg1551 <= ((8'ha0) != reg1522[(4'ha):(2'h2)]);
                      reg1552 <= {(~$signed((8'ha5)))};
                    end
                end
              reg1553 <= $signed($unsigned(((reg1485 ~^ reg1484) ?
                  reg1552 : forvar1490[(1'h0):(1'h0)])));
            end
          else
            begin
              for (forvar1533 = (1'h0); (forvar1533 < (2'h3)); forvar1533 = (forvar1533 + (1'h1)))
                begin
                  for (forvar1534 = (1'h0); (forvar1534 < (2'h3)); forvar1534 = (forvar1534 + (1'h1)))
                    begin
                      reg1535 <= ($unsigned((reg1522 <<< (reg1517 <<< reg1486))) * $unsigned((reg1487 ?
                          ((8'hb4) >>> reg1471) : {reg1511})));
                    end
                  if (reg1461[(2'h3):(1'h0)])
                    begin
                      reg1536 <= $unsigned(((|(reg1494 ?
                          reg1546 : (8'hb4))) ^~ $signed((reg1478 ~^ reg1455))));
                    end
                  else
                    begin
                      reg1536 <= $signed((&wire1453[(1'h1):(1'h1)]));
                      reg1537 <= ((((forvar1506 ? forvar1502 : reg1461) ?
                          forvar1482 : (forvar1548 ?
                              reg1456 : forvar1456)) < (reg1499[(2'h2):(1'h0)] > (^~forvar1514))) || (((reg1488 ?
                          reg1460 : reg1464) << {reg1494}) == (^(reg1468 ?
                          reg1470 : reg1487))));
                      reg1538 <= ((wire4[(3'h6):(1'h1)] ?
                          (~|$unsigned(reg1531)) : (reg1545[(3'h6):(1'h0)] ?
                              forvar1502[(3'h7):(3'h7)] : forvar1482[(4'he):(4'hb)])) != reg1532);
                      reg1539 <= $signed($signed($unsigned($unsigned(reg1459))));
                    end
                  for (forvar1540 = (1'h0); (forvar1540 < (2'h2)); forvar1540 = (forvar1540 + (1'h1)))
                    begin
                      reg1541 <= ($unsigned(reg1503[(4'h8):(1'h0)]) ?
                          reg1460[(2'h2):(1'h0)] : $unsigned(({wire1} ?
                              $signed(forvar1531) : reg1501[(3'h6):(1'h0)])));
                      reg1542 <= ($unsigned($unsigned($unsigned(forvar1485))) == ($signed($signed(wire0)) ?
                          (reg1501[(4'ha):(1'h1)] >= (forvar1538 ?
                              forvar1541 : (8'hb7))) : (forvar1524[(4'h9):(3'h4)] ^~ ((8'ha4) >> (8'haf)))));
                    end
                  for (forvar1543 = (1'h0); (forvar1543 < (2'h2)); forvar1543 = (forvar1543 + (1'h1)))
                    begin
                      reg1544 <= $unsigned($signed(reg1467));
                    end
                end
              for (forvar1545 = (1'h0); (forvar1545 < (2'h3)); forvar1545 = (forvar1545 + (1'h1)))
                begin
                  for (forvar1546 = (1'h0); (forvar1546 < (2'h2)); forvar1546 = (forvar1546 + (1'h1)))
                    begin
                      reg1547 <= ({(8'ha2)} ?
                          $signed((~|(reg1520 && (8'ha9)))) : reg1492[(1'h1):(1'h1)]);
                      reg1548 <= $signed(reg1488[(3'h4):(3'h4)]);
                      reg1549 <= (~|reg1503[(1'h0):(1'h0)]);
                      reg1550 <= reg1492[(3'h5):(3'h4)];
                    end
                  if ((~reg1491))
                    begin
                      reg1551 <= {reg1497};
                      reg1552 <= reg1536;
                    end
                  else
                    begin
                      reg1551 <= forvar1518;
                    end
                  reg1553 <= (&reg1491[(4'ha):(4'h9)]);
                  for (forvar1554 = (1'h0); (forvar1554 < (2'h3)); forvar1554 = (forvar1554 + (1'h1)))
                    begin
                      reg1555 <= ($signed((((8'ha4) & (8'ha4)) || forvar1502[(4'h8):(1'h0)])) <= $signed(forvar1543[(2'h2):(2'h2)]));
                      reg1556 <= $unsigned(($unsigned(wire5[(4'hb):(4'ha)]) ?
                          (|$signed(reg1485)) : forvar1456[(1'h1):(1'h1)]));
                    end
                end
              reg1557 <= $signed(($signed((reg1458 ? forvar1533 : reg1494)) ?
                  ($unsigned(reg1523) ?
                      $unsigned((8'hb5)) : (~forvar1531)) : ((reg1499 ?
                          reg1492 : reg1495) ?
                      (reg1530 ? reg1489 : reg1464) : $unsigned((8'haa)))));
            end
          if (wire4[(2'h3):(2'h3)])
            begin
              for (forvar1558 = (1'h0); (forvar1558 < (2'h2)); forvar1558 = (forvar1558 + (1'h1)))
                begin
                  for (forvar1559 = (1'h0); (forvar1559 < (1'h0)); forvar1559 = (forvar1559 + (1'h1)))
                    begin
                      reg1560 <= reg1455;
                      reg1561 <= ($signed(reg1457[(3'h4):(3'h4)]) >>> ((reg1536[(4'h8):(2'h2)] ^ reg1543) ?
                          $unsigned($unsigned(reg1485)) : $signed((forvar1550 ?
                              forvar1490 : reg1457))));
                      reg1562 <= (($signed($signed(reg1507)) ?
                          $signed({forvar1495}) : wire0) < ($unsigned((reg1488 >> reg1556)) ?
                          (((8'hb5) >>> forvar1559) ^~ (&reg1488)) : ($signed(reg1467) >= (forvar1485 ?
                              reg1468 : forvar1506))));
                    end
                  if (reg1550[(2'h2):(1'h1)])
                    begin
                      reg1563 <= forvar1546[(2'h2):(1'h0)];
                      reg1564 <= (($unsigned((reg1525 ? forvar1546 : reg1513)) ?
                              (~|$signed(forvar1455)) : (~|(reg1472 > wire4))) ?
                          ($signed(forvar1524[(4'h8):(3'h4)]) << reg1493) : forvar1510[(3'h4):(1'h0)]);
                      reg1565 <= ($signed(($signed(forvar1490) ?
                              $unsigned(reg1496) : forvar1501)) ?
                          $signed((8'haf)) : (~|reg1489));
                      reg1566 <= ((reg1456 >= {(reg1495 != reg1565)}) ?
                          $unsigned(((reg1502 & reg1565) | (reg1505 ?
                              forvar1546 : forvar1486))) : (-{(!reg1504)}));
                    end
                  else
                    begin
                      reg1563 <= forvar1461[(2'h2):(2'h2)];
                      reg1564 <= ((~|(reg1465[(2'h2):(1'h0)] < (forvar1456 != (8'ha4)))) << reg1455);
                    end
                  for (forvar1567 = (1'h0); (forvar1567 < (1'h1)); forvar1567 = (forvar1567 + (1'h1)))
                    begin
                      reg1568 <= (forvar1567[(1'h0):(1'h0)] ^ reg1521[(3'h4):(2'h3)]);
                      reg1569 <= $unsigned((|forvar1550[(2'h2):(1'h0)]));
                      reg1570 <= (8'hab);
                    end
                end
              if (reg1564[(4'ha):(2'h2)])
                begin
                  for (forvar1571 = (1'h0); (forvar1571 < (2'h3)); forvar1571 = (forvar1571 + (1'h1)))
                    begin
                      reg1572 <= ((reg1515 < $signed((forvar1543 ?
                              reg1527 : reg1495))) ?
                          {$unsigned((+reg1503))} : $unsigned(($unsigned(reg1540) | reg1477)));
                      reg1573 <= reg1486;
                      reg1574 <= (8'hab);
                    end
                  if ((($signed(forvar1476) ? $signed((8'h9c)) : {(&reg1498)}) ?
                      $signed((~forvar1540[(3'h5):(3'h4)])) : (~$signed(forvar1541[(1'h0):(1'h0)]))))
                    begin
                      reg1575 <= forvar1534;
                      reg1576 <= $signed((((~reg1456) ?
                          {reg1542} : reg1537[(4'h8):(4'h8)]) & ((wire1453 | reg1517) ?
                          $unsigned(reg1543) : $unsigned(forvar1545))));
                    end
                  else
                    begin
                      reg1575 <= {$signed({(reg1471 <<< reg1459)})};
                      reg1576 <= {reg1468};
                    end
                  for (forvar1577 = (1'h0); (forvar1577 < (2'h2)); forvar1577 = (forvar1577 + (1'h1)))
                    begin
                      reg1578 <= ($signed($signed({reg1563})) << ($unsigned((^~reg1500)) << {$unsigned(forvar1476)}));
                    end
                  reg1579 <= {{((reg1458 ? reg1546 : reg1469) ?
                              $signed(reg1465) : (-reg1530))}};
                end
              else
                begin
                  if ($unsigned(reg1469))
                    begin
                      reg1571 <= $unsigned(($unsigned((-(8'hb7))) ^~ ((wire1453 <<< reg1503) ?
                          forvar1506[(3'h6):(3'h4)] : {forvar1461})));
                      reg1572 <= (reg1532[(3'h7):(2'h2)] ?
                          reg1460 : (~&((reg1479 ?
                              reg1571 : (8'hb5)) + (^~reg1574))));
                    end
                  else
                    begin
                      reg1571 <= ((reg1561[(4'h8):(1'h1)] ?
                          reg1489[(1'h1):(1'h1)] : ($unsigned((8'hae)) ?
                              (reg1487 ?
                                  reg1546 : reg1574) : {forvar1518})) > $unsigned(($unsigned(reg1516) ?
                          (+reg1490) : $signed(reg1539))));
                    end
                  reg1573 <= $signed($signed(reg1546[(2'h3):(1'h0)]));
                end
            end
          else
            begin
              reg1558 <= reg1525;
              for (forvar1559 = (1'h0); (forvar1559 < (1'h1)); forvar1559 = (forvar1559 + (1'h1)))
                begin
                  for (forvar1560 = (1'h0); (forvar1560 < (2'h2)); forvar1560 = (forvar1560 + (1'h1)))
                    begin
                      reg1561 <= (8'hae);
                      reg1562 <= (~^(reg1461 >> {reg1576}));
                      reg1563 <= ($signed(((reg1530 ? reg1468 : reg1500) ?
                          ((8'ha1) ^~ reg1520) : reg1500[(1'h0):(1'h0)])) || reg1519);
                    end
                  if (forvar1514)
                    begin
                      reg1564 <= reg1527;
                    end
                  else
                    begin
                      reg1564 <= (|((&$unsigned(reg1481)) <<< forvar1501[(1'h0):(1'h0)]));
                      reg1565 <= wire5[(2'h2):(1'h1)];
                      reg1566 <= (($signed({forvar1560}) ?
                          ((~|(8'ha8)) <= (reg1538 ^ (8'hb1))) : (8'hab)) >> (((forvar1567 >= forvar1494) ~^ forvar1529[(4'hb):(1'h1)]) <= $signed(forvar1571[(3'h4):(2'h2)])));
                    end
                end
              if ((^$unsigned(forvar1472)))
                begin
                  for (forvar1567 = (1'h0); (forvar1567 < (2'h2)); forvar1567 = (forvar1567 + (1'h1)))
                    begin
                      reg1568 <= $signed((-(8'hae)));
                      reg1569 <= (reg1487[(1'h1):(1'h0)] || {$signed($unsigned(forvar1459))});
                      reg1570 <= reg1471[(1'h0):(1'h0)];
                      reg1571 <= $signed(((+(forvar1456 || wire1451)) ?
                          $unsigned(reg1505[(4'h9):(1'h0)]) : {(-reg1511)}));
                    end
                  for (forvar1572 = (1'h0); (forvar1572 < (1'h1)); forvar1572 = (forvar1572 + (1'h1)))
                    begin
                      reg1573 <= ($unsigned((+(reg1509 >>> forvar1456))) >= (($signed((8'hb6)) > (8'hab)) ?
                          reg1458 : forvar1548[(1'h0):(1'h0)]));
                      reg1574 <= $unsigned(($unsigned((reg1575 ?
                              (8'ha8) : reg1523)) ?
                          $signed((+reg1558)) : (+$unsigned(wire1))));
                      reg1575 <= ($signed(reg1504[(3'h6):(3'h4)]) ?
                          reg1488[(4'h9):(2'h2)] : forvar1506);
                      reg1576 <= reg1497[(1'h1):(1'h0)];
                    end
                  if ((~|$signed($unsigned(((8'ha9) - reg1526)))))
                    begin
                      reg1577 <= {(~(8'hb0))};
                      reg1578 <= {($unsigned((forvar1467 ?
                              reg1478 : (8'hb2))) < (^~$unsigned(forvar1541)))};
                    end
                  else
                    begin
                      reg1577 <= $signed({reg1556[(2'h3):(1'h0)]});
                      reg1578 <= ((reg1543 ?
                              wire1451[(4'he):(1'h0)] : $unsigned((~&(8'ha9)))) ?
                          {reg1507} : $signed({(forvar1577 ?
                                  reg1550 : reg1549)}));
                      reg1579 <= forvar1510;
                      reg1580 <= reg1530;
                    end
                  if (((|forvar1501[(1'h1):(1'h1)]) < $signed(((reg1458 ?
                      (8'hb2) : forvar1531) > reg1492[(3'h6):(1'h1)]))))
                    begin
                      reg1581 <= reg1517;
                      reg1582 <= reg1456[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg1581 <= reg1561;
                      reg1582 <= $signed($unsigned($signed($signed(reg1465))));
                    end
                end
              else
                begin
                  if ($signed((((wire1295 ? reg1551 : reg1508) ?
                      (forvar1559 == reg1535) : (forvar1454 ?
                          reg1473 : reg1485)) <= {$unsigned(reg1470)})))
                    begin
                      reg1567 <= {$unsigned(forvar1482)};
                      reg1568 <= ((+(&wire0)) && reg1458);
                      reg1569 <= {reg1461};
                    end
                  else
                    begin
                      reg1567 <= reg1539[(1'h0):(1'h0)];
                      reg1568 <= forvar1548;
                    end
                end
              for (forvar1583 = (1'h0); (forvar1583 < (1'h0)); forvar1583 = (forvar1583 + (1'h1)))
                begin
                  if ((reg1512 ?
                      reg1573 : ($unsigned($unsigned((8'hab))) ?
                          reg1509 : $signed($unsigned(reg1555)))))
                    begin
                      reg1584 <= $signed(reg1458[(4'h8):(4'h8)]);
                    end
                  else
                    begin
                      reg1584 <= reg1582[(3'h7):(1'h1)];
                    end
                  for (forvar1585 = (1'h0); (forvar1585 < (1'h1)); forvar1585 = (forvar1585 + (1'h1)))
                    begin
                      reg1586 <= (!$signed(({(8'h9c)} << reg1578)));
                      reg1587 <= ((&$signed($signed(reg1466))) ?
                          reg1457 : {((forvar1476 + reg1458) << reg1457)});
                      reg1588 <= {reg1478[(2'h3):(2'h2)]};
                      reg1589 <= $signed((!$signed((reg1525 ^~ (8'hb1)))));
                    end
                end
            end
          for (forvar1590 = (1'h0); (forvar1590 < (1'h1)); forvar1590 = (forvar1590 + (1'h1)))
            begin
              if (forvar1577)
                begin
                  if (reg1540)
                    begin
                      reg1591 <= (-reg1570[(4'hb):(4'h9)]);
                      reg1592 <= (^(reg1552[(3'h4):(1'h1)] ~^ reg1531));
                      reg1593 <= reg1512;
                    end
                  else
                    begin
                      reg1591 <= $unsigned((~^$unsigned(reg1486)));
                      reg1592 <= reg1579[(2'h2):(1'h1)];
                      reg1593 <= $signed(reg1491);
                    end
                end
              else
                begin
                  reg1591 <= $unsigned((reg1563 > $signed(((8'hb5) ?
                      reg1492 : reg1582))));
                  for (forvar1592 = (1'h0); (forvar1592 < (1'h1)); forvar1592 = (forvar1592 + (1'h1)))
                    begin
                      reg1593 <= reg1545;
                      reg1594 <= (reg1576 ?
                          ((&((8'ha7) + reg1546)) <<< (8'h9f)) : ($signed((~&reg1474)) ?
                              reg1552[(3'h5):(1'h1)] : $signed((forvar1459 ?
                                  forvar1533 : (8'h9c)))));
                    end
                  if (((((reg1478 ? forvar1529 : reg1478) ?
                          (forvar1518 >> reg1467) : (forvar1546 ^ reg1472)) != {$signed(forvar1548)}) ?
                      reg1511[(2'h2):(1'h1)] : (reg1508[(3'h6):(3'h4)] <<< wire1295[(4'hb):(2'h2)])))
                    begin
                      reg1595 <= $signed($signed(forvar1470));
                      reg1596 <= forvar1554[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg1595 <= (-(8'h9d));
                      reg1596 <= (^~(forvar1548[(2'h2):(1'h1)] ^~ reg1596));
                    end
                end
              for (forvar1597 = (1'h0); (forvar1597 < (2'h2)); forvar1597 = (forvar1597 + (1'h1)))
                begin
                  for (forvar1598 = (1'h0); (forvar1598 < (1'h0)); forvar1598 = (forvar1598 + (1'h1)))
                    begin
                      reg1599 <= reg1519;
                    end
                  for (forvar1600 = (1'h0); (forvar1600 < (1'h0)); forvar1600 = (forvar1600 + (1'h1)))
                    begin
                      reg1601 <= reg1511[(3'h7):(2'h3)];
                      reg1602 <= $unsigned({(~|$unsigned((8'ha4)))});
                    end
                  for (forvar1603 = (1'h0); (forvar1603 < (2'h3)); forvar1603 = (forvar1603 + (1'h1)))
                    begin
                      reg1604 <= ((~&({wire1451} ?
                          (reg1546 << reg1495) : (reg1511 && reg1595))) < reg1523[(4'ha):(4'h8)]);
                    end
                end
              if (reg1489[(4'hb):(4'h8)])
                begin
                  if ((reg1595 ?
                      ((reg1573 ?
                          reg1503[(3'h6):(2'h2)] : reg1498) & $unsigned($signed(reg1576))) : ({$signed(reg1501)} << (8'hb9))))
                    begin
                      reg1605 <= ({(reg1541[(1'h1):(1'h1)] ?
                                  $unsigned(forvar1538) : (reg1462 - forvar1585))} ?
                          reg1544 : (8'hb6));
                      reg1606 <= (^(~&forvar1482));
                      reg1607 <= (^~reg1591[(1'h1):(1'h1)]);
                    end
                  else
                    begin
                      reg1605 <= ((&($unsigned(reg1525) <= ((8'hb6) <= (8'hab)))) ?
                          (((reg1582 && reg1591) ?
                              (forvar1461 ?
                                  reg1538 : reg1545) : {forvar1455}) | (forvar1454 ?
                              $unsigned(reg1478) : $signed(forvar1559))) : {((-reg1591) ?
                                  reg1493 : (reg1472 + reg1572))});
                      reg1606 <= $unsigned(reg1588[(4'h9):(3'h6)]);
                    end
                  for (forvar1608 = (1'h0); (forvar1608 < (2'h2)); forvar1608 = (forvar1608 + (1'h1)))
                    begin
                      reg1609 <= ((($signed(reg1558) & forvar1454) <<< (+forvar1531)) ?
                          $unsigned((-(reg1516 ?
                              forvar1572 : wire6))) : $unsigned(($unsigned(reg1549) ?
                              $signed(forvar1485) : $unsigned(forvar1597))));
                      reg1610 <= $signed({($unsigned(reg1548) ?
                              forvar1499 : {reg1469})});
                      reg1611 <= (~|($unsigned(reg1538[(1'h1):(1'h1)]) ?
                          reg1567[(3'h4):(3'h4)] : (~|(reg1560 ?
                              reg1513 : reg1586))));
                    end
                end
              else
                begin
                  if ($signed(({$signed(reg1488)} + reg1571[(2'h3):(2'h3)])))
                    begin
                      reg1605 <= (-((forvar1558[(1'h0):(1'h0)] - (reg1463 && reg1594)) - $unsigned((~|reg1458))));
                      reg1606 <= reg1528;
                    end
                  else
                    begin
                      reg1605 <= (~&forvar1598[(3'h7):(3'h4)]);
                      reg1606 <= reg1464;
                    end
                end
              for (forvar1612 = (1'h0); (forvar1612 < (1'h0)); forvar1612 = (forvar1612 + (1'h1)))
                begin
                  for (forvar1613 = (1'h0); (forvar1613 < (1'h1)); forvar1613 = (forvar1613 + (1'h1)))
                    begin
                      reg1614 <= {((8'hac) ?
                              $unsigned(reg1602) : wire1451[(4'ha):(1'h1)])};
                      reg1615 <= reg1498;
                    end
                  for (forvar1616 = (1'h0); (forvar1616 < (1'h0)); forvar1616 = (forvar1616 + (1'h1)))
                    begin
                      reg1617 <= reg1572;
                    end
                end
            end
        end
    end
  assign wire1618 = (reg1548[(1'h1):(1'h0)] ?
                        $unsigned((forvar1483[(1'h1):(1'h0)] ?
                            reg1472 : (wire4 ?
                                reg1463 : reg1617))) : (!$signed({reg1564})));
  always
    @(posedge clk) begin
      if ($signed(reg1591[(3'h5):(3'h5)]))
        begin
          if ($signed((~|(^~(forvar1600 ? reg1460 : reg1609)))))
            begin
              for (forvar1619 = (1'h0); (forvar1619 < (1'h0)); forvar1619 = (forvar1619 + (1'h1)))
                begin
                  if ((~|$unsigned((8'hb5))))
                    begin
                      reg1620 <= (reg1582[(1'h0):(1'h0)] == reg1499);
                      reg1621 <= $signed($unsigned(reg1523[(4'hb):(4'h9)]));
                    end
                  else
                    begin
                      reg1620 <= $signed((~&($unsigned(forvar1467) ?
                          (8'haf) : (~|(8'hb7)))));
                    end
                end
              reg1622 <= {forvar1485[(3'h4):(2'h2)]};
              reg1623 <= reg1576;
              for (forvar1624 = (1'h0); (forvar1624 < (1'h1)); forvar1624 = (forvar1624 + (1'h1)))
                begin
                  for (forvar1625 = (1'h0); (forvar1625 < (1'h1)); forvar1625 = (forvar1625 + (1'h1)))
                    begin
                      reg1626 <= ((~&((reg1521 ?
                              reg1468 : reg1571) * reg1497[(1'h0):(1'h0)])) ?
                          reg1570[(4'hd):(3'h7)] : forvar1590[(2'h2):(1'h1)]);
                    end
                  for (forvar1627 = (1'h0); (forvar1627 < (1'h1)); forvar1627 = (forvar1627 + (1'h1)))
                    begin
                      reg1628 <= reg1526[(3'h6):(1'h1)];
                      reg1629 <= {reg1485[(4'hb):(2'h3)]};
                      reg1630 <= $signed($unsigned((reg1537 << $unsigned(reg1607))));
                      reg1631 <= $unsigned($signed(reg1504[(3'h5):(3'h4)]));
                    end
                end
            end
          else
            begin
              if (reg1515)
                begin
                  for (forvar1619 = (1'h0); (forvar1619 < (1'h1)); forvar1619 = (forvar1619 + (1'h1)))
                    begin
                      reg1620 <= ((^~((forvar1603 != (8'hb3)) ?
                              reg1474 : $signed(reg1477))) ?
                          forvar1524[(2'h3):(1'h1)] : (^((&reg1558) ?
                              $signed(reg1604) : $unsigned(reg1606))));
                    end
                  if (reg1592[(4'ha):(1'h1)])
                    begin
                      reg1621 <= $signed($unsigned(reg1460));
                    end
                  else
                    begin
                      reg1621 <= (reg1607[(2'h2):(2'h2)] << {((reg1606 ?
                                  (8'h9e) : forvar1459) ?
                              $signed(reg1495) : ((8'hb0) ?
                                  reg1499 : forvar1456))});
                      reg1622 <= reg1509[(1'h0):(1'h0)];
                    end
                  for (forvar1623 = (1'h0); (forvar1623 < (2'h3)); forvar1623 = (forvar1623 + (1'h1)))
                    begin
                      reg1624 <= $unsigned($unsigned($signed((^forvar1567))));
                      reg1625 <= $signed((|((8'hb9) ?
                          {reg1459} : (reg1546 ? wire1453 : (8'ha0)))));
                    end
                  for (forvar1626 = (1'h0); (forvar1626 < (1'h0)); forvar1626 = (forvar1626 + (1'h1)))
                    begin
                      reg1627 <= ($signed($unsigned((~|reg1551))) ?
                          ($signed({forvar1597}) * (8'hb3)) : {reg1565});
                      reg1628 <= ($unsigned(((-reg1520) * $signed(reg1573))) + (forvar1540 == ($unsigned(forvar1543) ?
                          reg1561[(2'h3):(2'h3)] : $unsigned(forvar1499))));
                      reg1629 <= ({$signed((forvar1623 ?
                                  reg1542 : forvar1603))} ?
                          $unsigned((((8'ha8) || (8'ha8)) - (^~forvar1626))) : $signed(({reg1460} ?
                              (forvar1540 << reg1542) : reg1556)));
                    end
                end
              else
                begin
                  for (forvar1619 = (1'h0); (forvar1619 < (1'h1)); forvar1619 = (forvar1619 + (1'h1)))
                    begin
                      reg1620 <= ({(~reg1500)} ?
                          (reg1550[(1'h1):(1'h0)] ?
                              ((reg1572 * reg1593) | {forvar1558}) : $unsigned(forvar1590[(2'h2):(2'h2)])) : ($unsigned((reg1623 && reg1489)) ?
                              {reg1466[(4'h9):(1'h1)]} : $unsigned((forvar1590 ?
                                  reg1570 : forvar1499))));
                      reg1621 <= $unsigned($signed(forvar1554[(3'h7):(1'h0)]));
                      reg1622 <= reg1541[(1'h0):(1'h0)];
                      reg1623 <= $signed(reg1525);
                    end
                  reg1624 <= $unsigned({reg1550[(1'h1):(1'h1)]});
                  if ((-(($signed(wire0) ? (^~reg1627) : {(8'hb2)}) ?
                      $signed((~&forvar1459)) : $signed($signed(reg1601)))))
                    begin
                      reg1625 <= reg1542;
                      reg1626 <= ({reg1467} >>> (reg1487[(1'h0):(1'h0)] ?
                          reg1470[(1'h1):(1'h0)] : reg1593));
                      reg1627 <= {$signed(((!reg1539) ?
                              ((8'h9c) - reg1604) : (reg1498 == forvar1501)))};
                    end
                  else
                    begin
                      reg1625 <= reg1631;
                      reg1626 <= (($signed($signed(reg1471)) ?
                              $signed((-forvar1472)) : {((8'h9f) >> forvar1548)}) ?
                          ((8'ha0) ?
                              ($signed(reg1543) && (|reg1459)) : $signed($unsigned(reg1520))) : (({wire1295} ^~ {(8'hb3)}) ?
                              reg1537[(3'h4):(3'h4)] : ((&wire3) ?
                                  {reg1621} : (8'hab))));
                    end
                end
              for (forvar1630 = (1'h0); (forvar1630 < (2'h2)); forvar1630 = (forvar1630 + (1'h1)))
                begin
                  for (forvar1631 = (1'h0); (forvar1631 < (1'h0)); forvar1631 = (forvar1631 + (1'h1)))
                    begin
                      reg1632 <= (~&(+((forvar1600 + reg1587) <= (reg1555 < reg1592))));
                    end
                  for (forvar1633 = (1'h0); (forvar1633 < (2'h2)); forvar1633 = (forvar1633 + (1'h1)))
                    begin
                      reg1634 <= ((&(reg1459 ~^ (^reg1564))) ?
                          (^~$unsigned(reg1558)) : ($unsigned((8'ha9)) ?
                              ($unsigned(reg1548) ~^ reg1491[(4'hc):(4'hc)]) : ((~&(8'hb4)) ?
                                  (reg1553 ~^ reg1464) : (8'hb6))));
                      reg1635 <= wire4;
                    end
                  for (forvar1636 = (1'h0); (forvar1636 < (1'h0)); forvar1636 = (forvar1636 + (1'h1)))
                    begin
                      reg1637 <= $signed((&(reg1605[(1'h0):(1'h0)] ?
                          (-forvar1502) : (wire1 ? reg1629 : (8'hb9)))));
                    end
                  if (reg1560)
                    begin
                      reg1638 <= $signed(forvar1633);
                    end
                  else
                    begin
                      reg1638 <= (reg1509 >= {$unsigned({reg1457})});
                      reg1639 <= ($signed(reg1572) ?
                          $unsigned((forvar1545[(2'h3):(1'h0)] & (8'haf))) : (reg1511 < (((8'h9f) ?
                              reg1577 : reg1635) != (reg1459 ?
                              wire6 : reg1582))));
                      reg1640 <= (reg1638[(3'h6):(2'h3)] * reg1570);
                    end
                end
              for (forvar1641 = (1'h0); (forvar1641 < (2'h3)); forvar1641 = (forvar1641 + (1'h1)))
                begin
                  for (forvar1642 = (1'h0); (forvar1642 < (1'h1)); forvar1642 = (forvar1642 + (1'h1)))
                    begin
                      reg1643 <= reg1614[(3'h5):(1'h0)];
                      reg1644 <= reg1553[(1'h0):(1'h0)];
                      reg1645 <= reg1545;
                      reg1646 <= $unsigned($unsigned((reg1640[(3'h7):(2'h2)] ?
                          (&reg1639) : $signed(wire5))));
                    end
                  if ((reg1563 ?
                      reg1458[(5'h10):(4'hd)] : reg1462[(3'h7):(3'h4)]))
                    begin
                      reg1647 <= (forvar1456 ?
                          $signed(reg1494[(2'h3):(2'h2)]) : forvar1546);
                      reg1648 <= (&forvar1623);
                      reg1649 <= $signed((forvar1501 == forvar1499[(3'h4):(1'h0)]));
                    end
                  else
                    begin
                      reg1647 <= forvar1630;
                      reg1648 <= reg1605[(2'h2):(1'h1)];
                    end
                  reg1650 <= (+($unsigned((8'ha9)) >>> (&$signed(forvar1540))));
                  if ({$signed((reg1553 >>> $unsigned(forvar1550)))})
                    begin
                      reg1651 <= (forvar1534[(2'h2):(1'h0)] << ($unsigned($signed((8'hb2))) ?
                          (forvar1456[(2'h2):(2'h2)] ?
                              $unsigned(reg1491) : $signed(wire1453)) : ($signed(forvar1540) ?
                              $unsigned(reg1459) : (~(8'ha0)))));
                    end
                  else
                    begin
                      reg1651 <= (((~^{reg1557}) ?
                              reg1581 : $signed({reg1538})) ?
                          (~|(|{(8'ha1)})) : (($unsigned((8'ha2)) ?
                                  forvar1495[(1'h1):(1'h1)] : (reg1635 + reg1546)) ?
                              $signed(((8'hb2) <= (8'haa))) : ((forvar1592 ?
                                      reg1592 : reg1565) ?
                                  (reg1548 ?
                                      reg1485 : reg1488) : forvar1459[(3'h7):(3'h7)])));
                    end
                end
              if (wire1451[(4'hf):(4'hb)])
                begin
                  if (forvar1636)
                    begin
                      reg1652 <= (&reg1609[(3'h4):(1'h0)]);
                    end
                  else
                    begin
                      reg1652 <= $signed((~^(reg1492 > {forvar1608})));
                      reg1653 <= (((reg1624[(1'h1):(1'h0)] ?
                          (+(8'haa)) : (reg1571 >>> forvar1624)) + reg1456[(1'h1):(1'h1)]) * $signed(reg1635[(3'h6):(1'h1)]));
                    end
                end
              else
                begin
                  if ((|forvar1559))
                    begin
                      reg1652 <= $unsigned({(8'hae)});
                    end
                  else
                    begin
                      reg1652 <= reg1632;
                      reg1653 <= reg1503;
                    end
                  reg1654 <= ($unsigned({(reg1487 ?
                          reg1582 : reg1485)}) >>> ((&{forvar1567}) ?
                      $unsigned(reg1606) : {(reg1599 >>> reg1543)}));
                  for (forvar1655 = (1'h0); (forvar1655 < (2'h2)); forvar1655 = (forvar1655 + (1'h1)))
                    begin
                      reg1656 <= $signed(forvar1560);
                      reg1657 <= (~&((reg1594 ? (8'hb2) : (|forvar1583)) ?
                          reg1484[(4'h8):(2'h2)] : {wire3}));
                      reg1658 <= wire5[(3'h7):(1'h0)];
                    end
                end
            end
        end
      else
        begin
          for (forvar1619 = (1'h0); (forvar1619 < (2'h3)); forvar1619 = (forvar1619 + (1'h1)))
            begin
              if (reg1539[(3'h5):(2'h3)])
                begin
                  if (((~&{(!reg1515)}) ?
                      {forvar1642[(5'h10):(3'h4)]} : (!$signed(((8'h9f) ?
                          reg1484 : reg1468)))))
                    begin
                      reg1620 <= ((8'ha1) ?
                          $unsigned(reg1601[(3'h7):(2'h2)]) : (&{$signed(wire1453)}));
                      reg1621 <= ((|(~(reg1548 ? reg1487 : forvar1597))) ?
                          $unsigned($unsigned($unsigned(reg1635))) : $signed((wire1618[(2'h3):(2'h3)] >> forvar1486)));
                      reg1622 <= $unsigned(reg1485[(4'ha):(1'h0)]);
                    end
                  else
                    begin
                      reg1620 <= ({reg1592} ?
                          (|(((8'ha2) && (8'hb8)) ?
                              forvar1567 : $unsigned(forvar1501))) : (~{reg1596[(5'h10):(4'ha)]}));
                      reg1621 <= forvar1534;
                      reg1622 <= (((&(reg1466 ? reg1644 : (8'hb6))) ?
                              forvar1616 : ((reg1466 != reg1654) == $signed(forvar1455))) ?
                          {$unsigned(reg1507)} : (($signed((8'ha1)) ^ (-reg1580)) ?
                              $unsigned((~reg1560)) : ({forvar1583} ?
                                  reg1634 : (reg1644 ? reg1484 : forvar1603))));
                      reg1623 <= forvar1548;
                    end
                  reg1624 <= (^(reg1535 != forvar1598[(3'h4):(2'h2)]));
                  if (($signed((+(~forvar1545))) + {reg1557[(3'h6):(2'h2)]}))
                    begin
                      reg1625 <= (~|(8'ha3));
                      reg1626 <= (+(&$signed((~&forvar1454))));
                      reg1627 <= ($signed((+(reg1593 < forvar1543))) > reg1615[(2'h2):(1'h0)]);
                      reg1628 <= ((8'ha2) ?
                          $unsigned(reg1563[(3'h4):(3'h4)]) : (8'ha7));
                    end
                  else
                    begin
                      reg1625 <= ((($signed(reg1584) ?
                              {reg1565} : {forvar1619}) ?
                          forvar1577 : reg1497) << reg1513[(4'ha):(4'h8)]);
                      reg1626 <= reg1611;
                    end
                end
              else
                begin
                  reg1620 <= (-$unsigned($unsigned((+reg1494))));
                end
              for (forvar1629 = (1'h0); (forvar1629 < (1'h0)); forvar1629 = (forvar1629 + (1'h1)))
                begin
                  for (forvar1630 = (1'h0); (forvar1630 < (1'h1)); forvar1630 = (forvar1630 + (1'h1)))
                    begin
                      reg1631 <= reg1460;
                      reg1632 <= forvar1592;
                    end
                  if (reg1635[(1'h1):(1'h0)])
                    begin
                      reg1633 <= ($signed(($signed((8'ha4)) ?
                              reg1471[(2'h2):(1'h1)] : (~^reg1464))) ?
                          (^(+(reg1561 ?
                              reg1480 : forvar1524))) : (((&(8'h9d)) ~^ reg1629[(1'h0):(1'h0)]) << (^~(reg1497 ?
                              reg1550 : reg1580))));
                      reg1634 <= $signed(($signed((reg1637 >>> forvar1559)) ?
                          (8'hb2) : ($unsigned(reg1617) << (reg1657 >>> reg1610))));
                      reg1635 <= forvar1486;
                      reg1636 <= $signed($signed($unsigned({reg1556})));
                    end
                  else
                    begin
                      reg1633 <= (!(($unsigned(reg1577) ?
                          (-reg1569) : forvar1494[(3'h6):(1'h0)]) < $signed((-reg1465))));
                      reg1634 <= forvar1545[(3'h6):(3'h6)];
                      reg1635 <= $signed($unsigned(reg1490));
                      reg1636 <= forvar1597[(2'h3):(2'h3)];
                    end
                  reg1637 <= forvar1476;
                end
              reg1638 <= ((((+reg1650) ^ $unsigned(forvar1624)) ?
                  $signed($signed(wire1)) : reg1523[(1'h1):(1'h0)]) + (^{reg1567[(2'h2):(1'h1)]}));
              if ((+(~&$unsigned((reg1503 ? reg1645 : reg1645)))))
                begin
                  for (forvar1639 = (1'h0); (forvar1639 < (1'h0)); forvar1639 = (forvar1639 + (1'h1)))
                    begin
                      reg1640 <= {$signed((&(reg1643 ? (8'h9f) : reg1521)))};
                      reg1641 <= $signed($signed(forvar1597[(1'h0):(1'h0)]));
                      reg1642 <= $unsigned((forvar1597[(2'h3):(2'h2)] ?
                          $signed($signed(reg1579)) : ({(8'hb8)} - $signed(reg1474))));
                    end
                end
              else
                begin
                  if ((~$signed((reg1517[(4'ha):(1'h0)] ?
                      $signed((8'hb4)) : (reg1586 + reg1465)))))
                    begin
                      reg1639 <= $signed((&({reg1541} <<< wire1453)));
                      reg1640 <= (&forvar1560[(2'h2):(2'h2)]);
                      reg1641 <= $signed($unsigned(reg1500));
                    end
                  else
                    begin
                      reg1639 <= (reg1637[(2'h2):(1'h1)] << $signed((reg1575 ?
                          (|forvar1630) : (+reg1488))));
                      reg1640 <= {forvar1533};
                      reg1641 <= (wire2 ?
                          reg1463 : (($unsigned(reg1516) ?
                              $signed(reg1464) : $signed(wire1295)) < wire1618[(1'h0):(1'h0)]));
                    end
                  if ((+reg1536[(4'ha):(4'h9)]))
                    begin
                      reg1642 <= (|$signed(reg1577[(1'h1):(1'h1)]));
                      reg1643 <= $signed(($unsigned((~reg1654)) ?
                          (reg1607[(4'hd):(4'hb)] >= reg1620) : {reg1479[(2'h2):(2'h2)]}));
                      reg1644 <= (8'h9d);
                      reg1645 <= $unsigned(({$signed(reg1561)} ^~ reg1540));
                    end
                  else
                    begin
                      reg1642 <= $unsigned((((reg1615 ~^ forvar1554) ^ forvar1554) ?
                          $unsigned((-(8'h9c))) : (8'hb3)));
                      reg1643 <= reg1499[(3'h7):(3'h6)];
                      reg1644 <= $unsigned((forvar1559[(2'h3):(1'h0)] ?
                          $unsigned((forvar1572 < (8'ha1))) : ((reg1464 > reg1605) ?
                              (8'ha1) : (reg1505 >= reg1503))));
                      reg1645 <= reg1575;
                    end
                  for (forvar1646 = (1'h0); (forvar1646 < (2'h3)); forvar1646 = (forvar1646 + (1'h1)))
                    begin
                      reg1647 <= ((reg1507[(2'h2):(1'h0)] ?
                          reg1628 : (reg1653[(4'h8):(1'h1)] ?
                              $signed(wire4) : forvar1470[(4'ha):(2'h2)])) != forvar1583);
                      reg1648 <= $signed(reg1555);
                      reg1649 <= (reg1573 ?
                          reg1624[(1'h0):(1'h0)] : forvar1608[(1'h1):(1'h1)]);
                      reg1650 <= reg1621;
                    end
                end
            end
          for (forvar1651 = (1'h0); (forvar1651 < (1'h0)); forvar1651 = (forvar1651 + (1'h1)))
            begin
              reg1652 <= reg1467;
            end
          if (reg1469)
            begin
              if ($signed((^forvar1613)))
                begin
                  for (forvar1653 = (1'h0); (forvar1653 < (1'h1)); forvar1653 = (forvar1653 + (1'h1)))
                    begin
                      reg1654 <= (((^~reg1485[(3'h7):(3'h4)]) ?
                          ((reg1632 ? reg1602 : forvar1567) ?
                              (~&reg1522) : forvar1653[(4'h8):(1'h1)]) : (|(reg1481 ?
                              forvar1456 : reg1624))) <= reg1650);
                      reg1655 <= ($signed((forvar1577[(1'h0):(1'h0)] ?
                          $signed(forvar1560) : forvar1608[(4'ha):(1'h0)])) ^ $unsigned(($unsigned(forvar1483) ?
                          reg1625[(2'h3):(1'h0)] : ((8'hb6) ?
                              reg1640 : reg1486))));
                      reg1656 <= ({reg1519[(3'h4):(2'h2)]} < (+$unsigned($signed(reg1563))));
                    end
                  for (forvar1657 = (1'h0); (forvar1657 < (2'h2)); forvar1657 = (forvar1657 + (1'h1)))
                    begin
                      reg1658 <= reg1468[(4'ha):(1'h1)];
                      reg1659 <= $unsigned(reg1527[(4'hd):(3'h5)]);
                      reg1660 <= forvar1572[(3'h7):(3'h4)];
                      reg1661 <= $signed(((8'ha8) ?
                          ((reg1545 ?
                              reg1622 : forvar1655) < (~&reg1548)) : $unsigned(forvar1583)));
                    end
                  for (forvar1662 = (1'h0); (forvar1662 < (2'h2)); forvar1662 = (forvar1662 + (1'h1)))
                    begin
                      reg1663 <= reg1528[(2'h3):(2'h3)];
                      reg1664 <= (8'hb8);
                    end
                end
              else
                begin
                  if ((((((8'hb4) ? reg1548 : forvar1550) ?
                          $unsigned(reg1577) : ((8'hb2) ?
                              reg1538 : forvar1558)) * $unsigned((forvar1494 ^~ reg1546))) ?
                      (((reg1638 ?
                          reg1485 : forvar1592) <= reg1537) ^~ (^$unsigned(reg1611))) : forvar1538))
                    begin
                      reg1653 <= $unsigned(reg1538[(3'h4):(2'h2)]);
                    end
                  else
                    begin
                      reg1653 <= (!reg1637[(2'h3):(1'h0)]);
                    end
                  reg1654 <= (^~reg1474[(1'h0):(1'h0)]);
                  if ((|(((8'ha0) || reg1477[(1'h0):(1'h0)]) != $unsigned(reg1550[(2'h2):(1'h1)]))))
                    begin
                      reg1655 <= reg1626[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1655 <= (forvar1624 ?
                          (+((forvar1470 ? forvar1558 : forvar1472) ?
                              reg1565[(3'h7):(2'h3)] : {reg1639})) : reg1457);
                      reg1656 <= ($signed(((|(8'had)) == (8'ha5))) ?
                          (reg1478[(1'h1):(1'h0)] > $unsigned((reg1546 ?
                              reg1644 : (8'ha9)))) : (((reg1577 ?
                                  reg1495 : forvar1655) != reg1591[(1'h0):(1'h0)]) ?
                              (forvar1545[(2'h3):(2'h3)] ?
                                  reg1551[(1'h0):(1'h0)] : reg1651) : {((8'ha6) ~^ reg1557)}));
                    end
                end
              reg1665 <= $unsigned(forvar1612);
              for (forvar1666 = (1'h0); (forvar1666 < (1'h1)); forvar1666 = (forvar1666 + (1'h1)))
                begin
                  for (forvar1667 = (1'h0); (forvar1667 < (2'h2)); forvar1667 = (forvar1667 + (1'h1)))
                    begin
                      reg1668 <= $unsigned(wire1618);
                      reg1669 <= (^~((wire6 < {reg1576}) - (reg1546[(2'h2):(2'h2)] < (^~reg1539))));
                      reg1670 <= reg1525;
                    end
                  for (forvar1671 = (1'h0); (forvar1671 < (1'h1)); forvar1671 = (forvar1671 + (1'h1)))
                    begin
                      reg1672 <= ($unsigned(($unsigned(wire0) << $signed(reg1643))) ?
                          forvar1608 : $signed({(reg1574 < reg1467)}));
                      reg1673 <= {((reg1633[(2'h3):(2'h2)] ?
                                  (^forvar1483) : $signed(forvar1558)) ?
                              (|$signed(forvar1483)) : (~(8'ha9)))};
                      reg1674 <= (~^$signed((8'ha8)));
                    end
                  if ($signed($unsigned({reg1481})))
                    begin
                      reg1675 <= {$signed($signed($unsigned(reg1643)))};
                    end
                  else
                    begin
                      reg1675 <= {$signed($unsigned($unsigned(reg1622)))};
                      reg1676 <= (forvar1501 ?
                          reg1480 : forvar1657[(4'he):(3'h5)]);
                      reg1677 <= reg1544[(2'h3):(2'h3)];
                    end
                  reg1678 <= {{{$unsigned((8'haa))}}};
                end
            end
          else
            begin
              if (forvar1482[(4'h9):(3'h6)])
                begin
                  for (forvar1653 = (1'h0); (forvar1653 < (1'h1)); forvar1653 = (forvar1653 + (1'h1)))
                    begin
                      reg1654 <= $signed((!{$signed((8'hac))}));
                    end
                  for (forvar1655 = (1'h0); (forvar1655 < (1'h0)); forvar1655 = (forvar1655 + (1'h1)))
                    begin
                      reg1656 <= $unsigned($unsigned(($signed(reg1563) ?
                          forvar1476[(3'h6):(3'h4)] : $signed(reg1577))));
                      reg1657 <= ($signed(reg1642) & {(+(reg1473 ?
                              reg1625 : reg1537))});
                      reg1658 <= (!reg1635[(3'h7):(3'h5)]);
                      reg1659 <= reg1595;
                    end
                  for (forvar1660 = (1'h0); (forvar1660 < (2'h3)); forvar1660 = (forvar1660 + (1'h1)))
                    begin
                      reg1661 <= reg1491;
                    end
                end
              else
                begin
                  reg1653 <= ($signed(reg1462[(3'h6):(1'h1)]) ?
                      $unsigned($signed($signed(forvar1636))) : ($unsigned($unsigned(reg1623)) ?
                          ((reg1500 <= (8'hb7)) ?
                              $unsigned((8'h9e)) : $signed((8'ha7))) : ($signed(reg1517) && (forvar1461 ?
                              reg1558 : reg1516))));
                  if ($unsigned((~^$signed($signed((8'ha3))))))
                    begin
                      reg1654 <= (^~(!(!(wire3 ^~ reg1611))));
                      reg1655 <= ({(forvar1631[(2'h3):(2'h2)] ?
                                  forvar1629 : (reg1512 + reg1496))} ?
                          ($signed($unsigned((8'ha1))) > (+(forvar1624 && reg1463))) : ($signed(((8'h9d) ~^ (8'hb5))) ?
                              (8'hb2) : ((^(8'ha0)) ?
                                  reg1548[(3'h7):(3'h5)] : (reg1522 >>> reg1644))));
                      reg1656 <= (!{$unsigned($unsigned(reg1635))});
                      reg1657 <= ((8'hb9) ?
                          reg1601 : ($signed($unsigned((8'h9d))) | {$unsigned(forvar1514)}));
                    end
                  else
                    begin
                      reg1654 <= (-(8'ha0));
                    end
                end
              if (reg1665[(2'h2):(1'h1)])
                begin
                  for (forvar1662 = (1'h0); (forvar1662 < (1'h1)); forvar1662 = (forvar1662 + (1'h1)))
                    begin
                      reg1663 <= (reg1659[(3'h6):(1'h1)] ?
                          (forvar1467 ?
                              ($signed(reg1574) == (wire0 ?
                                  wire3 : reg1460)) : (~^forvar1626)) : forvar1627[(1'h0):(1'h0)]);
                      reg1664 <= (reg1521[(1'h1):(1'h1)] >>> $signed($signed(((8'hae) | reg1481))));
                    end
                  reg1665 <= $unsigned($signed($signed(reg1650)));
                  reg1666 <= $signed(forvar1558);
                end
              else
                begin
                  for (forvar1662 = (1'h0); (forvar1662 < (1'h1)); forvar1662 = (forvar1662 + (1'h1)))
                    begin
                      reg1663 <= (^($unsigned((+(8'h9c))) ?
                          ($unsigned(reg1474) ?
                              $unsigned(reg1676) : reg1508) : reg1460));
                    end
                  for (forvar1664 = (1'h0); (forvar1664 < (2'h2)); forvar1664 = (forvar1664 + (1'h1)))
                    begin
                      reg1665 <= reg1551;
                      reg1666 <= (forvar1598 <= ((8'hb3) ?
                          $signed((reg1572 >> reg1470)) : ((8'ha5) >> $signed((8'hb0)))));
                      reg1667 <= ($signed((~reg1469[(3'h6):(3'h5)])) & $unsigned(($unsigned(forvar1541) || $signed(reg1579))));
                    end
                end
              for (forvar1668 = (1'h0); (forvar1668 < (1'h0)); forvar1668 = (forvar1668 + (1'h1)))
                begin
                  for (forvar1669 = (1'h0); (forvar1669 < (1'h1)); forvar1669 = (forvar1669 + (1'h1)))
                    begin
                      reg1670 <= $signed((reg1462 <= reg1644));
                    end
                  if ($unsigned((($signed((8'ha8)) ?
                      (forvar1455 ?
                          reg1551 : wire0) : $unsigned(reg1484)) & $unsigned({(8'haa)}))))
                    begin
                      reg1671 <= $unsigned($signed(forvar1482));
                    end
                  else
                    begin
                      reg1671 <= ($unsigned(reg1592[(4'h8):(4'h8)]) - ((^~$signed(reg1519)) <<< forvar1585));
                      reg1672 <= $unsigned((~((~forvar1501) ?
                          (forvar1558 && reg1579) : wire1295)));
                    end
                end
              if ($signed($unsigned($signed($signed(reg1486)))))
                begin
                  if ($signed(((reg1553[(1'h0):(1'h0)] ?
                          {(8'haa)} : forvar1624) ?
                      ((|forvar1608) > reg1660[(1'h0):(1'h0)]) : ((!reg1652) >> $unsigned(wire5)))))
                    begin
                      reg1673 <= forvar1612[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1673 <= ({(reg1648 & (|reg1511))} ?
                          reg1615[(1'h0):(1'h0)] : $signed($unsigned($signed(wire2))));
                      reg1674 <= (reg1567[(3'h4):(3'h4)] ? {reg1485} : (8'h9f));
                      reg1675 <= (($unsigned(((8'hac) <<< reg1562)) ?
                          {$signed(forvar1660)} : (forvar1629 ?
                              (reg1495 ?
                                  forvar1590 : reg1669) : reg1644)) - reg1570);
                    end
                  for (forvar1676 = (1'h0); (forvar1676 < (2'h3)); forvar1676 = (forvar1676 + (1'h1)))
                    begin
                      reg1677 <= $unsigned($unsigned(reg1564[(2'h2):(2'h2)]));
                      reg1678 <= forvar1624;
                      reg1679 <= ((^forvar1560) == {$unsigned(reg1490[(3'h7):(3'h6)])});
                      reg1680 <= ($signed({((8'hae) + reg1485)}) ?
                          reg1464[(3'h6):(3'h6)] : reg1512[(1'h0):(1'h0)]);
                    end
                end
              else
                begin
                  if ((($unsigned((forvar1541 ?
                          reg1658 : forvar1495)) & {(reg1504 >> forvar1600)}) ?
                      {({reg1652} ?
                              (reg1672 * reg1628) : $unsigned(reg1544))} : $signed($unsigned((forvar1529 & reg1543)))))
                    begin
                      reg1673 <= $unsigned(forvar1639[(3'h5):(1'h0)]);
                      reg1674 <= {(8'hb9)};
                      reg1675 <= $signed(reg1528);
                    end
                  else
                    begin
                      reg1673 <= ((($unsigned(forvar1613) ?
                          {reg1675} : (~^(8'ha3))) >> reg1593[(1'h0):(1'h0)]) <= (-$signed((&forvar1476))));
                      reg1674 <= $signed(($signed(((8'h9d) && reg1477)) ?
                          (~^$unsigned(reg1490)) : ($signed(reg1663) ?
                              $unsigned(forvar1538) : {reg1576})));
                    end
                  if ($unsigned({({reg1496} && $signed(reg1648))}))
                    begin
                      reg1676 <= {(-(reg1527[(3'h5):(2'h2)] ?
                              {reg1607} : $unsigned(reg1578)))};
                      reg1677 <= (forvar1538 ?
                          reg1640 : $unsigned((&(reg1650 ?
                              reg1679 : (8'ha6)))));
                    end
                  else
                    begin
                      reg1676 <= $signed((reg1669[(4'ha):(4'ha)] ?
                          reg1623 : reg1678));
                    end
                  reg1678 <= ((~^(8'hae)) && $unsigned((((8'hb7) <= reg1502) ?
                      (reg1652 >= reg1582) : forvar1624)));
                end
            end
          if ($signed($unsigned($unsigned((8'hba)))))
            begin
              for (forvar1681 = (1'h0); (forvar1681 < (2'h2)); forvar1681 = (forvar1681 + (1'h1)))
                begin
                  reg1682 <= (($unsigned((~&(8'h9c))) ?
                          reg1521[(3'h4):(2'h3)] : $unsigned(forvar1483[(2'h2):(1'h0)])) ?
                      (8'h9f) : (reg1498[(3'h5):(3'h4)] ?
                          forvar1485[(2'h3):(2'h2)] : (~(-reg1520))));
                  for (forvar1683 = (1'h0); (forvar1683 < (1'h0)); forvar1683 = (forvar1683 + (1'h1)))
                    begin
                      reg1684 <= $unsigned({reg1487});
                      reg1685 <= (wire1618[(4'ha):(1'h0)] ?
                          {reg1540[(3'h7):(3'h4)]} : $signed($unsigned(forvar1585[(2'h2):(2'h2)])));
                      reg1686 <= ($signed($unsigned(forvar1454[(4'ha):(3'h6)])) ?
                          forvar1461[(2'h2):(2'h2)] : reg1523[(4'hc):(3'h7)]);
                      reg1687 <= reg1607;
                    end
                  if (((((reg1492 >>> reg1566) ?
                      $signed(reg1566) : {reg1582}) && $signed((reg1485 ?
                      forvar1541 : reg1458))) == {reg1561[(4'h8):(1'h1)]}))
                    begin
                      reg1688 <= $unsigned(({(forvar1630 > reg1625)} ?
                          $signed($signed(reg1660)) : ($signed((8'hb3)) ?
                              (reg1684 ?
                                  forvar1455 : forvar1531) : (+reg1464))));
                      reg1689 <= (reg1517 ?
                          (((reg1573 ^~ reg1550) ?
                              $unsigned(reg1646) : (reg1523 ?
                                  reg1475 : (8'had))) ~^ (!(reg1646 <<< reg1528))) : forvar1625[(3'h5):(1'h0)]);
                      reg1690 <= $signed((reg1522[(3'h6):(2'h3)] ?
                          $signed((reg1488 ?
                              forvar1671 : reg1526)) : $unsigned((wire1 ?
                              forvar1472 : (8'ha5)))));
                      reg1691 <= $signed((((!reg1596) ?
                              reg1545[(3'h7):(2'h3)] : $signed(forvar1543)) ?
                          reg1493[(2'h2):(1'h0)] : (reg1532[(4'hb):(1'h0)] <<< forvar1506[(1'h0):(1'h0)])));
                    end
                  else
                    begin
                      reg1688 <= $unsigned((($signed(forvar1567) | forvar1613) ?
                          $unsigned($unsigned(reg1558)) : (8'h9c)));
                      reg1689 <= forvar1660[(4'hc):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar1681 = (1'h0); (forvar1681 < (2'h2)); forvar1681 = (forvar1681 + (1'h1)))
                begin
                  for (forvar1682 = (1'h0); (forvar1682 < (1'h1)); forvar1682 = (forvar1682 + (1'h1)))
                    begin
                      reg1683 <= reg1631;
                      reg1684 <= $signed($unsigned($unsigned((reg1686 ?
                          (8'hb5) : reg1595))));
                    end
                  for (forvar1685 = (1'h0); (forvar1685 < (1'h1)); forvar1685 = (forvar1685 + (1'h1)))
                    begin
                      reg1686 <= {(8'hb7)};
                    end
                end
            end
        end
      if ($unsigned(((8'hb0) ~^ (~|((8'hae) ? wire1618 : (8'haa))))))
        begin
          reg1692 <= ($signed($unsigned($signed(reg1676))) << (~|$signed($unsigned((8'ha0)))));
        end
      else
        begin
          reg1692 <= $unsigned((forvar1558 >= {$unsigned(forvar1624)}));
          for (forvar1693 = (1'h0); (forvar1693 < (2'h3)); forvar1693 = (forvar1693 + (1'h1)))
            begin
              for (forvar1694 = (1'h0); (forvar1694 < (1'h0)); forvar1694 = (forvar1694 + (1'h1)))
                begin
                  for (forvar1695 = (1'h0); (forvar1695 < (2'h3)); forvar1695 = (forvar1695 + (1'h1)))
                    begin
                      reg1696 <= (~(reg1596[(3'h7):(3'h6)] ?
                          $unsigned(reg1649) : forvar1467));
                      reg1697 <= reg1492;
                      reg1698 <= forvar1454[(1'h1):(1'h1)];
                      reg1699 <= $signed((~$signed(wire1453)));
                    end
                  if (reg1602)
                    begin
                      reg1700 <= forvar1624[(2'h3):(2'h2)];
                    end
                  else
                    begin
                      reg1700 <= wire1618;
                      reg1701 <= (((reg1682 ?
                              reg1527[(4'ha):(3'h4)] : {(8'ha7)}) << {reg1463[(2'h2):(1'h1)]}) ?
                          ({$signed(reg1620)} ?
                              reg1556[(3'h5):(1'h0)] : $signed((~|reg1473))) : (+(reg1511 ?
                              reg1668[(1'h1):(1'h0)] : (-forvar1619))));
                      reg1702 <= $signed({(8'hb1)});
                      reg1703 <= (~&{reg1509[(4'h9):(3'h4)]});
                    end
                end
              if (reg1620)
                begin
                  for (forvar1704 = (1'h0); (forvar1704 < (1'h0)); forvar1704 = (forvar1704 + (1'h1)))
                    begin
                      reg1705 <= $signed($signed({(^reg1666)}));
                    end
                  if (forvar1472)
                    begin
                      reg1706 <= $signed(({$signed(reg1651)} ?
                          (~$signed(reg1545)) : reg1630));
                    end
                  else
                    begin
                      reg1706 <= (~&$unsigned({$unsigned(reg1455)}));
                      reg1707 <= $signed(($unsigned((reg1685 ~^ reg1515)) <= ($signed(reg1584) ?
                          ((8'hb6) ?
                              (8'ha3) : reg1572) : reg1463[(1'h1):(1'h1)])));
                    end
                end
              else
                begin
                  reg1704 <= $unsigned(((!$signed(reg1470)) - {{(8'h9e)}}));
                  for (forvar1705 = (1'h0); (forvar1705 < (1'h0)); forvar1705 = (forvar1705 + (1'h1)))
                    begin
                      reg1706 <= (^((^~(reg1464 || (8'hba))) <<< $signed((reg1672 >= reg1532))));
                      reg1707 <= forvar1603[(2'h2):(1'h0)];
                    end
                  if (forvar1577)
                    begin
                      reg1708 <= {{reg1670}};
                      reg1709 <= {$unsigned(((reg1614 ? reg1469 : forvar1685) ?
                              (forvar1543 ?
                                  reg1682 : forvar1695) : ((8'hb3) * reg1540)))};
                      reg1710 <= $unsigned((|$unsigned((|reg1709))));
                      reg1711 <= $signed(((^(reg1644 ~^ reg1475)) && forvar1629[(3'h5):(2'h2)]));
                    end
                  else
                    begin
                      reg1708 <= ($unsigned(forvar1619[(1'h1):(1'h0)]) ?
                          reg1666 : (~$signed((reg1579 ? reg1596 : reg1464))));
                    end
                end
              for (forvar1712 = (1'h0); (forvar1712 < (2'h3)); forvar1712 = (forvar1712 + (1'h1)))
                begin
                  for (forvar1713 = (1'h0); (forvar1713 < (1'h1)); forvar1713 = (forvar1713 + (1'h1)))
                    begin
                      reg1714 <= {reg1528[(3'h5):(3'h4)]};
                      reg1715 <= $signed($unsigned(forvar1583[(3'h6):(2'h3)]));
                      reg1716 <= (($unsigned((reg1628 ?
                          reg1504 : (8'hb9))) + (reg1696 - (&reg1674))) & $signed((~^(reg1626 >>> reg1633))));
                      reg1717 <= (^((~&$signed(reg1520)) ?
                          {(~(8'hab))} : (&$signed(reg1635))));
                    end
                  if ((8'hba))
                    begin
                      reg1718 <= $unsigned(($signed((-reg1659)) * $signed($signed(forvar1577))));
                      reg1719 <= $unsigned(((&{reg1459}) ?
                          wire0[(3'h5):(1'h1)] : reg1659[(2'h3):(2'h3)]));
                      reg1720 <= (reg1611 ~^ forvar1585[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg1718 <= forvar1571[(3'h4):(1'h0)];
                      reg1719 <= $signed($signed({reg1464}));
                    end
                  for (forvar1721 = (1'h0); (forvar1721 < (1'h1)); forvar1721 = (forvar1721 + (1'h1)))
                    begin
                      reg1722 <= {reg1634[(4'h9):(3'h7)]};
                    end
                  if (($unsigned(reg1644) ? reg1593 : reg1480))
                    begin
                      reg1723 <= reg1602[(4'h8):(3'h5)];
                      reg1724 <= (!(((reg1557 ~^ (8'hb3)) + $unsigned(forvar1631)) < (~^$signed(reg1708))));
                    end
                  else
                    begin
                      reg1723 <= reg1675;
                      reg1724 <= $unsigned(forvar1567[(2'h2):(2'h2)]);
                      reg1725 <= (reg1639 ?
                          forvar1456[(1'h0):(1'h0)] : $unsigned((~{reg1714})));
                    end
                end
              reg1726 <= forvar1572[(1'h0):(1'h0)];
            end
          for (forvar1727 = (1'h0); (forvar1727 < (1'h0)); forvar1727 = (forvar1727 + (1'h1)))
            begin
              reg1728 <= (8'h9e);
              if ((+(+reg1544[(4'he):(3'h4)])))
                begin
                  reg1729 <= ((+((8'ha4) ?
                          (^~reg1645) : (forvar1529 >>> forvar1682))) ?
                      (wire2 ?
                          forvar1651[(2'h2):(1'h0)] : (&reg1488)) : (((reg1634 ?
                          forvar1671 : reg1649) >>> $signed(reg1667)) ^ (8'ha2)));
                end
              else
                begin
                  if (((((reg1630 ? reg1723 : reg1668) ?
                          ((8'hac) ? reg1552 : reg1671) : $unsigned((8'hb9))) ?
                      {(reg1564 <= reg1647)} : {(reg1710 >> reg1549)}) << (+forvar1534[(2'h3):(1'h1)])))
                    begin
                      reg1729 <= {($signed(reg1575[(4'ha):(3'h7)]) ?
                              (^(8'h9e)) : $signed($signed((8'hb4))))};
                      reg1730 <= $unsigned($unsigned($signed({reg1669})));
                      reg1731 <= $signed(reg1630);
                      reg1732 <= reg1731[(3'h6):(2'h2)];
                    end
                  else
                    begin
                      reg1729 <= $signed($signed($signed($signed((8'h9d)))));
                      reg1730 <= ({{(^reg1467)}} ?
                          (wire4[(4'ha):(2'h3)] ?
                              $signed($signed(reg1625)) : (reg1643 >> (8'hb3))) : (~&(~$unsigned(forvar1705))));
                    end
                  if (reg1492[(3'h6):(3'h6)])
                    begin
                      reg1733 <= $unsigned(($unsigned($unsigned(reg1528)) <<< $unsigned((!reg1701))));
                    end
                  else
                    begin
                      reg1733 <= $unsigned($signed(reg1471));
                    end
                end
            end
          if ($signed(((&forvar1627[(1'h0):(1'h0)]) <<< wire6[(4'ha):(3'h4)])))
            begin
              if ($signed(($unsigned((8'hae)) ?
                  $signed(forvar1713[(2'h2):(2'h2)]) : wire1618)))
                begin
                  for (forvar1734 = (1'h0); (forvar1734 < (2'h3)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= (^($unsigned($unsigned((8'ha9))) ?
                          reg1642 : $unsigned((-reg1711))));
                    end
                  for (forvar1736 = (1'h0); (forvar1736 < (1'h0)); forvar1736 = (forvar1736 + (1'h1)))
                    begin
                      reg1737 <= (+$unsigned(wire3));
                      reg1738 <= $unsigned(reg1472);
                      reg1739 <= (+(^forvar1506));
                      reg1740 <= reg1553[(3'h6):(3'h4)];
                    end
                  if (((reg1574[(2'h2):(1'h1)] - {reg1466}) ?
                      (+reg1587) : (reg1517 ? reg1546 : $unsigned({reg1571}))))
                    begin
                      reg1741 <= {$unsigned(((!reg1477) - ((8'hb4) ^ reg1474)))};
                      reg1742 <= (($unsigned((reg1551 >>> forvar1486)) ?
                              ($signed(forvar1495) ?
                                  reg1637[(2'h3):(2'h2)] : reg1703[(2'h3):(2'h3)]) : forvar1664[(1'h1):(1'h0)]) ?
                          (reg1679[(3'h7):(1'h0)] ?
                              (!$unsigned((8'haf))) : (|(reg1477 ?
                                  reg1717 : reg1717))) : reg1539);
                      reg1743 <= reg1455[(3'h6):(1'h0)];
                      reg1744 <= reg1684[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg1741 <= forvar1630[(1'h0):(1'h0)];
                      reg1742 <= ((reg1738[(4'h9):(3'h5)] ?
                          {(reg1696 ~^ reg1722)} : ((8'hae) << (reg1676 ?
                              (8'hb4) : forvar1727))) * ($signed(reg1553) ?
                          {reg1547} : $signed(forvar1664)));
                      reg1743 <= ((reg1607[(4'ha):(4'ha)] ?
                          ((~^reg1532) | $signed(reg1488)) : (+reg1467[(2'h2):(1'h1)])) != reg1478);
                      reg1744 <= $unsigned((8'h9d));
                    end
                  if (reg1550[(1'h1):(1'h1)])
                    begin
                      reg1745 <= $signed($unsigned(reg1733));
                      reg1746 <= ($unsigned((|((8'ha7) != reg1462))) ?
                          reg1604[(4'h8):(1'h1)] : $unsigned({reg1498[(1'h0):(1'h0)]}));
                      reg1747 <= $unsigned({reg1553});
                      reg1748 <= ({(forvar1608 ^ (reg1494 ^~ reg1547))} ?
                          ((+{reg1708}) ?
                              reg1560[(3'h5):(2'h2)] : $signed($unsigned(wire1618))) : forvar1510[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1745 <= ($signed(forvar1625) <<< $unsigned(reg1522[(3'h5):(3'h4)]));
                      reg1746 <= {(((reg1594 ?
                              (8'ha0) : (8'hb0)) >>> reg1683[(3'h5):(2'h3)]) ^~ ((reg1728 ?
                              reg1560 : reg1651) ~^ {forvar1600}))};
                    end
                end
              else
                begin
                  for (forvar1734 = (1'h0); (forvar1734 < (1'h1)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= (((+reg1627[(2'h2):(2'h2)]) ?
                              reg1638 : (+(reg1596 || forvar1608))) ?
                          reg1659[(3'h6):(3'h5)] : reg1680);
                    end
                  for (forvar1736 = (1'h0); (forvar1736 < (1'h0)); forvar1736 = (forvar1736 + (1'h1)))
                    begin
                      reg1737 <= ($unsigned(forvar1571[(2'h3):(1'h1)]) ?
                          {$signed($unsigned(reg1560))} : ($unsigned({reg1697}) ?
                              ((!reg1706) ?
                                  (forvar1518 * reg1622) : $unsigned(reg1617)) : (8'ha7)));
                      reg1738 <= ((&$unsigned($unsigned(forvar1660))) ?
                          (($unsigned((8'hb8)) ~^ $signed(reg1680)) && reg1711) : $unsigned($unsigned((reg1636 || reg1560))));
                      reg1739 <= (8'hb3);
                      reg1740 <= $signed(forvar1631[(4'he):(1'h1)]);
                    end
                  if (reg1737)
                    begin
                      reg1741 <= $signed($unsigned(reg1631));
                      reg1742 <= reg1488[(4'h8):(2'h2)];
                      reg1743 <= (8'ha4);
                    end
                  else
                    begin
                      reg1741 <= $unsigned(forvar1543);
                      reg1742 <= (forvar1630 > {$signed($unsigned(reg1669))});
                    end
                  for (forvar1744 = (1'h0); (forvar1744 < (1'h0)); forvar1744 = (forvar1744 + (1'h1)))
                    begin
                      reg1745 <= ({((reg1478 + reg1572) ?
                              forvar1486 : reg1706[(1'h1):(1'h1)])} || $signed(((reg1625 >> reg1471) ?
                          $unsigned(forvar1597) : forvar1499)));
                      reg1746 <= ({((~^reg1561) ?
                              $unsigned(reg1479) : (reg1550 >= reg1490))} >= ((&(reg1481 ?
                              (8'ha4) : (8'hac))) ?
                          (((8'ha9) >= forvar1630) <<< (8'ha9)) : (~$unsigned(reg1646))));
                      reg1747 <= reg1477;
                    end
                end
              if (((^(reg1492[(1'h1):(1'h1)] ~^ (forvar1626 && reg1722))) ?
                  $signed((^$unsigned(reg1515))) : reg1546[(1'h1):(1'h0)]))
                begin
                  if ($signed((~&((reg1602 ^ reg1586) < $unsigned(reg1508)))))
                    begin
                      reg1749 <= $unsigned(((reg1739[(2'h3):(2'h2)] | (8'ha8)) ?
                          reg1593 : (forvar1631[(3'h6):(1'h1)] ?
                              $unsigned((8'hb2)) : forvar1660[(3'h4):(1'h1)])));
                      reg1750 <= (~&$unsigned(reg1654));
                      reg1751 <= {$signed(forvar1713[(1'h0):(1'h0)])};
                    end
                  else
                    begin
                      reg1749 <= reg1686[(3'h4):(3'h4)];
                    end
                  for (forvar1752 = (1'h0); (forvar1752 < (1'h0)); forvar1752 = (forvar1752 + (1'h1)))
                    begin
                      reg1753 <= reg1654;
                      reg1754 <= ((&forvar1467) ?
                          $signed((!(reg1560 ?
                              (8'ha5) : forvar1612))) : ($signed($unsigned(reg1466)) + reg1730));
                    end
                  for (forvar1755 = (1'h0); (forvar1755 < (1'h1)); forvar1755 = (forvar1755 + (1'h1)))
                    begin
                      reg1756 <= $signed((reg1486[(1'h0):(1'h0)] ?
                          forvar1664 : ((reg1544 * reg1488) ?
                              reg1549[(4'he):(1'h1)] : (forvar1454 >= reg1676))));
                    end
                end
              else
                begin
                  reg1749 <= forvar1681;
                end
              for (forvar1757 = (1'h0); (forvar1757 < (2'h2)); forvar1757 = (forvar1757 + (1'h1)))
                begin
                  for (forvar1758 = (1'h0); (forvar1758 < (1'h1)); forvar1758 = (forvar1758 + (1'h1)))
                    begin
                      reg1759 <= reg1553;
                    end
                end
            end
          else
            begin
              if (({$unsigned((wire6 || reg1652))} & ($signed((+forvar1486)) ^~ reg1543)))
                begin
                  for (forvar1734 = (1'h0); (forvar1734 < (1'h1)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= {$unsigned(((reg1685 > wire1451) ^ $signed(forvar1461)))};
                      reg1736 <= $unsigned(reg1702);
                    end
                  if ((^reg1542[(4'hb):(1'h1)]))
                    begin
                      reg1737 <= (((|reg1725[(1'h0):(1'h0)]) && $signed($unsigned(reg1700))) ?
                          (8'hb5) : (~|$unsigned($unsigned(reg1461))));
                      reg1738 <= $unsigned((8'hb6));
                      reg1739 <= reg1586[(3'h6):(3'h6)];
                      reg1740 <= ((^reg1609) > $signed(((~&reg1678) ?
                          {reg1564} : (reg1574 ? reg1746 : reg1569))));
                    end
                  else
                    begin
                      reg1737 <= (forvar1681[(3'h6):(2'h2)] ~^ ({reg1491} ?
                          (forvar1454[(3'h6):(2'h3)] > (^(8'had))) : (8'h9e)));
                      reg1738 <= (((!$signed(reg1744)) + forvar1653[(1'h0):(1'h0)]) ^~ $signed(($unsigned(forvar1757) + (^~forvar1472))));
                    end
                  if ((&({{reg1666}} + (8'hb3))))
                    begin
                      reg1741 <= (~forvar1646[(2'h2):(2'h2)]);
                      reg1742 <= (+(({reg1668} ?
                              $signed((8'hb2)) : $signed((8'hb1))) ?
                          (((8'h9d) | reg1487) && forvar1467) : $unsigned($signed(reg1582))));
                      reg1743 <= $unsigned($unsigned($unsigned((!reg1469))));
                      reg1744 <= $unsigned((($signed(reg1671) ?
                              (reg1595 ~^ reg1507) : (reg1562 ~^ reg1660)) ?
                          (~^((8'hab) ? reg1688 : wire1295)) : reg1475));
                    end
                  else
                    begin
                      reg1741 <= {(+wire1618)};
                      reg1742 <= $unsigned($signed({(forvar1613 ?
                              (8'ha2) : reg1739)}));
                      reg1743 <= ($unsigned($signed((reg1723 ?
                              reg1702 : reg1637))) ?
                          ({reg1470[(2'h2):(2'h2)]} ~^ $unsigned((reg1539 ?
                              reg1541 : reg1498))) : ((^((8'hb9) == forvar1482)) ?
                              $unsigned($signed((8'hb5))) : (-{reg1725})));
                      reg1744 <= ($signed(reg1560[(3'h4):(1'h1)]) || (8'ha0));
                    end
                  if ($signed((reg1578[(4'ha):(1'h1)] ?
                      $unsigned({reg1677}) : ((reg1579 ~^ reg1623) | ((8'h9c) ?
                          reg1729 : reg1667)))))
                    begin
                      reg1745 <= (reg1494[(3'h6):(2'h2)] ?
                          {$unsigned($signed((8'haa)))} : reg1675[(4'h8):(3'h4)]);
                      reg1746 <= (8'hac);
                    end
                  else
                    begin
                      reg1745 <= ({$signed({wire0})} ?
                          forvar1531[(3'h6):(1'h0)] : $signed(((reg1480 ?
                              reg1564 : reg1623) != reg1463[(2'h2):(2'h2)])));
                      reg1746 <= (^(reg1747 || (forvar1633 >>> ((8'ha2) ?
                          (8'ha5) : reg1706))));
                      reg1747 <= $unsigned($unsigned((^~reg1747)));
                    end
                end
              else
                begin
                  for (forvar1734 = (1'h0); (forvar1734 < (1'h1)); forvar1734 = (forvar1734 + (1'h1)))
                    begin
                      reg1735 <= (^~($signed($unsigned(forvar1485)) ?
                          (!(!(8'hab))) : $unsigned(forvar1669)));
                      reg1736 <= reg1696[(2'h3):(1'h0)];
                      reg1737 <= ((reg1588 > (~^{forvar1585})) * $unsigned((+$unsigned(reg1516))));
                      reg1738 <= ($signed(($signed(reg1744) ?
                              $signed(reg1477) : $signed(reg1730))) ?
                          ($signed(forvar1550[(2'h2):(1'h1)]) && $signed($unsigned(forvar1651))) : ($signed($signed((8'ha5))) ^ {(+forvar1721)}));
                    end
                  for (forvar1739 = (1'h0); (forvar1739 < (1'h0)); forvar1739 = (forvar1739 + (1'h1)))
                    begin
                      reg1740 <= forvar1626;
                      reg1741 <= (&(+reg1569));
                      reg1742 <= $signed((reg1674 << $unsigned((reg1745 ?
                          forvar1651 : forvar1518))));
                      reg1743 <= (8'ha7);
                    end
                  if ({(reg1604 & (^{reg1742}))})
                    begin
                      reg1744 <= (reg1538[(2'h3):(1'h1)] << (^{{(8'hac)}}));
                    end
                  else
                    begin
                      reg1744 <= (($signed(reg1527) ?
                          ((reg1486 & forvar1631) ?
                              ((8'hba) ?
                                  forvar1633 : reg1697) : (reg1660 | reg1652)) : ((8'ha9) ?
                              (reg1740 > reg1697) : forvar1524)) && $signed($signed((reg1743 == reg1587))));
                      reg1745 <= (+reg1587[(3'h5):(1'h1)]);
                      reg1746 <= (8'hab);
                      reg1747 <= {(!reg1640[(3'h7):(3'h4)])};
                    end
                end
              for (forvar1748 = (1'h0); (forvar1748 < (2'h2)); forvar1748 = (forvar1748 + (1'h1)))
                begin
                  for (forvar1749 = (1'h0); (forvar1749 < (2'h3)); forvar1749 = (forvar1749 + (1'h1)))
                    begin
                      reg1750 <= (reg1661[(1'h0):(1'h0)] >>> {(~|(forvar1655 >>> forvar1739))});
                      reg1751 <= (-reg1644[(4'h8):(3'h4)]);
                    end
                  if (({{reg1678[(4'ha):(1'h1)]}} ?
                      ($unsigned((reg1710 ? forvar1472 : reg1543)) * {((8'hb0) ?
                              reg1759 : reg1720)}) : (reg1704[(4'h9):(1'h0)] ?
                          (forvar1755 ^~ (reg1670 ?
                              (8'haa) : forvar1538)) : $signed((-forvar1541)))))
                    begin
                      reg1752 <= reg1635;
                      reg1753 <= (~&$unsigned(forvar1548[(1'h1):(1'h1)]));
                    end
                  else
                    begin
                      reg1752 <= ($signed($unsigned($signed((8'hba)))) && $unsigned((~&$signed(reg1552))));
                      reg1753 <= {($unsigned((reg1663 ?
                              reg1703 : forvar1483)) != $unsigned($signed(reg1738)))};
                    end
                end
            end
        end
      if ({((!(reg1489 ^~ wire1)) ?
              (((8'ha1) ^ (8'hba)) ?
                  $unsigned((8'hb2)) : forvar1616) : reg1553[(2'h3):(1'h0)])})
        begin
          for (forvar1760 = (1'h0); (forvar1760 < (1'h1)); forvar1760 = (forvar1760 + (1'h1)))
            begin
              if (forvar1758[(2'h2):(2'h2)])
                begin
                  if ((8'h9d))
                    begin
                      reg1761 <= ((~^(^(reg1587 ? forvar1748 : reg1643))) ?
                          (|($unsigned(reg1566) ?
                              $unsigned(wire5) : (reg1710 * reg1552))) : (+($signed(forvar1598) < ((8'hb7) <<< (8'ha9)))));
                    end
                  else
                    begin
                      reg1761 <= $signed(reg1627);
                      reg1762 <= (forvar1623[(4'h9):(3'h5)] ?
                          ($signed($signed(reg1729)) + ((8'hb9) ?
                              {forvar1585} : (8'hb8))) : (8'h9d));
                      reg1763 <= ({forvar1749} ?
                          (forvar1592 ?
                              $signed(reg1634) : (~^(reg1647 ?
                                  (8'h9e) : (8'ha3)))) : (forvar1590[(1'h0):(1'h0)] & $signed((reg1610 != reg1522))));
                      reg1764 <= ($unsigned((~reg1480)) ?
                          reg1576[(1'h1):(1'h0)] : forvar1734);
                    end
                end
              else
                begin
                  for (forvar1761 = (1'h0); (forvar1761 < (1'h1)); forvar1761 = (forvar1761 + (1'h1)))
                    begin
                      reg1762 <= (reg1626[(1'h0):(1'h0)] ?
                          ($unsigned({reg1572}) ?
                              (~^forvar1467[(4'hb):(4'h9)]) : {{forvar1494}}) : ({((8'h9d) < reg1691)} + ((reg1733 || forvar1545) <<< {(8'h9c)})));
                      reg1763 <= $unsigned((~(&((8'hac) ?
                          reg1665 : forvar1636))));
                      reg1764 <= reg1545;
                    end
                  for (forvar1765 = (1'h0); (forvar1765 < (2'h2)); forvar1765 = (forvar1765 + (1'h1)))
                    begin
                      reg1766 <= (forvar1518[(3'h7):(3'h4)] ?
                          reg1748 : $signed($signed(reg1587[(2'h2):(2'h2)])));
                      reg1767 <= (^(~&(!(forvar1657 > (8'hb3)))));
                    end
                  for (forvar1768 = (1'h0); (forvar1768 < (2'h3)); forvar1768 = (forvar1768 + (1'h1)))
                    begin
                      reg1769 <= $signed({$unsigned(forvar1490[(4'ha):(2'h2)])});
                      reg1770 <= reg1635;
                      reg1771 <= (|reg1733[(4'hb):(1'h1)]);
                      reg1772 <= (~^$unsigned(((reg1566 ^ reg1532) ^~ forvar1657)));
                    end
                  reg1773 <= ((({(8'hb5)} >> reg1513) >> (((8'hb2) + reg1730) >> $unsigned(reg1763))) || ($unsigned(reg1665) == (&{reg1770})));
                end
            end
          if (reg1467)
            begin
              for (forvar1774 = (1'h0); (forvar1774 < (2'h3)); forvar1774 = (forvar1774 + (1'h1)))
                begin
                  for (forvar1775 = (1'h0); (forvar1775 < (1'h1)); forvar1775 = (forvar1775 + (1'h1)))
                    begin
                      reg1776 <= (-{(8'h9e)});
                    end
                  reg1777 <= ($signed($unsigned((!forvar1572))) ?
                      ($signed({reg1541}) & (~&(+reg1605))) : ((forvar1646 < $signed((8'hb0))) ?
                          $unsigned(reg1581[(3'h4):(1'h0)]) : reg1581[(1'h0):(1'h0)]));
                end
            end
          else
            begin
              if (((reg1495 == ((&(8'hb5)) != ((8'hb1) ?
                  reg1642 : reg1578))) >>> $signed(($signed(reg1566) ?
                  reg1572[(3'h4):(2'h2)] : forvar1624[(4'h9):(3'h4)]))))
                begin
                  if (((forvar1629 ?
                          forvar1704[(4'hc):(4'ha)] : reg1474[(1'h1):(1'h0)]) ?
                      reg1471 : ((8'hb4) ?
                          reg1605 : (+(reg1586 << forvar1538)))))
                    begin
                      reg1774 <= $signed(({(forvar1660 << reg1732)} ?
                          forvar1668[(4'h8):(3'h5)] : forvar1456));
                      reg1775 <= (~&(reg1753 ?
                          $signed((&reg1485)) : $signed(reg1741)));
                    end
                  else
                    begin
                      reg1774 <= $signed(forvar1749[(1'h1):(1'h0)]);
                      reg1775 <= {forvar1461};
                      reg1776 <= {$unsigned(forvar1727)};
                      reg1777 <= (reg1580 ?
                          reg1704[(4'hb):(4'hb)] : {((-forvar1571) ?
                                  (8'h9e) : $signed(reg1517))});
                    end
                  if (($signed((reg1630 ? {reg1745} : $unsigned(wire1))) ?
                      $signed(reg1574) : reg1488))
                    begin
                      reg1778 <= reg1469[(3'h5):(3'h5)];
                      reg1779 <= reg1573;
                      reg1780 <= $signed(forvar1524);
                      reg1781 <= $signed($signed($signed(reg1749)));
                    end
                  else
                    begin
                      reg1778 <= (-{$signed(forvar1583[(3'h7):(2'h2)])});
                      reg1779 <= ((reg1490 ^ $unsigned(reg1567[(2'h3):(1'h0)])) ?
                          (forvar1682 ?
                              $signed((^reg1700)) : $unsigned((!forvar1642))) : reg1545);
                      reg1780 <= (~^(($signed(reg1493) ?
                              ((8'ha7) ? reg1677 : reg1628) : (reg1589 ?
                                  reg1744 : reg1495)) ?
                          ((&(8'ha0)) ^~ (~reg1751)) : $unsigned((~|reg1665))));
                    end
                end
              else
                begin
                  for (forvar1774 = (1'h0); (forvar1774 < (2'h2)); forvar1774 = (forvar1774 + (1'h1)))
                    begin
                      reg1775 <= $unsigned($unsigned($unsigned((reg1656 >>> reg1689))));
                    end
                  for (forvar1776 = (1'h0); (forvar1776 < (1'h0)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 <= (({(reg1704 >> reg1593)} ?
                          ((reg1780 ?
                              reg1549 : reg1513) & $signed(reg1722)) : {reg1653}) + $unsigned((~&(reg1683 ?
                          reg1669 : reg1699))));
                      reg1778 <= ($signed(reg1728) ?
                          ((8'h9f) ?
                              ((reg1667 ^ wire1618) < reg1773[(3'h5):(3'h5)]) : $unsigned(((8'haa) ?
                                  reg1766 : forvar1669))) : forvar1748);
                      reg1779 <= (reg1568 ?
                          {((reg1601 == reg1703) || reg1638[(2'h3):(2'h3)])} : (8'haf));
                      reg1780 <= $unsigned(reg1743[(2'h2):(1'h1)]);
                    end
                  reg1781 <= (!((~|(reg1749 ?
                      forvar1662 : reg1488)) ^ forvar1752[(1'h0):(1'h0)]));
                  reg1782 <= ((~|reg1457[(2'h2):(1'h0)]) ?
                      $signed($unsigned((~^reg1521))) : reg1771);
                end
              if (reg1469)
                begin
                  reg1783 <= reg1540[(3'h7):(2'h2)];
                  if ((+{(~(^reg1565))}))
                    begin
                      reg1784 <= ($unsigned(reg1571) ?
                          (wire2[(4'h8):(3'h7)] != $unsigned((~|reg1697))) : (reg1485 + {$signed(reg1701)}));
                      reg1785 <= {reg1696};
                      reg1786 <= reg1556[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg1784 <= $signed(($unsigned((reg1560 << reg1756)) ?
                          (~^(forvar1501 ? forvar1585 : (8'h9e))) : (8'hac)));
                      reg1785 <= $signed(reg1653);
                      reg1786 <= $signed((((reg1704 ?
                          reg1470 : wire1453) <= (reg1644 ?
                          reg1577 : forvar1486)) << (~&(reg1715 != reg1547))));
                    end
                  for (forvar1787 = (1'h0); (forvar1787 < (1'h0)); forvar1787 = (forvar1787 + (1'h1)))
                    begin
                      reg1788 <= ((8'haf) ?
                          (forvar1752 ?
                              ($signed(forvar1727) * $unsigned(reg1690)) : $signed(forvar1554)) : $signed($unsigned(reg1573[(4'hb):(3'h7)])));
                      reg1789 <= $signed(reg1707[(2'h2):(2'h2)]);
                    end
                end
              else
                begin
                  for (forvar1783 = (1'h0); (forvar1783 < (1'h0)); forvar1783 = (forvar1783 + (1'h1)))
                    begin
                      reg1784 <= $signed($signed(forvar1597));
                    end
                end
              reg1790 <= $unsigned((reg1692[(1'h1):(1'h1)] <<< (~^reg1481[(3'h4):(1'h0)])));
              if ($signed((reg1724[(4'hb):(3'h5)] ?
                  $signed((forvar1486 == reg1709)) : (~|(reg1551 || reg1690)))))
                begin
                  if ((!$unsigned(forvar1626[(2'h3):(1'h1)])))
                    begin
                      reg1791 <= (8'haf);
                      reg1792 <= (~&reg1614);
                      reg1793 <= reg1747;
                    end
                  else
                    begin
                      reg1791 <= (($unsigned(reg1528[(4'hb):(3'h4)]) ?
                          (^((8'hac) <= reg1522)) : (reg1674 ?
                              reg1750[(4'h9):(3'h4)] : reg1532[(4'hb):(1'h1)])) ~^ $unsigned($unsigned($unsigned(reg1767))));
                    end
                  if (reg1732)
                    begin
                      reg1794 <= (^~(~((forvar1639 ?
                          forvar1598 : reg1620) < $unsigned((8'ha9)))));
                      reg1795 <= $signed(($signed((~reg1552)) == ((reg1606 != reg1747) & {reg1515})));
                      reg1796 <= ($signed({(^reg1750)}) | $unsigned(($unsigned(reg1581) ?
                          (8'ha1) : (+reg1479))));
                    end
                  else
                    begin
                      reg1794 <= (^reg1791);
                      reg1795 <= (reg1780[(1'h1):(1'h1)] <= reg1584);
                      reg1796 <= reg1614[(3'h7):(2'h2)];
                    end
                end
              else
                begin
                  for (forvar1791 = (1'h0); (forvar1791 < (2'h2)); forvar1791 = (forvar1791 + (1'h1)))
                    begin
                      reg1792 <= reg1541;
                      reg1793 <= {$signed(reg1703[(2'h3):(1'h1)])};
                      reg1794 <= (((-forvar1612) ?
                          ((reg1500 >> forvar1768) > reg1667[(3'h4):(2'h3)]) : forvar1559[(2'h3):(2'h2)]) == (($signed((8'hb1)) - $signed(forvar1655)) ?
                          $signed($unsigned(reg1742)) : $unsigned((|reg1642))));
                    end
                end
            end
          for (forvar1797 = (1'h0); (forvar1797 < (1'h0)); forvar1797 = (forvar1797 + (1'h1)))
            begin
              for (forvar1798 = (1'h0); (forvar1798 < (1'h0)); forvar1798 = (forvar1798 + (1'h1)))
                begin
                  if ((~^$unsigned($signed(((8'haf) ? reg1679 : reg1584)))))
                    begin
                      reg1799 <= (reg1794[(3'h4):(2'h3)] ?
                          (((-reg1794) | {reg1552}) + reg1467) : wire0[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg1799 <= $signed(reg1567[(1'h1):(1'h0)]);
                      reg1800 <= $signed((forvar1664 ?
                          $signed($signed(forvar1461)) : ($signed(reg1473) ?
                              (reg1499 ?
                                  forvar1727 : (8'h9e)) : reg1475[(2'h2):(1'h0)])));
                      reg1801 <= (^~(($unsigned(forvar1721) ?
                          ((8'haf) ?
                              (8'hb5) : reg1799) : (reg1733 | reg1546)) <= $signed((forvar1758 == reg1515))));
                      reg1802 <= forvar1567[(1'h1):(1'h0)];
                    end
                  reg1803 <= reg1475;
                  if (reg1570[(4'hc):(4'hb)])
                    begin
                      reg1804 <= ((reg1641[(4'he):(4'hd)] + reg1523[(3'h7):(1'h1)]) ?
                          (reg1462[(4'hf):(1'h1)] >= {reg1463[(2'h3):(2'h3)]}) : $signed($unsigned($unsigned(reg1527))));
                    end
                  else
                    begin
                      reg1804 <= $unsigned($signed((reg1580[(3'h7):(3'h4)] - ((8'had) < reg1674))));
                      reg1805 <= (((!{wire6}) ^~ $signed(forvar1548)) ?
                          (|((~^reg1791) ?
                              ((8'hac) ?
                                  reg1701 : reg1544) : (reg1754 - forvar1567))) : $signed((!{reg1517})));
                      reg1806 <= ({forvar1669} ?
                          forvar1783[(4'hb):(1'h0)] : ((~&{reg1526}) ~^ $unsigned((reg1609 ?
                              reg1747 : reg1730))));
                    end
                end
            end
        end
      else
        begin
          reg1760 <= (~|reg1658[(2'h2):(1'h0)]);
          for (forvar1761 = (1'h0); (forvar1761 < (2'h3)); forvar1761 = (forvar1761 + (1'h1)))
            begin
              for (forvar1762 = (1'h0); (forvar1762 < (1'h0)); forvar1762 = (forvar1762 + (1'h1)))
                begin
                  if ($signed(reg1486[(2'h2):(1'h0)]))
                    begin
                      reg1763 <= ((($signed(reg1689) ?
                              (reg1800 ?
                                  (8'hba) : forvar1482) : reg1764[(1'h1):(1'h1)]) ?
                          (forvar1518 ~^ reg1683[(3'h7):(3'h5)]) : (-(reg1460 != reg1735))) < $signed($signed($unsigned((8'ha5)))));
                      reg1764 <= (reg1552 ?
                          (~^$signed(((8'ha5) >>> (8'hb4)))) : reg1460[(1'h1):(1'h1)]);
                      reg1765 <= reg1509;
                    end
                  else
                    begin
                      reg1763 <= (+forvar1653);
                    end
                  for (forvar1766 = (1'h0); (forvar1766 < (1'h0)); forvar1766 = (forvar1766 + (1'h1)))
                    begin
                      reg1767 <= reg1707[(3'h5):(3'h4)];
                      reg1768 <= forvar1762;
                    end
                end
              for (forvar1769 = (1'h0); (forvar1769 < (1'h1)); forvar1769 = (forvar1769 + (1'h1)))
                begin
                  for (forvar1770 = (1'h0); (forvar1770 < (2'h2)); forvar1770 = (forvar1770 + (1'h1)))
                    begin
                      reg1771 <= ($signed({reg1511[(3'h5):(3'h4)]}) ~^ $signed(($signed(forvar1548) ?
                          $unsigned(reg1767) : reg1571)));
                      reg1772 <= ($unsigned($unsigned((reg1754 <<< (8'hb9)))) ?
                          (+reg1733) : forvar1761);
                      reg1773 <= forvar1639;
                      reg1774 <= $unsigned(((~$unsigned((8'had))) ?
                          (8'hba) : $unsigned($signed((8'ha6)))));
                    end
                end
              if (forvar1546[(1'h1):(1'h0)])
                begin
                  reg1775 <= $signed(reg1744[(1'h0):(1'h0)]);
                  for (forvar1776 = (1'h0); (forvar1776 < (2'h2)); forvar1776 = (forvar1776 + (1'h1)))
                    begin
                      reg1777 <= reg1783;
                      reg1778 <= $unsigned({($signed(reg1469) << $unsigned(forvar1483))});
                      reg1779 <= $unsigned(((-(^~forvar1755)) ?
                          $unsigned((reg1783 ?
                              wire6 : reg1677)) : $unsigned((reg1776 ?
                              reg1573 : reg1775))));
                      reg1780 <= ($unsigned($unsigned(forvar1546)) && (($unsigned(reg1473) >= $signed(reg1761)) ?
                          (^~$signed(reg1543)) : (reg1665 ?
                              reg1475 : (forvar1798 ? forvar1524 : reg1793))));
                    end
                  if ({$signed({forvar1518})})
                    begin
                      reg1781 <= $unsigned(wire1453);
                      reg1782 <= forvar1757;
                      reg1783 <= $signed((reg1640[(3'h7):(1'h0)] >> $signed((8'hb1))));
                      reg1784 <= $unsigned(forvar1600[(4'h8):(4'h8)]);
                    end
                  else
                    begin
                      reg1781 <= reg1663[(4'ha):(3'h7)];
                      reg1782 <= forvar1734[(3'h4):(2'h2)];
                      reg1783 <= reg1785;
                      reg1784 <= (~&(-(reg1542 >= reg1579)));
                    end
                  for (forvar1785 = (1'h0); (forvar1785 < (1'h0)); forvar1785 = (forvar1785 + (1'h1)))
                    begin
                      reg1786 <= reg1772[(1'h1):(1'h0)];
                      reg1787 <= (+((~&(reg1584 <= reg1562)) != {$signed(reg1750)}));
                      reg1788 <= (reg1751[(4'h8):(2'h3)] <<< ($signed(reg1601[(3'h7):(3'h4)]) * $unsigned($unsigned(reg1502))));
                    end
                end
              else
                begin
                  for (forvar1775 = (1'h0); (forvar1775 < (1'h0)); forvar1775 = (forvar1775 + (1'h1)))
                    begin
                      reg1776 <= $unsigned((+(8'haa)));
                      reg1777 <= (forvar1760 * ($signed((|reg1785)) ^ {((8'ha3) ?
                              forvar1761 : reg1637)}));
                      reg1778 <= reg1491;
                    end
                  if (reg1586)
                    begin
                      reg1779 <= reg1563[(3'h7):(1'h1)];
                      reg1780 <= reg1744;
                      reg1781 <= $signed(((8'h9f) ? {(+reg1557)} : reg1467));
                    end
                  else
                    begin
                      reg1779 <= forvar1454[(4'h9):(3'h5)];
                      reg1780 <= $signed(((~|{reg1639}) && forvar1669[(4'hb):(4'h8)]));
                    end
                  for (forvar1782 = (1'h0); (forvar1782 < (1'h0)); forvar1782 = (forvar1782 + (1'h1)))
                    begin
                      reg1783 <= (^$unsigned(((reg1610 ?
                          (8'ha6) : forvar1770) ^~ $unsigned((8'hb4)))));
                      reg1784 <= (reg1769 ?
                          (((forvar1459 ? reg1455 : reg1680) >> reg1570) ?
                              $signed(reg1570) : ((!reg1724) ?
                                  $unsigned(forvar1766) : $unsigned(forvar1518))) : reg1542[(4'h8):(3'h6)]);
                    end
                  for (forvar1785 = (1'h0); (forvar1785 < (1'h1)); forvar1785 = (forvar1785 + (1'h1)))
                    begin
                      reg1786 <= $signed((^(!reg1766[(2'h2):(1'h1)])));
                      reg1787 <= {forvar1571};
                    end
                end
            end
          if (reg1683[(1'h1):(1'h1)])
            begin
              reg1789 <= (8'h9e);
            end
          else
            begin
              if ((reg1724[(3'h5):(1'h1)] ?
                  reg1768 : (~|({reg1660} <<< {reg1586}))))
                begin
                  if (reg1502)
                    begin
                      reg1789 <= reg1654;
                      reg1790 <= $signed({{(forvar1752 != forvar1461)}});
                    end
                  else
                    begin
                      reg1789 <= reg1462[(4'he):(3'h5)];
                      reg1790 <= ($signed(($signed(reg1633) >= (reg1803 * reg1594))) * $unsigned((|((8'hb3) ?
                          reg1680 : reg1513))));
                      reg1791 <= {{(reg1638 ?
                                  (reg1570 <= reg1696) : ((8'h9f) ?
                                      reg1620 : forvar1541))}};
                      reg1792 <= $unsigned(($unsigned($unsigned((8'h9c))) ?
                          $unsigned((forvar1499 ?
                              (8'hb4) : (8'ha9))) : {forvar1755[(2'h2):(1'h1)]}));
                    end
                end
              else
                begin
                  reg1789 <= (~^{$unsigned(reg1682)});
                  reg1790 <= (($unsigned({forvar1577}) & forvar1736) && $unsigned(((reg1696 ~^ reg1711) ?
                      (reg1770 <= reg1555) : forvar1657)));
                  for (forvar1791 = (1'h0); (forvar1791 < (2'h3)); forvar1791 = (forvar1791 + (1'h1)))
                    begin
                      reg1792 <= (^(-$signed(forvar1791[(2'h3):(1'h1)])));
                      reg1793 <= reg1579[(2'h3):(2'h2)];
                      reg1794 <= {(reg1682 ? reg1487 : reg1607[(3'h5):(2'h3)])};
                    end
                end
            end
        end
    end
  assign wire1807 = $signed(forvar1744[(2'h2):(2'h2)]);
  assign wire1808 = $signed((~|(~&{(8'hb8)})));
  assign wire1809 = ({({reg1586} <= reg1546[(1'h0):(1'h0)])} ?
                        ((-reg1611) ?
                            ({(8'h9d)} ?
                                {reg1754} : $signed(forvar1585)) : reg1521) : (8'hb1));
  always
    @(posedge clk) begin
      for (forvar1810 = (1'h0); (forvar1810 < (1'h1)); forvar1810 = (forvar1810 + (1'h1)))
        begin
          for (forvar1811 = (1'h0); (forvar1811 < (1'h0)); forvar1811 = (forvar1811 + (1'h1)))
            begin
              if (forvar1762)
                begin
                  for (forvar1812 = (1'h0); (forvar1812 < (2'h3)); forvar1812 = (forvar1812 + (1'h1)))
                    begin
                      reg1813 <= forvar1653[(2'h3):(1'h0)];
                      reg1814 <= ($signed(reg1699) & $unsigned({(forvar1613 >= forvar1612)}));
                      reg1815 <= (forvar1755[(1'h1):(1'h0)] ?
                          ({{(8'haf)}} ?
                              {{reg1498}} : reg1629) : $signed(reg1814));
                      reg1816 <= {reg1800[(1'h0):(1'h0)]};
                    end
                  if (($unsigned($unsigned($unsigned(reg1480))) >> (reg1686[(3'h5):(1'h0)] >= reg1509[(3'h6):(2'h2)])))
                    begin
                      reg1817 <= reg1717[(3'h6):(2'h3)];
                      reg1818 <= (8'haa);
                    end
                  else
                    begin
                      reg1817 <= reg1532[(2'h3):(1'h0)];
                    end
                  for (forvar1819 = (1'h0); (forvar1819 < (1'h1)); forvar1819 = (forvar1819 + (1'h1)))
                    begin
                      reg1820 <= (!$signed((~^reg1806[(3'h5):(3'h5)])));
                      reg1821 <= {forvar1639};
                      reg1822 <= ((~reg1666) ?
                          (reg1577 < ($signed(reg1469) & (reg1627 | reg1736))) : ((~^(reg1651 || forvar1671)) ?
                              $unsigned(((8'hb8) ?
                                  forvar1485 : (8'haf))) : (~|reg1561[(4'h9):(3'h5)])));
                    end
                end
              else
                begin
                  for (forvar1812 = (1'h0); (forvar1812 < (2'h3)); forvar1812 = (forvar1812 + (1'h1)))
                    begin
                      reg1813 <= reg1485[(3'h6):(2'h3)];
                      reg1814 <= ((~^$unsigned((reg1574 ?
                          (8'h9d) : forvar1667))) <<< $signed(reg1487[(2'h3):(1'h0)]));
                    end
                end
              if ((~|(forvar1545[(3'h5):(2'h3)] ?
                  {$signed(forvar1666)} : reg1706)))
                begin
                  if ($unsigned(((+(8'hae)) ^~ (~^(forvar1603 >> forvar1671)))))
                    begin
                      reg1823 <= $unsigned({((~|reg1785) && (8'hac))});
                    end
                  else
                    begin
                      reg1823 <= ((&((~^reg1644) ?
                          $signed(forvar1470) : (reg1726 <= reg1486))) <= (($unsigned(reg1539) ?
                              forvar1612[(1'h0):(1'h0)] : (^reg1715)) ?
                          $unsigned(((8'h9d) ?
                              reg1773 : reg1774)) : (+(|reg1666))));
                      reg1824 <= ((~(~^(reg1458 ? reg1649 : reg1640))) ?
                          (((reg1520 && (8'hb4)) ?
                              forvar1736[(1'h1):(1'h1)] : forvar1550[(1'h1):(1'h0)]) >= $signed((reg1677 << reg1587))) : $signed($signed((reg1760 ?
                              forvar1791 : (8'ha0)))));
                    end
                end
              else
                begin
                  if (((8'ha1) <= {$unsigned($unsigned(wire3))}))
                    begin
                      reg1823 <= $unsigned((8'ha6));
                      reg1824 <= (reg1555 ? reg1504 : forvar1502);
                      reg1825 <= ((({reg1551} ?
                              (reg1686 ~^ reg1565) : (reg1528 != reg1636)) >= reg1551[(3'h4):(1'h0)]) ?
                          (reg1649 ?
                              reg1639[(4'hd):(3'h4)] : (|(~forvar1540))) : ($signed({(8'hb6)}) ?
                              ($unsigned(reg1699) ?
                                  reg1475 : $unsigned(reg1676)) : (^~(reg1792 >>> reg1466))));
                    end
                  else
                    begin
                      reg1823 <= (!(^$signed($unsigned(reg1787))));
                      reg1824 <= (reg1577 >> reg1509[(2'h3):(2'h2)]);
                      reg1825 <= $unsigned(forvar1762[(2'h2):(2'h2)]);
                      reg1826 <= (((-$signed(reg1639)) << $signed((reg1515 ?
                              reg1550 : reg1737))) ?
                          (!(forvar1705[(3'h5):(1'h1)] ?
                              reg1722 : $unsigned(reg1699))) : reg1658[(1'h1):(1'h1)]);
                    end
                end
              for (forvar1827 = (1'h0); (forvar1827 < (2'h2)); forvar1827 = (forvar1827 + (1'h1)))
                begin
                  for (forvar1828 = (1'h0); (forvar1828 < (2'h2)); forvar1828 = (forvar1828 + (1'h1)))
                    begin
                      reg1829 <= ({reg1657} > ((^reg1614[(1'h1):(1'h1)]) ?
                          $signed((&(8'ha2))) : ((8'hb9) ?
                              $signed((8'ha2)) : $unsigned(reg1645))));
                      reg1830 <= forvar1583;
                      reg1831 <= ($unsigned($signed((reg1592 ?
                          forvar1631 : reg1475))) ^ $unsigned(reg1550[(2'h2):(1'h1)]));
                    end
                  for (forvar1832 = (1'h0); (forvar1832 < (2'h2)); forvar1832 = (forvar1832 + (1'h1)))
                    begin
                      reg1833 <= ($signed($unsigned(reg1736[(3'h5):(1'h0)])) ?
                          (!reg1750) : ($signed($signed(reg1753)) ?
                              reg1766[(3'h4):(1'h1)] : (forvar1758[(3'h6):(2'h2)] && ((8'hb6) ?
                                  (8'ha0) : (8'haf)))));
                    end
                  if (((&$signed($unsigned(wire1451))) ?
                      reg1647[(2'h3):(1'h1)] : wire1809[(2'h2):(1'h1)]))
                    begin
                      reg1834 <= (-$unsigned((^(|reg1500))));
                      reg1835 <= (+(($unsigned(forvar1639) ?
                          reg1645 : {reg1555}) == ((reg1748 < (8'hb1)) ?
                          $signed(forvar1782) : reg1507[(4'h8):(2'h3)])));
                      reg1836 <= (8'had);
                      reg1837 <= (forvar1776[(2'h3):(1'h1)] ?
                          (((reg1586 ? reg1610 : (8'hb6)) ?
                              forvar1748 : $unsigned(reg1654)) <<< ((+forvar1470) ?
                              forvar1791[(2'h3):(1'h0)] : $unsigned(reg1471))) : (&$signed({reg1532})));
                    end
                  else
                    begin
                      reg1834 <= reg1648[(4'h8):(2'h3)];
                      reg1835 <= (|(-reg1628[(1'h0):(1'h0)]));
                    end
                end
              reg1838 <= (reg1530[(3'h7):(2'h3)] ?
                  (~|(reg1780[(1'h0):(1'h0)] ?
                      (reg1833 ?
                          reg1703 : reg1633) : $signed(reg1707))) : (^(forvar1755[(1'h0):(1'h0)] ?
                      ((8'hb1) ?
                          forvar1524 : reg1486) : (forvar1501 - forvar1470))));
            end
          if (reg1593)
            begin
              for (forvar1839 = (1'h0); (forvar1839 < (2'h2)); forvar1839 = (forvar1839 + (1'h1)))
                begin
                  reg1840 <= $signed(({reg1773} ?
                      ({forvar1529} ^ (reg1710 <= forvar1598)) : (8'ha1)));
                  for (forvar1841 = (1'h0); (forvar1841 < (2'h2)); forvar1841 = (forvar1841 + (1'h1)))
                    begin
                      reg1842 <= (reg1664[(2'h2):(1'h1)] ?
                          (-(((8'haf) ? reg1735 : forvar1712) || ((8'hb1) ?
                              reg1579 : reg1522))) : $signed(reg1637[(3'h7):(3'h6)]));
                      reg1843 <= (forvar1783[(4'h8):(3'h5)] - $signed($unsigned($unsigned(reg1656))));
                      reg1844 <= forvar1839;
                      reg1845 <= {((~&(|wire1809)) == $signed((reg1669 ?
                              reg1599 : reg1766)))};
                    end
                  reg1846 <= (&(reg1759 ~^ $signed({forvar1744})));
                end
              if (reg1515[(3'h4):(1'h0)])
                begin
                  if ((&(|(8'ha5))))
                    begin
                      reg1847 <= (~|((reg1660[(1'h0):(1'h0)] ?
                              reg1470[(2'h3):(1'h0)] : forvar1839[(2'h2):(1'h1)]) ?
                          (&(reg1825 ? reg1760 : (8'ha6))) : wire6));
                      reg1848 <= ((~&(8'h9d)) == ((8'h9e) <<< ($signed(forvar1598) ?
                          (reg1572 + (8'ha3)) : (reg1766 >> (8'hab)))));
                      reg1849 <= (&wire1453[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg1847 <= forvar1765;
                      reg1848 <= reg1621[(1'h0):(1'h0)];
                    end
                  for (forvar1850 = (1'h0); (forvar1850 < (2'h2)); forvar1850 = (forvar1850 + (1'h1)))
                    begin
                      reg1851 <= forvar1485;
                      reg1852 <= reg1647;
                      reg1853 <= $signed(((forvar1819 != (reg1606 * forvar1685)) ?
                          $unsigned(reg1792) : (reg1830 ~^ (-(8'ha4)))));
                      reg1854 <= $signed(forvar1768[(3'h5):(3'h5)]);
                    end
                end
              else
                begin
                  reg1847 <= ((^~($signed(reg1560) ?
                          {reg1526} : forvar1646[(4'hf):(4'hf)])) ?
                      (forvar1541 ?
                          {reg1455[(2'h3):(1'h1)]} : (~$signed(forvar1510))) : (^({forvar1758} - (|reg1480))));
                  if ((reg1718 + $signed(($unsigned(forvar1540) ?
                      (reg1795 ? (8'ha0) : reg1474) : ((8'ha2) ?
                          reg1684 : forvar1704)))))
                    begin
                      reg1848 <= (!reg1674);
                      reg1849 <= reg1563[(3'h4):(3'h4)];
                      reg1850 <= $signed(reg1777);
                      reg1851 <= reg1543[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg1848 <= (8'hb6);
                    end
                  for (forvar1852 = (1'h0); (forvar1852 < (1'h0)); forvar1852 = (forvar1852 + (1'h1)))
                    begin
                      reg1853 <= ((((|reg1465) ?
                          $signed(reg1829) : (8'h9c)) && reg1582) && reg1762);
                      reg1854 <= ($signed($unsigned(((8'had) ?
                          (8'ha4) : forvar1514))) + (forvar1482[(5'h10):(4'h8)] ?
                          ((reg1705 ?
                              reg1764 : (8'hb4)) >= reg1775[(3'h5):(2'h2)]) : $unsigned($unsigned((8'ha6)))));
                      reg1855 <= forvar1459;
                      reg1856 <= forvar1755[(1'h0):(1'h0)];
                    end
                  for (forvar1857 = (1'h0); (forvar1857 < (2'h2)); forvar1857 = (forvar1857 + (1'h1)))
                    begin
                      reg1858 <= reg1843[(3'h7):(2'h3)];
                    end
                end
              for (forvar1859 = (1'h0); (forvar1859 < (1'h0)); forvar1859 = (forvar1859 + (1'h1)))
                begin
                  for (forvar1860 = (1'h0); (forvar1860 < (2'h2)); forvar1860 = (forvar1860 + (1'h1)))
                    begin
                      reg1861 <= reg1622;
                      reg1862 <= reg1493[(2'h2):(1'h1)];
                      reg1863 <= (^(forvar1660[(3'h5):(2'h2)] <= $signed((reg1789 ?
                          forvar1736 : reg1668))));
                    end
                  for (forvar1864 = (1'h0); (forvar1864 < (2'h3)); forvar1864 = (forvar1864 + (1'h1)))
                    begin
                      reg1865 <= ((reg1744 ?
                          ((reg1690 ? (8'ha9) : forvar1752) ?
                              (reg1650 >>> reg1567) : (reg1728 ?
                                  (8'hae) : forvar1776)) : ($unsigned(reg1683) ?
                              $signed(forvar1613) : $signed(reg1717))) <<< ($unsigned((reg1552 ?
                              (8'haf) : forvar1662)) ?
                          reg1571 : {(forvar1482 ? reg1739 : reg1853)}));
                      reg1866 <= reg1496;
                      reg1867 <= ($unsigned(forvar1524[(2'h2):(1'h1)]) + (reg1729[(3'h4):(2'h2)] & {(reg1588 >= reg1767)}));
                      reg1868 <= {forvar1529};
                    end
                  reg1869 <= $signed($signed(reg1547[(4'h9):(4'h8)]));
                  for (forvar1870 = (1'h0); (forvar1870 < (1'h0)); forvar1870 = (forvar1870 + (1'h1)))
                    begin
                      reg1871 <= (~&$unsigned($unsigned($signed(reg1813))));
                      reg1872 <= $unsigned(($signed((&reg1719)) ?
                          reg1697[(3'h6):(3'h5)] : (|$unsigned(reg1724))));
                    end
                end
              for (forvar1873 = (1'h0); (forvar1873 < (2'h3)); forvar1873 = (forvar1873 + (1'h1)))
                begin
                  reg1874 <= (~|{$unsigned($unsigned(forvar1727))});
                  for (forvar1875 = (1'h0); (forvar1875 < (2'h3)); forvar1875 = (forvar1875 + (1'h1)))
                    begin
                      reg1876 <= (-(((^reg1663) ?
                          {forvar1785} : (reg1784 ?
                              reg1719 : forvar1683)) ^ (((8'hb2) ?
                          reg1697 : reg1546) ^~ ((8'h9c) + reg1848))));
                      reg1877 <= (($unsigned(reg1486[(1'h1):(1'h0)]) >>> (&$signed((8'hae)))) ^ $unsigned($unsigned(reg1516[(2'h2):(1'h0)])));
                    end
                end
            end
          else
            begin
              if ($unsigned(forvar1499[(3'h6):(1'h1)]))
                begin
                  if ($unsigned(($signed(reg1525[(2'h2):(2'h2)]) ^ $unsigned(reg1614[(3'h5):(1'h1)]))))
                    begin
                      reg1839 <= (($signed((reg1847 & forvar1510)) >> ($signed(forvar1873) || (reg1512 * forvar1827))) ?
                          $unsigned(forvar1502) : (((forvar1560 << forvar1577) ?
                              (reg1634 ?
                                  reg1668 : reg1599) : (^reg1540)) <= $signed((^reg1511))));
                      reg1840 <= reg1464;
                      reg1841 <= $signed((+$signed(((8'h9f) * forvar1721))));
                      reg1842 <= ((+($unsigned(reg1615) ?
                          (~|reg1463) : (-reg1509))) >> (((reg1837 ?
                              reg1508 : reg1709) >> reg1871) ?
                          (reg1796[(4'ha):(2'h3)] ?
                              reg1668[(4'h8):(2'h2)] : $signed(reg1650)) : forvar1752));
                    end
                  else
                    begin
                      reg1839 <= (reg1785[(3'h6):(1'h1)] << (!$unsigned($unsigned(forvar1641))));
                      reg1840 <= reg1656[(4'h9):(3'h7)];
                      reg1841 <= reg1731[(3'h6):(1'h0)];
                      reg1842 <= {$signed((~^$unsigned(forvar1630)))};
                    end
                  for (forvar1843 = (1'h0); (forvar1843 < (2'h3)); forvar1843 = (forvar1843 + (1'h1)))
                    begin
                      reg1844 <= {(((~&reg1741) || (forvar1762 ?
                                  reg1791 : reg1573)) ?
                              forvar1694 : reg1865[(3'h7):(3'h4)])};
                      reg1845 <= {{forvar1828}};
                    end
                end
              else
                begin
                  reg1839 <= $unsigned($signed((&$unsigned(reg1769))));
                  reg1840 <= $signed($signed(((~&forvar1534) ?
                      $signed(reg1667) : $unsigned(forvar1785))));
                end
              if ($signed($signed(((forvar1676 << forvar1860) ?
                  $unsigned(reg1467) : (8'ha2)))))
                begin
                  reg1846 <= ((reg1643[(1'h1):(1'h1)] && (^~(reg1760 < reg1697))) > $unsigned(reg1581));
                end
              else
                begin
                  if ($signed(({forvar1752[(2'h3):(1'h1)]} ?
                      (8'hab) : $signed(((8'ha3) <<< reg1492)))))
                    begin
                      reg1846 <= (((^$unsigned((8'h9f))) <= $signed(((8'hb2) ?
                              reg1749 : (8'hb7)))) ?
                          (&$unsigned(reg1677)) : $unsigned(reg1469[(2'h3):(1'h1)]));
                      reg1847 <= $signed(forvar1819[(3'h4):(2'h3)]);
                    end
                  else
                    begin
                      reg1846 <= reg1768;
                      reg1847 <= (^~{$unsigned($unsigned(reg1765))});
                      reg1848 <= forvar1873;
                    end
                  if (($unsigned($unsigned({(8'ha9)})) ?
                      (~^$unsigned($unsigned(reg1737))) : reg1690))
                    begin
                      reg1849 <= $unsigned((($unsigned(forvar1734) >>> reg1621[(2'h3):(2'h2)]) <= (^~$unsigned(reg1563))));
                      reg1850 <= (~&reg1831[(1'h0):(1'h0)]);
                      reg1851 <= reg1805;
                    end
                  else
                    begin
                      reg1849 <= $signed(((-(wire0 ? reg1508 : reg1457)) ?
                          (reg1756[(4'h9):(3'h7)] << (forvar1721 | reg1493)) : (-reg1592)));
                      reg1850 <= $signed(reg1547[(1'h1):(1'h1)]);
                      reg1851 <= {((((8'ha1) ?
                                  reg1647 : forvar1538) ^~ reg1689[(3'h4):(1'h0)]) ?
                              forvar1538[(1'h0):(1'h0)] : {forvar1454[(2'h3):(1'h1)]})};
                      reg1852 <= ($signed(forvar1518) != {((forvar1486 ?
                              reg1523 : reg1744) * reg1696[(1'h0):(1'h0)])});
                    end
                end
              reg1853 <= forvar1639;
            end
          for (forvar1878 = (1'h0); (forvar1878 < (2'h3)); forvar1878 = (forvar1878 + (1'h1)))
            begin
              for (forvar1879 = (1'h0); (forvar1879 < (1'h0)); forvar1879 = (forvar1879 + (1'h1)))
                begin
                  for (forvar1880 = (1'h0); (forvar1880 < (2'h3)); forvar1880 = (forvar1880 + (1'h1)))
                    begin
                      reg1881 <= wire4;
                      reg1882 <= (^~$signed(reg1540));
                    end
                end
            end
          for (forvar1883 = (1'h0); (forvar1883 < (2'h2)); forvar1883 = (forvar1883 + (1'h1)))
            begin
              for (forvar1884 = (1'h0); (forvar1884 < (2'h2)); forvar1884 = (forvar1884 + (1'h1)))
                begin
                  for (forvar1885 = (1'h0); (forvar1885 < (1'h1)); forvar1885 = (forvar1885 + (1'h1)))
                    begin
                      reg1886 <= $signed(reg1532[(3'h7):(3'h6)]);
                      reg1887 <= $unsigned(($unsigned($unsigned(forvar1748)) ?
                          ($signed(forvar1626) * {reg1622}) : reg1724[(3'h6):(3'h5)]));
                      reg1888 <= ((reg1513[(2'h2):(1'h1)] <<< reg1497[(2'h2):(1'h1)]) < reg1544);
                    end
                  if (($signed((reg1582 << (reg1570 == reg1477))) != $signed($unsigned(forvar1631))))
                    begin
                      reg1889 <= reg1786[(2'h2):(2'h2)];
                      reg1890 <= $signed((~^$unsigned({forvar1734})));
                      reg1891 <= ((reg1486[(2'h2):(1'h1)] ^ ((reg1699 >= forvar1682) && $signed(reg1715))) <= (reg1692 ?
                          reg1840[(4'hc):(2'h3)] : $signed($unsigned(forvar1758))));
                      reg1892 <= $unsigned($signed(reg1702));
                    end
                  else
                    begin
                      reg1889 <= (({$unsigned(forvar1533)} | $signed(((8'hac) || reg1592))) ?
                          ({(reg1565 ? forvar1755 : (8'had))} ?
                              $unsigned(((8'h9f) >>> reg1750)) : (^(reg1725 ?
                                  reg1771 : reg1572))) : reg1628[(1'h1):(1'h0)]);
                    end
                  reg1893 <= ((forvar1883[(3'h4):(2'h2)] ?
                      {reg1815} : (|(reg1813 & forvar1884))) <= $unsigned($unsigned((reg1570 != (8'hb8)))));
                end
              for (forvar1894 = (1'h0); (forvar1894 < (2'h3)); forvar1894 = (forvar1894 + (1'h1)))
                begin
                  for (forvar1895 = (1'h0); (forvar1895 < (1'h1)); forvar1895 = (forvar1895 + (1'h1)))
                    begin
                      reg1896 <= ((~wire3) ?
                          $unsigned(reg1699[(4'h9):(4'h8)]) : $unsigned((^~((8'ha4) <<< forvar1811))));
                      reg1897 <= forvar1776[(2'h3):(1'h1)];
                      reg1898 <= $signed($signed(({reg1740} & reg1578[(2'h3):(2'h2)])));
                    end
                end
              for (forvar1899 = (1'h0); (forvar1899 < (2'h3)); forvar1899 = (forvar1899 + (1'h1)))
                begin
                  reg1900 <= (reg1660 ~^ $signed(wire1618[(2'h2):(2'h2)]));
                  for (forvar1901 = (1'h0); (forvar1901 < (1'h1)); forvar1901 = (forvar1901 + (1'h1)))
                    begin
                      reg1902 <= (^~$signed(forvar1631));
                    end
                end
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1297  (y, clk, wire1302, wire1301, wire1300, wire1299, wire1298);
  output wire [(32'h60c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire1302;
  input wire signed [(3'h4):(1'h0)] wire1301;
  input wire signed [(5'h10):(1'h0)] wire1300;
  input wire signed [(4'ha):(1'h0)] wire1299;
  input wire signed [(3'h4):(1'h0)] wire1298;
  wire signed [(3'h7):(1'h0)] wire1450;
  wire [(4'hb):(1'h0)] wire1449;
  reg signed [(4'hd):(1'h0)] reg1448 = (1'h0);
  reg [(4'h9):(1'h0)] reg1447 = (1'h0);
  reg [(3'h7):(1'h0)] reg1440 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1437 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1431 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1442 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1446 = (1'h0);
  reg [(2'h3):(1'h0)] reg1445 = (1'h0);
  reg [(2'h2):(1'h0)] reg1444 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1443 = (1'h0);
  reg [(4'hc):(1'h0)] reg1442 = (1'h0);
  reg [(3'h6):(1'h0)] reg1441 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1440 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1439 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1432 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1438 = (1'h0);
  reg [(2'h3):(1'h0)] reg1437 = (1'h0);
  reg [(4'he):(1'h0)] reg1436 = (1'h0);
  reg [(4'hd):(1'h0)] reg1435 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1434 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1433 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1432 = (1'h0);
  reg [(4'hb):(1'h0)] reg1431 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1430 = (1'h0);
  reg [(3'h6):(1'h0)] reg1415 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1413 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1412 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1429 = (1'h0);
  reg [(2'h3):(1'h0)] reg1428 = (1'h0);
  reg [(3'h4):(1'h0)] reg1427 = (1'h0);
  reg [(3'h7):(1'h0)] reg1426 = (1'h0);
  reg [(4'ha):(1'h0)] reg1425 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1419 = (1'h0);
  reg [(4'he):(1'h0)] reg1424 = (1'h0);
  reg [(3'h6):(1'h0)] reg1423 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1422 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1421 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1420 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1419 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1418 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1417 = (1'h0);
  reg [(4'h9):(1'h0)] reg1416 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1415 = (1'h0);
  reg [(4'h8):(1'h0)] reg1414 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1413 = (1'h0);
  reg [(4'hf):(1'h0)] reg1412 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1411 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1410 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1409 = (1'h0);
  reg [(2'h3):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1407 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1406 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1405 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1404 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1403 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1402 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1401 = (1'h0);
  reg [(4'hf):(1'h0)] reg1400 = (1'h0);
  reg [(4'h8):(1'h0)] reg1399 = (1'h0);
  reg [(4'hd):(1'h0)] reg1398 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1397 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1396 = (1'h0);
  reg [(3'h4):(1'h0)] reg1395 = (1'h0);
  reg [(2'h3):(1'h0)] reg1394 = (1'h0);
  reg [(3'h4):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1392 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1391 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1390 = (1'h0);
  reg [(3'h7):(1'h0)] reg1389 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1388 = (1'h0);
  reg [(4'ha):(1'h0)] reg1387 = (1'h0);
  reg [(2'h2):(1'h0)] reg1386 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1385 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1384 = (1'h0);
  reg [(5'h10):(1'h0)] reg1383 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1382 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1381 = (1'h0);
  reg [(3'h6):(1'h0)] reg1380 = (1'h0);
  reg [(4'hb):(1'h0)] reg1379 = (1'h0);
  reg [(4'hd):(1'h0)] reg1378 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1377 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1376 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1375 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1374 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1373 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1372 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1371 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1370 = (1'h0);
  reg [(4'ha):(1'h0)] reg1369 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1368 = (1'h0);
  reg [(3'h4):(1'h0)] reg1367 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1364 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1357 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1354 = (1'h0);
  reg [(4'hd):(1'h0)] reg1361 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1353 = (1'h0);
  reg [(3'h7):(1'h0)] reg1351 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1349 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1366 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1365 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1364 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1363 = (1'h0);
  reg [(4'hc):(1'h0)] reg1362 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1361 = (1'h0);
  reg [(4'hc):(1'h0)] reg1360 = (1'h0);
  reg [(3'h7):(1'h0)] reg1359 = (1'h0);
  reg [(4'he):(1'h0)] reg1358 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1357 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1356 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1355 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1354 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1353 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1352 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1351 = (1'h0);
  reg [(2'h3):(1'h0)] reg1350 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1349 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1348 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1347 = (1'h0);
  reg [(3'h4):(1'h0)] reg1346 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1345 = (1'h0);
  reg [(4'hd):(1'h0)] reg1337 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1334 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1333 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1332 = (1'h0);
  reg [(4'h9):(1'h0)] reg1344 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1343 = (1'h0);
  reg [(5'h10):(1'h0)] reg1342 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1341 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1340 = (1'h0);
  reg [(4'hd):(1'h0)] reg1339 = (1'h0);
  reg [(3'h7):(1'h0)] reg1338 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1337 = (1'h0);
  reg [(4'h9):(1'h0)] reg1336 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1335 = (1'h0);
  reg [(3'h6):(1'h0)] reg1334 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1333 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1332 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1331 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1330 = (1'h0);
  reg [(3'h7):(1'h0)] reg1329 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1321 = (1'h0);
  reg [(4'ha):(1'h0)] reg1318 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1317 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1314 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1313 = (1'h0);
  reg [(3'h7):(1'h0)] reg1312 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1311 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1308 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1304 = (1'h0);
  reg [(4'hf):(1'h0)] reg1328 = (1'h0);
  reg [(4'h9):(1'h0)] reg1327 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1326 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1325 = (1'h0);
  reg [(4'h9):(1'h0)] reg1324 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1323 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1322 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1321 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1320 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1319 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1318 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1317 = (1'h0);
  reg [(4'he):(1'h0)] reg1316 = (1'h0);
  reg [(3'h5):(1'h0)] reg1315 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1314 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1313 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1312 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1311 = (1'h0);
  reg [(4'hb):(1'h0)] reg1310 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1309 = (1'h0);
  reg [(4'h9):(1'h0)] reg1308 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1307 = (1'h0);
  reg [(4'hd):(1'h0)] reg1306 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1305 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1304 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1303 = (1'h0);
  assign y = {wire1450,
                 wire1449,
                 reg1448,
                 reg1447,
                 reg1440,
                 forvar1437,
                 forvar1431,
                 forvar1442,
                 reg1446,
                 reg1445,
                 reg1444,
                 reg1443,
                 reg1442,
                 reg1441,
                 forvar1440,
                 reg1439,
                 reg1432,
                 reg1438,
                 reg1437,
                 reg1436,
                 reg1435,
                 reg1434,
                 reg1433,
                 forvar1432,
                 reg1431,
                 forvar1430,
                 reg1415,
                 forvar1413,
                 forvar1412,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 reg1425,
                 forvar1419,
                 reg1424,
                 reg1423,
                 reg1422,
                 reg1421,
                 reg1420,
                 reg1419,
                 reg1418,
                 reg1417,
                 reg1416,
                 forvar1415,
                 reg1414,
                 reg1413,
                 reg1412,
                 reg1411,
                 forvar1410,
                 reg1409,
                 reg1408,
                 reg1407,
                 forvar1406,
                 forvar1405,
                 forvar1404,
                 reg1403,
                 reg1402,
                 forvar1401,
                 reg1400,
                 reg1399,
                 reg1398,
                 forvar1397,
                 reg1396,
                 reg1395,
                 reg1394,
                 reg1393,
                 reg1392,
                 forvar1391,
                 reg1390,
                 reg1389,
                 reg1388,
                 reg1387,
                 reg1386,
                 forvar1385,
                 forvar1384,
                 reg1383,
                 forvar1382,
                 reg1381,
                 reg1380,
                 reg1379,
                 reg1378,
                 forvar1377,
                 reg1376,
                 reg1375,
                 reg1374,
                 reg1373,
                 forvar1372,
                 forvar1371,
                 forvar1370,
                 reg1369,
                 reg1368,
                 reg1367,
                 forvar1364,
                 reg1357,
                 reg1354,
                 reg1361,
                 reg1353,
                 reg1351,
                 forvar1349,
                 reg1366,
                 reg1365,
                 reg1364,
                 reg1363,
                 reg1362,
                 forvar1361,
                 reg1360,
                 reg1359,
                 reg1358,
                 forvar1357,
                 reg1356,
                 reg1355,
                 forvar1354,
                 forvar1353,
                 reg1352,
                 forvar1351,
                 reg1350,
                 reg1349,
                 reg1348,
                 forvar1347,
                 reg1346,
                 forvar1345,
                 reg1337,
                 forvar1334,
                 reg1333,
                 reg1332,
                 reg1344,
                 reg1343,
                 reg1342,
                 reg1341,
                 forvar1340,
                 reg1339,
                 reg1338,
                 forvar1337,
                 reg1336,
                 forvar1335,
                 reg1334,
                 forvar1333,
                 forvar1332,
                 forvar1331,
                 reg1330,
                 reg1329,
                 forvar1321,
                 reg1318,
                 forvar1317,
                 forvar1314,
                 reg1313,
                 reg1312,
                 forvar1311,
                 forvar1308,
                 forvar1304,
                 reg1328,
                 reg1327,
                 reg1326,
                 forvar1325,
                 reg1324,
                 reg1323,
                 reg1322,
                 reg1321,
                 reg1320,
                 reg1319,
                 forvar1318,
                 reg1317,
                 reg1316,
                 reg1315,
                 reg1314,
                 forvar1313,
                 forvar1312,
                 reg1311,
                 reg1310,
                 reg1309,
                 reg1308,
                 reg1307,
                 reg1306,
                 reg1305,
                 reg1304,
                 forvar1303,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar1303 = (1'h0); (forvar1303 < (1'h1)); forvar1303 = (forvar1303 + (1'h1)))
        begin
          if (wire1301[(2'h3):(2'h3)])
            begin
              reg1304 <= $unsigned($unsigned(wire1301[(1'h0):(1'h0)]));
              if ($signed(($signed(wire1298) ?
                  (!wire1300) : (wire1300 ^~ (forvar1303 ?
                      (8'hb2) : (8'ha5))))))
                begin
                  reg1305 <= {((~reg1304[(2'h2):(1'h0)]) + $signed((wire1299 != (8'ha9))))};
                  if ($signed(wire1302))
                    begin
                      reg1306 <= (^reg1305);
                      reg1307 <= $signed($unsigned(wire1301[(1'h0):(1'h0)]));
                      reg1308 <= ((($unsigned(reg1306) >= $signed(wire1299)) & $signed((~&reg1305))) ?
                          wire1298[(1'h0):(1'h0)] : (forvar1303 <<< (^$unsigned(wire1302))));
                      reg1309 <= (+(wire1299[(4'ha):(4'ha)] ?
                          (wire1301[(2'h2):(2'h2)] ?
                              wire1299[(4'ha):(3'h6)] : (&wire1299)) : reg1306[(4'hb):(4'hb)]));
                    end
                  else
                    begin
                      reg1306 <= (^(8'ha2));
                      reg1307 <= (($unsigned(wire1300) + (wire1300[(4'hd):(4'h8)] ?
                              (~&reg1304) : $unsigned(wire1300))) ?
                          $unsigned({$unsigned(wire1299)}) : (~(~^$signed((8'ha8)))));
                    end
                end
              else
                begin
                  reg1305 <= $signed(reg1307[(1'h1):(1'h1)]);
                  reg1306 <= $unsigned(reg1304);
                  if ($signed(reg1306[(1'h0):(1'h0)]))
                    begin
                      reg1307 <= (^reg1304[(1'h1):(1'h1)]);
                      reg1308 <= ((($unsigned((8'h9c)) << reg1304) ?
                              $signed(reg1307[(1'h1):(1'h0)]) : $unsigned(wire1301[(2'h3):(1'h0)])) ?
                          (~&(!((8'h9e) ?
                              reg1307 : reg1309))) : ({(|wire1300)} | reg1309[(2'h2):(2'h2)]));
                      reg1309 <= $unsigned((^$unsigned((wire1300 < wire1298))));
                      reg1310 <= (^~$signed(wire1300));
                    end
                  else
                    begin
                      reg1307 <= {$signed((|$unsigned(reg1309)))};
                    end
                  reg1311 <= ((|((wire1298 ? wire1299 : wire1300) ?
                          (reg1305 || (8'h9f)) : wire1298[(2'h2):(1'h1)])) ?
                      ({wire1300[(1'h1):(1'h0)]} ?
                          ($signed(wire1298) == (wire1302 ?
                              (8'hab) : wire1299)) : ((reg1308 != wire1300) * reg1306)) : wire1302[(2'h3):(1'h0)]);
                end
              for (forvar1312 = (1'h0); (forvar1312 < (2'h2)); forvar1312 = (forvar1312 + (1'h1)))
                begin
                  for (forvar1313 = (1'h0); (forvar1313 < (1'h0)); forvar1313 = (forvar1313 + (1'h1)))
                    begin
                      reg1314 <= {{{(|(8'hb7))}}};
                      reg1315 <= reg1306;
                      reg1316 <= {$signed((+((8'ha3) ? reg1311 : reg1314)))};
                      reg1317 <= (((reg1311 ^~ (~^reg1307)) > wire1301[(2'h3):(2'h2)]) >= ((!reg1304) ?
                          ((reg1310 ? wire1298 : reg1308) ?
                              reg1304 : (8'hb8)) : (reg1308 > reg1304[(1'h0):(1'h0)])));
                    end
                  for (forvar1318 = (1'h0); (forvar1318 < (2'h2)); forvar1318 = (forvar1318 + (1'h1)))
                    begin
                      reg1319 <= (reg1304 ?
                          {wire1298} : $signed({(forvar1303 * wire1298)}));
                      reg1320 <= $signed((8'hb3));
                      reg1321 <= (reg1317[(1'h1):(1'h0)] | reg1310[(4'ha):(3'h5)]);
                      reg1322 <= forvar1318[(2'h2):(1'h0)];
                    end
                  if (reg1307[(1'h0):(1'h0)])
                    begin
                      reg1323 <= $unsigned($signed(($unsigned((8'hb5)) ?
                          reg1314[(2'h2):(1'h1)] : (reg1314 >> (8'ha7)))));
                    end
                  else
                    begin
                      reg1323 <= reg1314;
                      reg1324 <= reg1315;
                    end
                  for (forvar1325 = (1'h0); (forvar1325 < (1'h0)); forvar1325 = (forvar1325 + (1'h1)))
                    begin
                      reg1326 <= ($unsigned((-$unsigned(reg1309))) ?
                          ($signed((reg1319 ~^ reg1322)) > $signed((~^forvar1303))) : (((reg1323 ?
                                  reg1316 : forvar1303) ^~ (~|reg1315)) ?
                              $unsigned((reg1323 & reg1324)) : (((8'ha6) ?
                                  forvar1318 : wire1301) || (~reg1306))));
                      reg1327 <= ((~((~(8'h9e)) | $unsigned(forvar1312))) <<< (8'h9c));
                      reg1328 <= (wire1302 || $signed($unsigned((!(8'hac)))));
                    end
                end
            end
          else
            begin
              for (forvar1304 = (1'h0); (forvar1304 < (1'h1)); forvar1304 = (forvar1304 + (1'h1)))
                begin
                  if (((((reg1314 <<< reg1324) ^ reg1308) ?
                      reg1327[(2'h3):(2'h3)] : (reg1305[(2'h2):(1'h1)] ?
                          (reg1320 ^ wire1299) : (+forvar1312))) ^~ {$signed((reg1328 ?
                          (8'h9f) : (8'haa)))}))
                    begin
                      reg1305 <= (8'hae);
                      reg1306 <= (8'ha7);
                      reg1307 <= wire1298[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1305 <= (reg1316[(4'hb):(1'h0)] < $signed($signed(reg1317)));
                    end
                  for (forvar1308 = (1'h0); (forvar1308 < (1'h0)); forvar1308 = (forvar1308 + (1'h1)))
                    begin
                      reg1309 <= $unsigned(reg1316);
                    end
                end
              reg1310 <= $unsigned(({forvar1318} << (((8'hb2) >>> (8'haa)) ^ (forvar1325 <= reg1308))));
              if (($signed((|forvar1313)) ?
                  (((-reg1324) ?
                      {reg1310} : (^reg1315)) * $signed($unsigned(wire1300))) : (~|reg1309)))
                begin
                  for (forvar1311 = (1'h0); (forvar1311 < (1'h0)); forvar1311 = (forvar1311 + (1'h1)))
                    begin
                      reg1312 <= ($signed((~&reg1307[(2'h2):(1'h0)])) + ($unsigned((reg1327 ?
                          reg1305 : forvar1303)) & ((&reg1328) || wire1298)));
                      reg1313 <= (+wire1299[(1'h1):(1'h0)]);
                    end
                  for (forvar1314 = (1'h0); (forvar1314 < (1'h1)); forvar1314 = (forvar1314 + (1'h1)))
                    begin
                      reg1315 <= (-(~((~^reg1305) << (8'h9f))));
                    end
                  reg1316 <= {$signed(($signed(forvar1311) - reg1321))};
                end
              else
                begin
                  if ((reg1316 ?
                      ((forvar1303[(4'hc):(4'hc)] <= (8'ha4)) >>> reg1308[(3'h7):(2'h2)]) : $signed($unsigned((forvar1314 ?
                          reg1322 : forvar1318)))))
                    begin
                      reg1311 <= (^~($signed(forvar1308) ?
                          forvar1304 : $signed($unsigned(wire1301))));
                    end
                  else
                    begin
                      reg1311 <= reg1311[(2'h2):(1'h0)];
                      reg1312 <= $signed($signed(($unsigned((8'ha5)) ?
                          $signed(reg1323) : (~^reg1309))));
                      reg1313 <= (reg1314[(1'h1):(1'h1)] ?
                          forvar1308 : wire1301);
                      reg1314 <= $signed(reg1313[(3'h7):(3'h5)]);
                    end
                  if (reg1310)
                    begin
                      reg1315 <= forvar1318;
                      reg1316 <= forvar1325;
                    end
                  else
                    begin
                      reg1315 <= wire1298;
                      reg1316 <= (^~$signed(wire1302));
                    end
                  for (forvar1317 = (1'h0); (forvar1317 < (1'h0)); forvar1317 = (forvar1317 + (1'h1)))
                    begin
                      reg1318 <= reg1309;
                      reg1319 <= $unsigned((~^((reg1306 > reg1314) <= $signed(reg1311))));
                      reg1320 <= reg1318[(3'h5):(1'h0)];
                    end
                  for (forvar1321 = (1'h0); (forvar1321 < (2'h3)); forvar1321 = (forvar1321 + (1'h1)))
                    begin
                      reg1322 <= $signed(reg1323);
                    end
                end
            end
          reg1329 <= forvar1321[(1'h1):(1'h1)];
          reg1330 <= (8'hab);
        end
      for (forvar1331 = (1'h0); (forvar1331 < (2'h3)); forvar1331 = (forvar1331 + (1'h1)))
        begin
          if ((!(!(^$unsigned(wire1299)))))
            begin
              for (forvar1332 = (1'h0); (forvar1332 < (1'h1)); forvar1332 = (forvar1332 + (1'h1)))
                begin
                  for (forvar1333 = (1'h0); (forvar1333 < (2'h2)); forvar1333 = (forvar1333 + (1'h1)))
                    begin
                      reg1334 <= (reg1312 && {forvar1317[(4'hc):(3'h6)]});
                    end
                  for (forvar1335 = (1'h0); (forvar1335 < (1'h0)); forvar1335 = (forvar1335 + (1'h1)))
                    begin
                      reg1336 <= $unsigned($unsigned($unsigned((8'h9f))));
                    end
                  for (forvar1337 = (1'h0); (forvar1337 < (1'h1)); forvar1337 = (forvar1337 + (1'h1)))
                    begin
                      reg1338 <= (~^($unsigned(reg1319[(2'h2):(1'h0)]) ^ {$signed(reg1315)}));
                      reg1339 <= $signed((((forvar1325 ~^ forvar1331) ?
                              forvar1321[(1'h1):(1'h1)] : reg1309) ?
                          (((8'ha1) ? forvar1313 : wire1298) ?
                              (~^reg1309) : (reg1330 ?
                                  reg1322 : wire1301)) : (forvar1304 << (wire1300 < reg1315))));
                    end
                  for (forvar1340 = (1'h0); (forvar1340 < (1'h0)); forvar1340 = (forvar1340 + (1'h1)))
                    begin
                      reg1341 <= (reg1309 ?
                          $signed((~|$signed(reg1314))) : ($signed((reg1329 ?
                              forvar1318 : forvar1313)) >> {$signed((8'h9c))}));
                      reg1342 <= ($signed(reg1322[(1'h0):(1'h0)]) ?
                          wire1300[(4'he):(4'h8)] : forvar1311[(1'h1):(1'h1)]);
                      reg1343 <= {$unsigned($signed($signed(reg1339)))};
                    end
                end
              reg1344 <= $signed(({reg1320} & reg1342));
            end
          else
            begin
              reg1332 <= (forvar1331 ?
                  (($signed(reg1329) ?
                      reg1324[(1'h0):(1'h0)] : {forvar1312}) ~^ ($signed(reg1328) ?
                      (forvar1313 ^~ reg1318) : (reg1344 - (8'ha3)))) : $unsigned($signed($signed(reg1323))));
              reg1333 <= reg1334[(1'h1):(1'h0)];
              for (forvar1334 = (1'h0); (forvar1334 < (2'h3)); forvar1334 = (forvar1334 + (1'h1)))
                begin
                  for (forvar1335 = (1'h0); (forvar1335 < (2'h3)); forvar1335 = (forvar1335 + (1'h1)))
                    begin
                      reg1336 <= $signed((!($signed(forvar1333) ?
                          ((8'h9c) & (8'hb0)) : (&forvar1335))));
                    end
                  if (((reg1304[(1'h1):(1'h0)] ?
                      reg1341[(1'h0):(1'h0)] : reg1304[(1'h1):(1'h1)]) >= reg1320[(1'h0):(1'h0)]))
                    begin
                      reg1337 <= reg1314[(1'h0):(1'h0)];
                      reg1338 <= reg1343;
                      reg1339 <= (reg1337 ?
                          $unsigned({{wire1298}}) : reg1318[(4'h9):(3'h7)]);
                    end
                  else
                    begin
                      reg1337 <= {(|$unsigned($unsigned((8'hb1))))};
                      reg1338 <= $signed($unsigned(reg1315));
                      reg1339 <= $unsigned(reg1338[(2'h2):(1'h1)]);
                    end
                  for (forvar1340 = (1'h0); (forvar1340 < (1'h1)); forvar1340 = (forvar1340 + (1'h1)))
                    begin
                      reg1341 <= (forvar1314 ?
                          ((|(reg1339 ? forvar1311 : (8'hb7))) ?
                              reg1314[(1'h1):(1'h1)] : ((reg1315 ?
                                      wire1300 : wire1302) ?
                                  ((8'hba) <= reg1316) : forvar1333[(1'h0):(1'h0)])) : (+((reg1326 & forvar1303) != forvar1334[(3'h5):(3'h5)])));
                      reg1342 <= (8'hb1);
                    end
                end
            end
          for (forvar1345 = (1'h0); (forvar1345 < (1'h0)); forvar1345 = (forvar1345 + (1'h1)))
            begin
              reg1346 <= $signed($signed($signed($signed(reg1316))));
              for (forvar1347 = (1'h0); (forvar1347 < (1'h1)); forvar1347 = (forvar1347 + (1'h1)))
                begin
                  reg1348 <= $unsigned((|$signed($unsigned(reg1326))));
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed($unsigned($signed(reg1310))))
        begin
          reg1349 <= forvar1303[(1'h1):(1'h0)];
          reg1350 <= reg1346[(2'h3):(2'h3)];
          for (forvar1351 = (1'h0); (forvar1351 < (2'h3)); forvar1351 = (forvar1351 + (1'h1)))
            begin
              reg1352 <= (~^reg1329[(1'h0):(1'h0)]);
              for (forvar1353 = (1'h0); (forvar1353 < (1'h1)); forvar1353 = (forvar1353 + (1'h1)))
                begin
                  for (forvar1354 = (1'h0); (forvar1354 < (1'h1)); forvar1354 = (forvar1354 + (1'h1)))
                    begin
                      reg1355 <= (reg1333[(2'h3):(1'h1)] ?
                          $unsigned(($signed(reg1338) && $unsigned(reg1307))) : $signed((forvar1317 ?
                              wire1300[(4'h9):(3'h5)] : $signed(forvar1321))));
                      reg1356 <= $signed(($signed((forvar1337 * reg1349)) && reg1322));
                    end
                end
              for (forvar1357 = (1'h0); (forvar1357 < (2'h3)); forvar1357 = (forvar1357 + (1'h1)))
                begin
                  if ((forvar1334[(3'h4):(3'h4)] ?
                      ((^~$unsigned(reg1312)) >= forvar1311) : (reg1323 ?
                          ((&(8'hb8)) ^ (~&(8'hae))) : ($unsigned((8'h9e)) ?
                              $unsigned(reg1342) : reg1305[(2'h2):(2'h2)]))))
                    begin
                      reg1358 <= reg1330[(1'h1):(1'h1)];
                      reg1359 <= ((((forvar1331 >= (8'hb4)) >= $unsigned(reg1314)) && $signed(forvar1347)) >= $unsigned($signed($unsigned((8'h9e)))));
                    end
                  else
                    begin
                      reg1358 <= $unsigned(($signed(forvar1312[(1'h1):(1'h0)]) + $signed(reg1338)));
                      reg1359 <= (^~reg1308[(2'h3):(2'h2)]);
                      reg1360 <= reg1346;
                    end
                  for (forvar1361 = (1'h0); (forvar1361 < (1'h0)); forvar1361 = (forvar1361 + (1'h1)))
                    begin
                      reg1362 <= $signed(reg1327[(3'h7):(3'h4)]);
                      reg1363 <= ($unsigned((reg1305[(3'h5):(3'h4)] >= reg1310[(1'h1):(1'h0)])) ?
                          $signed({(~&reg1350)}) : ($signed($unsigned(reg1362)) + (!$signed(reg1307))));
                      reg1364 <= forvar1340;
                      reg1365 <= $signed({$signed(reg1343)});
                    end
                  reg1366 <= reg1349[(2'h3):(1'h1)];
                end
            end
        end
      else
        begin
          if ($signed(((|(&reg1348)) & reg1337[(4'hb):(3'h4)])))
            begin
              for (forvar1349 = (1'h0); (forvar1349 < (2'h2)); forvar1349 = (forvar1349 + (1'h1)))
                begin
                  if ((!reg1305))
                    begin
                      reg1350 <= $signed(((reg1356 >>> (|reg1326)) <= {forvar1325[(2'h3):(1'h0)]}));
                      reg1351 <= (|($signed({(8'hb0)}) >= reg1339[(3'h7):(1'h0)]));
                      reg1352 <= (reg1346[(3'h4):(1'h0)] ?
                          {((forvar1334 ?
                                  reg1346 : reg1342) != (forvar1354 ~^ reg1329))} : (^forvar1331));
                    end
                  else
                    begin
                      reg1350 <= ($unsigned(((reg1337 ? forvar1345 : (8'hb5)) ?
                              (forvar1357 && reg1320) : {forvar1333})) ?
                          (forvar1303 || reg1342[(1'h1):(1'h0)]) : (!(((8'hba) <= reg1312) > (reg1306 ?
                              (8'ha6) : reg1344))));
                      reg1351 <= ((-($unsigned(forvar1331) ?
                              ((8'ha9) ^ forvar1334) : ((8'ha5) >>> forvar1333))) ?
                          (~|(((8'h9f) <= (8'hb9)) ?
                              (+reg1309) : ((8'hb0) ?
                                  forvar1353 : reg1336))) : ($signed((&forvar1354)) ?
                              (reg1318 >= reg1350) : $signed((^reg1349))));
                      reg1352 <= reg1328;
                      reg1353 <= $unsigned((+(!forvar1304)));
                    end
                end
              if ((~|forvar1333[(1'h1):(1'h1)]))
                begin
                  for (forvar1354 = (1'h0); (forvar1354 < (2'h2)); forvar1354 = (forvar1354 + (1'h1)))
                    begin
                      reg1355 <= ($unsigned(forvar1332) ?
                          (+$unsigned(reg1342)) : (forvar1313 ~^ $signed(reg1351)));
                    end
                  reg1356 <= wire1301;
                  for (forvar1357 = (1'h0); (forvar1357 < (1'h1)); forvar1357 = (forvar1357 + (1'h1)))
                    begin
                      reg1358 <= ($unsigned($signed(reg1320[(2'h2):(1'h1)])) ?
                          ($unsigned(reg1323[(1'h1):(1'h1)]) << ((8'ha6) ?
                              (forvar1312 - (8'hac)) : (wire1300 ?
                                  reg1338 : reg1304))) : $unsigned(((~forvar1331) << $signed((8'hb5)))));
                      reg1359 <= {$unsigned((reg1339[(3'h7):(2'h2)] ?
                              $signed(reg1348) : (reg1364 << forvar1354)))};
                      reg1360 <= ((8'ha7) ?
                          ($unsigned(forvar1331) >> forvar1325) : reg1315);
                    end
                  reg1361 <= (($signed((reg1366 ?
                      reg1348 : forvar1340)) >= ((8'ha1) ?
                      forvar1303[(4'h8):(3'h6)] : $signed(forvar1325))) & $signed(((forvar1314 ?
                          reg1313 : reg1349) ?
                      forvar1304[(4'h8):(1'h1)] : reg1356[(3'h5):(2'h3)])));
                end
              else
                begin
                  reg1354 <= (~reg1320);
                  reg1355 <= (((+$unsigned(forvar1333)) ?
                          ($unsigned(reg1332) ~^ reg1309) : ({(8'hb6)} & forvar1314)) ?
                      reg1354[(2'h2):(1'h1)] : (reg1305 ~^ {(+reg1364)}));
                  if (reg1327)
                    begin
                      reg1356 <= ($unsigned(((reg1328 ? reg1353 : reg1338) ?
                          $signed((8'ha0)) : (|(8'ha3)))) && (+(reg1315[(1'h1):(1'h1)] ?
                          (reg1307 ? reg1320 : reg1308) : (reg1308 ?
                              forvar1313 : (8'ha0)))));
                      reg1357 <= (($signed(((8'h9c) ? reg1305 : reg1308)) ?
                              reg1312 : {(reg1304 ? reg1358 : reg1319)}) ?
                          $unsigned((!(reg1359 ?
                              forvar1354 : (8'ha4)))) : reg1346[(1'h0):(1'h0)]);
                      reg1358 <= $signed($signed(((+forvar1317) | {reg1352})));
                      reg1359 <= ((|reg1358) >>> $unsigned(forvar1312[(1'h1):(1'h0)]));
                    end
                  else
                    begin
                      reg1356 <= reg1339;
                    end
                  if (reg1307[(1'h1):(1'h1)])
                    begin
                      reg1360 <= forvar1331;
                    end
                  else
                    begin
                      reg1360 <= (((|$signed(wire1300)) <= reg1353) <= $signed($unsigned($signed(forvar1303))));
                      reg1361 <= $unsigned($unsigned($signed(((8'hac) ?
                          forvar1311 : reg1315))));
                      reg1362 <= $signed(((reg1330[(2'h3):(1'h0)] ?
                              reg1362[(4'hc):(4'h9)] : wire1298) ?
                          reg1365 : $signed($unsigned((8'hb0)))));
                      reg1363 <= (+(reg1364 ? forvar1335 : forvar1304));
                    end
                end
              for (forvar1364 = (1'h0); (forvar1364 < (2'h3)); forvar1364 = (forvar1364 + (1'h1)))
                begin
                  reg1365 <= reg1312;
                  if (((^~reg1346[(1'h0):(1'h0)]) ?
                      $signed($unsigned($signed(reg1321))) : {$signed($unsigned(reg1350))}))
                    begin
                      reg1366 <= (|reg1365[(2'h2):(1'h0)]);
                      reg1367 <= $unsigned($signed(({forvar1353} + reg1315)));
                      reg1368 <= ({((!reg1365) > (reg1304 ?
                                  forvar1321 : forvar1334))} ?
                          (reg1333 <<< $signed((-reg1328))) : $unsigned(reg1334));
                      reg1369 <= forvar1303[(3'h4):(1'h0)];
                    end
                  else
                    begin
                      reg1366 <= reg1313;
                      reg1367 <= $signed($unsigned(((reg1338 ?
                              forvar1331 : wire1302) ?
                          ((8'had) ^ (8'hb2)) : $unsigned(reg1322))));
                      reg1368 <= $signed(((-reg1332) ?
                          reg1338 : reg1369[(3'h7):(3'h5)]));
                    end
                end
            end
          else
            begin
              if (reg1310[(1'h1):(1'h1)])
                begin
                  reg1349 <= ((&(forvar1361[(4'hc):(3'h7)] | (reg1360 & forvar1311))) & $signed($unsigned($unsigned(wire1300))));
                  reg1350 <= (($unsigned($signed(forvar1347)) ?
                      (wire1301 >>> (8'hb4)) : (8'hab)) << reg1317);
                  if ($signed((|$signed((!(8'h9e))))))
                    begin
                      reg1351 <= {(~|(~|(+(8'ha6))))};
                      reg1352 <= (forvar1345[(4'hf):(2'h2)] ?
                          reg1308 : {{(|reg1309)}});
                      reg1353 <= (&((8'ha5) & (reg1367[(2'h2):(1'h0)] <<< {reg1319})));
                      reg1354 <= forvar1332[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg1351 <= $signed($signed(reg1305[(2'h2):(1'h0)]));
                      reg1352 <= (reg1306 | (reg1359[(1'h1):(1'h1)] & $unsigned((forvar1325 ?
                          forvar1313 : forvar1318))));
                    end
                end
              else
                begin
                  for (forvar1349 = (1'h0); (forvar1349 < (2'h2)); forvar1349 = (forvar1349 + (1'h1)))
                    begin
                      reg1350 <= forvar1351;
                      reg1351 <= (^($unsigned($unsigned(forvar1321)) >> {$unsigned((8'h9e))}));
                    end
                  if ((~|$signed((8'hab))))
                    begin
                      reg1352 <= (!(forvar1334 ^~ (-forvar1333)));
                    end
                  else
                    begin
                      reg1352 <= forvar1354[(2'h3):(2'h3)];
                      reg1353 <= forvar1349;
                      reg1354 <= reg1313[(1'h1):(1'h0)];
                    end
                end
              reg1355 <= $signed(((forvar1335 ?
                      $signed(reg1315) : $signed(reg1311)) ?
                  forvar1308 : {(8'ha0)}));
            end
          for (forvar1370 = (1'h0); (forvar1370 < (1'h0)); forvar1370 = (forvar1370 + (1'h1)))
            begin
              for (forvar1371 = (1'h0); (forvar1371 < (1'h1)); forvar1371 = (forvar1371 + (1'h1)))
                begin
                  for (forvar1372 = (1'h0); (forvar1372 < (2'h3)); forvar1372 = (forvar1372 + (1'h1)))
                    begin
                      reg1373 <= $unsigned(reg1308);
                      reg1374 <= ((wire1299 ?
                          (wire1298 != wire1302[(1'h1):(1'h0)]) : ($signed(reg1336) ?
                              $unsigned((8'ha2)) : (reg1327 ?
                                  reg1320 : reg1355))) && $signed(($signed(reg1323) ?
                          reg1342[(4'ha):(2'h2)] : (8'hb2))));
                      reg1375 <= reg1355;
                      reg1376 <= (&((|forvar1321) ?
                          {(^reg1361)} : (((8'hb0) >= (8'ha4)) + {(8'hb0)})));
                    end
                  for (forvar1377 = (1'h0); (forvar1377 < (2'h2)); forvar1377 = (forvar1377 + (1'h1)))
                    begin
                      reg1378 <= (((reg1343 ?
                              (|forvar1312) : $signed((8'hb5))) ~^ ($unsigned(reg1348) - {(8'hb1)})) ?
                          reg1357 : $unsigned({{wire1298}}));
                      reg1379 <= {forvar1334};
                      reg1380 <= reg1308[(3'h5):(3'h4)];
                      reg1381 <= reg1341[(1'h1):(1'h0)];
                    end
                  for (forvar1382 = (1'h0); (forvar1382 < (1'h0)); forvar1382 = (forvar1382 + (1'h1)))
                    begin
                      reg1383 <= ($signed(((reg1313 ? reg1356 : reg1309) ?
                          reg1311[(4'h8):(1'h0)] : $unsigned(forvar1371))) <<< (+(-(wire1300 != (8'hb6)))));
                    end
                end
              for (forvar1384 = (1'h0); (forvar1384 < (2'h2)); forvar1384 = (forvar1384 + (1'h1)))
                begin
                  for (forvar1385 = (1'h0); (forvar1385 < (2'h3)); forvar1385 = (forvar1385 + (1'h1)))
                    begin
                      reg1386 <= reg1350[(1'h0):(1'h0)];
                    end
                  if ($unsigned(reg1348[(2'h2):(1'h0)]))
                    begin
                      reg1387 <= $unsigned(((reg1386 ?
                              reg1321 : (forvar1321 - reg1354)) ?
                          reg1375 : {(reg1367 ? reg1361 : (8'hac))}));
                      reg1388 <= (|(forvar1345 ?
                          (^~{(8'ha6)}) : {$unsigned(reg1322)}));
                      reg1389 <= (reg1364[(1'h1):(1'h0)] && $unsigned({(reg1321 ?
                              forvar1321 : reg1307)}));
                    end
                  else
                    begin
                      reg1387 <= $unsigned((reg1342 <<< (8'h9e)));
                      reg1388 <= reg1320[(2'h2):(1'h1)];
                      reg1389 <= {(+(~^forvar1331))};
                      reg1390 <= $signed(reg1336[(1'h0):(1'h0)]);
                    end
                end
              for (forvar1391 = (1'h0); (forvar1391 < (2'h2)); forvar1391 = (forvar1391 + (1'h1)))
                begin
                  if ({$signed(({reg1332} ?
                          (~|forvar1331) : (reg1338 && reg1358)))})
                    begin
                      reg1392 <= (^~$signed({(~reg1379)}));
                      reg1393 <= $signed(forvar1331);
                    end
                  else
                    begin
                      reg1392 <= reg1317[(1'h0):(1'h0)];
                      reg1393 <= ((~$signed($unsigned(reg1334))) ?
                          (~forvar1304[(3'h4):(2'h2)]) : $unsigned(reg1307[(1'h1):(1'h0)]));
                    end
                  if ($signed($signed($unsigned((reg1365 ^ forvar1318)))))
                    begin
                      reg1394 <= (reg1388[(3'h5):(3'h5)] << $signed(($unsigned((8'ha3)) <<< $unsigned(reg1360))));
                      reg1395 <= {forvar1337};
                    end
                  else
                    begin
                      reg1394 <= (forvar1377 ? reg1392 : {wire1302});
                      reg1395 <= $signed(($unsigned(((8'hb5) ~^ reg1333)) ?
                          ((forvar1377 ? forvar1337 : forvar1340) ?
                              ((8'h9c) ^~ reg1342) : (!forvar1340)) : {((8'ha9) ?
                                  reg1336 : reg1352)}));
                      reg1396 <= forvar1351[(4'he):(4'h9)];
                    end
                  for (forvar1397 = (1'h0); (forvar1397 < (2'h2)); forvar1397 = (forvar1397 + (1'h1)))
                    begin
                      reg1398 <= ($unsigned(reg1359) ?
                          {(reg1351 ^~ (reg1310 ?
                                  reg1380 : reg1328))} : $unsigned(reg1365));
                      reg1399 <= $unsigned(reg1318);
                      reg1400 <= ((((forvar1361 < reg1338) & (reg1359 ?
                          reg1348 : reg1308)) * forvar1391[(4'ha):(3'h6)]) << (($unsigned(reg1307) + (forvar1353 != reg1343)) >>> $unsigned((8'ha1))));
                    end
                  for (forvar1401 = (1'h0); (forvar1401 < (1'h0)); forvar1401 = (forvar1401 + (1'h1)))
                    begin
                      reg1402 <= ((~|((-(8'ha1)) & (reg1346 || forvar1382))) ~^ $unsigned(reg1313[(2'h2):(1'h1)]));
                    end
                end
              reg1403 <= {(^$signed(wire1298))};
            end
          for (forvar1404 = (1'h0); (forvar1404 < (1'h0)); forvar1404 = (forvar1404 + (1'h1)))
            begin
              for (forvar1405 = (1'h0); (forvar1405 < (1'h0)); forvar1405 = (forvar1405 + (1'h1)))
                begin
                  for (forvar1406 = (1'h0); (forvar1406 < (1'h0)); forvar1406 = (forvar1406 + (1'h1)))
                    begin
                      reg1407 <= (($unsigned({forvar1311}) ?
                          (8'ha1) : ($unsigned(reg1376) ?
                              $unsigned(forvar1340) : $unsigned(reg1358))) >= $unsigned((!(^~(8'h9c)))));
                      reg1408 <= $signed(reg1308[(2'h2):(1'h1)]);
                    end
                end
              reg1409 <= forvar1357[(3'h7):(3'h5)];
              for (forvar1410 = (1'h0); (forvar1410 < (1'h1)); forvar1410 = (forvar1410 + (1'h1)))
                begin
                  if (reg1309)
                    begin
                      reg1411 <= {$unsigned((^$unsigned(reg1349)))};
                    end
                  else
                    begin
                      reg1411 <= (($unsigned({reg1394}) + forvar1404) | reg1338[(1'h1):(1'h0)]);
                    end
                end
            end
          if (((reg1315[(2'h2):(1'h1)] ?
              (reg1307[(2'h2):(1'h0)] ?
                  $signed(reg1313) : (-forvar1353)) : forvar1345[(4'h8):(3'h5)]) * {(reg1394[(1'h0):(1'h0)] ?
                  (!reg1368) : {reg1358})}))
            begin
              if ($unsigned(reg1355))
                begin
                  if ($signed(({forvar1410} ? {$signed(reg1379)} : forvar1318)))
                    begin
                      reg1412 <= $unsigned((^~{forvar1333}));
                      reg1413 <= $signed(reg1352[(3'h7):(1'h1)]);
                    end
                  else
                    begin
                      reg1412 <= reg1362[(3'h4):(1'h1)];
                      reg1413 <= $unsigned($signed((~&reg1409)));
                    end
                  reg1414 <= (({reg1376[(2'h2):(2'h2)]} ?
                          forvar1317 : {(8'ha7)}) ?
                      $signed($signed((^~reg1316))) : (|{forvar1331}));
                  for (forvar1415 = (1'h0); (forvar1415 < (1'h1)); forvar1415 = (forvar1415 + (1'h1)))
                    begin
                      reg1416 <= (+$unsigned(($unsigned(forvar1347) > (-reg1360))));
                      reg1417 <= $signed({reg1330[(1'h0):(1'h0)]});
                    end
                end
              else
                begin
                  reg1412 <= reg1339;
                  reg1413 <= (forvar1332[(2'h2):(2'h2)] << reg1366[(1'h0):(1'h0)]);
                end
              reg1418 <= {({(~^reg1316)} || reg1350)};
              if (((~|((reg1417 ? reg1398 : forvar1406) ?
                      reg1320[(1'h1):(1'h0)] : forvar1404)) ?
                  reg1417 : (~reg1334[(3'h4):(3'h4)])))
                begin
                  reg1419 <= reg1408[(2'h3):(1'h1)];
                  reg1420 <= ((!({reg1388} >= $unsigned((8'had)))) + ($signed(reg1351) != $signed(((8'ha1) == reg1310))));
                  if (((((~(8'hba)) ~^ (reg1369 ? reg1400 : (8'ha1))) ?
                      ((reg1408 >= (8'ha0)) ?
                          reg1356[(2'h2):(1'h0)] : ((8'hab) ?
                              (8'had) : wire1302)) : ($signed(reg1414) > (~|reg1373))) << reg1419))
                    begin
                      reg1421 <= (~^{(^~$unsigned((8'ha5)))});
                      reg1422 <= (($unsigned($signed(reg1395)) ^ reg1386[(1'h0):(1'h0)]) ?
                          ({(-(8'h9e))} ?
                              $unsigned($unsigned((8'hb7))) : $signed((reg1418 ?
                                  forvar1371 : reg1322))) : $signed(reg1368[(4'hc):(4'h9)]));
                    end
                  else
                    begin
                      reg1421 <= reg1338;
                      reg1422 <= reg1312[(2'h2):(1'h1)];
                      reg1423 <= (reg1306[(3'h7):(3'h4)] || (&(reg1329[(1'h0):(1'h0)] && (8'ha7))));
                      reg1424 <= reg1308[(1'h0):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar1419 = (1'h0); (forvar1419 < (2'h2)); forvar1419 = (forvar1419 + (1'h1)))
                    begin
                      reg1420 <= $unsigned(forvar1335);
                      reg1421 <= reg1307[(2'h2):(1'h0)];
                    end
                  if ((reg1366[(3'h4):(1'h1)] ?
                      {$signed((-forvar1314))} : (((reg1374 && reg1422) << $unsigned(forvar1313)) && $unsigned($signed((8'ha9))))))
                    begin
                      reg1422 <= $signed((~^{((8'haa) << (8'ha5))}));
                      reg1423 <= (forvar1357[(3'h4):(2'h2)] ?
                          (^(^$signed((8'hac)))) : forvar1321);
                      reg1424 <= ((|((reg1319 ?
                              reg1387 : reg1313) > (^(8'hb1)))) ?
                          reg1396 : {((forvar1340 >> reg1319) ?
                                  reg1361 : $unsigned(forvar1314))});
                      reg1425 <= reg1393[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1422 <= wire1301[(2'h3):(1'h0)];
                      reg1423 <= reg1376;
                      reg1424 <= {{(((8'haa) ?
                                  forvar1333 : reg1316) >>> $signed(forvar1304))}};
                      reg1425 <= {reg1311};
                    end
                  if ($signed({$unsigned((reg1358 ? reg1368 : reg1358))}))
                    begin
                      reg1426 <= (~^forvar1331[(3'h5):(3'h4)]);
                    end
                  else
                    begin
                      reg1426 <= (|{($unsigned(reg1414) ?
                              (^reg1369) : (&forvar1325))});
                      reg1427 <= (8'ha1);
                      reg1428 <= forvar1318;
                      reg1429 <= $signed(((^~forvar1405[(2'h3):(1'h0)]) <= reg1309[(3'h5):(2'h2)]));
                    end
                end
            end
          else
            begin
              for (forvar1412 = (1'h0); (forvar1412 < (2'h3)); forvar1412 = (forvar1412 + (1'h1)))
                begin
                  for (forvar1413 = (1'h0); (forvar1413 < (1'h1)); forvar1413 = (forvar1413 + (1'h1)))
                    begin
                      reg1414 <= ({(~|((8'hb5) > reg1308))} < (~^$unsigned(reg1379)));
                    end
                  reg1415 <= $unsigned(($unsigned($signed(reg1379)) ?
                      reg1378[(2'h2):(1'h0)] : (8'hac)));
                end
            end
        end
      for (forvar1430 = (1'h0); (forvar1430 < (1'h1)); forvar1430 = (forvar1430 + (1'h1)))
        begin
          if (reg1400)
            begin
              if ($signed(reg1398))
                begin
                  reg1431 <= reg1337[(3'h4):(1'h0)];
                  for (forvar1432 = (1'h0); (forvar1432 < (1'h0)); forvar1432 = (forvar1432 + (1'h1)))
                    begin
                      reg1433 <= (~^{($unsigned(forvar1397) ?
                              $unsigned(reg1321) : forvar1334[(3'h5):(2'h2)])});
                    end
                  if (reg1392)
                    begin
                      reg1434 <= $unsigned(((wire1298 ?
                          (|reg1305) : forvar1412) <= ((forvar1312 ~^ forvar1337) || {forvar1412})));
                    end
                  else
                    begin
                      reg1434 <= ($unsigned($signed({forvar1405})) <= (|reg1321));
                      reg1435 <= reg1383[(3'h6):(2'h2)];
                      reg1436 <= $signed(((reg1350[(1'h0):(1'h0)] ?
                          reg1318 : (&reg1407)) <= {reg1327[(1'h0):(1'h0)]}));
                      reg1437 <= $unsigned(({(+reg1369)} ?
                          $unsigned({forvar1415}) : ({forvar1353} - $unsigned((8'h9d)))));
                    end
                  reg1438 <= $signed(reg1366);
                end
              else
                begin
                  if ((8'ha6))
                    begin
                      reg1431 <= $unsigned(wire1301);
                      reg1432 <= forvar1325[(3'h6):(1'h1)];
                      reg1433 <= ($signed({reg1394[(2'h3):(2'h3)]}) ?
                          $unsigned(reg1431[(1'h0):(1'h0)]) : $signed($unsigned($unsigned(reg1337))));
                      reg1434 <= (|reg1421);
                    end
                  else
                    begin
                      reg1431 <= {$signed((forvar1345 ^ $unsigned((8'h9e))))};
                      reg1432 <= reg1352[(2'h3):(2'h3)];
                    end
                end
              reg1439 <= (8'had);
              for (forvar1440 = (1'h0); (forvar1440 < (2'h2)); forvar1440 = (forvar1440 + (1'h1)))
                begin
                  reg1441 <= (((|(reg1332 ? reg1364 : wire1300)) ?
                      (8'haf) : (~&((8'ha9) || (8'hac)))) ^~ reg1316);
                end
              if ((+reg1376))
                begin
                  reg1442 <= {(~&{(forvar1314 ? reg1439 : reg1339)})};
                  if (forvar1382)
                    begin
                      reg1443 <= $unsigned({$signed((reg1339 - (8'haf)))});
                      reg1444 <= (forvar1405[(1'h0):(1'h0)] - (reg1428 ^ reg1358[(4'h8):(2'h3)]));
                      reg1445 <= reg1413[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1443 <= forvar1333;
                      reg1444 <= {(((reg1428 ? reg1409 : (8'h9f)) ?
                                  (reg1402 * reg1339) : (!reg1356)) ?
                              reg1431[(2'h3):(2'h2)] : reg1304[(2'h2):(2'h2)])};
                      reg1445 <= forvar1432;
                      reg1446 <= reg1434;
                    end
                end
              else
                begin
                  for (forvar1442 = (1'h0); (forvar1442 < (2'h2)); forvar1442 = (forvar1442 + (1'h1)))
                    begin
                      reg1443 <= (((((8'ha5) ?
                          reg1431 : reg1400) || reg1396[(2'h3):(1'h1)]) || (&(reg1438 ?
                          reg1434 : reg1381))) < $unsigned($signed($unsigned(reg1334))));
                      reg1444 <= $signed((+$signed(reg1317)));
                      reg1445 <= {reg1355};
                      reg1446 <= reg1436[(1'h0):(1'h0)];
                    end
                end
            end
          else
            begin
              for (forvar1431 = (1'h0); (forvar1431 < (1'h1)); forvar1431 = (forvar1431 + (1'h1)))
                begin
                  if ($unsigned(reg1351[(3'h6):(3'h6)]))
                    begin
                      reg1432 <= (|$signed($unsigned((&reg1321))));
                      reg1433 <= $unsigned($unsigned(reg1386));
                    end
                  else
                    begin
                      reg1432 <= reg1307[(1'h0):(1'h0)];
                      reg1433 <= (~&($unsigned($unsigned(reg1329)) ?
                          $unsigned((reg1375 ?
                              reg1415 : (8'ha4))) : reg1421[(4'h9):(3'h7)]));
                      reg1434 <= {{reg1357[(1'h1):(1'h0)]}};
                      reg1435 <= $signed((|forvar1321[(1'h1):(1'h1)]));
                    end
                  reg1436 <= {{reg1351}};
                end
              if ((~|reg1304))
                begin
                  for (forvar1437 = (1'h0); (forvar1437 < (2'h2)); forvar1437 = (forvar1437 + (1'h1)))
                    begin
                      reg1438 <= reg1351[(1'h1):(1'h1)];
                      reg1439 <= reg1425[(1'h0):(1'h0)];
                      reg1440 <= $unsigned($signed((~(forvar1440 <<< reg1425))));
                      reg1441 <= reg1310[(3'h5):(2'h2)];
                    end
                  for (forvar1442 = (1'h0); (forvar1442 < (2'h3)); forvar1442 = (forvar1442 + (1'h1)))
                    begin
                      reg1443 <= $unsigned($signed($unsigned((forvar1437 ^~ reg1336))));
                      reg1444 <= (8'ha4);
                    end
                end
              else
                begin
                  for (forvar1437 = (1'h0); (forvar1437 < (2'h2)); forvar1437 = (forvar1437 + (1'h1)))
                    begin
                      reg1438 <= ({$unsigned($signed(reg1329))} ?
                          ((forvar1442[(3'h4):(2'h3)] ?
                              forvar1312[(2'h3):(2'h3)] : reg1441[(3'h6):(3'h6)]) >>> wire1298[(1'h0):(1'h0)]) : ((~|{reg1381}) <= $signed(forvar1382)));
                      reg1439 <= (reg1342 ?
                          {(|forvar1332[(1'h1):(1'h0)])} : reg1321[(1'h1):(1'h0)]);
                    end
                  if (($unsigned((^(8'hae))) <= $unsigned({reg1425})))
                    begin
                      reg1440 <= (8'ha6);
                      reg1441 <= $unsigned($signed($unsigned(reg1383)));
                      reg1442 <= forvar1332[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1440 <= ({reg1437[(2'h2):(1'h0)]} ?
                          ((~^$signed(reg1380)) ?
                              forvar1308 : reg1383) : (((forvar1377 ?
                                  reg1326 : forvar1340) < {(8'hb3)}) ?
                              ($signed(reg1348) * {reg1407}) : $signed(reg1356[(1'h1):(1'h0)])));
                      reg1441 <= (($unsigned((forvar1311 ?
                              reg1320 : reg1441)) >> $signed(forvar1405)) ?
                          (~((-forvar1325) ?
                              (reg1424 ?
                                  (8'hac) : reg1378) : reg1353)) : ({forvar1331[(4'hc):(1'h1)]} ?
                              (&(~^(8'hb0))) : ($signed(reg1326) != reg1398[(4'hb):(3'h5)])));
                      reg1442 <= (!({(reg1334 ~^ reg1324)} ?
                          $signed((~^forvar1413)) : reg1319));
                      reg1443 <= reg1412[(4'he):(4'h8)];
                    end
                end
              reg1445 <= forvar1432;
              reg1446 <= (~&reg1338[(3'h5):(3'h4)]);
            end
          reg1447 <= forvar1314[(1'h1):(1'h0)];
          reg1448 <= ({$unsigned(forvar1317[(3'h7):(3'h7)])} >> (reg1412[(3'h5):(3'h4)] ?
              reg1324[(2'h3):(1'h0)] : reg1306[(2'h3):(2'h3)]));
        end
    end
  assign wire1449 = $unsigned($signed(reg1333[(3'h4):(1'h1)]));
  assign wire1450 = reg1346;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7  (y, clk, wire8, wire9, wire10, wire11, wire12);
  output wire [(32'h1875):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire8;
  input wire [(4'ha):(1'h0)] wire9;
  input wire signed [(4'hc):(1'h0)] wire10;
  input wire [(4'hb):(1'h0)] wire11;
  input wire signed [(4'hf):(1'h0)] wire12;
  wire signed [(2'h2):(1'h0)] wire1294;
  reg signed [(4'ha):(1'h0)] reg1293 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1292 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1291 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1290 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1289 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1288 = (1'h0);
  reg [(3'h4):(1'h0)] reg1287 = (1'h0);
  reg [(4'hc):(1'h0)] reg1286 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1285 = (1'h0);
  reg [(3'h5):(1'h0)] reg1284 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1283 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1282 = (1'h0);
  reg [(4'hd):(1'h0)] reg1279 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1278 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1275 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1274 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1282 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1281 = (1'h0);
  reg [(4'hb):(1'h0)] reg1280 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1279 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1278 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1277 = (1'h0);
  reg [(4'hf):(1'h0)] reg1276 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1275 = (1'h0);
  reg [(4'hf):(1'h0)] reg1274 = (1'h0);
  reg [(4'he):(1'h0)] reg1273 = (1'h0);
  reg [(2'h3):(1'h0)] reg1272 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1271 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1270 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1269 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1268 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1267 = (1'h0);
  reg [(4'hc):(1'h0)] reg1266 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1265 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1264 = (1'h0);
  reg [(4'he):(1'h0)] reg1262 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1261 = (1'h0);
  reg [(2'h2):(1'h0)] reg1264 = (1'h0);
  reg [(3'h4):(1'h0)] reg1263 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1262 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1261 = (1'h0);
  reg [(5'h10):(1'h0)] reg1258 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1260 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1259 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1258 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1257 = (1'h0);
  reg [(3'h6):(1'h0)] reg1256 = (1'h0);
  reg [(3'h7):(1'h0)] reg1253 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1251 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1248 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1245 = (1'h0);
  reg [(5'h10):(1'h0)] reg1255 = (1'h0);
  reg [(2'h3):(1'h0)] reg1254 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1253 = (1'h0);
  reg [(3'h4):(1'h0)] reg1252 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1251 = (1'h0);
  reg [(4'hf):(1'h0)] reg1250 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1249 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1248 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1247 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1246 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1245 = (1'h0);
  reg [(3'h5):(1'h0)] reg1244 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1243 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1242 = (1'h0);
  reg [(3'h4):(1'h0)] reg1241 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1240 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1201 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1236 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1235 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1231 = (1'h0);
  reg [(2'h3):(1'h0)] reg1239 = (1'h0);
  reg [(5'h10):(1'h0)] reg1238 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1237 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1236 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1235 = (1'h0);
  reg [(5'h10):(1'h0)] reg1234 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1233 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1232 = (1'h0);
  reg [(4'hd):(1'h0)] reg1231 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1230 = (1'h0);
  reg [(3'h5):(1'h0)] reg1229 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1228 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1226 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1223 = (1'h0);
  reg [(5'h10):(1'h0)] reg1227 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1226 = (1'h0);
  reg [(3'h4):(1'h0)] reg1225 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1224 = (1'h0);
  reg [(4'hb):(1'h0)] reg1223 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1222 = (1'h0);
  reg [(3'h7):(1'h0)] reg1221 = (1'h0);
  reg [(4'h8):(1'h0)] reg1220 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1219 = (1'h0);
  reg [(3'h5):(1'h0)] reg1218 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1217 = (1'h0);
  reg [(3'h4):(1'h0)] reg1216 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1215 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1214 = (1'h0);
  reg [(3'h4):(1'h0)] reg1213 = (1'h0);
  reg [(4'hc):(1'h0)] reg1212 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1211 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1210 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1209 = (1'h0);
  reg [(4'he):(1'h0)] forvar1208 = (1'h0);
  reg [(4'h9):(1'h0)] reg1200 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1199 = (1'h0);
  reg [(3'h7):(1'h0)] reg1207 = (1'h0);
  reg [(3'h4):(1'h0)] reg1206 = (1'h0);
  reg [(4'he):(1'h0)] reg1205 = (1'h0);
  reg [(4'he):(1'h0)] reg1204 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1203 = (1'h0);
  reg [(3'h6):(1'h0)] reg1202 = (1'h0);
  reg [(4'hb):(1'h0)] reg1201 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1200 = (1'h0);
  reg [(3'h7):(1'h0)] reg1199 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1198 = (1'h0);
  reg [(4'ha):(1'h0)] reg1197 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1196 = (1'h0);
  reg [(2'h2):(1'h0)] reg1195 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1194 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1193 = (1'h0);
  reg [(2'h3):(1'h0)] reg1192 = (1'h0);
  reg [(3'h4):(1'h0)] reg1191 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1190 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1189 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1188 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1187 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1186 = (1'h0);
  reg [(2'h2):(1'h0)] reg1185 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1184 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1183 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1182 = (1'h0);
  reg [(4'ha):(1'h0)] reg1181 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1180 = (1'h0);
  reg [(4'he):(1'h0)] forvar1179 = (1'h0);
  reg [(4'he):(1'h0)] reg1178 = (1'h0);
  reg [(2'h3):(1'h0)] reg1177 = (1'h0);
  reg [(5'h10):(1'h0)] reg1176 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1175 = (1'h0);
  reg [(4'h9):(1'h0)] reg1174 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1173 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1172 = (1'h0);
  reg [(4'h9):(1'h0)] reg1171 = (1'h0);
  reg [(4'h9):(1'h0)] reg1170 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1169 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1168 = (1'h0);
  reg [(4'ha):(1'h0)] reg1167 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1166 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1165 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1164 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1163 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1162 = (1'h0);
  reg [(4'hc):(1'h0)] reg1166 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1165 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1164 = (1'h0);
  reg [(2'h3):(1'h0)] reg1163 = (1'h0);
  reg [(3'h6):(1'h0)] reg1162 = (1'h0);
  reg [(4'hf):(1'h0)] reg1135 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1136 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1161 = (1'h0);
  reg [(3'h6):(1'h0)] reg1160 = (1'h0);
  reg [(4'hf):(1'h0)] reg1159 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1158 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1157 = (1'h0);
  reg [(4'hc):(1'h0)] reg1156 = (1'h0);
  reg [(4'h9):(1'h0)] reg1155 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1154 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1152 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1151 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1149 = (1'h0);
  reg [(4'hb):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1149 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1148 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1147 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1146 = (1'h0);
  reg [(3'h7):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1144 = (1'h0);
  reg [(5'h10):(1'h0)] reg1143 = (1'h0);
  reg [(4'hf):(1'h0)] reg1142 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1141 = (1'h0);
  reg [(3'h6):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1139 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1138 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1137 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1136 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1135 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1130 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1129 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1123 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1118 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1114 = (1'h0);
  reg [(5'h10):(1'h0)] reg1134 = (1'h0);
  reg [(3'h5):(1'h0)] reg1133 = (1'h0);
  reg [(2'h3):(1'h0)] reg1132 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1131 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1130 = (1'h0);
  reg [(3'h6):(1'h0)] reg1129 = (1'h0);
  reg [(3'h5):(1'h0)] reg1128 = (1'h0);
  reg [(2'h2):(1'h0)] reg1127 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1125 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1120 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1117 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1115 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1113 = (1'h0);
  reg [(4'hf):(1'h0)] reg1109 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1106 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1101 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1100 = (1'h0);
  reg [(3'h7):(1'h0)] reg1098 = (1'h0);
  reg [(4'h8):(1'h0)] reg1090 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1099 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1097 = (1'h0);
  reg [(4'hf):(1'h0)] reg1092 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1126 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1125 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1124 = (1'h0);
  reg [(4'h9):(1'h0)] reg1123 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1122 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1120 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1119 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1116 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1112 = (1'h0);
  reg [(4'hd):(1'h0)] reg1118 = (1'h0);
  reg [(3'h4):(1'h0)] reg1117 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1116 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1115 = (1'h0);
  reg [(4'hb):(1'h0)] reg1114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1113 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1112 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1111 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1110 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1109 = (1'h0);
  reg [(2'h2):(1'h0)] reg1108 = (1'h0);
  reg [(4'hf):(1'h0)] reg1107 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1106 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1105 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1104 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1103 = (1'h0);
  reg [(4'h8):(1'h0)] reg1102 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1101 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1100 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1099 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1098 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1097 = (1'h0);
  reg [(4'hb):(1'h0)] reg1096 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1095 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1094 = (1'h0);
  reg [(4'he):(1'h0)] reg1093 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1092 = (1'h0);
  reg [(3'h7):(1'h0)] reg1091 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1090 = (1'h0);
  reg [(4'hb):(1'h0)] reg1089 = (1'h0);
  reg [(4'hf):(1'h0)] reg1088 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1087 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1086 = (1'h0);
  reg [(4'ha):(1'h0)] reg1085 = (1'h0);
  reg [(4'hb):(1'h0)] reg1084 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1083 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1082 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1081 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1080 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1079 = (1'h0);
  reg [(4'ha):(1'h0)] reg1078 = (1'h0);
  reg [(4'hb):(1'h0)] reg1077 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1076 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1075 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1074 = (1'h0);
  reg [(4'he):(1'h0)] forvar1073 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1072 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1071 = (1'h0);
  reg [(5'h10):(1'h0)] reg1070 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1069 = (1'h0);
  reg [(4'hf):(1'h0)] reg1067 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1066 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1062 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1059 = (1'h0);
  reg [(4'he):(1'h0)] reg1058 = (1'h0);
  reg [(4'hd):(1'h0)] reg1057 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1052 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1051 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1050 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1068 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1067 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1066 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1065 = (1'h0);
  reg [(4'hc):(1'h0)] reg1064 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1063 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1062 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1061 = (1'h0);
  reg [(4'hd):(1'h0)] reg1060 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1059 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1058 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1057 = (1'h0);
  reg [(3'h7):(1'h0)] reg1056 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1054 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1049 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1048 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1045 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1055 = (1'h0);
  reg [(4'hf):(1'h0)] reg1054 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1053 = (1'h0);
  reg [(4'hc):(1'h0)] reg1052 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1051 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1050 = (1'h0);
  reg [(4'h8):(1'h0)] reg1049 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1048 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1047 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1046 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1045 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1044 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1043 = (1'h0);
  reg [(4'hf):(1'h0)] reg1042 = (1'h0);
  reg [(3'h5):(1'h0)] reg1041 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1040 = (1'h0);
  reg [(5'h10):(1'h0)] reg1039 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1038 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1037 = (1'h0);
  reg [(2'h2):(1'h0)] reg1036 = (1'h0);
  reg [(3'h5):(1'h0)] reg1035 = (1'h0);
  reg [(4'h9):(1'h0)] reg1034 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1033 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1032 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1031 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1030 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1020 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1028 = (1'h0);
  reg [(4'h8):(1'h0)] reg1027 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1026 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1025 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1024 = (1'h0);
  reg [(3'h4):(1'h0)] reg1023 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1022 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1021 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1020 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1019 = (1'h0);
  reg [(3'h4):(1'h0)] reg1013 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1011 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1008 = (1'h0);
  reg [(2'h2):(1'h0)] reg1007 = (1'h0);
  reg [(2'h2):(1'h0)] reg1004 = (1'h0);
  reg [(3'h5):(1'h0)] reg1000 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg999 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1018 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1017 = (1'h0);
  reg [(4'ha):(1'h0)] reg1016 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1015 = (1'h0);
  reg [(2'h3):(1'h0)] reg1014 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1013 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1012 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1011 = (1'h0);
  reg [(4'h8):(1'h0)] reg1010 = (1'h0);
  reg [(4'h9):(1'h0)] reg1009 = (1'h0);
  reg [(4'hb):(1'h0)] reg1008 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1007 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1006 = (1'h0);
  reg [(4'hf):(1'h0)] reg1005 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1004 = (1'h0);
  reg [(3'h7):(1'h0)] reg1003 = (1'h0);
  reg [(2'h3):(1'h0)] reg1002 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1001 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1000 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar999 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar998 = (1'h0);
  reg [(3'h5):(1'h0)] reg997 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg996 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar995 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar994 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar960 = (1'h0);
  reg [(4'h8):(1'h0)] reg963 = (1'h0);
  reg [(4'h9):(1'h0)] reg959 = (1'h0);
  reg signed [(4'he):(1'h0)] reg993 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar989 = (1'h0);
  reg [(3'h7):(1'h0)] reg984 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg992 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg991 = (1'h0);
  reg [(3'h5):(1'h0)] reg990 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg989 = (1'h0);
  reg [(4'h8):(1'h0)] reg988 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg987 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg986 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg985 = (1'h0);
  reg [(3'h5):(1'h0)] forvar984 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg982 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg983 = (1'h0);
  reg [(2'h3):(1'h0)] forvar982 = (1'h0);
  reg [(3'h5):(1'h0)] reg981 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg980 = (1'h0);
  reg [(3'h4):(1'h0)] reg979 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg978 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg977 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg976 = (1'h0);
  reg [(3'h5):(1'h0)] reg975 = (1'h0);
  reg [(5'h10):(1'h0)] reg974 = (1'h0);
  reg [(4'he):(1'h0)] reg973 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg972 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg971 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar970 = (1'h0);
  reg [(2'h3):(1'h0)] forvar969 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg968 = (1'h0);
  reg [(2'h2):(1'h0)] reg967 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg966 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg965 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg964 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar963 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg962 = (1'h0);
  reg [(5'h10):(1'h0)] reg961 = (1'h0);
  reg [(3'h6):(1'h0)] reg960 = (1'h0);
  reg [(4'h9):(1'h0)] forvar959 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg958 = (1'h0);
  reg [(4'h9):(1'h0)] forvar949 = (1'h0);
  reg [(5'h10):(1'h0)] reg957 = (1'h0);
  reg [(2'h3):(1'h0)] reg956 = (1'h0);
  reg [(4'he):(1'h0)] reg955 = (1'h0);
  reg [(4'h9):(1'h0)] forvar954 = (1'h0);
  reg [(3'h5):(1'h0)] reg953 = (1'h0);
  reg [(4'hd):(1'h0)] reg952 = (1'h0);
  reg [(4'hd):(1'h0)] reg951 = (1'h0);
  reg [(3'h6):(1'h0)] reg950 = (1'h0);
  reg [(2'h3):(1'h0)] reg949 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg948 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg947 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg946 = (1'h0);
  reg [(4'hf):(1'h0)] forvar945 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg945 = (1'h0);
  reg [(2'h2):(1'h0)] reg919 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg944 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg943 = (1'h0);
  reg [(3'h5):(1'h0)] reg942 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg941 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg940 = (1'h0);
  reg [(4'he):(1'h0)] reg939 = (1'h0);
  reg [(3'h6):(1'h0)] reg938 = (1'h0);
  reg [(2'h2):(1'h0)] forvar937 = (1'h0);
  reg [(3'h5):(1'h0)] reg936 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg935 = (1'h0);
  reg signed [(4'he):(1'h0)] reg934 = (1'h0);
  reg [(5'h10):(1'h0)] reg933 = (1'h0);
  reg [(2'h2):(1'h0)] forvar932 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg931 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar930 = (1'h0);
  reg [(5'h10):(1'h0)] forvar929 = (1'h0);
  reg [(3'h5):(1'h0)] reg928 = (1'h0);
  reg [(4'hd):(1'h0)] reg927 = (1'h0);
  reg [(3'h4):(1'h0)] reg926 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg925 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg924 = (1'h0);
  reg [(4'hb):(1'h0)] reg923 = (1'h0);
  reg [(4'hb):(1'h0)] forvar922 = (1'h0);
  reg [(4'ha):(1'h0)] reg921 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar920 = (1'h0);
  reg [(2'h2):(1'h0)] forvar919 = (1'h0);
  reg [(3'h5):(1'h0)] reg918 = (1'h0);
  reg signed [(4'he):(1'h0)] reg917 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg916 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar915 = (1'h0);
  reg [(4'hc):(1'h0)] reg914 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg913 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg912 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg911 = (1'h0);
  reg [(4'h9):(1'h0)] reg910 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg909 = (1'h0);
  reg [(4'hf):(1'h0)] reg908 = (1'h0);
  reg [(4'hf):(1'h0)] forvar907 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg906 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg903 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar899 = (1'h0);
  reg [(4'ha):(1'h0)] forvar896 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg905 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg904 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar903 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg902 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg901 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg900 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg899 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar898 = (1'h0);
  reg [(2'h2):(1'h0)] reg897 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg895 = (1'h0);
  reg [(4'hb):(1'h0)] reg898 = (1'h0);
  reg [(4'ha):(1'h0)] forvar897 = (1'h0);
  reg [(3'h7):(1'h0)] reg896 = (1'h0);
  reg [(5'h10):(1'h0)] forvar895 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg894 = (1'h0);
  reg [(5'h10):(1'h0)] reg893 = (1'h0);
  reg [(3'h5):(1'h0)] reg892 = (1'h0);
  reg [(2'h3):(1'h0)] reg891 = (1'h0);
  reg [(4'ha):(1'h0)] forvar890 = (1'h0);
  reg [(4'hc):(1'h0)] reg889 = (1'h0);
  reg [(4'h9):(1'h0)] forvar888 = (1'h0);
  reg [(3'h6):(1'h0)] reg887 = (1'h0);
  reg [(4'ha):(1'h0)] reg886 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar885 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar884 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg875 = (1'h0);
  reg [(4'hf):(1'h0)] forvar873 = (1'h0);
  reg [(4'hf):(1'h0)] reg883 = (1'h0);
  reg [(4'ha):(1'h0)] reg882 = (1'h0);
  reg [(4'hf):(1'h0)] reg881 = (1'h0);
  reg [(4'h8):(1'h0)] reg880 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar879 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg878 = (1'h0);
  reg [(4'h8):(1'h0)] reg877 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg876 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar875 = (1'h0);
  reg [(3'h5):(1'h0)] reg874 = (1'h0);
  reg [(4'hd):(1'h0)] reg873 = (1'h0);
  reg [(4'h9):(1'h0)] reg872 = (1'h0);
  reg [(2'h3):(1'h0)] reg871 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg870 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg869 = (1'h0);
  reg [(4'hf):(1'h0)] reg868 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar867 = (1'h0);
  reg [(4'h8):(1'h0)] reg866 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg865 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar864 = (1'h0);
  reg signed [(4'he):(1'h0)] reg863 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg864 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar863 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar862 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg853 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg861 = (1'h0);
  reg [(4'ha):(1'h0)] reg860 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg859 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar858 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg857 = (1'h0);
  reg [(4'h9):(1'h0)] reg856 = (1'h0);
  reg [(2'h3):(1'h0)] reg855 = (1'h0);
  reg [(3'h4):(1'h0)] reg854 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar853 = (1'h0);
  reg [(4'hb):(1'h0)] reg852 = (1'h0);
  reg [(2'h2):(1'h0)] reg851 = (1'h0);
  reg [(3'h4):(1'h0)] reg850 = (1'h0);
  reg [(4'he):(1'h0)] reg849 = (1'h0);
  reg [(3'h6):(1'h0)] forvar848 = (1'h0);
  reg [(3'h5):(1'h0)] reg847 = (1'h0);
  reg [(4'he):(1'h0)] forvar846 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar845 = (1'h0);
  reg [(3'h5):(1'h0)] forvar844 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg843 = (1'h0);
  reg [(4'he):(1'h0)] reg842 = (1'h0);
  reg [(4'hf):(1'h0)] forvar841 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar840 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg830 = (1'h0);
  reg [(3'h6):(1'h0)] forvar827 = (1'h0);
  reg [(4'hd):(1'h0)] reg839 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar838 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg837 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg836 = (1'h0);
  reg [(3'h7):(1'h0)] reg835 = (1'h0);
  reg [(4'ha):(1'h0)] reg834 = (1'h0);
  reg [(4'ha):(1'h0)] reg833 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg832 = (1'h0);
  reg signed [(4'he):(1'h0)] reg831 = (1'h0);
  reg [(2'h2):(1'h0)] forvar830 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg829 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg828 = (1'h0);
  reg [(4'hc):(1'h0)] reg827 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg826 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar825 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg824 = (1'h0);
  reg [(4'hb):(1'h0)] reg823 = (1'h0);
  reg [(4'he):(1'h0)] reg822 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg821 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg820 = (1'h0);
  reg [(2'h2):(1'h0)] reg819 = (1'h0);
  reg [(2'h2):(1'h0)] forvar818 = (1'h0);
  reg [(2'h2):(1'h0)] reg817 = (1'h0);
  reg [(2'h2):(1'h0)] reg816 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg815 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg814 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar813 = (1'h0);
  reg [(4'hf):(1'h0)] forvar812 = (1'h0);
  reg [(4'hf):(1'h0)] forvar811 = (1'h0);
  reg [(3'h7):(1'h0)] forvar810 = (1'h0);
  reg [(4'hf):(1'h0)] reg809 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg808 = (1'h0);
  reg [(3'h7):(1'h0)] reg807 = (1'h0);
  reg [(4'ha):(1'h0)] reg806 = (1'h0);
  reg [(4'h9):(1'h0)] reg805 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg804 = (1'h0);
  reg [(3'h7):(1'h0)] reg803 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar802 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg801 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar800 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar799 = (1'h0);
  reg [(3'h5):(1'h0)] reg798 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg797 = (1'h0);
  reg [(4'h9):(1'h0)] reg796 = (1'h0);
  reg [(4'he):(1'h0)] reg795 = (1'h0);
  reg [(4'hd):(1'h0)] forvar794 = (1'h0);
  reg [(3'h6):(1'h0)] forvar793 = (1'h0);
  reg [(5'h10):(1'h0)] forvar792 = (1'h0);
  reg [(4'he):(1'h0)] reg791 = (1'h0);
  reg [(2'h2):(1'h0)] forvar790 = (1'h0);
  reg [(2'h3):(1'h0)] reg789 = (1'h0);
  reg [(3'h6):(1'h0)] forvar788 = (1'h0);
  reg [(3'h7):(1'h0)] reg787 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg786 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg785 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg784 = (1'h0);
  reg [(4'h9):(1'h0)] reg783 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg782 = (1'h0);
  reg [(4'hc):(1'h0)] reg781 = (1'h0);
  reg [(3'h6):(1'h0)] forvar780 = (1'h0);
  reg signed [(4'he):(1'h0)] reg779 = (1'h0);
  reg [(4'h9):(1'h0)] reg778 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar777 = (1'h0);
  reg [(4'hb):(1'h0)] forvar776 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg775 = (1'h0);
  reg [(3'h4):(1'h0)] reg774 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg773 = (1'h0);
  reg [(4'hc):(1'h0)] reg772 = (1'h0);
  reg [(4'h8):(1'h0)] reg771 = (1'h0);
  reg [(3'h6):(1'h0)] reg770 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg769 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar768 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg767 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar763 = (1'h0);
  reg [(4'hc):(1'h0)] reg766 = (1'h0);
  reg [(3'h7):(1'h0)] reg765 = (1'h0);
  reg [(4'h9):(1'h0)] reg764 = (1'h0);
  reg [(4'ha):(1'h0)] reg763 = (1'h0);
  reg [(4'ha):(1'h0)] reg751 = (1'h0);
  reg [(2'h3):(1'h0)] reg762 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg761 = (1'h0);
  reg [(4'h9):(1'h0)] forvar760 = (1'h0);
  reg [(4'h9):(1'h0)] reg759 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg758 = (1'h0);
  reg signed [(4'he):(1'h0)] reg757 = (1'h0);
  reg [(4'hd):(1'h0)] reg756 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg755 = (1'h0);
  reg [(4'hd):(1'h0)] reg754 = (1'h0);
  reg [(4'h9):(1'h0)] reg753 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg752 = (1'h0);
  reg [(4'he):(1'h0)] forvar751 = (1'h0);
  reg signed [(4'he):(1'h0)] reg750 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg749 = (1'h0);
  reg [(4'h9):(1'h0)] reg748 = (1'h0);
  reg [(4'hf):(1'h0)] forvar747 = (1'h0);
  reg [(3'h6):(1'h0)] reg725 = (1'h0);
  reg [(2'h2):(1'h0)] forvar724 = (1'h0);
  reg [(2'h2):(1'h0)] forvar723 = (1'h0);
  reg [(2'h3):(1'h0)] forvar718 = (1'h0);
  reg [(4'hf):(1'h0)] reg713 = (1'h0);
  reg [(3'h4):(1'h0)] forvar711 = (1'h0);
  reg [(2'h2):(1'h0)] forvar704 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg746 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar745 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg744 = (1'h0);
  reg [(2'h3):(1'h0)] reg743 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg742 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg741 = (1'h0);
  reg [(3'h5):(1'h0)] forvar740 = (1'h0);
  reg [(4'hb):(1'h0)] reg739 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar738 = (1'h0);
  reg [(3'h4):(1'h0)] forvar737 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg736 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg734 = (1'h0);
  reg [(4'h9):(1'h0)] forvar733 = (1'h0);
  reg [(3'h7):(1'h0)] reg729 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar727 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg735 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar734 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg733 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg732 = (1'h0);
  reg [(4'hb):(1'h0)] reg731 = (1'h0);
  reg signed [(4'he):(1'h0)] reg730 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar729 = (1'h0);
  reg [(3'h4):(1'h0)] reg728 = (1'h0);
  reg [(3'h4):(1'h0)] reg727 = (1'h0);
  reg [(4'ha):(1'h0)] reg726 = (1'h0);
  reg [(4'ha):(1'h0)] forvar725 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg724 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg723 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg722 = (1'h0);
  reg [(4'h9):(1'h0)] reg721 = (1'h0);
  reg [(2'h3):(1'h0)] reg720 = (1'h0);
  reg [(3'h7):(1'h0)] reg719 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg718 = (1'h0);
  reg [(3'h6):(1'h0)] reg717 = (1'h0);
  reg [(3'h7):(1'h0)] reg716 = (1'h0);
  reg [(3'h7):(1'h0)] reg715 = (1'h0);
  reg [(3'h4):(1'h0)] reg714 = (1'h0);
  reg [(4'h8):(1'h0)] forvar713 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg712 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar708 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg711 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg710 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg703 = (1'h0);
  reg [(4'h8):(1'h0)] reg705 = (1'h0);
  reg [(3'h6):(1'h0)] reg709 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg708 = (1'h0);
  reg [(4'hb):(1'h0)] reg707 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg706 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar705 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg704 = (1'h0);
  reg [(3'h6):(1'h0)] forvar703 = (1'h0);
  wire [(5'h10):(1'h0)] wire13;
  wire signed [(4'h8):(1'h0)] wire14;
  wire signed [(4'hb):(1'h0)] wire701;
  assign y = {wire1294,
                 reg1293,
                 forvar1292,
                 reg1291,
                 reg1290,
                 forvar1289,
                 reg1288,
                 reg1287,
                 reg1286,
                 forvar1285,
                 reg1284,
                 reg1283,
                 forvar1282,
                 reg1279,
                 forvar1278,
                 reg1275,
                 forvar1274,
                 reg1282,
                 reg1281,
                 reg1280,
                 forvar1279,
                 reg1278,
                 reg1277,
                 reg1276,
                 forvar1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 forvar1271,
                 reg1270,
                 forvar1269,
                 reg1268,
                 reg1267,
                 reg1266,
                 reg1265,
                 forvar1264,
                 reg1262,
                 forvar1261,
                 reg1264,
                 reg1263,
                 forvar1262,
                 reg1261,
                 reg1258,
                 reg1260,
                 reg1259,
                 forvar1258,
                 reg1257,
                 reg1256,
                 reg1253,
                 forvar1251,
                 reg1248,
                 forvar1245,
                 reg1255,
                 reg1254,
                 forvar1253,
                 reg1252,
                 reg1251,
                 reg1250,
                 reg1249,
                 forvar1248,
                 reg1247,
                 reg1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 forvar1242,
                 reg1241,
                 forvar1240,
                 forvar1201,
                 reg1236,
                 forvar1235,
                 forvar1231,
                 reg1239,
                 reg1238,
                 reg1237,
                 forvar1236,
                 reg1235,
                 reg1234,
                 reg1233,
                 reg1232,
                 reg1231,
                 reg1230,
                 reg1229,
                 reg1228,
                 forvar1226,
                 forvar1223,
                 reg1227,
                 reg1226,
                 reg1225,
                 reg1224,
                 reg1223,
                 reg1222,
                 reg1221,
                 reg1220,
                 forvar1219,
                 reg1218,
                 reg1217,
                 reg1216,
                 reg1215,
                 forvar1214,
                 reg1213,
                 reg1212,
                 reg1211,
                 reg1210,
                 reg1209,
                 forvar1208,
                 reg1200,
                 forvar1199,
                 reg1207,
                 reg1206,
                 reg1205,
                 reg1204,
                 reg1203,
                 reg1202,
                 reg1201,
                 forvar1200,
                 reg1199,
                 reg1198,
                 reg1197,
                 forvar1196,
                 reg1195,
                 forvar1194,
                 reg1193,
                 reg1192,
                 reg1191,
                 reg1190,
                 forvar1189,
                 forvar1188,
                 forvar1187,
                 reg1186,
                 reg1185,
                 forvar1184,
                 reg1183,
                 reg1182,
                 reg1181,
                 reg1180,
                 forvar1179,
                 reg1178,
                 reg1177,
                 reg1176,
                 forvar1175,
                 reg1174,
                 reg1173,
                 forvar1172,
                 reg1171,
                 reg1170,
                 forvar1169,
                 forvar1168,
                 reg1167,
                 forvar1166,
                 reg1165,
                 reg1164,
                 forvar1163,
                 forvar1162,
                 reg1166,
                 forvar1165,
                 forvar1164,
                 reg1163,
                 reg1162,
                 reg1135,
                 reg1136,
                 reg1161,
                 reg1160,
                 reg1159,
                 forvar1158,
                 reg1157,
                 reg1156,
                 reg1155,
                 reg1154,
                 forvar1153,
                 reg1152,
                 reg1151,
                 reg1149,
                 reg1150,
                 forvar1149,
                 reg1148,
                 forvar1147,
                 reg1146,
                 reg1145,
                 reg1144,
                 reg1143,
                 reg1142,
                 reg1141,
                 reg1140,
                 reg1139,
                 reg1138,
                 reg1137,
                 forvar1136,
                 forvar1135,
                 forvar1130,
                 forvar1129,
                 forvar1123,
                 forvar1118,
                 forvar1114,
                 reg1134,
                 reg1133,
                 reg1132,
                 reg1131,
                 reg1130,
                 reg1129,
                 reg1128,
                 reg1127,
                 forvar1125,
                 forvar1120,
                 forvar1117,
                 forvar1115,
                 forvar1113,
                 reg1109,
                 reg1106,
                 reg1101,
                 forvar1100,
                 reg1098,
                 reg1090,
                 reg1099,
                 reg1097,
                 reg1092,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1123,
                 reg1122,
                 reg1121,
                 reg1120,
                 reg1119,
                 forvar1116,
                 reg1112,
                 reg1118,
                 reg1117,
                 reg1116,
                 reg1115,
                 reg1114,
                 reg1113,
                 forvar1112,
                 reg1111,
                 forvar1110,
                 forvar1109,
                 reg1108,
                 reg1107,
                 forvar1106,
                 reg1105,
                 reg1104,
                 reg1103,
                 reg1102,
                 forvar1101,
                 reg1100,
                 forvar1099,
                 forvar1098,
                 forvar1097,
                 reg1096,
                 reg1095,
                 reg1094,
                 reg1093,
                 forvar1092,
                 reg1091,
                 forvar1090,
                 reg1089,
                 reg1088,
                 reg1087,
                 forvar1086,
                 reg1085,
                 reg1084,
                 reg1083,
                 reg1082,
                 forvar1081,
                 forvar1080,
                 reg1079,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1075,
                 forvar1074,
                 forvar1073,
                 forvar1072,
                 reg1071,
                 reg1070,
                 forvar1069,
                 reg1067,
                 forvar1066,
                 forvar1062,
                 forvar1059,
                 reg1058,
                 reg1057,
                 forvar1052,
                 reg1051,
                 forvar1050,
                 reg1068,
                 forvar1067,
                 reg1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 forvar1058,
                 forvar1057,
                 reg1056,
                 forvar1054,
                 forvar1049,
                 reg1048,
                 forvar1045,
                 reg1055,
                 reg1054,
                 reg1053,
                 reg1052,
                 forvar1051,
                 reg1050,
                 reg1049,
                 forvar1048,
                 reg1047,
                 reg1046,
                 reg1045,
                 reg1044,
                 forvar1043,
                 reg1042,
                 reg1041,
                 reg1040,
                 reg1039,
                 forvar1038,
                 forvar1037,
                 reg1036,
                 reg1035,
                 reg1034,
                 reg1033,
                 forvar1032,
                 forvar1031,
                 forvar1030,
                 reg1020,
                 reg1029,
                 reg1028,
                 reg1027,
                 reg1026,
                 reg1025,
                 forvar1024,
                 reg1023,
                 reg1022,
                 reg1021,
                 forvar1020,
                 forvar1019,
                 reg1013,
                 forvar1011,
                 forvar1008,
                 reg1007,
                 reg1004,
                 reg1000,
                 reg999,
                 reg1018,
                 reg1017,
                 reg1016,
                 reg1015,
                 reg1014,
                 forvar1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1009,
                 reg1008,
                 forvar1007,
                 reg1006,
                 reg1005,
                 forvar1004,
                 reg1003,
                 reg1002,
                 reg1001,
                 forvar1000,
                 forvar999,
                 forvar998,
                 reg997,
                 reg996,
                 forvar995,
                 forvar994,
                 forvar960,
                 reg963,
                 reg959,
                 reg993,
                 forvar989,
                 reg984,
                 reg992,
                 reg991,
                 reg990,
                 reg989,
                 reg988,
                 reg987,
                 reg986,
                 reg985,
                 forvar984,
                 reg982,
                 reg983,
                 forvar982,
                 reg981,
                 reg980,
                 reg979,
                 reg978,
                 reg977,
                 reg976,
                 reg975,
                 reg974,
                 reg973,
                 reg972,
                 reg971,
                 forvar970,
                 forvar969,
                 reg968,
                 reg967,
                 reg966,
                 reg965,
                 reg964,
                 forvar963,
                 reg962,
                 reg961,
                 reg960,
                 forvar959,
                 reg958,
                 forvar949,
                 reg957,
                 reg956,
                 reg955,
                 forvar954,
                 reg953,
                 reg952,
                 reg951,
                 reg950,
                 reg949,
                 reg948,
                 reg947,
                 reg946,
                 forvar945,
                 reg945,
                 reg919,
                 reg944,
                 reg943,
                 reg942,
                 reg941,
                 reg940,
                 reg939,
                 reg938,
                 forvar937,
                 reg936,
                 reg935,
                 reg934,
                 reg933,
                 forvar932,
                 reg931,
                 forvar930,
                 forvar929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg923,
                 forvar922,
                 reg921,
                 forvar920,
                 forvar919,
                 reg918,
                 reg917,
                 reg916,
                 forvar915,
                 reg914,
                 reg913,
                 reg912,
                 reg911,
                 reg910,
                 reg909,
                 reg908,
                 forvar907,
                 reg906,
                 reg903,
                 forvar899,
                 forvar896,
                 reg905,
                 reg904,
                 forvar903,
                 reg902,
                 reg901,
                 reg900,
                 reg899,
                 forvar898,
                 reg897,
                 reg895,
                 reg898,
                 forvar897,
                 reg896,
                 forvar895,
                 reg894,
                 reg893,
                 reg892,
                 reg891,
                 forvar890,
                 reg889,
                 forvar888,
                 reg887,
                 reg886,
                 forvar885,
                 forvar884,
                 reg875,
                 forvar873,
                 reg883,
                 reg882,
                 reg881,
                 reg880,
                 forvar879,
                 reg878,
                 reg877,
                 reg876,
                 forvar875,
                 reg874,
                 reg873,
                 reg872,
                 reg871,
                 reg870,
                 reg869,
                 reg868,
                 forvar867,
                 reg866,
                 reg865,
                 forvar864,
                 reg863,
                 reg864,
                 forvar863,
                 forvar862,
                 reg853,
                 reg861,
                 reg860,
                 reg859,
                 forvar858,
                 reg857,
                 reg856,
                 reg855,
                 reg854,
                 forvar853,
                 reg852,
                 reg851,
                 reg850,
                 reg849,
                 forvar848,
                 reg847,
                 forvar846,
                 forvar845,
                 forvar844,
                 reg843,
                 reg842,
                 forvar841,
                 forvar840,
                 reg830,
                 forvar827,
                 reg839,
                 forvar838,
                 reg837,
                 reg836,
                 reg835,
                 reg834,
                 reg833,
                 reg832,
                 reg831,
                 forvar830,
                 reg829,
                 reg828,
                 reg827,
                 reg826,
                 forvar825,
                 reg824,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 forvar818,
                 reg817,
                 reg816,
                 reg815,
                 reg814,
                 forvar813,
                 forvar812,
                 forvar811,
                 forvar810,
                 reg809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 forvar802,
                 reg801,
                 forvar800,
                 forvar799,
                 reg798,
                 reg797,
                 reg796,
                 reg795,
                 forvar794,
                 forvar793,
                 forvar792,
                 reg791,
                 forvar790,
                 reg789,
                 forvar788,
                 reg787,
                 reg786,
                 reg785,
                 reg784,
                 reg783,
                 reg782,
                 reg781,
                 forvar780,
                 reg779,
                 reg778,
                 forvar777,
                 forvar776,
                 reg775,
                 reg774,
                 reg773,
                 reg772,
                 reg771,
                 reg770,
                 reg769,
                 forvar768,
                 reg767,
                 forvar763,
                 reg766,
                 reg765,
                 reg764,
                 reg763,
                 reg751,
                 reg762,
                 reg761,
                 forvar760,
                 reg759,
                 reg758,
                 reg757,
                 reg756,
                 reg755,
                 reg754,
                 reg753,
                 reg752,
                 forvar751,
                 reg750,
                 reg749,
                 reg748,
                 forvar747,
                 reg725,
                 forvar724,
                 forvar723,
                 forvar718,
                 reg713,
                 forvar711,
                 forvar704,
                 reg746,
                 forvar745,
                 reg744,
                 reg743,
                 reg742,
                 reg741,
                 forvar740,
                 reg739,
                 forvar738,
                 forvar737,
                 reg736,
                 reg734,
                 forvar733,
                 reg729,
                 forvar727,
                 reg735,
                 forvar734,
                 reg733,
                 reg732,
                 reg731,
                 reg730,
                 forvar729,
                 reg728,
                 reg727,
                 reg726,
                 forvar725,
                 reg724,
                 reg723,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 reg714,
                 forvar713,
                 reg712,
                 forvar708,
                 reg711,
                 reg710,
                 reg703,
                 reg705,
                 reg709,
                 reg708,
                 reg707,
                 reg706,
                 forvar705,
                 reg704,
                 forvar703,
                 wire13,
                 wire14,
                 wire701,
                 (1'h0)};
  assign wire13 = ({wire9} ^~ (&(((8'hb0) < wire8) <= wire10[(3'h7):(1'h1)])));
  assign wire14 = ($signed($signed($unsigned((8'ha2)))) < ((~|(8'h9f)) ^~ $unsigned((wire11 ?
                      wire12 : wire8))));
  module15 modinst702 (.clk(clk), .wire20(wire11), .y(wire701), .wire17(wire14), .wire19(wire13), .wire16(wire12), .wire18(wire8));
  always
    @(posedge clk) begin
      if ((~(~|({(8'ha8)} + wire12))))
        begin
          if (wire13[(3'h4):(3'h4)])
            begin
              for (forvar703 = (1'h0); (forvar703 < (2'h2)); forvar703 = (forvar703 + (1'h1)))
                begin
                  reg704 <= (($unsigned(wire10[(1'h1):(1'h0)]) ?
                      (8'hba) : wire701[(1'h1):(1'h1)]) - (^wire701));
                end
              for (forvar705 = (1'h0); (forvar705 < (1'h1)); forvar705 = (forvar705 + (1'h1)))
                begin
                  reg706 <= wire701[(3'h6):(2'h2)];
                  reg707 <= (~(reg704 ? wire701 : ((~^wire9) < wire701)));
                  if (((((wire9 ?
                      wire9 : wire11) > wire8) ^ (~$signed(wire12))) >>> $unsigned((~|$unsigned(wire12)))))
                    begin
                      reg708 <= (8'hb8);
                      reg709 <= reg708[(4'he):(4'h8)];
                    end
                  else
                    begin
                      reg708 <= wire12[(3'h5):(3'h5)];
                      reg709 <= $signed(($signed($signed(forvar705)) - ($unsigned(wire12) ?
                          $unsigned(wire8) : (reg704 ? reg704 : wire8))));
                    end
                end
            end
          else
            begin
              if ($signed($unsigned(wire14)))
                begin
                  for (forvar703 = (1'h0); (forvar703 < (1'h1)); forvar703 = (forvar703 + (1'h1)))
                    begin
                      reg704 <= $signed((^~$signed((wire9 + wire9))));
                      reg705 <= ((($signed(reg704) ?
                          reg708 : wire10[(4'hc):(1'h1)]) >> ((|forvar705) || (wire701 ?
                          reg706 : forvar705))) >> forvar703[(3'h5):(3'h4)]);
                    end
                end
              else
                begin
                  if (wire12)
                    begin
                      reg703 <= $signed({((~reg706) ?
                              (wire701 ? wire14 : reg707) : (^~forvar705))});
                    end
                  else
                    begin
                      reg703 <= wire12;
                      reg704 <= (reg706 ?
                          $unsigned((&((8'hb7) ?
                              wire13 : reg703))) : (~|reg705[(3'h5):(3'h4)]));
                      reg705 <= (~&forvar705);
                      reg706 <= (($unsigned((^(8'h9e))) >= (~$unsigned(wire11))) >>> reg706);
                    end
                  if ($unsigned((($unsigned(wire701) || (reg707 < reg708)) > ({forvar705} ?
                      reg703 : wire12[(3'h5):(1'h1)]))))
                    begin
                      reg707 <= (reg708[(3'h5):(1'h0)] ?
                          (wire12[(1'h0):(1'h0)] ?
                              (8'h9d) : (&reg704[(1'h0):(1'h0)])) : $unsigned((~&$unsigned(wire9))));
                      reg708 <= wire9;
                    end
                  else
                    begin
                      reg707 <= forvar703[(3'h4):(2'h2)];
                      reg708 <= (&(8'ha0));
                      reg709 <= $unsigned((-(^~reg705[(2'h2):(2'h2)])));
                      reg710 <= ($signed($signed(forvar705)) == $signed(($signed(wire11) << reg705[(2'h3):(2'h3)])));
                    end
                end
              reg711 <= ((^~(reg708[(1'h1):(1'h0)] ?
                  $signed(reg703) : reg704[(3'h4):(3'h4)])) << $signed(reg710[(4'h9):(4'h8)]));
            end
        end
      else
        begin
          if (reg711)
            begin
              for (forvar703 = (1'h0); (forvar703 < (1'h1)); forvar703 = (forvar703 + (1'h1)))
                begin
                  if ($unsigned((($signed(reg704) ?
                          (~reg711) : reg705[(1'h0):(1'h0)]) ?
                      reg703 : $signed(reg705[(4'h8):(2'h2)]))))
                    begin
                      reg704 <= $unsigned((wire13 ^~ ((reg704 ?
                          (8'ha7) : reg710) + (reg711 << reg707))));
                      reg705 <= $signed(reg708[(4'h8):(3'h6)]);
                      reg706 <= (|($unsigned((-wire701)) < {reg709}));
                      reg707 <= ((reg710 - $unsigned((^~wire14))) == (reg711 ?
                          $signed({wire10}) : ($unsigned(reg704) ?
                              (reg709 ? (8'h9c) : reg709) : (~(8'ha1)))));
                    end
                  else
                    begin
                      reg704 <= forvar705;
                      reg705 <= (wire10 & (-((wire14 ? wire14 : wire9) ?
                          $unsigned((8'hba)) : (wire12 ? reg704 : (8'ha9)))));
                    end
                end
              for (forvar708 = (1'h0); (forvar708 < (2'h3)); forvar708 = (forvar708 + (1'h1)))
                begin
                  if (wire9)
                    begin
                      reg709 <= ((8'hb0) ?
                          (~^$unsigned((-reg705))) : (wire11 >>> $unsigned($unsigned(reg708))));
                      reg710 <= (reg706[(2'h2):(2'h2)] ~^ ($signed((8'ha8)) ?
                          $unsigned(((8'hb0) ?
                              reg711 : reg703)) : $unsigned(wire12[(4'hb):(3'h5)])));
                      reg711 <= ($signed((~(reg708 ?
                          forvar705 : reg711))) && reg703[(2'h2):(2'h2)]);
                      reg712 <= (-reg706[(1'h0):(1'h0)]);
                    end
                  else
                    begin
                      reg709 <= (|((^~$unsigned(wire11)) ^~ ((+reg706) ?
                          (&reg706) : (wire10 ? wire11 : wire9))));
                    end
                  for (forvar713 = (1'h0); (forvar713 < (2'h3)); forvar713 = (forvar713 + (1'h1)))
                    begin
                      reg714 <= $signed(reg704);
                      reg715 <= (-$signed($signed($unsigned(wire14))));
                      reg716 <= ({{((8'h9d) <<< wire13)}} > {reg708[(4'hc):(2'h3)]});
                      reg717 <= reg706[(3'h4):(1'h1)];
                    end
                  if ($signed(((-(+reg709)) ?
                      {reg715} : $signed((reg711 ? (8'hb8) : wire9)))))
                    begin
                      reg718 <= (&wire10[(4'h9):(2'h3)]);
                      reg719 <= (~|$signed(wire13[(4'hd):(4'hc)]));
                      reg720 <= reg717;
                    end
                  else
                    begin
                      reg718 <= (~|$signed(forvar705[(2'h3):(1'h0)]));
                      reg719 <= ({reg714} && $signed($signed({reg714})));
                    end
                  if (wire701[(1'h0):(1'h0)])
                    begin
                      reg721 <= $unsigned($signed((8'ha7)));
                      reg722 <= $unsigned(reg717[(2'h2):(1'h1)]);
                      reg723 <= reg718;
                      reg724 <= reg721;
                    end
                  else
                    begin
                      reg721 <= $signed({$signed(((8'ha3) ? reg723 : reg708))});
                      reg722 <= ({($unsigned(reg721) ?
                              reg722 : $signed(reg721))} >>> reg703[(2'h2):(1'h0)]);
                    end
                end
              if (($signed(($signed(reg720) < {(8'ha5)})) ?
                  ((reg709[(3'h4):(3'h4)] >= $signed(reg716)) ?
                      (reg723 >> (reg719 ?
                          wire12 : reg707)) : wire12[(4'hb):(3'h5)]) : (((-wire13) || (reg723 ?
                      (8'hb9) : forvar708)) * {(-reg712)})))
                begin
                  for (forvar725 = (1'h0); (forvar725 < (2'h3)); forvar725 = (forvar725 + (1'h1)))
                    begin
                      reg726 <= {$unsigned(((wire8 ?
                              reg716 : (8'ha0)) & wire8))};
                      reg727 <= (^~(((reg722 > (8'had)) & (~&reg716)) ?
                          (8'hb0) : (~{reg724})));
                      reg728 <= $unsigned($signed($unsigned((reg706 ?
                          wire701 : reg726))));
                    end
                  for (forvar729 = (1'h0); (forvar729 < (1'h1)); forvar729 = (forvar729 + (1'h1)))
                    begin
                      reg730 <= $signed((reg721[(2'h3):(2'h3)] ?
                          (~^$signed(reg716)) : ({reg718} ?
                              reg712[(1'h0):(1'h0)] : reg703[(2'h3):(1'h1)])));
                      reg731 <= $unsigned($signed(wire9));
                      reg732 <= ($signed(reg719[(2'h3):(1'h1)]) ?
                          $signed(($signed(wire13) ?
                              (wire11 ?
                                  wire13 : forvar703) : $unsigned(forvar705))) : forvar725);
                      reg733 <= $signed((~^({reg706} ^~ {forvar703})));
                    end
                  for (forvar734 = (1'h0); (forvar734 < (2'h3)); forvar734 = (forvar734 + (1'h1)))
                    begin
                      reg735 <= $signed(reg711);
                    end
                end
              else
                begin
                  for (forvar725 = (1'h0); (forvar725 < (2'h3)); forvar725 = (forvar725 + (1'h1)))
                    begin
                      reg726 <= (~$unsigned($unsigned({(8'hb1)})));
                    end
                  for (forvar727 = (1'h0); (forvar727 < (2'h3)); forvar727 = (forvar727 + (1'h1)))
                    begin
                      reg728 <= $signed($signed(forvar725[(4'ha):(2'h2)]));
                    end
                  if ($signed($unsigned(forvar705[(1'h1):(1'h0)])))
                    begin
                      reg729 <= reg708;
                      reg730 <= (8'ha8);
                      reg731 <= reg705;
                      reg732 <= (forvar734 ?
                          ($unsigned((wire9 ?
                              (8'hb4) : (8'had))) + (~&(wire12 > reg726))) : ($signed(reg735) ?
                              $signed($unsigned(reg716)) : $signed((-reg721))));
                    end
                  else
                    begin
                      reg729 <= reg711[(4'h8):(3'h6)];
                    end
                  for (forvar733 = (1'h0); (forvar733 < (2'h3)); forvar733 = (forvar733 + (1'h1)))
                    begin
                      reg734 <= {reg722[(2'h2):(1'h0)]};
                      reg735 <= (|forvar703);
                      reg736 <= (reg714 ? reg719 : forvar705);
                    end
                end
              for (forvar737 = (1'h0); (forvar737 < (2'h3)); forvar737 = (forvar737 + (1'h1)))
                begin
                  for (forvar738 = (1'h0); (forvar738 < (1'h0)); forvar738 = (forvar738 + (1'h1)))
                    begin
                      reg739 <= (~$unsigned($signed($signed(reg716))));
                    end
                  for (forvar740 = (1'h0); (forvar740 < (2'h2)); forvar740 = (forvar740 + (1'h1)))
                    begin
                      reg741 <= $signed($signed($signed((!(8'ha4)))));
                      reg742 <= reg714;
                      reg743 <= (~((forvar727 ?
                              (forvar729 * forvar734) : wire701[(3'h5):(3'h4)]) ?
                          (~|forvar705[(3'h4):(1'h0)]) : $signed((|reg723))));
                      reg744 <= {(reg730[(1'h0):(1'h0)] <<< $unsigned(((8'hb4) <= forvar737)))};
                    end
                  for (forvar745 = (1'h0); (forvar745 < (2'h2)); forvar745 = (forvar745 + (1'h1)))
                    begin
                      reg746 <= ((+$unsigned(((8'hba) & reg708))) ?
                          reg703[(1'h1):(1'h1)] : ({{reg733}} * {$signed(forvar703)}));
                    end
                end
            end
          else
            begin
              for (forvar703 = (1'h0); (forvar703 < (1'h0)); forvar703 = (forvar703 + (1'h1)))
                begin
                  for (forvar704 = (1'h0); (forvar704 < (2'h3)); forvar704 = (forvar704 + (1'h1)))
                    begin
                      reg705 <= $signed((reg707 ?
                          reg721 : $unsigned(reg723[(4'h8):(1'h0)])));
                      reg706 <= $unsigned($signed({reg718[(3'h4):(1'h1)]}));
                      reg707 <= {(reg735[(2'h3):(1'h0)] ?
                              reg732 : reg730[(1'h0):(1'h0)])};
                    end
                  if ($signed(reg735))
                    begin
                      reg708 <= $unsigned($signed($unsigned((reg726 ?
                          wire14 : (8'hb7)))));
                    end
                  else
                    begin
                      reg708 <= {($unsigned((reg708 ?
                              wire10 : forvar725)) ^~ $signed((~|reg717)))};
                      reg709 <= reg709;
                      reg710 <= reg734;
                    end
                end
              if ({reg722[(1'h0):(1'h0)]})
                begin
                  for (forvar711 = (1'h0); (forvar711 < (1'h1)); forvar711 = (forvar711 + (1'h1)))
                    begin
                      reg712 <= ({((~^reg724) ?
                                  forvar705[(1'h0):(1'h0)] : reg734)} ?
                          wire12 : (~&({(8'ha7)} > (^~wire13))));
                      reg713 <= $signed((forvar737[(2'h2):(1'h0)] - ((reg722 ?
                          reg739 : reg717) + $unsigned(forvar745))));
                    end
                end
              else
                begin
                  for (forvar711 = (1'h0); (forvar711 < (1'h1)); forvar711 = (forvar711 + (1'h1)))
                    begin
                      reg712 <= {$unsigned((!reg718))};
                      reg713 <= $unsigned(reg729[(3'h7):(3'h4)]);
                    end
                  if (((8'ha9) ?
                      $signed(((^reg727) ?
                          {reg724} : {reg744})) : forvar705[(3'h5):(2'h3)]))
                    begin
                      reg714 <= forvar713[(1'h1):(1'h0)];
                      reg715 <= $signed(($signed($signed(reg727)) ?
                          reg724[(2'h3):(2'h3)] : $signed((!reg732))));
                      reg716 <= $signed(forvar711[(1'h1):(1'h0)]);
                      reg717 <= {$unsigned($unsigned((!forvar738)))};
                    end
                  else
                    begin
                      reg714 <= (&$signed({(reg714 + reg746)}));
                      reg715 <= $signed(($unsigned(((8'h9d) ?
                              reg746 : reg705)) ?
                          ($signed(forvar704) || (reg703 << reg733)) : $unsigned((wire12 ^~ reg735))));
                    end
                  for (forvar718 = (1'h0); (forvar718 < (1'h0)); forvar718 = (forvar718 + (1'h1)))
                    begin
                      reg719 <= $unsigned((|reg719[(3'h7):(1'h0)]));
                      reg720 <= (~|$unsigned((+(forvar727 && reg717))));
                      reg721 <= $signed({(&{(8'h9c)})});
                      reg722 <= {$signed(reg709)};
                    end
                end
              for (forvar723 = (1'h0); (forvar723 < (2'h2)); forvar723 = (forvar723 + (1'h1)))
                begin
                  for (forvar724 = (1'h0); (forvar724 < (2'h3)); forvar724 = (forvar724 + (1'h1)))
                    begin
                      reg725 <= {(^reg704[(3'h4):(2'h3)])};
                    end
                  reg726 <= $signed($unsigned(reg732));
                  if ($unsigned((8'h9e)))
                    begin
                      reg727 <= $signed(forvar723[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg727 <= $signed({((forvar740 ? reg720 : forvar734) ?
                              (reg735 ?
                                  reg721 : forvar737) : $signed(reg726))});
                      reg728 <= reg713[(3'h7):(3'h6)];
                    end
                  for (forvar729 = (1'h0); (forvar729 < (1'h1)); forvar729 = (forvar729 + (1'h1)))
                    begin
                      reg730 <= (!{((reg716 ?
                              (8'hb3) : reg721) + $signed(reg720))});
                      reg731 <= forvar711[(2'h2):(1'h1)];
                      reg732 <= forvar713;
                      reg733 <= $unsigned({((reg730 ? reg736 : reg707) ?
                              $signed(reg743) : $unsigned(wire13))});
                    end
                end
            end
          for (forvar747 = (1'h0); (forvar747 < (1'h0)); forvar747 = (forvar747 + (1'h1)))
            begin
              if (forvar718)
                begin
                  if ($unsigned(((^$signed(reg727)) ?
                      (reg716[(1'h1):(1'h1)] == (~|reg744)) : ($unsigned(reg705) - reg713))))
                    begin
                      reg748 <= $signed((((|reg744) <<< (forvar745 <<< (8'hba))) == (~|(forvar725 ?
                          reg739 : wire12))));
                      reg749 <= {{$signed((reg708 ? forvar737 : wire11))}};
                    end
                  else
                    begin
                      reg748 <= forvar718[(1'h0):(1'h0)];
                      reg749 <= ($signed($signed($unsigned(reg748))) ?
                          $signed(((wire11 ? (8'haa) : reg709) ?
                              $signed((8'ha6)) : wire11[(3'h4):(2'h2)])) : (((reg720 ?
                                  forvar723 : reg731) == (!reg714)) ?
                              reg710 : ($signed(wire14) != ((8'ha5) && reg733))));
                      reg750 <= $unsigned((+{$signed(wire13)}));
                    end
                  for (forvar751 = (1'h0); (forvar751 < (2'h3)); forvar751 = (forvar751 + (1'h1)))
                    begin
                      reg752 <= reg708[(3'h4):(2'h2)];
                      reg753 <= reg723;
                      reg754 <= $signed({reg722});
                      reg755 <= (wire8 || forvar747[(2'h2):(1'h0)]);
                    end
                  if (($signed(reg705) ? reg733[(4'hb):(4'hb)] : forvar733))
                    begin
                      reg756 <= forvar711[(3'h4):(1'h0)];
                      reg757 <= $signed(($unsigned((8'h9c)) ?
                          ((reg753 ^~ reg726) && (forvar727 ?
                              forvar734 : wire11)) : ((~^reg733) ?
                              reg703[(1'h1):(1'h1)] : $signed(wire14))));
                    end
                  else
                    begin
                      reg756 <= (~|reg708);
                      reg757 <= $unsigned((reg707 ?
                          forvar703[(3'h6):(2'h2)] : reg704));
                      reg758 <= $unsigned(reg734);
                      reg759 <= {$unsigned((!$signed(reg749)))};
                    end
                  for (forvar760 = (1'h0); (forvar760 < (1'h1)); forvar760 = (forvar760 + (1'h1)))
                    begin
                      reg761 <= (&(|(+$unsigned(wire701))));
                      reg762 <= (~&$signed((|reg735)));
                    end
                end
              else
                begin
                  if (forvar705)
                    begin
                      reg748 <= ($signed(reg710[(3'h5):(3'h4)]) | ((reg744[(3'h4):(2'h3)] >>> ((8'hb4) ?
                          reg735 : reg762)) <<< forvar708[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg748 <= (-forvar725[(2'h3):(1'h1)]);
                      reg749 <= forvar734;
                      reg750 <= (~&reg733);
                      reg751 <= ((~$unsigned(reg753[(1'h0):(1'h0)])) << ((forvar718[(1'h0):(1'h0)] == reg756[(4'ha):(2'h2)]) + $signed(reg761[(2'h3):(2'h3)])));
                    end
                end
              if ({($unsigned(reg724) ? {wire13} : reg711)})
                begin
                  if ($unsigned((($signed(reg723) ?
                      (&reg721) : (reg757 ?
                          reg717 : forvar724)) & {reg727[(2'h2):(1'h0)]})))
                    begin
                      reg763 <= reg751[(2'h2):(1'h1)];
                      reg764 <= $signed((((forvar708 >>> forvar725) || (reg731 || forvar727)) ?
                          ((reg730 ^ reg733) >= reg757) : $signed($unsigned(forvar708))));
                    end
                  else
                    begin
                      reg763 <= ((|$unsigned({reg715})) >= $unsigned($unsigned(reg715)));
                      reg764 <= reg751;
                      reg765 <= ((8'hb2) ?
                          reg729 : (($signed(reg757) >= (+reg752)) >= $unsigned(forvar713)));
                      reg766 <= $unsigned((reg744 ?
                          (+$unsigned((8'had))) : (8'hb3)));
                    end
                end
              else
                begin
                  for (forvar763 = (1'h0); (forvar763 < (2'h2)); forvar763 = (forvar763 + (1'h1)))
                    begin
                      reg764 <= (^(((^reg728) ?
                          forvar760 : (!reg750)) * ((reg766 ?
                          (8'hb8) : reg765) ~^ $unsigned(reg705))));
                      reg765 <= reg729[(3'h5):(2'h3)];
                      reg766 <= $signed({reg755});
                      reg767 <= {$unsigned(($unsigned(reg763) > (reg746 ?
                              (8'h9c) : reg707)))};
                    end
                  for (forvar768 = (1'h0); (forvar768 < (1'h1)); forvar768 = (forvar768 + (1'h1)))
                    begin
                      reg769 <= (reg718 || ((~(8'hb6)) ?
                          $unsigned((|reg706)) : reg704));
                      reg770 <= (+(+(+(~|reg758))));
                    end
                  if ((reg725[(2'h3):(1'h1)] || reg756[(4'hc):(4'hb)]))
                    begin
                      reg771 <= forvar763[(2'h3):(1'h1)];
                    end
                  else
                    begin
                      reg771 <= {{$unsigned({(8'haf)})}};
                    end
                  if (((forvar725[(4'ha):(3'h7)] << forvar729) ?
                      forvar729[(4'hc):(1'h1)] : reg726))
                    begin
                      reg772 <= (forvar747[(4'he):(3'h6)] ? reg728 : wire11);
                      reg773 <= $signed(($unsigned(wire11[(4'h8):(3'h5)]) ?
                          $unsigned(forvar704) : (~^{reg706})));
                      reg774 <= reg705;
                    end
                  else
                    begin
                      reg772 <= $unsigned(reg709[(1'h1):(1'h0)]);
                      reg773 <= (({{(8'ha5)}} ? $signed(reg707) : (8'ha9)) ?
                          (reg772 | {$unsigned(forvar740)}) : (forvar704 == $signed($signed(reg709))));
                      reg774 <= reg709;
                      reg775 <= (!{(~|((8'hab) ? reg728 : reg731))});
                    end
                end
              for (forvar776 = (1'h0); (forvar776 < (2'h2)); forvar776 = (forvar776 + (1'h1)))
                begin
                  for (forvar777 = (1'h0); (forvar777 < (2'h3)); forvar777 = (forvar777 + (1'h1)))
                    begin
                      reg778 <= reg742;
                      reg779 <= $unsigned(reg769[(2'h2):(1'h0)]);
                    end
                  for (forvar780 = (1'h0); (forvar780 < (1'h1)); forvar780 = (forvar780 + (1'h1)))
                    begin
                      reg781 <= {$unsigned($signed((~&forvar733)))};
                      reg782 <= (!((8'hb4) >> ((reg763 << reg723) ?
                          (forvar724 * wire701) : reg748[(1'h1):(1'h1)])));
                      reg783 <= $unsigned(((~^$unsigned((8'hb4))) ?
                          $signed($unsigned(reg717)) : reg770[(2'h2):(2'h2)]));
                    end
                  if (((8'ha2) ?
                      (reg769 <<< (reg705[(2'h2):(1'h1)] + (reg748 ?
                          reg727 : reg770))) : $signed($unsigned((^reg713)))))
                    begin
                      reg784 <= forvar705;
                      reg785 <= reg711[(3'h4):(2'h2)];
                      reg786 <= $signed(($signed((~^forvar705)) ?
                          (reg759[(1'h1):(1'h1)] ?
                              (reg767 >>> forvar713) : reg708[(1'h1):(1'h0)]) : (((8'ha4) + (8'had)) ?
                              wire14[(3'h4):(1'h0)] : forvar747)));
                    end
                  else
                    begin
                      reg784 <= (!(8'hb8));
                      reg785 <= $unsigned((reg762 || ((wire9 && reg748) ?
                          (^~reg786) : reg719[(2'h3):(1'h0)])));
                      reg786 <= forvar723;
                      reg787 <= $signed($unsigned(reg762));
                    end
                  for (forvar788 = (1'h0); (forvar788 < (2'h2)); forvar788 = (forvar788 + (1'h1)))
                    begin
                      reg789 <= (^$unsigned($signed(forvar705[(1'h0):(1'h0)])));
                    end
                end
            end
          for (forvar790 = (1'h0); (forvar790 < (1'h0)); forvar790 = (forvar790 + (1'h1)))
            begin
              reg791 <= ((reg785[(3'h5):(1'h1)] != reg764[(4'h9):(3'h4)]) ?
                  ($unsigned((&(8'hba))) ^~ forvar727[(1'h1):(1'h1)]) : (-$unsigned({forvar780})));
            end
          for (forvar792 = (1'h0); (forvar792 < (1'h0)); forvar792 = (forvar792 + (1'h1)))
            begin
              for (forvar793 = (1'h0); (forvar793 < (2'h3)); forvar793 = (forvar793 + (1'h1)))
                begin
                  for (forvar794 = (1'h0); (forvar794 < (2'h3)); forvar794 = (forvar794 + (1'h1)))
                    begin
                      reg795 <= $signed($unsigned(($unsigned(reg718) >>> reg779[(4'he):(4'hd)])));
                      reg796 <= $unsigned($unsigned(((~&reg734) * $signed((8'h9c)))));
                      reg797 <= reg754;
                    end
                end
              reg798 <= ($signed(reg791[(4'ha):(3'h7)]) ?
                  (((8'hb2) ^ ((8'ha3) + reg766)) ?
                      $unsigned(reg731[(4'hb):(2'h3)]) : $unsigned({reg771})) : ({(~|reg754)} ^~ $unsigned($signed((8'h9c)))));
              for (forvar799 = (1'h0); (forvar799 < (1'h0)); forvar799 = (forvar799 + (1'h1)))
                begin
                  for (forvar800 = (1'h0); (forvar800 < (2'h2)); forvar800 = (forvar800 + (1'h1)))
                    begin
                      reg801 <= (^(^$signed((reg785 > (8'h9e)))));
                    end
                  for (forvar802 = (1'h0); (forvar802 < (1'h1)); forvar802 = (forvar802 + (1'h1)))
                    begin
                      reg803 <= reg754[(4'h9):(2'h2)];
                    end
                  if ($unsigned($unsigned((reg762[(1'h1):(1'h1)] ?
                      forvar780[(3'h6):(3'h4)] : $signed(reg744)))))
                    begin
                      reg804 <= $unsigned((((^forvar729) ?
                          (-reg785) : (!forvar776)) | reg711));
                      reg805 <= (^$unsigned(({reg724} ?
                          (|reg765) : (reg766 >= reg730))));
                      reg806 <= $signed(((~^(reg718 ?
                          forvar802 : reg789)) ^~ (reg773 >> (reg719 << reg706))));
                      reg807 <= {({(forvar792 ?
                                  reg706 : forvar723)} > {((8'ha7) >>> forvar740)})};
                    end
                  else
                    begin
                      reg804 <= (|({((8'haa) >>> (8'ha4))} ?
                          $unsigned((+reg770)) : $unsigned(reg735)));
                      reg805 <= (^reg722);
                      reg806 <= ((~$unsigned((~forvar723))) ?
                          $signed($unsigned($signed(reg767))) : $unsigned((8'h9c)));
                      reg807 <= (wire14[(1'h0):(1'h0)] < (($signed(reg757) ~^ $unsigned(wire9)) ?
                          ($signed(reg749) ?
                              (~^reg710) : (8'hb5)) : {$signed(reg803)}));
                    end
                  if ((8'haa))
                    begin
                      reg808 <= ($signed($signed($signed(reg774))) && forvar711[(2'h3):(1'h1)]);
                    end
                  else
                    begin
                      reg808 <= reg746[(3'h4):(3'h4)];
                      reg809 <= reg765;
                    end
                end
            end
        end
      for (forvar810 = (1'h0); (forvar810 < (2'h2)); forvar810 = (forvar810 + (1'h1)))
        begin
          for (forvar811 = (1'h0); (forvar811 < (1'h1)); forvar811 = (forvar811 + (1'h1)))
            begin
              for (forvar812 = (1'h0); (forvar812 < (1'h1)); forvar812 = (forvar812 + (1'h1)))
                begin
                  for (forvar813 = (1'h0); (forvar813 < (2'h2)); forvar813 = (forvar813 + (1'h1)))
                    begin
                      reg814 <= (&{(forvar738 * (~&reg753))});
                      reg815 <= {reg805};
                      reg816 <= {$unsigned($signed($unsigned(wire14)))};
                      reg817 <= (($signed(forvar780) ?
                          ($unsigned(forvar811) ?
                              $unsigned(reg718) : (|reg709)) : ((forvar711 >>> reg713) & (forvar792 >>> forvar780))) - ({(forvar740 << forvar763)} > {$unsigned(reg728)}));
                    end
                  for (forvar818 = (1'h0); (forvar818 < (1'h0)); forvar818 = (forvar818 + (1'h1)))
                    begin
                      reg819 <= $signed(forvar703);
                      reg820 <= $unsigned((wire14[(3'h7):(3'h4)] ?
                          $unsigned((8'ha2)) : reg718));
                    end
                  if ((reg752[(1'h1):(1'h1)] ? reg705[(3'h6):(1'h0)] : reg726))
                    begin
                      reg821 <= (reg774[(3'h4):(2'h2)] ?
                          forvar818[(1'h1):(1'h1)] : $unsigned((reg717[(2'h2):(2'h2)] ?
                              $unsigned(reg735) : (~^reg713))));
                      reg822 <= reg732[(4'ha):(2'h2)];
                      reg823 <= $signed(reg706[(1'h1):(1'h0)]);
                      reg824 <= ($signed((^~$unsigned(reg796))) ?
                          $signed($signed((|(8'hb8)))) : (8'haa));
                    end
                  else
                    begin
                      reg821 <= $unsigned(($unsigned((reg822 ~^ forvar776)) & reg803[(3'h5):(2'h3)]));
                      reg822 <= ((reg717[(2'h3):(2'h3)] ?
                              reg750 : $unsigned((reg806 && (8'hae)))) ?
                          $unsigned({(~^reg711)}) : (reg783[(4'h8):(4'h8)] <= ($unsigned((8'hac)) >>> (reg766 ?
                              forvar792 : reg763))));
                      reg823 <= $unsigned(reg784);
                      reg824 <= {((!((8'h9d) ? (8'hb5) : forvar723)) ?
                              ($signed(reg757) ~^ (^~reg733)) : (reg771[(1'h1):(1'h1)] ?
                                  $unsigned((8'ha5)) : (|forvar768)))};
                    end
                end
              if ($unsigned((reg816[(2'h2):(2'h2)] ?
                  reg765[(3'h5):(1'h1)] : $signed((wire10 ? reg757 : reg729)))))
                begin
                  for (forvar825 = (1'h0); (forvar825 < (1'h0)); forvar825 = (forvar825 + (1'h1)))
                    begin
                      reg826 <= $signed($unsigned(reg770));
                      reg827 <= forvar813[(3'h6):(3'h4)];
                      reg828 <= $unsigned(reg751[(1'h0):(1'h0)]);
                      reg829 <= (forvar734[(3'h6):(3'h5)] ?
                          reg809[(4'he):(4'h9)] : reg749[(1'h1):(1'h0)]);
                    end
                  for (forvar830 = (1'h0); (forvar830 < (2'h2)); forvar830 = (forvar830 + (1'h1)))
                    begin
                      reg831 <= (((|$signed(reg784)) ?
                          $signed($unsigned(wire8)) : (8'hb2)) == (!forvar705[(1'h0):(1'h0)]));
                      reg832 <= $unsigned(reg712[(2'h3):(1'h0)]);
                      reg833 <= wire9;
                      reg834 <= reg723[(2'h3):(2'h3)];
                    end
                  if ($unsigned(reg805))
                    begin
                      reg835 <= {$signed(({forvar737} ? (8'hb2) : {wire10}))};
                      reg836 <= reg823;
                      reg837 <= (|$unsigned(({forvar777} <<< (reg715 ?
                          forvar792 : reg732))));
                    end
                  else
                    begin
                      reg835 <= ({{reg732[(4'hc):(2'h3)]}} ?
                          (~(reg770[(3'h6):(1'h0)] ?
                              (reg835 ? reg775 : reg789) : (reg786 ?
                                  (8'ha0) : forvar723))) : $signed((&(reg836 && reg764))));
                      reg836 <= {{(8'haf)}};
                      reg837 <= $unsigned(reg736);
                    end
                  for (forvar838 = (1'h0); (forvar838 < (2'h3)); forvar838 = (forvar838 + (1'h1)))
                    begin
                      reg839 <= reg796[(4'h9):(3'h5)];
                    end
                end
              else
                begin
                  for (forvar825 = (1'h0); (forvar825 < (1'h0)); forvar825 = (forvar825 + (1'h1)))
                    begin
                      reg826 <= forvar703;
                    end
                  for (forvar827 = (1'h0); (forvar827 < (2'h2)); forvar827 = (forvar827 + (1'h1)))
                    begin
                      reg828 <= $signed($signed($signed((reg751 ?
                          reg758 : reg782))));
                      reg829 <= $unsigned(($unsigned({reg815}) ?
                          $signed(reg814[(1'h0):(1'h0)]) : ({reg774} ?
                              $unsigned(forvar812) : {forvar713})));
                      reg830 <= ($signed((forvar725 ?
                          $unsigned((8'haa)) : (reg712 + (8'ha6)))) > (($unsigned(reg730) <= (!reg808)) ?
                          (reg728 && ((8'ha8) == forvar733)) : $unsigned($unsigned(reg834))));
                      reg831 <= ((-(wire14 ^ $signed((8'ha2)))) < $signed($signed({reg727})));
                    end
                end
              for (forvar840 = (1'h0); (forvar840 < (1'h0)); forvar840 = (forvar840 + (1'h1)))
                begin
                  for (forvar841 = (1'h0); (forvar841 < (2'h3)); forvar841 = (forvar841 + (1'h1)))
                    begin
                      reg842 <= (^~$signed(((reg721 >= forvar745) ?
                          reg770 : (reg839 ? reg833 : (8'ha2)))));
                      reg843 <= $signed(reg728);
                    end
                end
            end
        end
      for (forvar844 = (1'h0); (forvar844 < (1'h1)); forvar844 = (forvar844 + (1'h1)))
        begin
          if (reg762)
            begin
              for (forvar845 = (1'h0); (forvar845 < (2'h2)); forvar845 = (forvar845 + (1'h1)))
                begin
                  for (forvar846 = (1'h0); (forvar846 < (2'h2)); forvar846 = (forvar846 + (1'h1)))
                    begin
                      reg847 <= (wire10 ?
                          $unsigned($signed(reg733[(1'h0):(1'h0)])) : forvar788[(2'h3):(2'h2)]);
                    end
                end
              for (forvar848 = (1'h0); (forvar848 < (1'h0)); forvar848 = (forvar848 + (1'h1)))
                begin
                  if (reg771[(2'h2):(2'h2)])
                    begin
                      reg849 <= reg753[(2'h3):(1'h1)];
                      reg850 <= (^$unsigned($signed((forvar848 <<< reg827))));
                      reg851 <= (8'hac);
                      reg852 <= {reg820[(3'h5):(2'h3)]};
                    end
                  else
                    begin
                      reg849 <= (~|$signed(reg850));
                      reg850 <= (8'ha1);
                      reg851 <= $unsigned(($signed(wire8) >> {$unsigned(reg730)}));
                      reg852 <= forvar727;
                    end
                  for (forvar853 = (1'h0); (forvar853 < (1'h0)); forvar853 = (forvar853 + (1'h1)))
                    begin
                      reg854 <= (((^(forvar734 ?
                          reg727 : (8'hb2))) ^ (+(|reg823))) == (((reg710 ?
                                  (8'ha9) : forvar737) ?
                              forvar790[(1'h0):(1'h0)] : reg817) ?
                          $signed((forvar800 <<< forvar734)) : (reg712[(1'h0):(1'h0)] ?
                              (forvar760 >>> reg749) : $unsigned((8'hb4)))));
                      reg855 <= (reg762[(2'h2):(1'h0)] ?
                          $unsigned(forvar745[(2'h3):(2'h2)]) : ({{(8'haa)}} >= reg803[(2'h2):(1'h1)]));
                    end
                  if ({$signed((8'hb3))})
                    begin
                      reg856 <= $unsigned(reg766);
                    end
                  else
                    begin
                      reg856 <= $signed((|forvar727));
                      reg857 <= ($signed(((reg806 ? reg820 : forvar840) ?
                          (|reg807) : wire9)) >>> ($unsigned($signed(reg772)) ^ reg721[(2'h2):(2'h2)]));
                    end
                  for (forvar858 = (1'h0); (forvar858 < (1'h0)); forvar858 = (forvar858 + (1'h1)))
                    begin
                      reg859 <= (^~(8'hb4));
                      reg860 <= $unsigned(reg766);
                    end
                end
              reg861 <= $signed($signed($unsigned((!reg765))));
            end
          else
            begin
              for (forvar845 = (1'h0); (forvar845 < (1'h1)); forvar845 = (forvar845 + (1'h1)))
                begin
                  for (forvar846 = (1'h0); (forvar846 < (2'h3)); forvar846 = (forvar846 + (1'h1)))
                    begin
                      reg847 <= {{(reg773 * reg787)}};
                    end
                  for (forvar848 = (1'h0); (forvar848 < (1'h1)); forvar848 = (forvar848 + (1'h1)))
                    begin
                      reg849 <= $signed(reg726[(2'h2):(2'h2)]);
                      reg850 <= ({((^reg789) ?
                                  wire8[(3'h7):(2'h3)] : (reg724 ?
                                      reg707 : reg850))} ?
                          reg798 : reg774[(2'h2):(2'h2)]);
                    end
                  if ({{reg779}})
                    begin
                      reg851 <= {$unsigned(reg711)};
                      reg852 <= ((-(~|forvar763)) ? reg769 : reg827);
                    end
                  else
                    begin
                      reg851 <= $signed((($signed(forvar723) == reg835) ?
                          (reg835 ?
                              $signed(wire9) : reg855[(2'h3):(1'h1)]) : reg801[(3'h5):(3'h5)]));
                      reg852 <= $unsigned((~$signed({reg720})));
                      reg853 <= $signed((forvar760[(3'h4):(2'h3)] ?
                          (((8'ha0) ? reg769 : forvar812) ?
                              $signed(reg771) : reg843) : ((reg791 ?
                              forvar844 : reg823) ^ $unsigned(forvar802))));
                      reg854 <= reg756[(2'h3):(1'h1)];
                    end
                end
              reg855 <= forvar727[(1'h1):(1'h1)];
            end
          for (forvar862 = (1'h0); (forvar862 < (1'h1)); forvar862 = (forvar862 + (1'h1)))
            begin
              if (reg826)
                begin
                  for (forvar863 = (1'h0); (forvar863 < (1'h1)); forvar863 = (forvar863 + (1'h1)))
                    begin
                      reg864 <= ($signed($unsigned((forvar713 || reg796))) - $unsigned(reg754));
                    end
                end
              else
                begin
                  reg863 <= $signed($unsigned($signed((forvar827 != (8'hb5)))));
                  for (forvar864 = (1'h0); (forvar864 < (2'h2)); forvar864 = (forvar864 + (1'h1)))
                    begin
                      reg865 <= reg739[(3'h4):(3'h4)];
                    end
                  reg866 <= $signed({$signed($signed(wire701))});
                  for (forvar867 = (1'h0); (forvar867 < (2'h2)); forvar867 = (forvar867 + (1'h1)))
                    begin
                      reg868 <= $unsigned(forvar776[(1'h1):(1'h1)]);
                      reg869 <= (&forvar848[(3'h6):(3'h6)]);
                    end
                end
              if (reg761[(1'h0):(1'h0)])
                begin
                  if ({(((reg711 ? reg706 : forvar813) ?
                          $unsigned(forvar802) : (~forvar705)) | ((reg789 <= reg823) > (reg820 >> forvar760)))})
                    begin
                      reg870 <= (8'hb2);
                      reg871 <= (reg797 ~^ $signed((8'ha7)));
                      reg872 <= reg851[(1'h0):(1'h0)];
                      reg873 <= $signed($signed(reg798));
                    end
                  else
                    begin
                      reg870 <= {{((reg864 ? reg759 : reg787) ?
                                  reg826 : (forvar827 ? wire9 : reg750))}};
                      reg871 <= $unsigned({$signed((forvar813 ?
                              forvar718 : forvar845))});
                    end
                  reg874 <= reg869[(4'ha):(1'h1)];
                  for (forvar875 = (1'h0); (forvar875 < (2'h3)); forvar875 = (forvar875 + (1'h1)))
                    begin
                      reg876 <= (reg773[(2'h2):(1'h1)] ?
                          ((8'hac) - $signed((forvar799 > (8'ha5)))) : $unsigned(reg850[(2'h2):(1'h1)]));
                      reg877 <= forvar840;
                      reg878 <= (&((!(reg861 ?
                          (8'haf) : (8'hba))) & reg754[(2'h3):(1'h1)]));
                    end
                  for (forvar879 = (1'h0); (forvar879 < (1'h0)); forvar879 = (forvar879 + (1'h1)))
                    begin
                      reg880 <= (^~(^~((reg820 ? reg744 : reg851) != (8'h9e))));
                      reg881 <= forvar848[(1'h1):(1'h1)];
                      reg882 <= ($signed((((8'had) <= reg860) * (wire10 ?
                              (8'hb3) : reg815))) ?
                          (($signed(reg861) ?
                                  forvar723[(1'h1):(1'h1)] : $signed((8'ha2))) ?
                              reg833[(1'h0):(1'h0)] : forvar729[(2'h3):(1'h0)]) : (8'h9e));
                      reg883 <= {(8'hab)};
                    end
                end
              else
                begin
                  reg870 <= ($signed(($unsigned((8'ha1)) ?
                      reg869[(4'h8):(1'h0)] : (reg713 ?
                          reg859 : forvar812))) >>> reg852[(3'h7):(1'h0)]);
                  if ($signed(reg785[(1'h0):(1'h0)]))
                    begin
                      reg871 <= {$unsigned(($signed(wire14) ?
                              forvar867 : ((8'hb8) ? reg772 : reg732)))};
                    end
                  else
                    begin
                      reg871 <= ($signed(((reg721 != reg808) ?
                          reg708 : (reg731 ?
                              reg826 : reg703))) == (reg798 & $signed({forvar800})));
                      reg872 <= ($signed(reg826[(2'h3):(1'h1)]) - {reg711});
                    end
                  for (forvar873 = (1'h0); (forvar873 < (2'h2)); forvar873 = (forvar873 + (1'h1)))
                    begin
                      reg874 <= reg781[(1'h0):(1'h0)];
                      reg875 <= (+((((8'ha7) ? reg859 : (8'h9d)) ?
                              reg855 : $unsigned(reg771)) ?
                          $unsigned($signed(forvar793)) : (~(8'ha7))));
                    end
                end
              for (forvar884 = (1'h0); (forvar884 < (2'h3)); forvar884 = (forvar884 + (1'h1)))
                begin
                  for (forvar885 = (1'h0); (forvar885 < (1'h0)); forvar885 = (forvar885 + (1'h1)))
                    begin
                      reg886 <= {reg805};
                      reg887 <= (^~$unsigned({(-reg703)}));
                    end
                  for (forvar888 = (1'h0); (forvar888 < (1'h0)); forvar888 = (forvar888 + (1'h1)))
                    begin
                      reg889 <= ({((^~forvar723) >= (reg763 ?
                              reg722 : forvar751))} + (^~(^~$unsigned(reg872))));
                    end
                  for (forvar890 = (1'h0); (forvar890 < (2'h3)); forvar890 = (forvar890 + (1'h1)))
                    begin
                      reg891 <= $unsigned(((~|reg856[(1'h1):(1'h0)]) ?
                          ($signed(reg865) ?
                              {reg847} : (reg835 ?
                                  reg816 : (8'hb6))) : (~reg878[(1'h1):(1'h0)])));
                      reg892 <= (($signed((^~reg727)) <<< reg761[(2'h3):(1'h0)]) ?
                          reg705 : wire10);
                      reg893 <= forvar733[(3'h6):(3'h6)];
                      reg894 <= ($signed((reg861 + ((8'hac) ?
                              wire701 : (8'ha0)))) ?
                          $unsigned({forvar863}) : {(~^reg787[(1'h0):(1'h0)])});
                    end
                end
            end
        end
      if (reg847)
        begin
          if ($signed((-(8'hb3))))
            begin
              if ($signed((|wire11)))
                begin
                  for (forvar895 = (1'h0); (forvar895 < (1'h1)); forvar895 = (forvar895 + (1'h1)))
                    begin
                      reg896 <= $unsigned({$signed($signed((8'hb8)))});
                    end
                  for (forvar897 = (1'h0); (forvar897 < (1'h1)); forvar897 = (forvar897 + (1'h1)))
                    begin
                      reg898 <= (reg756[(4'hd):(4'hd)] ?
                          ($signed((reg834 * forvar885)) ?
                              $unsigned({reg801}) : reg791[(3'h5):(3'h4)]) : reg824[(4'he):(4'hb)]);
                    end
                end
              else
                begin
                  if ($unsigned((~|reg789)))
                    begin
                      reg895 <= reg779[(2'h2):(1'h0)];
                    end
                  else
                    begin
                      reg895 <= reg876[(3'h7):(3'h5)];
                      reg896 <= reg871;
                      reg897 <= forvar811;
                    end
                  for (forvar898 = (1'h0); (forvar898 < (2'h2)); forvar898 = (forvar898 + (1'h1)))
                    begin
                      reg899 <= forvar768[(2'h2):(1'h0)];
                      reg900 <= reg828;
                      reg901 <= ({reg824} >> wire701);
                      reg902 <= $signed((&(&forvar884)));
                    end
                  for (forvar903 = (1'h0); (forvar903 < (2'h3)); forvar903 = (forvar903 + (1'h1)))
                    begin
                      reg904 <= ((($unsigned(reg717) ^~ forvar776) <<< $signed((forvar760 ?
                              wire14 : reg870))) ?
                          ($unsigned(reg827) ?
                              reg744[(1'h1):(1'h1)] : forvar846) : reg765[(2'h2):(1'h0)]);
                      reg905 <= {$unsigned(reg863)};
                    end
                end
            end
          else
            begin
              reg895 <= (8'hb0);
              for (forvar896 = (1'h0); (forvar896 < (1'h0)); forvar896 = (forvar896 + (1'h1)))
                begin
                  for (forvar897 = (1'h0); (forvar897 < (1'h1)); forvar897 = (forvar897 + (1'h1)))
                    begin
                      reg898 <= (~^(((-reg714) ?
                              {reg728} : (reg784 ? reg781 : reg850)) ?
                          ($signed(forvar863) ?
                              $unsigned(reg748) : $signed(reg865)) : (forvar812 ?
                              reg829 : forvar885)));
                    end
                  for (forvar899 = (1'h0); (forvar899 < (2'h2)); forvar899 = (forvar899 + (1'h1)))
                    begin
                      reg900 <= ($unsigned({$unsigned(reg742)}) >> $signed(($unsigned(reg863) || {forvar780})));
                      reg901 <= $signed(((forvar863 ~^ reg872[(3'h4):(1'h0)]) ?
                          $unsigned($signed(reg803)) : $signed(reg823[(1'h0):(1'h0)])));
                      reg902 <= reg783[(3'h5):(2'h2)];
                      reg903 <= $unsigned({reg806});
                    end
                end
            end
        end
      else
        begin
          if ((({reg723} <<< forvar704) ?
              (reg820[(3'h7):(1'h0)] << reg786[(1'h0):(1'h0)]) : ((forvar713[(2'h3):(2'h3)] ?
                      (reg746 ? reg898 : reg707) : $unsigned(forvar863)) ?
                  (~^(-reg875)) : (reg847[(2'h3):(1'h1)] != $signed(reg895)))))
            begin
              reg895 <= (8'h9c);
              if (reg772)
                begin
                  if ($unsigned($signed($signed($signed(forvar841)))))
                    begin
                      reg896 <= {$unsigned((~&(^(8'ha1))))};
                      reg897 <= (^~(-(forvar705 ?
                          (-reg736) : $signed(forvar737))));
                      reg898 <= ($unsigned($signed((&(8'hb2)))) ^ (!((reg758 || forvar818) + $signed((8'ha1)))));
                    end
                  else
                    begin
                      reg896 <= forvar725[(2'h2):(1'h1)];
                      reg897 <= (^~(~|($unsigned((8'ha4)) ?
                          (reg751 ? (8'h9c) : (8'had)) : $unsigned((8'ha2)))));
                      reg898 <= (!forvar813);
                    end
                  for (forvar899 = (1'h0); (forvar899 < (2'h2)); forvar899 = (forvar899 + (1'h1)))
                    begin
                      reg900 <= {((8'hb4) ?
                              ((^~reg732) ?
                                  reg887[(3'h4):(3'h4)] : {reg808}) : ($signed(reg775) ?
                                  reg806[(3'h4):(1'h1)] : $unsigned(forvar780)))};
                      reg901 <= {$signed($unsigned(reg898))};
                      reg902 <= $signed((&$unsigned((reg804 <= reg873))));
                    end
                end
              else
                begin
                  if (forvar760)
                    begin
                      reg896 <= ($unsigned(({reg898} ?
                          (forvar862 == reg713) : (~^reg843))) | reg847);
                    end
                  else
                    begin
                      reg896 <= reg878[(4'h8):(2'h3)];
                      reg897 <= $signed((-$signed((reg731 <= reg769))));
                      reg898 <= (!(+(+$signed(forvar838))));
                    end
                  reg899 <= (wire9[(1'h1):(1'h1)] ~^ ((~(&(8'haa))) && reg895[(4'h8):(3'h4)]));
                  reg900 <= $signed(reg828[(3'h7):(2'h3)]);
                  reg901 <= reg741[(1'h0):(1'h0)];
                end
            end
          else
            begin
              for (forvar895 = (1'h0); (forvar895 < (2'h2)); forvar895 = (forvar895 + (1'h1)))
                begin
                  if ((((8'ha2) ?
                      {$signed(reg883)} : ($signed(reg715) || (reg886 != reg708))) ^ {(8'ha5)}))
                    begin
                      reg896 <= ({reg781[(1'h0):(1'h0)]} || {($unsigned(reg827) >>> {reg720})});
                      reg897 <= $signed(reg860);
                      reg898 <= ((((forvar794 + reg843) ?
                                  forvar794[(3'h4):(1'h1)] : (~|reg705)) ?
                              ($signed(reg905) ?
                                  (forvar708 ~^ reg891) : $signed(reg826)) : ({reg847} == (reg746 == wire12))) ?
                          (8'hb4) : $unsigned($unsigned((reg764 ?
                              forvar751 : reg717))));
                    end
                  else
                    begin
                      reg896 <= $signed(forvar713[(3'h4):(2'h2)]);
                      reg897 <= ((!{((8'had) <<< forvar813)}) & $unsigned(forvar718[(2'h2):(1'h1)]));
                    end
                  if (($signed((reg836 ? ((8'ha6) <= reg742) : reg863)) ?
                      $unsigned($unsigned((forvar800 ?
                          (8'hac) : forvar885))) : ((!(^~forvar903)) ^ (^(reg757 ?
                          reg886 : reg781)))))
                    begin
                      reg899 <= reg855[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg899 <= (((reg876[(4'h8):(3'h4)] ~^ (forvar729 ?
                              reg891 : reg831)) ~^ reg849) ?
                          $signed(reg791[(4'hc):(2'h3)]) : reg753);
                      reg900 <= forvar705;
                      reg901 <= $unsigned($unsigned($unsigned((+reg763))));
                      reg902 <= (((-forvar848[(2'h2):(2'h2)]) ^ ($signed(reg795) ?
                          (reg708 >>> forvar777) : (reg767 ?
                              wire11 : reg723))) && ((~^$signed((8'hb7))) ?
                          ((reg901 ? reg889 : reg871) ~^ ((8'ha0) ?
                              reg805 : reg832)) : $unsigned($unsigned(reg852))));
                    end
                end
              for (forvar903 = (1'h0); (forvar903 < (2'h2)); forvar903 = (forvar903 + (1'h1)))
                begin
                  if (((~&$signed(reg815[(1'h0):(1'h0)])) ?
                      reg869 : (((forvar858 ? (8'ha4) : reg765) ?
                          (reg873 ? forvar825 : reg809) : (reg878 ?
                              reg713 : reg716)) >> (&{reg764}))))
                    begin
                      reg904 <= reg716;
                      reg905 <= ($unsigned(($unsigned(reg817) - $signed((8'ha6)))) ?
                          $signed(($signed(reg772) && $signed(reg787))) : $unsigned(($unsigned(reg895) <= $unsigned((8'hb6)))));
                      reg906 <= reg716[(2'h2):(2'h2)];
                    end
                  else
                    begin
                      reg904 <= (~|(~&(&(wire10 ? (8'ha8) : (8'hab)))));
                    end
                end
              if (reg826[(3'h6):(2'h3)])
                begin
                  for (forvar907 = (1'h0); (forvar907 < (1'h1)); forvar907 = (forvar907 + (1'h1)))
                    begin
                      reg908 <= $signed((forvar888 < $signed(reg743)));
                      reg909 <= reg856[(3'h6):(2'h2)];
                      reg910 <= reg870;
                    end
                  reg911 <= $unsigned(reg808);
                end
              else
                begin
                  for (forvar907 = (1'h0); (forvar907 < (1'h0)); forvar907 = (forvar907 + (1'h1)))
                    begin
                      reg908 <= $signed(((reg824 && forvar737[(1'h1):(1'h0)]) == reg730[(4'he):(1'h1)]));
                      reg909 <= (forvar751 >= reg712);
                      reg910 <= (($signed(reg754[(4'h8):(3'h5)]) ?
                              $signed((|(8'hae))) : (-(reg755 ^~ (8'ha7)))) ?
                          (~^({forvar879} > (reg806 >> reg798))) : ({(~forvar718)} ?
                              (8'ha6) : (~^$unsigned(reg821))));
                    end
                  if ((~^$unsigned($signed((reg730 ? reg900 : forvar725)))))
                    begin
                      reg911 <= ({{reg782[(4'h9):(4'h8)]}} >> (reg822 - $signed((forvar840 ?
                          reg746 : reg847))));
                      reg912 <= (~((forvar827 - $signed(reg911)) >= $signed($unsigned(reg843))));
                      reg913 <= (~|$unsigned((8'hac)));
                    end
                  else
                    begin
                      reg911 <= (reg849 ^~ $signed($unsigned(forvar751)));
                      reg912 <= reg869;
                      reg913 <= $signed(reg900);
                      reg914 <= {({$unsigned(forvar777)} >> ((wire701 * reg857) ?
                              {(8'h9c)} : forvar841[(4'h9):(2'h3)]))};
                    end
                  for (forvar915 = (1'h0); (forvar915 < (1'h0)); forvar915 = (forvar915 + (1'h1)))
                    begin
                      reg916 <= (&reg761[(3'h4):(2'h2)]);
                      reg917 <= $signed(reg764);
                      reg918 <= reg849;
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      if (forvar718)
        begin
          for (forvar919 = (1'h0); (forvar919 < (1'h0)); forvar919 = (forvar919 + (1'h1)))
            begin
              for (forvar920 = (1'h0); (forvar920 < (1'h1)); forvar920 = (forvar920 + (1'h1)))
                begin
                  reg921 <= (~(reg798[(3'h5):(2'h3)] ?
                      $unsigned(forvar841) : (8'ha6)));
                  for (forvar922 = (1'h0); (forvar922 < (2'h3)); forvar922 = (forvar922 + (1'h1)))
                    begin
                      reg923 <= ((reg772 != forvar899[(3'h4):(2'h3)]) + $signed(({(8'hb2)} * forvar763[(1'h0):(1'h0)])));
                      reg924 <= (!reg910);
                    end
                  if ($signed((reg713 ?
                      ({reg750} ? (!reg904) : {reg801}) : ((reg723 ?
                          reg906 : reg774) | (8'h9d)))))
                    begin
                      reg925 <= $signed((wire701[(2'h3):(2'h2)] >= {reg717[(1'h0):(1'h0)]}));
                    end
                  else
                    begin
                      reg925 <= {forvar740[(2'h3):(2'h2)]};
                      reg926 <= $signed({($unsigned(reg894) - forvar846)});
                      reg927 <= (~^{reg755[(2'h2):(2'h2)]});
                      reg928 <= ($signed((forvar863[(4'h9):(1'h0)] == (reg905 ?
                          reg829 : reg805))) & (^$signed((reg724 ?
                          (8'ha7) : forvar811))));
                    end
                end
              for (forvar929 = (1'h0); (forvar929 < (1'h1)); forvar929 = (forvar929 + (1'h1)))
                begin
                  for (forvar930 = (1'h0); (forvar930 < (1'h0)); forvar930 = (forvar930 + (1'h1)))
                    begin
                      reg931 <= reg906;
                    end
                end
              for (forvar932 = (1'h0); (forvar932 < (1'h1)); forvar932 = (forvar932 + (1'h1)))
                begin
                  if ($signed($unsigned($signed($signed(reg926)))))
                    begin
                      reg933 <= (($unsigned(reg913[(4'h9):(3'h7)]) ~^ ($signed(forvar930) << reg820[(1'h0):(1'h0)])) <<< (|$unsigned(reg823[(4'ha):(3'h5)])));
                      reg934 <= reg839;
                      reg935 <= {$signed((8'ha5))};
                      reg936 <= $unsigned((-({reg918} ?
                          reg733 : $unsigned((8'hb3)))));
                    end
                  else
                    begin
                      reg933 <= (~(~|((forvar799 ? forvar737 : reg755) ?
                          $signed(reg775) : ((8'hb5) <= forvar737))));
                      reg934 <= $unsigned(reg913[(2'h3):(2'h2)]);
                    end
                  for (forvar937 = (1'h0); (forvar937 < (1'h0)); forvar937 = (forvar937 + (1'h1)))
                    begin
                      reg938 <= {($unsigned({forvar704}) >> ((wire701 ?
                              forvar747 : reg820) ^ {wire13}))};
                      reg939 <= ($signed($signed((reg761 ?
                          reg791 : reg731))) * forvar825);
                      reg940 <= {(({reg791} ?
                              reg923[(3'h6):(3'h4)] : (reg853 & reg868)) * (8'hb6))};
                    end
                  if (reg708[(3'h5):(2'h2)])
                    begin
                      reg941 <= {(reg708 ? reg859 : reg729[(3'h7):(1'h0)])};
                      reg942 <= forvar788[(3'h6):(1'h0)];
                      reg943 <= $unsigned($signed(forvar713[(2'h2):(2'h2)]));
                      reg944 <= $unsigned($unsigned(forvar811));
                    end
                  else
                    begin
                      reg941 <= reg843[(4'h9):(3'h5)];
                    end
                end
            end
        end
      else
        begin
          reg919 <= (((reg916 & (forvar895 ? reg924 : reg868)) ?
              ((reg921 ? reg721 : reg801) < reg771) : ($unsigned(reg914) ?
                  $unsigned(reg766) : $signed((8'hb6)))) ^ reg748[(2'h3):(2'h3)]);
        end
      if ((reg933[(2'h3):(1'h0)] ? (-(^(reg938 >> forvar790))) : reg767))
        begin
          reg945 <= ($signed(($signed(reg717) ?
              (reg850 ? (8'ha1) : reg914) : reg717[(1'h0):(1'h0)])) != reg779);
        end
      else
        begin
          for (forvar945 = (1'h0); (forvar945 < (1'h1)); forvar945 = (forvar945 + (1'h1)))
            begin
              if ($signed((^(forvar827[(2'h2):(1'h1)] >> forvar897[(3'h4):(2'h2)]))))
                begin
                  if (((((^forvar827) ? (~reg815) : (~forvar768)) ?
                          ((~&(8'ha2)) ?
                              forvar708 : $unsigned(reg829)) : $unsigned((reg795 * forvar825))) ?
                      ($unsigned({reg854}) >> $unsigned((forvar740 == reg897))) : $unsigned(forvar895[(4'he):(1'h1)])))
                    begin
                      reg946 <= (forvar793 << {(~&$signed((8'hb4)))});
                      reg947 <= $unsigned((forvar723[(1'h1):(1'h1)] || {reg749}));
                      reg948 <= reg771;
                    end
                  else
                    begin
                      reg946 <= (|(8'hac));
                      reg947 <= ((^(~^(~^reg765))) ?
                          reg893 : $signed(((forvar922 >> (8'hb8)) > (&reg714))));
                      reg948 <= $signed((~&$unsigned(reg863[(3'h5):(1'h1)])));
                    end
                end
              else
                begin
                  reg946 <= (reg854[(1'h1):(1'h1)] ?
                      $unsigned(((!reg783) ?
                          {forvar793} : (forvar879 ?
                              reg849 : forvar810))) : forvar793);
                end
              if (($signed({$signed(reg773)}) * (8'ha8)))
                begin
                  reg949 <= {reg853[(2'h2):(1'h1)]};
                  if (($unsigned(((8'hb7) ?
                      reg705[(3'h5):(3'h4)] : forvar848[(2'h2):(2'h2)])) + (-($unsigned(reg878) ?
                      (~|reg748) : {wire10}))))
                    begin
                      reg950 <= $unsigned({$unsigned(reg889[(3'h4):(1'h1)])});
                      reg951 <= $signed((((reg880 == reg944) != forvar864) >>> ($unsigned((8'hab)) - $signed(forvar800))));
                      reg952 <= {$signed(reg733[(4'hf):(4'hd)])};
                      reg953 <= forvar858;
                    end
                  else
                    begin
                      reg950 <= (((reg798[(2'h2):(2'h2)] ?
                              reg735[(3'h7):(3'h5)] : $signed((8'hb8))) != $signed(((8'haf) ?
                              reg787 : reg753))) ?
                          reg939 : {($unsigned(forvar738) ? (8'haa) : reg944)});
                    end
                  for (forvar954 = (1'h0); (forvar954 < (1'h1)); forvar954 = (forvar954 + (1'h1)))
                    begin
                      reg955 <= $unsigned(forvar915);
                      reg956 <= (($unsigned((~&reg756)) ?
                          {reg876} : (^reg798)) << ({forvar776[(3'h7):(1'h1)]} && forvar888[(1'h1):(1'h1)]));
                      reg957 <= $signed(reg744[(2'h3):(2'h3)]);
                    end
                end
              else
                begin
                  for (forvar949 = (1'h0); (forvar949 < (2'h3)); forvar949 = (forvar949 + (1'h1)))
                    begin
                      reg950 <= reg832[(1'h0):(1'h0)];
                    end
                end
              reg958 <= (-(~reg746));
            end
          if (reg893[(4'he):(3'h4)])
            begin
              for (forvar959 = (1'h0); (forvar959 < (1'h0)); forvar959 = (forvar959 + (1'h1)))
                begin
                  if (({{reg816[(2'h2):(1'h0)]}} ^~ $unsigned(({(8'hb0)} & $signed(forvar838)))))
                    begin
                      reg960 <= (reg943 ?
                          (|((~&forvar793) - (reg905 ?
                              (8'hba) : (8'hb0)))) : (reg851 ?
                              reg751[(4'h8):(2'h3)] : ($signed(reg871) ^ (forvar920 ^ forvar780))));
                      reg961 <= $unsigned((reg720 ?
                          $unsigned(reg896) : $signed($unsigned(reg815))));
                      reg962 <= $signed($unsigned(($signed(reg742) >> (wire10 >> reg779))));
                    end
                  else
                    begin
                      reg960 <= reg934;
                      reg961 <= (+(~$unsigned(forvar919[(2'h2):(1'h1)])));
                    end
                  for (forvar963 = (1'h0); (forvar963 < (2'h2)); forvar963 = (forvar963 + (1'h1)))
                    begin
                      reg964 <= {$unsigned(forvar838)};
                      reg965 <= ($unsigned((&(reg832 ?
                          (8'h9e) : (8'h9e)))) == ($unsigned((+reg899)) ?
                          $signed((~^(8'hb5))) : ({reg715} >> (reg831 ?
                              reg891 : (8'hb2)))));
                      reg966 <= $signed((((forvar838 - (8'ha8)) ?
                          forvar932 : $unsigned((8'hba))) & $unsigned($unsigned(reg952))));
                      reg967 <= $unsigned(reg940);
                    end
                  reg968 <= $unsigned($unsigned(reg817));
                end
              for (forvar969 = (1'h0); (forvar969 < (1'h0)); forvar969 = (forvar969 + (1'h1)))
                begin
                  for (forvar970 = (1'h0); (forvar970 < (1'h0)); forvar970 = (forvar970 + (1'h1)))
                    begin
                      reg971 <= forvar845;
                      reg972 <= {$unsigned((!reg712))};
                      reg973 <= $unsigned($unsigned($signed({reg785})));
                    end
                  if (($signed({(reg769 * reg972)}) ?
                      (($unsigned((8'hba)) ?
                              $unsigned(forvar922) : (reg910 <= reg917)) ?
                          (|$unsigned(reg804)) : forvar896) : ((&(reg949 ?
                              reg866 : reg710)) ?
                          {(reg829 * reg943)} : reg854[(1'h1):(1'h0)])))
                    begin
                      reg974 <= reg769[(4'h8):(4'h8)];
                      reg975 <= $unsigned($signed(reg855[(2'h3):(1'h1)]));
                      reg976 <= (~^reg869[(4'h8):(4'h8)]);
                    end
                  else
                    begin
                      reg974 <= $signed(($signed({reg880}) >> reg713));
                      reg975 <= reg804;
                      reg976 <= $unsigned((^reg965[(1'h1):(1'h0)]));
                    end
                  reg977 <= forvar895[(1'h1):(1'h1)];
                  if (((((&wire13) ^ (wire13 > forvar704)) != $signed(reg900[(4'h9):(2'h2)])) >= reg831))
                    begin
                      reg978 <= $unsigned((^~(~&(wire8 ? (8'had) : reg952))));
                      reg979 <= (reg866 != reg887);
                      reg980 <= reg856[(1'h0):(1'h0)];
                      reg981 <= $unsigned(forvar768[(4'hf):(3'h7)]);
                    end
                  else
                    begin
                      reg978 <= (&(forvar788[(2'h3):(1'h1)] & $unsigned((forvar810 ?
                          (8'hb2) : reg949))));
                      reg979 <= {reg775};
                      reg980 <= (!(({forvar818} | (!forvar930)) ?
                          reg839 : ((reg736 ?
                              forvar723 : reg927) - (reg729 - reg952))));
                    end
                end
              if ((|reg949[(2'h2):(1'h0)]))
                begin
                  for (forvar982 = (1'h0); (forvar982 < (1'h0)); forvar982 = (forvar982 + (1'h1)))
                    begin
                      reg983 <= (~|reg746);
                    end
                end
              else
                begin
                  reg982 <= $unsigned($unsigned(($signed(reg957) && reg707[(4'h8):(3'h5)])));
                end
              if ($signed((reg878[(3'h5):(3'h5)] ?
                  forvar800[(4'ha):(4'h9)] : ($signed(reg979) && (reg834 <<< (8'ha1))))))
                begin
                  for (forvar984 = (1'h0); (forvar984 < (1'h1)); forvar984 = (forvar984 + (1'h1)))
                    begin
                      reg985 <= {(+(forvar777[(3'h6):(3'h6)] ?
                              forvar963[(3'h7):(2'h3)] : {forvar780}))};
                      reg986 <= {reg927[(1'h0):(1'h0)]};
                      reg987 <= $unsigned($signed(($unsigned(reg809) * reg957)));
                      reg988 <= (forvar740 ?
                          $signed(((forvar760 ^~ forvar959) ?
                              reg918[(3'h4):(1'h1)] : $signed(forvar738))) : {{$unsigned(forvar802)}});
                    end
                  if ((reg925 >>> $unsigned({(reg877 | reg831)})))
                    begin
                      reg989 <= (forvar945[(3'h4):(2'h3)] <= reg785[(1'h1):(1'h0)]);
                      reg990 <= reg725;
                      reg991 <= (8'hb9);
                      reg992 <= ((($signed(reg735) ?
                              $signed(forvar793) : reg971[(3'h6):(3'h4)]) ?
                          $unsigned({reg807}) : $unsigned((reg814 && forvar858))) - $signed(reg983[(2'h2):(1'h0)]));
                    end
                  else
                    begin
                      reg989 <= $signed($unsigned(forvar954[(1'h0):(1'h0)]));
                    end
                end
              else
                begin
                  if (((reg820 ?
                      $signed((forvar704 ?
                          reg770 : (8'ha2))) : (reg770[(2'h3):(1'h0)] != {reg839})) + $unsigned(((forvar873 ?
                      reg814 : forvar788) ^~ $unsigned((8'hba))))))
                    begin
                      reg984 <= $unsigned($unsigned((^(reg975 ?
                          reg834 : reg882))));
                      reg985 <= ($unsigned({forvar862[(3'h4):(1'h0)]}) || reg989[(3'h5):(1'h0)]);
                      reg986 <= $unsigned(forvar884);
                    end
                  else
                    begin
                      reg984 <= $signed((~(&(8'ha5))));
                    end
                  reg987 <= reg897;
                  reg988 <= $signed(($signed(forvar729) >= reg726[(1'h0):(1'h0)]));
                  for (forvar989 = (1'h0); (forvar989 < (1'h1)); forvar989 = (forvar989 + (1'h1)))
                    begin
                      reg990 <= $signed($unsigned(reg936[(1'h1):(1'h0)]));
                      reg991 <= (({(reg728 ~^ forvar718)} & {((8'haa) | forvar903)}) != (!reg720[(2'h2):(1'h0)]));
                      reg992 <= (reg779 ?
                          {reg831} : {(+reg874[(3'h4):(2'h3)])});
                      reg993 <= forvar776;
                    end
                end
            end
          else
            begin
              reg959 <= $unsigned((8'hb5));
              if ((reg781[(3'h4):(2'h2)] ? forvar790 : reg778[(4'h8):(4'h8)]))
                begin
                  if (({$unsigned({(8'hb5)})} ?
                      $signed({reg896[(2'h3):(2'h2)]}) : reg755[(3'h4):(2'h3)]))
                    begin
                      reg960 <= reg723[(2'h3):(2'h2)];
                      reg961 <= (8'h9e);
                      reg962 <= $unsigned($signed(($signed(reg864) ~^ forvar724[(1'h1):(1'h1)])));
                      reg963 <= reg839[(2'h3):(2'h3)];
                    end
                  else
                    begin
                      reg960 <= $unsigned((!$unsigned(reg953)));
                    end
                  if ((($unsigned($unsigned(forvar799)) ?
                          ($unsigned(forvar949) == reg957[(4'he):(3'h7)]) : $unsigned($unsigned(reg916))) ?
                      $signed(($signed(reg927) && forvar841)) : (^({reg878} << ((8'ha2) + reg928)))))
                    begin
                      reg964 <= reg735;
                      reg965 <= $unsigned(wire14[(2'h2):(1'h1)]);
                      reg966 <= $signed((^~$signed((wire11 ?
                          reg764 : reg759))));
                      reg967 <= forvar734[(4'he):(3'h6)];
                    end
                  else
                    begin
                      reg964 <= ($signed($unsigned($unsigned(forvar879))) & reg765[(1'h1):(1'h0)]);
                    end
                end
              else
                begin
                  for (forvar960 = (1'h0); (forvar960 < (1'h1)); forvar960 = (forvar960 + (1'h1)))
                    begin
                      reg961 <= {reg961[(4'he):(4'h9)]};
                      reg962 <= reg770[(1'h0):(1'h0)];
                      reg963 <= reg763;
                      reg964 <= $unsigned($unsigned($signed($signed((8'h9e)))));
                    end
                end
            end
          for (forvar994 = (1'h0); (forvar994 < (1'h1)); forvar994 = (forvar994 + (1'h1)))
            begin
              for (forvar995 = (1'h0); (forvar995 < (1'h1)); forvar995 = (forvar995 + (1'h1)))
                begin
                  reg996 <= {reg758[(1'h0):(1'h0)]};
                  reg997 <= (~|((^(~|reg866)) ?
                      ({forvar705} ?
                          reg771[(1'h1):(1'h1)] : forvar963) : ((~^(8'hb2)) * {reg961})));
                end
            end
        end
      for (forvar998 = (1'h0); (forvar998 < (1'h1)); forvar998 = (forvar998 + (1'h1)))
        begin
          if (reg964)
            begin
              for (forvar999 = (1'h0); (forvar999 < (2'h2)); forvar999 = (forvar999 + (1'h1)))
                begin
                  for (forvar1000 = (1'h0); (forvar1000 < (1'h1)); forvar1000 = (forvar1000 + (1'h1)))
                    begin
                      reg1001 <= {(~(8'hb7))};
                      reg1002 <= ((^~forvar740) <<< reg814);
                      reg1003 <= (reg887[(2'h3):(2'h2)] <= reg795[(2'h3):(2'h3)]);
                    end
                  for (forvar1004 = (1'h0); (forvar1004 < (1'h1)); forvar1004 = (forvar1004 + (1'h1)))
                    begin
                      reg1005 <= (reg980 >= (^~$signed((~&(8'haf)))));
                    end
                end
              reg1006 <= ($signed(({(8'h9f)} ?
                  ((8'haf) ?
                      forvar845 : forvar718) : reg947[(3'h7):(1'h0)])) << reg972[(1'h0):(1'h0)]);
              for (forvar1007 = (1'h0); (forvar1007 < (1'h1)); forvar1007 = (forvar1007 + (1'h1)))
                begin
                  reg1008 <= (8'ha1);
                  if ($signed($signed(forvar825)))
                    begin
                      reg1009 <= $unsigned(reg807[(3'h7):(3'h6)]);
                    end
                  else
                    begin
                      reg1009 <= $signed((($signed(forvar929) ?
                              $unsigned(reg948) : (forvar713 | forvar915)) ?
                          (reg816 || $signed(reg839)) : {wire14[(4'h8):(2'h3)]}));
                      reg1010 <= reg928[(1'h0):(1'h0)];
                      reg1011 <= $unsigned((reg981[(3'h4):(3'h4)] ?
                          {$unsigned(forvar896)} : $unsigned(((8'hb7) ?
                              wire8 : reg852))));
                      reg1012 <= $unsigned($unsigned(($unsigned((8'h9c)) ?
                          {reg707} : reg960)));
                    end
                  for (forvar1013 = (1'h0); (forvar1013 < (2'h3)); forvar1013 = (forvar1013 + (1'h1)))
                    begin
                      reg1014 <= $signed($signed((+$unsigned(reg983))));
                      reg1015 <= $signed($signed($unsigned((~forvar800))));
                      reg1016 <= (8'hb1);
                      reg1017 <= $unsigned($signed({(&reg874)}));
                    end
                end
              reg1018 <= $unsigned(((~|(reg988 ?
                  (8'ha7) : (8'hb1))) != ((|reg735) << (^~reg975))));
            end
          else
            begin
              reg999 <= reg819[(1'h1):(1'h1)];
              if ((-(reg803[(2'h3):(2'h3)] ? (+(~(8'ha6))) : $signed((8'ha8)))))
                begin
                  if ((-((8'hac) ?
                      reg707[(2'h2):(1'h1)] : forvar984[(1'h0):(1'h0)])))
                    begin
                      reg1000 <= $unsigned(reg912);
                    end
                  else
                    begin
                      reg1000 <= (!$signed($unsigned($unsigned(reg821))));
                      reg1001 <= $unsigned(((((8'ha6) != reg863) ?
                              $signed(reg1015) : $signed(reg993)) ?
                          $signed((reg732 ? (8'ha4) : reg842)) : {(reg997 ?
                                  reg854 : reg752)}));
                    end
                end
              else
                begin
                  if ($unsigned((reg758[(1'h0):(1'h0)] <<< ((&(8'hb3)) == (reg971 ?
                      reg880 : (8'hb5))))))
                    begin
                      reg1000 <= ($unsigned((~|$signed((8'hb5)))) ?
                          ($unsigned($signed(forvar994)) * reg986) : $signed((^~(forvar888 ?
                              forvar1007 : reg748))));
                      reg1001 <= reg727;
                      reg1002 <= $signed(reg1011[(3'h4):(1'h1)]);
                      reg1003 <= {$signed($signed({forvar867}))};
                    end
                  else
                    begin
                      reg1000 <= reg710[(2'h2):(2'h2)];
                      reg1001 <= $unsigned((~&forvar810));
                      reg1002 <= $signed(($unsigned({reg829}) ?
                          (~|$unsigned((8'hb9))) : $signed(wire11)));
                    end
                  if (reg771)
                    begin
                      reg1004 <= (!$signed($unsigned((reg916 - reg769))));
                      reg1005 <= $signed({$unsigned((8'hae))});
                      reg1006 <= ($signed((~&(reg787 ^ reg832))) ~^ $unsigned(forvar903[(1'h1):(1'h0)]));
                      reg1007 <= (reg952[(3'h7):(3'h5)] || ($signed((^~forvar932)) > reg1018));
                    end
                  else
                    begin
                      reg1004 <= ($unsigned(($unsigned(reg806) ~^ $unsigned(forvar999))) ?
                          $unsigned(wire14) : ((forvar737 >> {forvar794}) << $unsigned($signed(reg958))));
                      reg1005 <= (~^(~|reg988[(2'h2):(1'h1)]));
                    end
                end
              if ($unsigned(reg1014[(2'h3):(1'h1)]))
                begin
                  reg1008 <= reg721;
                end
              else
                begin
                  for (forvar1008 = (1'h0); (forvar1008 < (2'h2)); forvar1008 = (forvar1008 + (1'h1)))
                    begin
                      reg1009 <= (~&{(reg866 ?
                              (~reg982) : reg917[(3'h4):(3'h4)])});
                      reg1010 <= $unsigned({reg752[(3'h6):(2'h3)]});
                    end
                  for (forvar1011 = (1'h0); (forvar1011 < (2'h3)); forvar1011 = (forvar1011 + (1'h1)))
                    begin
                      reg1012 <= reg786[(1'h0):(1'h0)];
                      reg1013 <= ((~^$signed((+reg938))) ?
                          reg834 : ($unsigned((reg971 ?
                              reg953 : reg999)) > (|forvar915)));
                    end
                end
            end
          for (forvar1019 = (1'h0); (forvar1019 < (2'h2)); forvar1019 = (forvar1019 + (1'h1)))
            begin
              if ($unsigned(($unsigned((wire11 & reg904)) ?
                  reg772[(4'hc):(2'h3)] : reg843)))
                begin
                  for (forvar1020 = (1'h0); (forvar1020 < (1'h1)); forvar1020 = (forvar1020 + (1'h1)))
                    begin
                      reg1021 <= (~|$signed({$unsigned(reg759)}));
                      reg1022 <= {$unsigned($unsigned((reg853 >> forvar888)))};
                      reg1023 <= ((((^~reg833) ?
                          reg756 : forvar895[(4'hc):(4'ha)]) != $signed(reg868)) ^ (8'hb6));
                    end
                  for (forvar1024 = (1'h0); (forvar1024 < (2'h2)); forvar1024 = (forvar1024 + (1'h1)))
                    begin
                      reg1025 <= (((forvar885 > $signed(reg789)) ?
                              (~^reg968) : ((~&reg941) ?
                                  (~&reg719) : (reg847 ? (8'h9f) : reg828))) ?
                          reg883 : ($unsigned((reg964 & reg985)) - forvar888));
                    end
                  if ($unsigned($unsigned(($signed(reg975) & $unsigned(reg839)))))
                    begin
                      reg1026 <= (|((reg1023[(3'h4):(1'h1)] ?
                              $unsigned(reg955) : {forvar734}) ?
                          {((8'hb7) > forvar885)} : ((forvar793 ?
                              (8'ha3) : reg749) >>> $unsigned(reg724))));
                    end
                  else
                    begin
                      reg1026 <= reg873;
                      reg1027 <= ((~&(!{forvar1011})) ?
                          (&forvar1008[(2'h2):(1'h0)]) : forvar1019[(2'h3):(2'h2)]);
                      reg1028 <= forvar995;
                      reg1029 <= reg911;
                    end
                end
              else
                begin
                  if ($unsigned((reg732 ?
                      ((~reg787) <<< (8'hb6)) : $signed({forvar838}))))
                    begin
                      reg1020 <= (-reg951);
                      reg1021 <= $signed(reg1011[(3'h7):(2'h3)]);
                      reg1022 <= reg990[(2'h3):(1'h1)];
                      reg1023 <= $signed(($unsigned(wire9) ?
                          reg758 : (reg704 << forvar929[(2'h2):(1'h1)])));
                    end
                  else
                    begin
                      reg1020 <= (~forvar937);
                      reg1021 <= reg751;
                      reg1022 <= ((reg1003 ?
                          $unsigned((8'hb8)) : reg953) ^ $unsigned($signed((reg938 && (8'hba)))));
                    end
                  for (forvar1024 = (1'h0); (forvar1024 < (2'h2)); forvar1024 = (forvar1024 + (1'h1)))
                    begin
                      reg1025 <= ($unsigned($signed((forvar875 == reg895))) >= $unsigned($unsigned(((8'haf) ?
                          reg781 : forvar747))));
                      reg1026 <= $unsigned(reg1005[(4'hd):(2'h2)]);
                    end
                  if ((|$unsigned(($unsigned(reg717) ^~ forvar920))))
                    begin
                      reg1027 <= {((forvar844 ^~ reg966[(4'hd):(3'h4)]) <= ((reg872 == reg941) ?
                              ((8'h9c) ^~ reg786) : (reg983 || (8'hae))))};
                    end
                  else
                    begin
                      reg1027 <= (~reg727[(2'h3):(1'h1)]);
                      reg1028 <= forvar897[(4'h8):(1'h1)];
                      reg1029 <= ((reg986[(4'h9):(3'h5)] ?
                              $signed($signed((8'haa))) : $unsigned($signed(forvar919))) ?
                          {forvar811[(3'h7):(2'h3)]} : $unsigned(forvar776[(3'h5):(2'h2)]));
                    end
                end
            end
          for (forvar1030 = (1'h0); (forvar1030 < (2'h3)); forvar1030 = (forvar1030 + (1'h1)))
            begin
              for (forvar1031 = (1'h0); (forvar1031 < (2'h3)); forvar1031 = (forvar1031 + (1'h1)))
                begin
                  for (forvar1032 = (1'h0); (forvar1032 < (2'h3)); forvar1032 = (forvar1032 + (1'h1)))
                    begin
                      reg1033 <= (((reg819[(1'h0):(1'h0)] ?
                                  (-reg827) : (|forvar959)) ?
                              (8'ha3) : $unsigned((reg894 ?
                                  reg1009 : forvar727))) ?
                          forvar885 : (8'hac));
                      reg1034 <= ((^reg748[(3'h7):(1'h1)]) ?
                          reg966 : reg957[(4'h9):(3'h7)]);
                      reg1035 <= reg865[(1'h0):(1'h0)];
                    end
                end
              reg1036 <= ((forvar790[(2'h2):(1'h0)] <= ((+(8'hb4)) == $signed(reg916))) ?
                  {(&reg766[(4'h9):(4'h8)])} : reg714[(1'h0):(1'h0)]);
              for (forvar1037 = (1'h0); (forvar1037 < (2'h3)); forvar1037 = (forvar1037 + (1'h1)))
                begin
                  for (forvar1038 = (1'h0); (forvar1038 < (2'h2)); forvar1038 = (forvar1038 + (1'h1)))
                    begin
                      reg1039 <= $unsigned($signed({(^~reg1002)}));
                      reg1040 <= (~(reg814[(1'h1):(1'h1)] ?
                          reg944 : forvar1013[(3'h7):(2'h3)]));
                      reg1041 <= $signed($signed(reg911));
                      reg1042 <= (reg987[(4'h8):(3'h5)] ?
                          reg781[(3'h4):(1'h1)] : {$signed((&(8'hb9)))});
                    end
                end
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1043 = (1'h0); (forvar1043 < (1'h0)); forvar1043 = (forvar1043 + (1'h1)))
        begin
          if (wire14[(2'h3):(2'h3)])
            begin
              reg1044 <= (reg1015[(4'he):(1'h0)] ?
                  (^((forvar1037 ? (8'hac) : reg749) ?
                      forvar853[(2'h3):(1'h0)] : $unsigned(reg791))) : $signed($signed(forvar1043)));
              if ($unsigned($unsigned($unsigned((-reg1036)))))
                begin
                  if ((^$signed(({forvar959} || forvar713))))
                    begin
                      reg1045 <= ((+(^~$unsigned(reg750))) << ((wire10[(2'h3):(2'h3)] ?
                          reg997 : reg900[(3'h5):(1'h1)]) >= $signed($signed(reg826))));
                      reg1046 <= ((reg964[(1'h0):(1'h0)] ?
                              (~^(reg719 | (8'ha1))) : (&$signed(reg1029))) ?
                          reg796 : reg1023[(2'h3):(2'h3)]);
                    end
                  else
                    begin
                      reg1045 <= forvar810[(3'h4):(1'h1)];
                      reg1046 <= (~|forvar724[(1'h0):(1'h0)]);
                      reg1047 <= forvar1032[(1'h1):(1'h0)];
                    end
                  for (forvar1048 = (1'h0); (forvar1048 < (1'h1)); forvar1048 = (forvar1048 + (1'h1)))
                    begin
                      reg1049 <= $signed(reg899[(1'h1):(1'h1)]);
                      reg1050 <= $unsigned(reg1023[(2'h2):(2'h2)]);
                    end
                  for (forvar1051 = (1'h0); (forvar1051 < (1'h1)); forvar1051 = (forvar1051 + (1'h1)))
                    begin
                      reg1052 <= (^$signed(reg775[(3'h4):(2'h2)]));
                      reg1053 <= (^reg807);
                      reg1054 <= $unsigned(({forvar1004} != ($signed(reg779) ?
                          (reg796 ? reg865 : (8'hb8)) : (reg785 ?
                              reg721 : (8'hb3)))));
                      reg1055 <= (((reg983[(2'h2):(1'h0)] ?
                              (^~reg987) : reg1005[(1'h0):(1'h0)]) ?
                          {(+(8'hae))} : ((forvar845 ? forvar705 : reg716) ?
                              $signed(reg821) : (forvar1030 || (8'hab)))) <<< $signed(((8'ha4) ?
                          $unsigned(forvar813) : (forvar737 >>> (8'hac)))));
                    end
                end
              else
                begin
                  for (forvar1045 = (1'h0); (forvar1045 < (2'h2)); forvar1045 = (forvar1045 + (1'h1)))
                    begin
                      reg1046 <= {($unsigned((^~forvar949)) ?
                              $unsigned(forvar994[(4'ha):(2'h3)]) : reg960)};
                      reg1047 <= ($unsigned((8'hb6)) ?
                          {$unsigned($unsigned((8'hac)))} : $signed($unsigned({reg895})));
                      reg1048 <= forvar989;
                    end
                  for (forvar1049 = (1'h0); (forvar1049 < (2'h3)); forvar1049 = (forvar1049 + (1'h1)))
                    begin
                      reg1050 <= (reg892 ?
                          ($unsigned((~|wire10)) ?
                              reg991 : forvar838[(4'h8):(3'h7)]) : (^~($unsigned(reg982) ?
                              (~&reg936) : (|reg758))));
                    end
                  for (forvar1051 = (1'h0); (forvar1051 < (2'h2)); forvar1051 = (forvar1051 + (1'h1)))
                    begin
                      reg1052 <= {$signed(reg711[(4'hb):(1'h0)])};
                      reg1053 <= (^~(forvar907 ?
                          forvar745 : {forvar984[(3'h4):(2'h2)]}));
                    end
                  for (forvar1054 = (1'h0); (forvar1054 < (1'h0)); forvar1054 = (forvar1054 + (1'h1)))
                    begin
                      reg1055 <= ((~&reg903) ?
                          {(+reg782)} : reg1007[(1'h0):(1'h0)]);
                    end
                end
              reg1056 <= ((!(^{reg950})) ?
                  reg743[(2'h2):(1'h1)] : reg722[(2'h3):(2'h3)]);
              for (forvar1057 = (1'h0); (forvar1057 < (1'h0)); forvar1057 = (forvar1057 + (1'h1)))
                begin
                  for (forvar1058 = (1'h0); (forvar1058 < (1'h1)); forvar1058 = (forvar1058 + (1'h1)))
                    begin
                      reg1059 <= $unsigned(($unsigned((reg972 >= forvar799)) ?
                          (^~$signed(reg1002)) : reg960));
                      reg1060 <= forvar827;
                      reg1061 <= (((~|(reg821 ?
                          reg731 : forvar777)) - reg963) == {((&reg856) ?
                              $signed(reg891) : (reg872 ? reg843 : reg973))});
                      reg1062 <= (~&reg781);
                    end
                  if ($unsigned((forvar810[(3'h7):(1'h0)] ?
                      $signed((reg765 >>> forvar853)) : (~^(&(8'hb5))))))
                    begin
                      reg1063 <= reg860[(3'h6):(1'h0)];
                      reg1064 <= $signed({$signed($signed(reg814))});
                    end
                  else
                    begin
                      reg1063 <= $unsigned(reg934);
                      reg1064 <= reg770;
                    end
                  if (forvar960)
                    begin
                      reg1065 <= (-$signed((reg893[(4'h9):(4'h9)] <<< $unsigned(reg926))));
                      reg1066 <= ($signed(((~^reg910) > $signed(reg953))) << (reg948 ?
                          reg856 : $unsigned($signed(reg1062))));
                    end
                  else
                    begin
                      reg1065 <= forvar873;
                    end
                  for (forvar1067 = (1'h0); (forvar1067 < (1'h0)); forvar1067 = (forvar1067 + (1'h1)))
                    begin
                      reg1068 <= reg850;
                    end
                end
            end
          else
            begin
              if (forvar930)
                begin
                  reg1044 <= forvar725;
                  for (forvar1045 = (1'h0); (forvar1045 < (2'h2)); forvar1045 = (forvar1045 + (1'h1)))
                    begin
                      reg1046 <= (reg720[(2'h2):(1'h0)] ?
                          $unsigned((8'hb3)) : reg730);
                      reg1047 <= $signed((($unsigned(forvar708) ?
                              {reg1049} : {(8'hba)}) ?
                          ((forvar846 ^ forvar733) + reg886[(3'h6):(2'h2)]) : reg958[(4'hc):(4'h8)]));
                      reg1048 <= (($signed({(8'hb9)}) ?
                          ($unsigned(forvar711) ?
                              $unsigned((8'hb3)) : (forvar846 != reg903)) : reg1008[(3'h6):(3'h5)]) < forvar1008[(1'h1):(1'h1)]);
                      reg1049 <= forvar768;
                    end
                end
              else
                begin
                  reg1044 <= {$unsigned(reg923)};
                end
              for (forvar1050 = (1'h0); (forvar1050 < (1'h1)); forvar1050 = (forvar1050 + (1'h1)))
                begin
                  reg1051 <= ((reg857[(4'h8):(2'h2)] ?
                          (~^{reg744}) : $unsigned((reg723 ?
                              forvar740 : reg886))) ?
                      $signed(reg911) : {forvar945});
                  for (forvar1052 = (1'h0); (forvar1052 < (2'h2)); forvar1052 = (forvar1052 + (1'h1)))
                    begin
                      reg1053 <= {((~|(~(8'hb9))) << {reg774[(1'h0):(1'h0)]})};
                    end
                  if (((+({forvar875} == forvar802)) == ((8'hae) - {(reg712 > forvar812)})))
                    begin
                      reg1054 <= (reg773 || $unsigned($unsigned($unsigned(reg1003))));
                    end
                  else
                    begin
                      reg1054 <= reg948[(3'h4):(2'h3)];
                      reg1055 <= {((forvar1030[(4'ha):(4'ha)] ?
                                  reg765 : (reg971 + forvar863)) ?
                              reg865[(2'h2):(2'h2)] : forvar919)};
                      reg1056 <= (8'hba);
                      reg1057 <= $unsigned($signed((+$signed(reg1015))));
                    end
                end
              if ((~((reg905[(2'h2):(2'h2)] ?
                  (reg986 ?
                      forvar711 : forvar848) : (+reg944)) + forvar954[(3'h6):(1'h1)])))
                begin
                  reg1058 <= $unsigned((+$signed(reg826)));
                  for (forvar1059 = (1'h0); (forvar1059 < (2'h3)); forvar1059 = (forvar1059 + (1'h1)))
                    begin
                      reg1060 <= (reg804[(3'h4):(2'h3)] ? (8'ha5) : reg1035);
                      reg1061 <= reg819;
                      reg1062 <= $signed(((forvar858[(3'h7):(3'h5)] ?
                          forvar776[(1'h1):(1'h1)] : reg750[(4'he):(3'h5)]) | $signed((reg763 >>> reg763))));
                      reg1063 <= ($signed(($signed(reg1003) ?
                          (8'h9f) : (reg883 >>> reg804))) * (reg722[(2'h3):(2'h2)] != reg883));
                    end
                  reg1064 <= (~&forvar999[(2'h2):(1'h0)]);
                end
              else
                begin
                  if ({(($signed(reg754) <<< $signed(reg839)) ?
                          forvar1019 : ((reg859 ? reg892 : (8'ha8)) ?
                              $signed((8'ha5)) : $signed((8'ha7))))})
                    begin
                      reg1058 <= $signed($signed(reg1039[(3'h5):(2'h2)]));
                      reg1059 <= (forvar999[(1'h0):(1'h0)] || reg753);
                    end
                  else
                    begin
                      reg1058 <= $unsigned((((reg942 ? (8'hb3) : forvar802) ?
                              $unsigned(forvar845) : forvar724[(1'h0):(1'h0)]) ?
                          reg828[(1'h1):(1'h0)] : ({reg967} ^ $signed((8'hb7)))));
                      reg1059 <= (reg1016[(3'h7):(3'h6)] <= (8'hb2));
                      reg1060 <= (($unsigned(reg789[(1'h0):(1'h0)]) ?
                          reg703[(1'h0):(1'h0)] : reg889) >= forvar1031[(3'h6):(3'h4)]);
                      reg1061 <= reg1053[(3'h4):(2'h3)];
                    end
                  for (forvar1062 = (1'h0); (forvar1062 < (1'h1)); forvar1062 = (forvar1062 + (1'h1)))
                    begin
                      reg1063 <= reg931[(3'h7):(1'h1)];
                      reg1064 <= {reg855[(1'h0):(1'h0)]};
                      reg1065 <= $unsigned(reg955[(3'h6):(3'h4)]);
                    end
                  for (forvar1066 = (1'h0); (forvar1066 < (1'h1)); forvar1066 = (forvar1066 + (1'h1)))
                    begin
                      reg1067 <= (8'h9d);
                      reg1068 <= reg817;
                    end
                  for (forvar1069 = (1'h0); (forvar1069 < (2'h2)); forvar1069 = (forvar1069 + (1'h1)))
                    begin
                      reg1070 <= (|$signed($signed(reg1065[(3'h7):(3'h6)])));
                      reg1071 <= $signed((($unsigned(reg895) ?
                          $unsigned(forvar896) : $unsigned(reg1029)) >> $unsigned(forvar1032)));
                    end
                end
            end
          for (forvar1072 = (1'h0); (forvar1072 < (2'h2)); forvar1072 = (forvar1072 + (1'h1)))
            begin
              for (forvar1073 = (1'h0); (forvar1073 < (1'h1)); forvar1073 = (forvar1073 + (1'h1)))
                begin
                  for (forvar1074 = (1'h0); (forvar1074 < (2'h2)); forvar1074 = (forvar1074 + (1'h1)))
                    begin
                      reg1075 <= forvar841[(2'h2):(1'h1)];
                    end
                  reg1076 <= (((reg889[(3'h5):(3'h5)] + $unsigned(reg759)) ?
                          $signed((8'hb7)) : ((reg946 ?
                              reg870 : reg931) <= $unsigned(reg832))) ?
                      $signed($unsigned((~|reg753))) : (~|((+reg898) ?
                          forvar1069 : forvar1043[(3'h6):(3'h5)])));
                  reg1077 <= (|reg917[(2'h3):(2'h3)]);
                end
              reg1078 <= {($unsigned($signed(forvar1008)) ?
                      (((8'hba) ?
                          forvar724 : reg710) + reg1033[(2'h2):(2'h2)]) : ((-reg972) ?
                          {reg836} : {reg984}))};
              reg1079 <= $unsigned($unsigned(((reg795 >>> reg1010) | (reg986 ?
                  reg774 : forvar1024))));
              for (forvar1080 = (1'h0); (forvar1080 < (1'h1)); forvar1080 = (forvar1080 + (1'h1)))
                begin
                  for (forvar1081 = (1'h0); (forvar1081 < (1'h1)); forvar1081 = (forvar1081 + (1'h1)))
                    begin
                      reg1082 <= ((|((reg973 ?
                          forvar794 : (8'haa)) != ((8'h9e) | reg1071))) >> ({reg863[(4'hc):(2'h2)]} ?
                          reg765 : $signed($unsigned(reg945))));
                      reg1083 <= ((($signed(reg908) ?
                              forvar989 : (reg814 & forvar760)) ?
                          (reg942[(3'h5):(3'h4)] ?
                              $unsigned(reg718) : reg743) : reg783) > ((-(+wire9)) ?
                          ($signed(reg880) ?
                              $signed(reg1035) : (8'ha2)) : (~^{(8'hb8)})));
                      reg1084 <= (~&($signed((reg1045 ?
                          reg815 : forvar1031)) ^ $unsigned(reg751[(3'h7):(1'h0)])));
                      reg1085 <= reg893[(2'h3):(1'h1)];
                    end
                  for (forvar1086 = (1'h0); (forvar1086 < (1'h1)); forvar1086 = (forvar1086 + (1'h1)))
                    begin
                      reg1087 <= forvar969;
                      reg1088 <= $unsigned(($unsigned((-reg967)) ?
                          (!(8'haa)) : ((&reg734) & (reg987 ?
                              reg857 : reg834))));
                    end
                end
            end
          reg1089 <= (reg909 ^ $signed(reg801));
        end
      if ($unsigned($signed($unsigned($signed(forvar885)))))
        begin
          for (forvar1090 = (1'h0); (forvar1090 < (2'h2)); forvar1090 = (forvar1090 + (1'h1)))
            begin
              reg1091 <= ($unsigned($signed((reg847 ~^ forvar737))) ?
                  ((forvar888[(4'h8):(3'h4)] ^ reg1008) + (^~((8'ha2) ?
                      reg1005 : forvar1013))) : $unsigned(reg1087[(4'he):(4'ha)]));
              for (forvar1092 = (1'h0); (forvar1092 < (2'h3)); forvar1092 = (forvar1092 + (1'h1)))
                begin
                  if ((((&reg752[(1'h0):(1'h0)]) * (reg918 - $unsigned(wire14))) ?
                      reg1066[(4'h9):(3'h5)] : (~&((~&wire8) ?
                          forvar844 : (reg1079 && (8'ha1))))))
                    begin
                      reg1093 <= reg923;
                      reg1094 <= $unsigned($unsigned((-$unsigned(reg843))));
                      reg1095 <= {reg826[(4'hb):(3'h6)]};
                      reg1096 <= ((^~reg801) ?
                          wire14[(3'h5):(2'h2)] : forvar1090);
                    end
                  else
                    begin
                      reg1093 <= (^~((|{reg863}) <<< (^~{reg1095})));
                    end
                end
            end
          for (forvar1097 = (1'h0); (forvar1097 < (1'h1)); forvar1097 = (forvar1097 + (1'h1)))
            begin
              for (forvar1098 = (1'h0); (forvar1098 < (1'h1)); forvar1098 = (forvar1098 + (1'h1)))
                begin
                  for (forvar1099 = (1'h0); (forvar1099 < (2'h2)); forvar1099 = (forvar1099 + (1'h1)))
                    begin
                      reg1100 <= ($unsigned((~{reg1058})) ?
                          $unsigned(forvar780) : reg1048);
                    end
                  for (forvar1101 = (1'h0); (forvar1101 < (2'h3)); forvar1101 = (forvar1101 + (1'h1)))
                    begin
                      reg1102 <= $unsigned({reg710});
                      reg1103 <= forvar1080;
                      reg1104 <= reg1049[(2'h3):(1'h0)];
                      reg1105 <= $unsigned(({(reg831 <<< forvar1081)} ?
                          $signed((reg710 <= reg1093)) : (reg732[(4'hb):(3'h6)] ?
                              {reg1021} : (forvar840 == reg704))));
                    end
                  for (forvar1106 = (1'h0); (forvar1106 < (2'h3)); forvar1106 = (forvar1106 + (1'h1)))
                    begin
                      reg1107 <= reg815[(1'h0):(1'h0)];
                    end
                end
              reg1108 <= forvar725[(3'h4):(1'h0)];
              for (forvar1109 = (1'h0); (forvar1109 < (1'h1)); forvar1109 = (forvar1109 + (1'h1)))
                begin
                  for (forvar1110 = (1'h0); (forvar1110 < (2'h2)); forvar1110 = (forvar1110 + (1'h1)))
                    begin
                      reg1111 <= ($unsigned($unsigned(reg834)) ?
                          (($signed(forvar1032) ?
                                  $unsigned(reg1028) : reg834[(3'h4):(3'h4)]) ?
                              reg910 : (8'ha8)) : (^(forvar1097 ?
                              $unsigned(reg902) : $unsigned(forvar1057))));
                    end
                end
              if ($unsigned(reg829[(4'ha):(1'h0)]))
                begin
                  for (forvar1112 = (1'h0); (forvar1112 < (2'h2)); forvar1112 = (forvar1112 + (1'h1)))
                    begin
                      reg1113 <= (($unsigned(forvar998[(3'h4):(3'h4)]) ?
                              reg1083 : $signed($unsigned(reg899))) ?
                          (~^$unsigned(reg869)) : {($unsigned(forvar1032) ?
                                  {reg707} : reg830[(2'h3):(2'h2)])});
                      reg1114 <= {$unsigned((reg984 || (8'ha4)))};
                      reg1115 <= reg873;
                      reg1116 <= ($unsigned(reg722[(1'h1):(1'h1)]) - (~&((|forvar879) ?
                          $unsigned(forvar853) : $signed(reg1087))));
                    end
                  if ({({forvar867[(3'h6):(1'h0)]} ?
                          ((reg795 & forvar711) ?
                              (reg850 + reg851) : forvar969) : reg956)})
                    begin
                      reg1117 <= {(reg1111[(3'h6):(3'h4)] << ((forvar1074 || forvar1051) ?
                              $unsigned((8'hb4)) : $unsigned(reg1039)))};
                      reg1118 <= {(~&reg786)};
                    end
                  else
                    begin
                      reg1117 <= {{(forvar984[(1'h1):(1'h0)] ?
                                  (reg875 ? reg897 : (8'ha1)) : (reg772 ?
                                      reg764 : reg1044))}};
                      reg1118 <= (8'hab);
                    end
                end
              else
                begin
                  if ($signed(reg851[(1'h0):(1'h0)]))
                    begin
                      reg1112 <= (~$unsigned((^~$unsigned(reg847))));
                    end
                  else
                    begin
                      reg1112 <= ((((reg1026 > wire12) == (forvar1024 ~^ forvar896)) >> {(reg805 ?
                              (8'ha1) : forvar895)}) >> (~$unsigned($signed(reg761))));
                      reg1113 <= ((-(|{reg973})) ?
                          $signed(({forvar713} ?
                              (!(8'ha3)) : reg866[(1'h1):(1'h1)])) : (reg1046[(4'h8):(3'h7)] - forvar1008[(1'h1):(1'h1)]));
                      reg1114 <= {reg974[(4'hc):(4'hb)]};
                      reg1115 <= (&{{reg1026[(3'h6):(2'h3)]}});
                    end
                  for (forvar1116 = (1'h0); (forvar1116 < (2'h3)); forvar1116 = (forvar1116 + (1'h1)))
                    begin
                      reg1117 <= reg769[(4'h8):(3'h7)];
                      reg1118 <= reg852;
                      reg1119 <= (|$unsigned((&$signed((8'h9c)))));
                      reg1120 <= reg786[(1'h1):(1'h0)];
                    end
                  if ($unsigned($unsigned($signed((reg1039 ?
                      reg1001 : reg984)))))
                    begin
                      reg1121 <= {(-(forvar1097 >= $signed((8'hb9))))};
                    end
                  else
                    begin
                      reg1121 <= (reg1035 >> ($unsigned(((8'hb0) << reg990)) ?
                          ((~(8'ha4)) ?
                              forvar982[(1'h1):(1'h1)] : (~forvar827)) : $unsigned((reg709 ?
                              forvar922 : reg730))));
                      reg1122 <= (~|(((8'haa) == (|(8'ha4))) && $signed((reg712 ?
                          reg847 : reg900))));
                      reg1123 <= (8'h9d);
                    end
                  if ($signed(forvar799))
                    begin
                      reg1124 <= (((~&{reg1007}) >> ($signed(reg707) ?
                              (~&forvar825) : {reg965})) ?
                          reg897 : ((+reg752[(3'h6):(2'h3)]) == $unsigned((forvar737 * reg1049))));
                      reg1125 <= {$unsigned($unsigned(forvar1069))};
                      reg1126 <= forvar919;
                    end
                  else
                    begin
                      reg1124 <= forvar846;
                      reg1125 <= $unsigned(reg904[(2'h3):(2'h2)]);
                      reg1126 <= ((+(forvar1109 << $signed(forvar888))) ?
                          reg891[(1'h1):(1'h1)] : (reg987 ?
                              ((reg955 < (8'h9e)) ?
                                  reg860 : (wire8 >> (8'ha8))) : forvar1013));
                    end
                end
            end
        end
      else
        begin
          if (($unsigned(($unsigned(reg719) * {forvar1112})) ?
              reg909[(1'h0):(1'h0)] : (+$signed($signed(reg1039)))))
            begin
              for (forvar1090 = (1'h0); (forvar1090 < (1'h0)); forvar1090 = (forvar1090 + (1'h1)))
                begin
                  if (forvar794[(2'h3):(1'h1)])
                    begin
                      reg1091 <= forvar830;
                    end
                  else
                    begin
                      reg1091 <= reg1029[(1'h1):(1'h0)];
                      reg1092 <= ((8'ha1) ?
                          reg1057 : {$signed(forvar705[(3'h7):(1'h0)])});
                      reg1093 <= (!reg1070[(3'h5):(2'h2)]);
                    end
                  if ({{reg1042}})
                    begin
                      reg1094 <= reg1079;
                    end
                  else
                    begin
                      reg1094 <= $signed($unsigned(((forvar999 ?
                          (8'hb7) : reg830) >>> reg1021)));
                      reg1095 <= (reg783 && $unsigned(((&forvar844) >>> $signed((8'h9f)))));
                      reg1096 <= $unsigned(($signed(reg725[(2'h3):(2'h2)]) <<< forvar885));
                      reg1097 <= reg1076[(1'h0):(1'h0)];
                    end
                  for (forvar1098 = (1'h0); (forvar1098 < (2'h2)); forvar1098 = (forvar1098 + (1'h1)))
                    begin
                      reg1099 <= $signed(reg938);
                    end
                end
            end
          else
            begin
              reg1090 <= forvar989;
              if ((~|forvar724))
                begin
                  reg1091 <= $unsigned((~|{$signed(reg816)}));
                end
              else
                begin
                  if (reg724[(2'h2):(1'h0)])
                    begin
                      reg1091 <= reg1115[(1'h1):(1'h0)];
                    end
                  else
                    begin
                      reg1091 <= (reg853 >> $unsigned($signed((reg1112 <= reg1055))));
                    end
                  for (forvar1092 = (1'h0); (forvar1092 < (1'h1)); forvar1092 = (forvar1092 + (1'h1)))
                    begin
                      reg1093 <= {($unsigned(((8'hb3) ? reg757 : forvar800)) ?
                              (^~$signed(forvar777)) : ($unsigned(forvar919) >= reg1116))};
                      reg1094 <= reg1036[(1'h0):(1'h0)];
                      reg1095 <= (~forvar729);
                      reg1096 <= $unsigned(reg750);
                    end
                end
              if ($unsigned($unsigned($unsigned(reg1078[(1'h1):(1'h0)]))))
                begin
                  reg1097 <= reg806[(3'h4):(3'h4)];
                  reg1098 <= $unsigned($unsigned($unsigned($signed(reg923))));
                  reg1099 <= reg944[(1'h0):(1'h0)];
                  for (forvar1100 = (1'h0); (forvar1100 < (2'h2)); forvar1100 = (forvar1100 + (1'h1)))
                    begin
                      reg1101 <= ($signed((^~reg958)) + {$signed(((8'h9d) >> (8'ha4)))});
                      reg1102 <= {(^~{$unsigned(reg979)})};
                      reg1103 <= $unsigned($signed((^reg1094[(4'h8):(4'h8)])));
                      reg1104 <= $unsigned((^$signed(forvar853)));
                    end
                end
              else
                begin
                  if ($signed((!(~^((8'h9e) ? reg965 : reg1117)))))
                    begin
                      reg1097 <= (($signed(reg909) << $signed(reg1067[(1'h0):(1'h0)])) ?
                          $signed(reg1091[(1'h0):(1'h0)]) : reg852);
                      reg1098 <= $unsigned({{{reg938}}});
                      reg1099 <= $signed((^~{$unsigned(reg831)}));
                      reg1100 <= ($signed($unsigned({reg1017})) ?
                          reg806 : ((!(~^forvar733)) >>> reg755[(3'h4):(2'h2)]));
                    end
                  else
                    begin
                      reg1097 <= reg999;
                      reg1098 <= $signed({(~&$signed(reg881))});
                    end
                  for (forvar1101 = (1'h0); (forvar1101 < (2'h3)); forvar1101 = (forvar1101 + (1'h1)))
                    begin
                      reg1102 <= $signed($unsigned($unsigned($unsigned(forvar1013))));
                    end
                  if ($signed(reg782))
                    begin
                      reg1103 <= $unsigned(reg743);
                      reg1104 <= (^~forvar929);
                      reg1105 <= reg756;
                    end
                  else
                    begin
                      reg1103 <= $unsigned((|{(reg939 ? reg761 : reg1023)}));
                      reg1104 <= ((&{(8'hab)}) ?
                          {reg821} : ($signed((reg996 != reg1062)) ?
                              reg926 : (reg1023[(1'h1):(1'h0)] ?
                                  {reg842} : $unsigned(reg826))));
                      reg1105 <= reg1029;
                    end
                end
              if (reg911)
                begin
                  if ($signed((&(reg934[(2'h2):(2'h2)] >= reg927[(1'h0):(1'h0)]))))
                    begin
                      reg1106 <= $signed($signed(($unsigned(forvar1067) * {reg1049})));
                    end
                  else
                    begin
                      reg1106 <= (($signed((reg787 != (8'ha4))) ?
                          {(^(8'ha6))} : $unsigned($unsigned(reg939))) <<< (8'hab));
                      reg1107 <= $signed(reg707);
                      reg1108 <= $unsigned((+{reg912}));
                      reg1109 <= $signed(({$unsigned(reg1053)} ?
                          {$signed(reg706)} : (!$unsigned(forvar1049))));
                    end
                  for (forvar1110 = (1'h0); (forvar1110 < (1'h0)); forvar1110 = (forvar1110 + (1'h1)))
                    begin
                      reg1111 <= (!(8'hab));
                      reg1112 <= (~&((((8'hb1) ? wire10 : reg754) ?
                              (reg952 ?
                                  forvar875 : reg1079) : $unsigned(reg863)) ?
                          (reg843 ?
                              (~|forvar945) : $signed((8'hba))) : {reg987[(4'hb):(2'h3)]}));
                    end
                end
              else
                begin
                  if ($signed(reg869[(4'h8):(3'h4)]))
                    begin
                      reg1106 <= forvar1101;
                    end
                  else
                    begin
                      reg1106 <= $unsigned(($signed($unsigned(forvar903)) ?
                          reg720[(2'h3):(1'h1)] : forvar799[(4'h8):(4'h8)]));
                    end
                  reg1107 <= (reg909 && (8'had));
                end
            end
          if ($unsigned({{(forvar959 ^ (8'h9e))}}))
            begin
              for (forvar1113 = (1'h0); (forvar1113 < (2'h3)); forvar1113 = (forvar1113 + (1'h1)))
                begin
                  reg1114 <= $signed(reg823[(4'h9):(1'h0)]);
                  for (forvar1115 = (1'h0); (forvar1115 < (1'h0)); forvar1115 = (forvar1115 + (1'h1)))
                    begin
                      reg1116 <= ((+$signed($signed(reg714))) <= $signed($signed({wire10})));
                    end
                  for (forvar1117 = (1'h0); (forvar1117 < (2'h3)); forvar1117 = (forvar1117 + (1'h1)))
                    begin
                      reg1118 <= reg903[(2'h3):(1'h1)];
                      reg1119 <= $unsigned(reg789);
                    end
                  for (forvar1120 = (1'h0); (forvar1120 < (2'h3)); forvar1120 = (forvar1120 + (1'h1)))
                    begin
                      reg1121 <= forvar790[(2'h2):(2'h2)];
                      reg1122 <= forvar884;
                      reg1123 <= ($unsigned((reg964 ?
                          reg732 : {reg822})) <<< reg821[(2'h3):(2'h2)]);
                    end
                end
              reg1124 <= $unsigned(forvar1004[(1'h1):(1'h1)]);
              if ($unsigned(reg779[(3'h6):(1'h1)]))
                begin
                  for (forvar1125 = (1'h0); (forvar1125 < (1'h0)); forvar1125 = (forvar1125 + (1'h1)))
                    begin
                      reg1126 <= (reg751[(4'ha):(2'h3)] >> $signed(((reg990 ?
                              reg938 : (8'hb9)) ?
                          $signed(reg784) : $signed(reg1048))));
                      reg1127 <= ((forvar734[(3'h5):(1'h0)] - wire11[(4'h9):(3'h4)]) ?
                          (($unsigned((8'ha8)) * $signed(forvar862)) ^ (reg831 ?
                              $unsigned(reg758) : reg826[(4'h8):(3'h7)])) : (+(^~reg839[(3'h6):(3'h5)])));
                      reg1128 <= $unsigned($unsigned(reg989));
                    end
                  reg1129 <= reg980[(2'h2):(1'h0)];
                end
              else
                begin
                  reg1125 <= $unsigned(($signed((forvar1081 << reg1059)) ?
                      forvar708[(3'h5):(2'h2)] : ((reg870 ^~ reg718) >> (forvar1020 ?
                          (8'ha0) : reg897))));
                  if ((^~$unsigned((~|(&reg975)))))
                    begin
                      reg1126 <= forvar790;
                      reg1127 <= $unsigned((^~$signed((^reg1011))));
                      reg1128 <= forvar1109[(2'h3):(1'h0)];
                      reg1129 <= reg814[(1'h1):(1'h1)];
                    end
                  else
                    begin
                      reg1126 <= forvar862;
                      reg1127 <= $unsigned((^{reg1050}));
                    end
                  if ($unsigned((^~forvar1066[(3'h5):(2'h2)])))
                    begin
                      reg1130 <= (wire701 ?
                          forvar846 : (!$unsigned((~^forvar703))));
                    end
                  else
                    begin
                      reg1130 <= {(8'hb2)};
                      reg1131 <= {({reg729[(3'h6):(1'h0)]} >> forvar995[(4'hc):(3'h4)])};
                      reg1132 <= (~reg853);
                      reg1133 <= {(~^forvar848[(2'h2):(2'h2)])};
                    end
                  reg1134 <= ($signed($unsigned((reg798 ?
                      forvar885 : reg943))) || forvar884[(3'h4):(2'h2)]);
                end
            end
          else
            begin
              for (forvar1113 = (1'h0); (forvar1113 < (1'h0)); forvar1113 = (forvar1113 + (1'h1)))
                begin
                  for (forvar1114 = (1'h0); (forvar1114 < (1'h0)); forvar1114 = (forvar1114 + (1'h1)))
                    begin
                      reg1115 <= forvar747;
                    end
                  for (forvar1116 = (1'h0); (forvar1116 < (2'h3)); forvar1116 = (forvar1116 + (1'h1)))
                    begin
                      reg1117 <= $signed((reg1003 ?
                          (~{reg865}) : reg1058[(4'hc):(1'h1)]));
                    end
                end
              for (forvar1118 = (1'h0); (forvar1118 < (2'h2)); forvar1118 = (forvar1118 + (1'h1)))
                begin
                  if (reg744[(1'h0):(1'h0)])
                    begin
                      reg1119 <= reg1085[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg1119 <= ((reg1116[(2'h3):(1'h0)] <<< $unsigned((reg939 ?
                              reg925 : forvar984))) ?
                          ($unsigned((forvar989 >> reg927)) ?
                              $signed($signed(reg861)) : reg732) : (!((reg735 & reg755) ?
                              $unsigned(forvar725) : (^reg733))));
                      reg1120 <= ((~$unsigned({reg1105})) ?
                          $signed((8'hb1)) : $signed({reg791}));
                      reg1121 <= ($signed(reg944[(4'ha):(4'h8)]) && forvar800);
                      reg1122 <= $unsigned($signed({(forvar727 == forvar838)}));
                    end
                  for (forvar1123 = (1'h0); (forvar1123 < (1'h0)); forvar1123 = (forvar1123 + (1'h1)))
                    begin
                      reg1124 <= $unsigned({{(reg870 ? reg962 : reg1088)}});
                    end
                  if (($unsigned(reg1101) ? wire9 : $signed(reg808)))
                    begin
                      reg1125 <= reg1042;
                      reg1126 <= (reg767 & (~&reg957[(4'ha):(4'ha)]));
                    end
                  else
                    begin
                      reg1125 <= (~^$signed((reg1090[(1'h1):(1'h1)] ?
                          (forvar792 | reg726) : $signed(reg1089))));
                      reg1126 <= ($unsigned($unsigned({reg963})) ?
                          ($unsigned($signed((8'hae))) <= {((8'haf) ?
                                  reg842 : reg761)}) : $unsigned((8'hba)));
                      reg1127 <= {wire13};
                      reg1128 <= (($unsigned($unsigned(reg849)) ^~ (^reg1079[(4'h9):(4'h9)])) << ((~&(reg766 ?
                          (8'hb3) : reg901)) << (&reg961[(4'hd):(1'h0)])));
                    end
                end
              for (forvar1129 = (1'h0); (forvar1129 < (1'h1)); forvar1129 = (forvar1129 + (1'h1)))
                begin
                  for (forvar1130 = (1'h0); (forvar1130 < (2'h2)); forvar1130 = (forvar1130 + (1'h1)))
                    begin
                      reg1131 <= (~$signed(($signed(reg1099) - $unsigned(reg1130))));
                      reg1132 <= (reg826[(4'he):(4'h8)] ?
                          $signed(((!reg916) ?
                              (reg955 ?
                                  reg1133 : (8'h9f)) : reg1060)) : (($signed(reg1105) | reg965[(2'h2):(2'h2)]) ?
                              ($signed((8'hac)) ?
                                  (^~reg797) : $unsigned(reg755)) : reg940[(1'h1):(1'h0)]));
                      reg1133 <= reg988[(1'h0):(1'h0)];
                    end
                end
            end
        end
      if ((((~^reg731) ?
          $signed((8'ha2)) : reg1116[(4'ha):(2'h3)]) != $unsigned(reg1066[(2'h2):(1'h1)])))
        begin
          for (forvar1135 = (1'h0); (forvar1135 < (1'h0)); forvar1135 = (forvar1135 + (1'h1)))
            begin
              for (forvar1136 = (1'h0); (forvar1136 < (1'h1)); forvar1136 = (forvar1136 + (1'h1)))
                begin
                  reg1137 <= $unsigned(reg711[(4'hb):(1'h0)]);
                  if ($unsigned(reg824))
                    begin
                      reg1138 <= $unsigned($signed($unsigned(reg1049)));
                      reg1139 <= $unsigned((forvar963[(3'h5):(2'h2)] * reg819));
                    end
                  else
                    begin
                      reg1138 <= {$unsigned(reg870[(2'h3):(1'h0)])};
                      reg1139 <= (forvar1118[(4'h8):(3'h4)] < reg739);
                      reg1140 <= (({wire13[(2'h2):(1'h1)]} << $unsigned($unsigned(reg931))) ?
                          ($signed(forvar1090[(4'hb):(3'h6)]) ~^ reg1022[(3'h4):(2'h2)]) : $signed(($unsigned(reg711) ?
                              (forvar1048 || (8'hb6)) : (reg719 ?
                                  reg918 : reg1128))));
                    end
                  if (reg933[(3'h7):(2'h2)])
                    begin
                      reg1141 <= reg940[(3'h6):(1'h1)];
                    end
                  else
                    begin
                      reg1141 <= $unsigned((^reg756[(4'hc):(3'h4)]));
                      reg1142 <= (^reg1070[(2'h2):(1'h1)]);
                      reg1143 <= $signed((reg886 ?
                          (8'haa) : $unsigned(reg709)));
                      reg1144 <= (forvar890[(3'h6):(2'h3)] ?
                          $unsigned($unsigned((reg1040 ?
                              (8'haa) : reg1040))) : ($unsigned($signed(reg851)) ^~ forvar919));
                    end
                  if (({(~&(^reg1058))} == (!$signed((^~wire12)))))
                    begin
                      reg1145 <= reg918;
                      reg1146 <= $signed(($unsigned((~reg778)) & $unsigned({(8'hb9)})));
                    end
                  else
                    begin
                      reg1145 <= {$unsigned($unsigned((forvar1086 * reg988)))};
                    end
                end
              for (forvar1147 = (1'h0); (forvar1147 < (2'h2)); forvar1147 = (forvar1147 + (1'h1)))
                begin
                  reg1148 <= forvar945[(3'h6):(2'h2)];
                end
              if ($signed((^~reg1035)))
                begin
                  for (forvar1149 = (1'h0); (forvar1149 < (1'h1)); forvar1149 = (forvar1149 + (1'h1)))
                    begin
                      reg1150 <= {(reg861 == $signed(reg764[(3'h6):(2'h2)]))};
                    end
                end
              else
                begin
                  reg1149 <= reg703[(1'h1):(1'h0)];
                  if ((^~reg1111))
                    begin
                      reg1150 <= (((8'hb8) >>> reg1041) ?
                          reg726[(2'h3):(2'h3)] : (~&$signed($unsigned((8'hb9)))));
                      reg1151 <= (^~(^$signed((reg851 != reg900))));
                    end
                  else
                    begin
                      reg1150 <= forvar740[(3'h5):(2'h2)];
                      reg1151 <= $signed((8'h9e));
                      reg1152 <= ((+forvar1024[(4'h8):(4'h8)]) ?
                          (~|{(reg876 ? reg795 : reg981)}) : $unsigned(reg837));
                    end
                  for (forvar1153 = (1'h0); (forvar1153 < (1'h0)); forvar1153 = (forvar1153 + (1'h1)))
                    begin
                      reg1154 <= $unsigned(forvar982[(2'h3):(1'h0)]);
                      reg1155 <= ($unsigned(reg1000) << forvar1125);
                      reg1156 <= reg997[(1'h0):(1'h0)];
                      reg1157 <= reg905;
                    end
                  for (forvar1158 = (1'h0); (forvar1158 < (1'h0)); forvar1158 = (forvar1158 + (1'h1)))
                    begin
                      reg1159 <= $signed($signed(($unsigned(reg1006) ?
                          forvar875 : {reg789})));
                      reg1160 <= reg913[(4'hb):(3'h4)];
                      reg1161 <= ({reg1005} | $signed($unsigned(forvar777[(2'h3):(1'h0)])));
                    end
                end
            end
        end
      else
        begin
          if (reg710)
            begin
              for (forvar1135 = (1'h0); (forvar1135 < (1'h1)); forvar1135 = (forvar1135 + (1'h1)))
                begin
                  reg1136 <= reg769[(3'h6):(3'h4)];
                  if ({$unsigned((|$signed((8'ha7))))})
                    begin
                      reg1137 <= (~&((8'h9f) ?
                          $signed(reg831[(1'h0):(1'h0)]) : $signed(forvar729)));
                      reg1138 <= reg893;
                      reg1139 <= reg823;
                      reg1140 <= $signed($signed($unsigned(forvar723[(2'h2):(1'h0)])));
                    end
                  else
                    begin
                      reg1137 <= $unsigned(($signed(forvar818[(1'h0):(1'h0)]) ^~ reg1059[(3'h7):(2'h2)]));
                      reg1138 <= reg927[(2'h3):(1'h1)];
                      reg1139 <= (reg1028 || $unsigned($unsigned((reg1116 || reg1100))));
                      reg1140 <= $signed((reg785 * $signed((reg945 - forvar1050))));
                    end
                end
            end
          else
            begin
              if (($unsigned((forvar897[(2'h2):(1'h0)] <<< $signed(reg1012))) <= {forvar763}))
                begin
                  if (reg1091)
                    begin
                      reg1135 <= ($signed($unsigned((forvar793 ~^ reg1049))) ?
                          (~^((forvar1125 ~^ reg1106) ?
                              reg1108 : (forvar776 ?
                                  reg710 : forvar790))) : forvar1136[(4'hd):(2'h3)]);
                      reg1136 <= (reg868[(4'ha):(4'h8)] || reg948[(2'h3):(1'h1)]);
                      reg1137 <= (reg877[(3'h7):(1'h0)] ^ $unsigned(($signed(reg1144) != $unsigned(reg727))));
                    end
                  else
                    begin
                      reg1135 <= $unsigned(($signed((reg983 ?
                          (8'h9c) : reg1035)) + $signed($signed(reg749))));
                      reg1136 <= (reg979 >> ((reg831 ?
                          forvar1114[(3'h4):(3'h4)] : $unsigned(reg1006)) & ((~reg1152) ?
                          (^~forvar1125) : ((8'hae) + forvar999))));
                      reg1137 <= forvar768[(2'h3):(2'h2)];
                    end
                end
              else
                begin
                  if ((reg861[(1'h1):(1'h0)] ?
                      (+reg836) : $signed(($unsigned(reg905) ?
                          $signed(forvar1072) : $signed(reg955)))))
                    begin
                      reg1135 <= reg741[(3'h7):(3'h5)];
                      reg1136 <= ((reg824 < ($signed(reg814) ?
                          reg952 : forvar729)) * (reg868 & (^~(+forvar1115))));
                      reg1137 <= (~&$signed($unsigned($unsigned(forvar963))));
                      reg1138 <= $unsigned((($unsigned(reg1076) ?
                              {reg973} : reg1161) ?
                          ((8'hab) >>> $unsigned(reg803)) : (-(forvar1007 - reg1006))));
                    end
                  else
                    begin
                      reg1135 <= $signed($signed(forvar725));
                      reg1136 <= ((~|reg1000[(1'h1):(1'h0)]) || $signed($unsigned(reg1028)));
                      reg1137 <= reg731;
                    end
                  reg1139 <= $unsigned(($signed(reg955) <<< ($signed(reg823) - (reg866 ?
                      reg934 : reg933))));
                  if ($signed($signed((!forvar718))))
                    begin
                      reg1140 <= (($signed($signed(reg1048)) ?
                              forvar724[(1'h1):(1'h1)] : $unsigned($unsigned(forvar920))) ?
                          $unsigned(($signed(reg806) < forvar848[(2'h2):(1'h0)])) : ($signed((forvar989 ?
                                  forvar1098 : reg710)) ?
                              (&(reg861 && forvar813)) : $unsigned({reg918})));
                      reg1141 <= (+$unsigned(((~^reg822) & ((8'ha4) <<< forvar922))));
                    end
                  else
                    begin
                      reg1140 <= (reg1009[(1'h0):(1'h0)] ?
                          ({$signed(reg924)} ?
                              $signed(reg1014[(1'h0):(1'h0)]) : $unsigned((forvar794 ?
                                  reg1137 : reg1149))) : reg767[(2'h2):(2'h2)]);
                      reg1141 <= wire13[(2'h2):(1'h0)];
                    end
                end
            end
          reg1142 <= forvar800;
          reg1143 <= $signed(reg1136);
          reg1144 <= (~wire701[(4'ha):(3'h7)]);
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(reg1087[(4'hc):(4'hb)]))
        begin
          reg1162 <= {$unsigned(($unsigned(forvar768) ?
                  reg1068 : (~^forvar864)))};
          if ((reg1095 ?
              ((8'had) ?
                  reg1022 : (reg822 ?
                      forvar724 : $signed(reg914))) : $unsigned({reg1089[(2'h2):(1'h1)]})))
            begin
              reg1163 <= $unsigned($signed({(+reg1109)}));
              for (forvar1164 = (1'h0); (forvar1164 < (2'h3)); forvar1164 = (forvar1164 + (1'h1)))
                begin
                  for (forvar1165 = (1'h0); (forvar1165 < (2'h3)); forvar1165 = (forvar1165 + (1'h1)))
                    begin
                      reg1166 <= $signed((((-reg1151) ?
                              (reg928 ?
                                  reg964 : forvar777) : reg899[(1'h0):(1'h0)]) ?
                          (&(forvar884 ?
                              (8'ha8) : wire13)) : reg955[(2'h3):(1'h0)]));
                    end
                end
            end
          else
            begin
              reg1163 <= (-reg1025[(4'he):(4'he)]);
            end
        end
      else
        begin
          for (forvar1162 = (1'h0); (forvar1162 < (1'h1)); forvar1162 = (forvar1162 + (1'h1)))
            begin
              for (forvar1163 = (1'h0); (forvar1163 < (1'h0)); forvar1163 = (forvar1163 + (1'h1)))
                begin
                  if ($unsigned(forvar1117[(3'h4):(2'h2)]))
                    begin
                      reg1164 <= $signed({{(reg926 << reg859)}});
                    end
                  else
                    begin
                      reg1164 <= (^($unsigned((~(8'hb0))) < (^(reg904 ~^ reg828))));
                      reg1165 <= (($unsigned($signed(forvar1019)) > forvar1052) ?
                          ({(reg949 || reg936)} <= (|$signed(reg1057))) : reg873[(1'h0):(1'h0)]);
                    end
                  for (forvar1166 = (1'h0); (forvar1166 < (1'h1)); forvar1166 = (forvar1166 + (1'h1)))
                    begin
                      reg1167 <= ((((-reg988) ?
                                  $signed(forvar733) : $unsigned(reg1108)) ?
                              {forvar845} : ((~&(8'ha9)) ?
                                  {reg1152} : (reg1027 >> reg1127))) ?
                          reg814[(1'h0):(1'h0)] : ($unsigned((reg1166 ?
                                  reg1125 : reg996)) ?
                              $signed(reg808[(4'hf):(3'h6)]) : $signed(reg902[(4'h8):(3'h5)])));
                    end
                end
              for (forvar1168 = (1'h0); (forvar1168 < (1'h1)); forvar1168 = (forvar1168 + (1'h1)))
                begin
                  for (forvar1169 = (1'h0); (forvar1169 < (1'h1)); forvar1169 = (forvar1169 + (1'h1)))
                    begin
                      reg1170 <= reg1132[(2'h2):(1'h1)];
                      reg1171 <= $unsigned(reg764[(3'h5):(3'h4)]);
                    end
                  for (forvar1172 = (1'h0); (forvar1172 < (1'h0)); forvar1172 = (forvar1172 + (1'h1)))
                    begin
                      reg1173 <= {{{((8'hb6) ? reg1064 : reg720)}}};
                      reg1174 <= $signed(($unsigned((forvar903 ?
                          reg1160 : forvar1153)) >> (|$unsigned(reg976))));
                    end
                end
              for (forvar1175 = (1'h0); (forvar1175 < (1'h1)); forvar1175 = (forvar1175 + (1'h1)))
                begin
                  if ($unsigned(reg1144))
                    begin
                      reg1176 <= $unsigned($signed(forvar1090));
                      reg1177 <= $unsigned((8'hb0));
                      reg1178 <= ((($unsigned(reg783) ?
                              $signed(forvar811) : (~^reg1083)) ?
                          reg914[(4'h9):(3'h4)] : reg767[(1'h0):(1'h0)]) && {forvar1000});
                    end
                  else
                    begin
                      reg1176 <= (~|((reg1174 ? reg1111 : $signed(forvar897)) ?
                          ((+reg912) ~^ $unsigned(reg770)) : (reg1071[(3'h4):(1'h0)] ~^ $unsigned(reg1102))));
                      reg1177 <= $signed((reg1053[(2'h2):(1'h0)] ?
                          $signed((!reg951)) : $signed((wire9 != (8'h9c)))));
                      reg1178 <= ((^{(-forvar884)}) ?
                          forvar1136 : (!forvar818[(1'h1):(1'h0)]));
                    end
                  for (forvar1179 = (1'h0); (forvar1179 < (2'h3)); forvar1179 = (forvar1179 + (1'h1)))
                    begin
                      reg1180 <= $signed($unsigned(({reg824} && reg853)));
                      reg1181 <= $signed(((reg742[(3'h4):(1'h0)] <= (reg746 < forvar998)) ?
                          reg827[(2'h3):(1'h1)] : $unsigned((forvar703 ?
                              forvar1038 : reg719))));
                      reg1182 <= reg1070[(4'hd):(4'hc)];
                    end
                end
              reg1183 <= $unsigned((reg1046 ^ ($signed((8'h9d)) ?
                  $unsigned(reg1155) : $unsigned(reg830))));
            end
        end
      for (forvar1184 = (1'h0); (forvar1184 < (2'h3)); forvar1184 = (forvar1184 + (1'h1)))
        begin
          reg1185 <= reg783;
          reg1186 <= $signed($unsigned($signed((reg1018 ?
              forvar1059 : (8'hb2)))));
          for (forvar1187 = (1'h0); (forvar1187 < (1'h1)); forvar1187 = (forvar1187 + (1'h1)))
            begin
              for (forvar1188 = (1'h0); (forvar1188 < (1'h1)); forvar1188 = (forvar1188 + (1'h1)))
                begin
                  for (forvar1189 = (1'h0); (forvar1189 < (1'h1)); forvar1189 = (forvar1189 + (1'h1)))
                    begin
                      reg1190 <= $signed($signed(reg1060));
                      reg1191 <= (-($signed((~reg1111)) ?
                          (~|reg1152) : reg1128));
                      reg1192 <= ($unsigned((|reg1063[(2'h3):(2'h2)])) ~^ forvar998);
                    end
                  reg1193 <= (~|$unsigned({(!reg709)}));
                end
              for (forvar1194 = (1'h0); (forvar1194 < (1'h0)); forvar1194 = (forvar1194 + (1'h1)))
                begin
                  reg1195 <= $signed({$signed({forvar1038})});
                  for (forvar1196 = (1'h0); (forvar1196 < (1'h1)); forvar1196 = (forvar1196 + (1'h1)))
                    begin
                      reg1197 <= (-forvar873[(4'h9):(4'h9)]);
                      reg1198 <= $signed((($signed(forvar723) ^ reg859) ?
                          ({forvar998} != $signed((8'hb6))) : ({forvar711} ?
                              reg1027[(2'h3):(2'h3)] : (^reg938))));
                    end
                end
            end
          if ($signed($signed($signed(forvar907[(2'h2):(2'h2)]))))
            begin
              if (($unsigned(reg1039) ?
                  ((~^(reg773 ? reg1101 : reg1078)) ?
                      $unsigned($unsigned(reg1142)) : $unsigned((~reg1107))) : {forvar1020}))
                begin
                  reg1199 <= reg1106;
                  for (forvar1200 = (1'h0); (forvar1200 < (1'h0)); forvar1200 = (forvar1200 + (1'h1)))
                    begin
                      reg1201 <= (reg717[(3'h4):(1'h1)] >= reg968);
                      reg1202 <= (8'h9d);
                    end
                  reg1203 <= $signed(((reg1060[(4'hd):(2'h3)] ^~ (reg874 ?
                          reg903 : reg733)) ?
                      ($signed(reg774) || (forvar1101 ?
                          forvar1011 : wire10)) : ($unsigned(forvar1130) || ((8'hb2) ?
                          (8'h9f) : forvar1057))));
                  if ((((!reg953) || (!forvar1163)) ^~ (((^reg1070) | reg1198) ?
                      (-$unsigned(reg931)) : $signed((reg707 ?
                          forvar1049 : reg1144)))))
                    begin
                      reg1204 <= (forvar1116[(3'h4):(3'h4)] + (!(reg828[(2'h3):(1'h1)] ?
                          forvar1162[(3'h6):(3'h4)] : reg1186[(4'hd):(1'h1)])));
                      reg1205 <= reg735[(4'hc):(1'h1)];
                      reg1206 <= ($signed(forvar725) - (((^reg883) ?
                              reg1082[(2'h3):(1'h0)] : $unsigned((8'ha7))) ?
                          $unsigned($unsigned(reg757)) : reg1070[(3'h4):(2'h3)]));
                    end
                  else
                    begin
                      reg1204 <= {$signed({$signed(reg767)})};
                      reg1205 <= reg952[(2'h2):(1'h0)];
                      reg1206 <= reg769[(1'h1):(1'h1)];
                      reg1207 <= forvar1099[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar1199 = (1'h0); (forvar1199 < (2'h3)); forvar1199 = (forvar1199 + (1'h1)))
                    begin
                      reg1200 <= reg1108[(1'h0):(1'h0)];
                      reg1201 <= $unsigned($signed($unsigned(reg712[(1'h1):(1'h0)])));
                    end
                end
              for (forvar1208 = (1'h0); (forvar1208 < (2'h2)); forvar1208 = (forvar1208 + (1'h1)))
                begin
                  if ({{$signed((~^reg1173))}})
                    begin
                      reg1209 <= (&reg1010[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg1209 <= forvar711;
                      reg1210 <= $unsigned((($signed((8'ha5)) ?
                          (~(8'h9c)) : (-reg1133)) > ($unsigned((8'ha0)) ?
                          forvar845[(4'h9):(2'h3)] : {forvar1004})));
                      reg1211 <= forvar844[(1'h0):(1'h0)];
                      reg1212 <= (reg1050 ?
                          $unsigned(((^~reg1029) >= ((8'ha1) ?
                              wire9 : reg1036))) : (!(&{reg1011})));
                    end
                  reg1213 <= (($unsigned((reg1162 ? reg957 : (8'hb1))) ?
                          reg1118 : (8'ha0)) ?
                      {((8'h9d) ?
                              reg1017[(4'h8):(3'h6)] : (reg758 * (8'hb6)))} : (($signed(reg1173) * (reg952 - reg1010)) ?
                          $unsigned(reg981) : reg911[(2'h2):(1'h1)]));
                  for (forvar1214 = (1'h0); (forvar1214 < (2'h3)); forvar1214 = (forvar1214 + (1'h1)))
                    begin
                      reg1215 <= reg741;
                      reg1216 <= $signed(forvar1032);
                      reg1217 <= (~$signed($unsigned((reg1000 >= forvar1208))));
                      reg1218 <= (^~(-($signed((8'haa)) << (forvar959 ?
                          reg886 : reg806))));
                    end
                  for (forvar1219 = (1'h0); (forvar1219 < (2'h3)); forvar1219 = (forvar1219 + (1'h1)))
                    begin
                      reg1220 <= $signed({$signed({reg871})});
                      reg1221 <= $signed(forvar1208[(3'h6):(2'h2)]);
                      reg1222 <= $signed(reg1202[(1'h0):(1'h0)]);
                    end
                end
              if ((~^reg805[(2'h3):(1'h1)]))
                begin
                  if (($unsigned({{reg1163}}) ?
                      ($signed({forvar989}) ?
                          forvar1114 : {$unsigned(reg819)}) : (~^((reg1220 ?
                          reg834 : forvar725) ~^ (&reg1018)))))
                    begin
                      reg1223 <= reg703;
                      reg1224 <= (reg706[(2'h3):(1'h1)] ?
                          (|(((8'ha0) >> reg1180) <= (reg849 || forvar1020))) : reg902[(3'h6):(2'h3)]);
                    end
                  else
                    begin
                      reg1223 <= (($unsigned(reg1181[(3'h6):(2'h3)]) ?
                          $signed((!reg875)) : $unsigned((reg976 <= reg989))) <= (^$signed($unsigned(reg1106))));
                    end
                  if ($signed(forvar1031[(4'h8):(2'h2)]))
                    begin
                      reg1225 <= (^~$unsigned($signed(forvar863)));
                      reg1226 <= (-(^$unsigned((reg917 ? reg1108 : (8'had)))));
                      reg1227 <= {({(|reg924)} > reg925[(2'h2):(2'h2)])};
                    end
                  else
                    begin
                      reg1225 <= $unsigned(forvar1011);
                      reg1226 <= $unsigned((reg908 ?
                          (|(~^forvar1118)) : $unsigned($signed(forvar1165))));
                    end
                end
              else
                begin
                  for (forvar1223 = (1'h0); (forvar1223 < (1'h0)); forvar1223 = (forvar1223 + (1'h1)))
                    begin
                      reg1224 <= forvar888;
                      reg1225 <= ((~&reg1161) == ($unsigned({reg1191}) ?
                          ((forvar724 ^ forvar1054) ?
                              reg940 : (reg729 ^ reg754)) : ((reg782 ?
                              (8'ha8) : reg923) | {reg889})));
                    end
                  for (forvar1226 = (1'h0); (forvar1226 < (2'h2)); forvar1226 = (forvar1226 + (1'h1)))
                    begin
                      reg1227 <= $signed(reg1078[(2'h2):(2'h2)]);
                      reg1228 <= (forvar1045 ^ reg752);
                      reg1229 <= reg774;
                      reg1230 <= $signed($unsigned((|(8'hb4))));
                    end
                end
              if (reg758[(2'h2):(1'h1)])
                begin
                  if (((&(reg830 ^~ (-forvar845))) ?
                      $signed(({reg987} - (reg785 ?
                          (8'hab) : forvar1116))) : (~(+reg1058))))
                    begin
                      reg1231 <= ((|{(forvar1223 ? reg1109 : reg906)}) ?
                          forvar1098 : reg1193[(4'h8):(4'h8)]);
                      reg1232 <= $unsigned(({reg1011} * $unsigned(reg741[(3'h5):(3'h4)])));
                      reg1233 <= reg887[(3'h5):(3'h4)];
                    end
                  else
                    begin
                      reg1231 <= (!forvar827[(2'h2):(2'h2)]);
                      reg1232 <= ($unsigned($signed($signed(reg1113))) - $signed(forvar812));
                      reg1233 <= forvar907;
                      reg1234 <= $signed(($unsigned(forvar1092) ?
                          ((forvar1125 >= reg1101) || {reg849}) : ((!forvar1074) <<< (reg779 > reg755))));
                    end
                  reg1235 <= (reg864[(1'h0):(1'h0)] ?
                      reg1161[(1'h0):(1'h0)] : (|{$unsigned(reg964)}));
                  for (forvar1236 = (1'h0); (forvar1236 < (2'h3)); forvar1236 = (forvar1236 + (1'h1)))
                    begin
                      reg1237 <= forvar818;
                      reg1238 <= {($unsigned($unsigned(reg1016)) << $signed($signed(reg857)))};
                      reg1239 <= $signed($unsigned(($unsigned(reg783) ?
                          forvar873[(1'h1):(1'h0)] : reg1207[(3'h4):(1'h0)])));
                    end
                end
              else
                begin
                  for (forvar1231 = (1'h0); (forvar1231 < (1'h0)); forvar1231 = (forvar1231 + (1'h1)))
                    begin
                      reg1232 <= (~(!$unsigned((8'h9c))));
                      reg1233 <= reg1076[(3'h5):(1'h1)];
                      reg1234 <= (!$unsigned(reg1093));
                    end
                  for (forvar1235 = (1'h0); (forvar1235 < (1'h1)); forvar1235 = (forvar1235 + (1'h1)))
                    begin
                      reg1236 <= (forvar1165 ?
                          (forvar1072 <= reg961[(4'ha):(1'h0)]) : (~&$unsigned((forvar932 ?
                              reg880 : reg1195))));
                      reg1237 <= (~&$unsigned({$signed((8'ha4))}));
                      reg1238 <= $signed((~&reg808[(1'h0):(1'h0)]));
                    end
                end
            end
          else
            begin
              reg1199 <= $signed(($unsigned((reg984 << reg1177)) ?
                  ((~&reg1227) <= $unsigned(reg1095)) : reg1001));
              if (reg946)
                begin
                  for (forvar1200 = (1'h0); (forvar1200 < (2'h3)); forvar1200 = (forvar1200 + (1'h1)))
                    begin
                      reg1201 <= reg949[(2'h2):(1'h1)];
                      reg1202 <= reg971[(3'h4):(1'h1)];
                    end
                end
              else
                begin
                  reg1200 <= reg1201[(2'h2):(2'h2)];
                  for (forvar1201 = (1'h0); (forvar1201 < (1'h0)); forvar1201 = (forvar1201 + (1'h1)))
                    begin
                      reg1202 <= ($signed((-$unsigned(reg1097))) ?
                          forvar738 : (((~reg817) || (&reg1003)) >= $unsigned((reg828 ?
                              reg901 : reg947))));
                      reg1203 <= (($signed($unsigned(reg977)) ?
                          forvar790[(1'h1):(1'h0)] : ($signed(forvar794) ^~ reg1079[(4'hc):(1'h0)])) <<< $unsigned(((forvar794 ?
                              forvar920 : reg1059) ?
                          reg755[(3'h6):(1'h0)] : (reg1015 >>> reg863))));
                    end
                  reg1204 <= (reg1045 ?
                      (reg705[(1'h0):(1'h0)] && ((8'hb2) ?
                          {forvar1099} : {wire10})) : $unsigned(reg832));
                  if ($unsigned(reg977))
                    begin
                      reg1205 <= (^~$unsigned($signed($unsigned((8'h9d)))));
                      reg1206 <= $signed($signed((~^forvar1153[(1'h1):(1'h0)])));
                    end
                  else
                    begin
                      reg1205 <= $unsigned(((~^(reg973 >>> forvar959)) + {((8'hba) < forvar825)}));
                    end
                end
            end
        end
      for (forvar1240 = (1'h0); (forvar1240 < (2'h3)); forvar1240 = (forvar1240 + (1'h1)))
        begin
          reg1241 <= (+$signed({$signed((8'hb9))}));
          if ($unsigned((|$signed(((8'ha9) ~^ reg850)))))
            begin
              if ({((reg921 ~^ reg1155) ?
                      $unsigned($signed((8'ha7))) : {reg770[(3'h6):(2'h2)]})})
                begin
                  for (forvar1242 = (1'h0); (forvar1242 < (1'h0)); forvar1242 = (forvar1242 + (1'h1)))
                    begin
                      reg1243 <= $unsigned(((~(reg975 ?
                          forvar840 : reg786)) << $signed(reg710[(3'h4):(2'h2)])));
                    end
                  reg1244 <= (&reg898);
                end
              else
                begin
                  for (forvar1242 = (1'h0); (forvar1242 < (1'h1)); forvar1242 = (forvar1242 + (1'h1)))
                    begin
                      reg1243 <= $unsigned(({(8'hb4)} ?
                          $signed(((8'ha7) ?
                              reg894 : forvar920)) : (reg733[(4'h9):(4'h9)] ?
                              (reg1132 + forvar1226) : ((8'ha6) <<< reg1089))));
                    end
                  reg1244 <= {$signed((^~(reg982 | reg997)))};
                end
              if ($signed((|({reg742} * forvar1147))))
                begin
                  if ((&((~^(reg832 >>> reg1041)) & (~|$signed(reg1053)))))
                    begin
                      reg1245 <= {(forvar1057 ?
                              forvar1100 : {$signed(reg1035)})};
                    end
                  else
                    begin
                      reg1245 <= reg1197[(4'ha):(1'h0)];
                      reg1246 <= reg709;
                      reg1247 <= $signed(reg782[(3'h4):(1'h1)]);
                    end
                  for (forvar1248 = (1'h0); (forvar1248 < (1'h0)); forvar1248 = (forvar1248 + (1'h1)))
                    begin
                      reg1249 <= (((reg1107 ?
                          ((8'ha3) ^~ reg1212) : $signed(forvar863)) <<< reg1015) == $unsigned($unsigned((^reg973))));
                      reg1250 <= $signed($unsigned(($unsigned(reg1079) ?
                          (forvar711 ?
                              forvar853 : reg834) : forvar838[(4'he):(4'hb)])));
                      reg1251 <= {{(!(|(8'haa)))}};
                      reg1252 <= $signed(((8'ha9) ?
                          $signed(reg987) : (|reg1193[(1'h1):(1'h1)])));
                    end
                  for (forvar1253 = (1'h0); (forvar1253 < (2'h3)); forvar1253 = (forvar1253 + (1'h1)))
                    begin
                      reg1254 <= $unsigned($unsigned(($signed(forvar890) ^~ {reg1046})));
                      reg1255 <= $unsigned($signed((forvar737 ?
                          reg1192 : reg764)));
                    end
                end
              else
                begin
                  for (forvar1245 = (1'h0); (forvar1245 < (1'h0)); forvar1245 = (forvar1245 + (1'h1)))
                    begin
                      reg1246 <= reg918;
                      reg1247 <= (-(reg1107 | $signed(reg923)));
                      reg1248 <= $signed($signed(wire11));
                    end
                  if ((reg1228[(2'h3):(2'h3)] ?
                      ($unsigned((forvar959 * (8'ha7))) ^~ forvar1113) : ({(reg971 >= forvar1175)} | ((+reg1215) ?
                          $signed(reg1134) : {(8'hb1)}))))
                    begin
                      reg1249 <= (8'haf);
                      reg1250 <= reg1000[(1'h0):(1'h0)];
                      reg1251 <= reg1230;
                    end
                  else
                    begin
                      reg1249 <= (~^($signed($signed(reg767)) ?
                          ((!forvar1099) + ((8'h9e) ?
                              (8'hab) : forvar763)) : (reg1156[(3'h5):(2'h3)] ?
                              (~^reg1003) : (forvar1090 ? (8'ha9) : (8'hb8)))));
                      reg1250 <= forvar1032;
                    end
                  reg1252 <= (~^forvar802);
                  for (forvar1253 = (1'h0); (forvar1253 < (1'h0)); forvar1253 = (forvar1253 + (1'h1)))
                    begin
                      reg1254 <= $unsigned((forvar1106 < ((reg1135 == reg852) ?
                          reg829 : $unsigned(reg943))));
                      reg1255 <= reg918[(3'h5):(3'h4)];
                    end
                end
            end
          else
            begin
              for (forvar1242 = (1'h0); (forvar1242 < (1'h1)); forvar1242 = (forvar1242 + (1'h1)))
                begin
                  reg1243 <= ((&$unsigned({reg1216})) ?
                      $signed((+(forvar1253 ?
                          forvar1109 : (8'hac)))) : ((((8'hb2) ?
                                  reg809 : reg865) ?
                              {forvar1072} : (forvar776 * (8'ha0))) ?
                          forvar1112 : (((8'hae) & reg897) < reg826[(4'he):(1'h0)])));
                  if ($signed($unsigned(((&(8'hb8)) < (reg1106 | reg1097)))))
                    begin
                      reg1244 <= (|{($unsigned(reg902) ?
                              reg856[(4'h9):(3'h4)] : forvar885)});
                      reg1245 <= ($signed($unsigned(reg786[(1'h0):(1'h0)])) >>> reg1145);
                      reg1246 <= $signed((~((forvar738 ~^ forvar1226) ?
                          reg1078 : $signed((8'ha9)))));
                      reg1247 <= $unsigned({$signed({forvar813})});
                    end
                  else
                    begin
                      reg1244 <= $signed($signed(reg1144));
                      reg1245 <= $signed(forvar711);
                      reg1246 <= $unsigned({forvar960[(1'h0):(1'h0)]});
                      reg1247 <= $signed(forvar949);
                    end
                end
              for (forvar1248 = (1'h0); (forvar1248 < (2'h3)); forvar1248 = (forvar1248 + (1'h1)))
                begin
                  reg1249 <= {($signed($unsigned((8'hb0))) ?
                          $signed(((8'had) ?
                              reg1068 : reg1018)) : reg847[(1'h0):(1'h0)])};
                  reg1250 <= (reg837[(2'h2):(1'h0)] ?
                      (~^{(forvar1242 ?
                              reg980 : reg774)}) : $signed((((8'hae) <= reg1062) == reg1220[(3'h4):(2'h2)])));
                  for (forvar1251 = (1'h0); (forvar1251 < (2'h3)); forvar1251 = (forvar1251 + (1'h1)))
                    begin
                      reg1252 <= {$unsigned($unsigned((reg849 ?
                              reg730 : reg830)))};
                      reg1253 <= $unsigned(({(forvar907 ?
                                  forvar1069 : reg1111)} ?
                          $unsigned($signed(forvar734)) : reg909[(3'h5):(1'h0)]));
                      reg1254 <= (((reg1248 == reg1165) ?
                              (forvar793 ?
                                  (reg854 ^ (8'hb7)) : (reg1075 ?
                                      forvar737 : (8'hb4))) : $signed({forvar776})) ?
                          $unsigned(((8'ha8) ?
                              $unsigned(forvar897) : {reg1157})) : (&reg1047[(2'h2):(2'h2)]));
                    end
                  if (forvar708[(3'h7):(1'h1)])
                    begin
                      reg1255 <= (reg881[(4'hd):(3'h4)] || reg966[(4'hb):(2'h3)]);
                      reg1256 <= {(reg950[(3'h5):(3'h5)] * $unsigned((^~reg1071)))};
                      reg1257 <= ((((reg1137 != forvar790) ?
                          (forvar984 ?
                              (8'hb5) : reg1062) : forvar1038[(3'h5):(1'h1)]) || reg1028) ^~ (8'hba));
                    end
                  else
                    begin
                      reg1255 <= (~|$unsigned(((&reg1167) || (reg1062 ?
                          reg1140 : forvar812))));
                      reg1256 <= ($signed(($signed(reg725) <<< (8'h9c))) << (!reg980[(1'h0):(1'h0)]));
                    end
                end
              if (reg1125)
                begin
                  for (forvar1258 = (1'h0); (forvar1258 < (1'h1)); forvar1258 = (forvar1258 + (1'h1)))
                    begin
                      reg1259 <= $signed((reg827 ?
                          $unsigned($unsigned(reg852)) : ((|reg910) ?
                              (8'hb5) : {forvar1149})));
                    end
                  reg1260 <= (forvar1069[(1'h0):(1'h0)] >>> (~^$unsigned((forvar825 ?
                      reg774 : (8'hb4)))));
                end
              else
                begin
                  if ((~&$signed((~|(~forvar1168)))))
                    begin
                      reg1258 <= ($signed(reg795) ?
                          $unsigned((^~reg963)) : (|((reg1025 && reg736) > {reg1112})));
                      reg1259 <= (~((reg1156 ?
                          reg1160 : $signed(reg946)) ~^ $unsigned(reg1079[(3'h6):(3'h4)])));
                      reg1260 <= ({(reg1114[(1'h1):(1'h1)] <= (~&reg1096))} ?
                          (~{reg714[(1'h1):(1'h0)]}) : $signed(reg806[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg1258 <= ((-$unsigned(reg898[(4'h8):(1'h0)])) ?
                          forvar1045[(2'h2):(2'h2)] : ($signed(forvar1169[(2'h3):(1'h0)]) ?
                              ((reg874 ? (8'hb4) : reg1022) ?
                                  ((8'hb0) <= reg1083) : reg1106) : (reg990[(2'h3):(2'h3)] & reg783)));
                    end
                end
            end
          if ((~^reg868))
            begin
              reg1261 <= $unsigned(forvar998);
              if (reg1053)
                begin
                  for (forvar1262 = (1'h0); (forvar1262 < (1'h0)); forvar1262 = (forvar1262 + (1'h1)))
                    begin
                      reg1263 <= $unsigned($signed($unsigned(reg733[(2'h3):(1'h0)])));
                      reg1264 <= forvar895[(3'h7):(3'h7)];
                    end
                end
              else
                begin
                  for (forvar1262 = (1'h0); (forvar1262 < (2'h2)); forvar1262 = (forvar1262 + (1'h1)))
                    begin
                      reg1263 <= $signed((^{$signed(reg861)}));
                      reg1264 <= {forvar922};
                    end
                end
            end
          else
            begin
              for (forvar1261 = (1'h0); (forvar1261 < (2'h2)); forvar1261 = (forvar1261 + (1'h1)))
                begin
                  if (reg1250[(4'he):(2'h2)])
                    begin
                      reg1262 <= {$unsigned(((~&forvar788) == forvar1258[(3'h4):(2'h2)]))};
                      reg1263 <= (reg1052[(4'hc):(3'h5)] ~^ ((~&reg936) ?
                          reg787[(1'h1):(1'h1)] : reg741));
                    end
                  else
                    begin
                      reg1262 <= reg942;
                      reg1263 <= reg704[(1'h0):(1'h0)];
                    end
                  for (forvar1264 = (1'h0); (forvar1264 < (2'h3)); forvar1264 = (forvar1264 + (1'h1)))
                    begin
                      reg1265 <= $unsigned($signed($signed($unsigned(forvar1067))));
                      reg1266 <= reg1051[(2'h3):(2'h3)];
                      reg1267 <= {$unsigned($signed($signed(forvar838)))};
                      reg1268 <= $signed(forvar1162[(3'h7):(1'h0)]);
                    end
                  for (forvar1269 = (1'h0); (forvar1269 < (1'h1)); forvar1269 = (forvar1269 + (1'h1)))
                    begin
                      reg1270 <= ($signed(((-reg887) ?
                              $signed(forvar1072) : $unsigned((8'ha4)))) ?
                          $signed(reg1057) : {reg1092});
                    end
                  for (forvar1271 = (1'h0); (forvar1271 < (1'h0)); forvar1271 = (forvar1271 + (1'h1)))
                    begin
                      reg1272 <= forvar1166[(2'h2):(1'h0)];
                      reg1273 <= (^reg805[(3'h5):(1'h0)]);
                    end
                end
              if (reg961[(3'h6):(2'h2)])
                begin
                  reg1274 <= reg980[(1'h1):(1'h1)];
                  for (forvar1275 = (1'h0); (forvar1275 < (2'h3)); forvar1275 = (forvar1275 + (1'h1)))
                    begin
                      reg1276 <= forvar932;
                      reg1277 <= (reg789 ?
                          $unsigned($unsigned((forvar1219 ?
                              reg1002 : (8'hb4)))) : reg1017[(2'h3):(1'h1)]);
                      reg1278 <= $signed((~^reg1178));
                    end
                  for (forvar1279 = (1'h0); (forvar1279 < (2'h3)); forvar1279 = (forvar1279 + (1'h1)))
                    begin
                      reg1280 <= ($unsigned($unsigned($signed(reg1167))) < {forvar899});
                      reg1281 <= $signed(forvar1011[(2'h3):(2'h3)]);
                      reg1282 <= ({(~|(reg1000 <<< forvar984))} ?
                          ($signed(reg984[(2'h2):(1'h0)]) ?
                              ((^forvar995) ?
                                  (forvar999 ?
                                      reg1259 : reg904) : {reg1226}) : forvar1062[(3'h5):(2'h3)]) : $unsigned(reg1180));
                    end
                end
              else
                begin
                  for (forvar1274 = (1'h0); (forvar1274 < (2'h2)); forvar1274 = (forvar1274 + (1'h1)))
                    begin
                      reg1275 <= (reg895 > $unsigned((^(forvar1223 ?
                          reg757 : forvar1214))));
                    end
                  if ((-(~|$unsigned($unsigned(reg989)))))
                    begin
                      reg1276 <= ($signed(((forvar1129 ~^ reg1185) == reg1275[(3'h7):(1'h0)])) ?
                          {$signed((^reg1100))} : (!{(|(8'hae))}));
                    end
                  else
                    begin
                      reg1276 <= forvar711[(2'h3):(1'h0)];
                      reg1277 <= $signed(forvar1019);
                    end
                  for (forvar1278 = (1'h0); (forvar1278 < (2'h3)); forvar1278 = (forvar1278 + (1'h1)))
                    begin
                      reg1279 <= $signed(($unsigned((reg1130 - reg1186)) ?
                          {$unsigned(reg765)} : $signed($unsigned(forvar963))));
                      reg1280 <= reg1157;
                      reg1281 <= $unsigned(forvar1274);
                    end
                  for (forvar1282 = (1'h0); (forvar1282 < (2'h3)); forvar1282 = (forvar1282 + (1'h1)))
                    begin
                      reg1283 <= $unsigned(forvar841[(4'hf):(4'hc)]);
                    end
                end
              reg1284 <= (~reg1250[(4'ha):(4'ha)]);
              for (forvar1285 = (1'h0); (forvar1285 < (2'h3)); forvar1285 = (forvar1285 + (1'h1)))
                begin
                  if (($signed(reg865[(2'h2):(1'h0)]) + reg836))
                    begin
                      reg1286 <= reg752;
                      reg1287 <= {$unsigned($signed($signed(forvar896)))};
                      reg1288 <= {({forvar867[(2'h2):(1'h1)]} < {reg883})};
                    end
                  else
                    begin
                      reg1286 <= reg875;
                      reg1287 <= {(-(~&(reg926 & (8'h9e))))};
                    end
                  for (forvar1289 = (1'h0); (forvar1289 < (2'h2)); forvar1289 = (forvar1289 + (1'h1)))
                    begin
                      reg1290 <= reg1207;
                      reg1291 <= ($signed(({(8'hb8)} ?
                          (~&reg1204) : (reg1277 ?
                              (8'hab) : reg938))) * $unsigned((+$signed((8'hb9)))));
                    end
                  for (forvar1292 = (1'h0); (forvar1292 < (1'h1)); forvar1292 = (forvar1292 + (1'h1)))
                    begin
                      reg1293 <= ({($signed(forvar768) ?
                                  (reg1199 ^ reg919) : reg1237)} ?
                          (reg1145[(2'h3):(2'h3)] ?
                              reg963[(4'h8):(4'h8)] : reg861[(1'h1):(1'h1)]) : $signed(reg960));
                    end
                end
            end
        end
    end
  assign wire1294 = wire8;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module15
#( parameter param700 = (!(~&(((8'ha4) ? (8'hb4) : (8'hb7)) ? ((8'hba) ? (8'had) : (8'hb7)) : ((8'h9d) << (8'ha2))))) )
(y, clk, wire20, wire19, wire18, wire17, wire16);
  output wire [(32'hbe0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire20;
  input wire signed [(5'h10):(1'h0)] wire19;
  input wire [(4'hc):(1'h0)] wire18;
  input wire signed [(3'h6):(1'h0)] wire17;
  input wire signed [(4'hf):(1'h0)] wire16;
  reg [(4'hd):(1'h0)] reg699 = (1'h0);
  reg [(5'h10):(1'h0)] reg698 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg697 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg696 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg695 = (1'h0);
  reg [(3'h5):(1'h0)] reg694 = (1'h0);
  reg [(4'hf):(1'h0)] reg693 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg692 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg691 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg690 = (1'h0);
  reg [(5'h10):(1'h0)] reg689 = (1'h0);
  reg [(2'h3):(1'h0)] forvar688 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg687 = (1'h0);
  reg [(4'h8):(1'h0)] forvar686 = (1'h0);
  reg [(3'h5):(1'h0)] forvar685 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg684 = (1'h0);
  reg [(5'h10):(1'h0)] reg683 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg682 = (1'h0);
  reg [(2'h3):(1'h0)] reg681 = (1'h0);
  reg [(4'hd):(1'h0)] forvar680 = (1'h0);
  reg [(4'hd):(1'h0)] reg679 = (1'h0);
  reg [(3'h4):(1'h0)] reg678 = (1'h0);
  reg [(4'he):(1'h0)] reg677 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg676 = (1'h0);
  reg [(2'h2):(1'h0)] reg675 = (1'h0);
  reg signed [(4'he):(1'h0)] reg674 = (1'h0);
  reg [(3'h7):(1'h0)] reg673 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg672 = (1'h0);
  reg [(5'h10):(1'h0)] forvar671 = (1'h0);
  reg [(3'h6):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar669 = (1'h0);
  reg [(4'hc):(1'h0)] reg662 = (1'h0);
  reg [(4'he):(1'h0)] forvar659 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg658 = (1'h0);
  reg [(4'hd):(1'h0)] forvar657 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar647 = (1'h0);
  reg [(4'h9):(1'h0)] forvar642 = (1'h0);
  reg [(4'he):(1'h0)] forvar650 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar649 = (1'h0);
  reg [(4'h9):(1'h0)] forvar645 = (1'h0);
  reg [(2'h2):(1'h0)] reg637 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg646 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg651 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar643 = (1'h0);
  reg [(3'h5):(1'h0)] forvar638 = (1'h0);
  reg [(4'hb):(1'h0)] reg668 = (1'h0);
  reg [(4'h8):(1'h0)] reg667 = (1'h0);
  reg [(2'h2):(1'h0)] reg666 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar665 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg664 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg663 = (1'h0);
  reg [(4'hd):(1'h0)] forvar662 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg661 = (1'h0);
  reg [(2'h3):(1'h0)] reg660 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg659 = (1'h0);
  reg [(4'h8):(1'h0)] forvar658 = (1'h0);
  reg [(4'hc):(1'h0)] reg657 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar656 = (1'h0);
  reg [(4'hd):(1'h0)] reg655 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg654 = (1'h0);
  reg [(5'h10):(1'h0)] reg653 = (1'h0);
  reg [(4'ha):(1'h0)] reg652 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar651 = (1'h0);
  reg [(4'hc):(1'h0)] reg650 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg649 = (1'h0);
  reg [(4'h9):(1'h0)] reg648 = (1'h0);
  reg [(4'h8):(1'h0)] reg647 = (1'h0);
  reg [(4'hf):(1'h0)] forvar646 = (1'h0);
  reg [(2'h2):(1'h0)] reg645 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg644 = (1'h0);
  reg [(4'hb):(1'h0)] reg643 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg642 = (1'h0);
  reg [(4'ha):(1'h0)] reg641 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg640 = (1'h0);
  reg [(2'h2):(1'h0)] reg639 = (1'h0);
  reg [(3'h6):(1'h0)] reg638 = (1'h0);
  reg [(4'ha):(1'h0)] forvar637 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg636 = (1'h0);
  reg [(4'hc):(1'h0)] reg635 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg634 = (1'h0);
  reg [(4'h8):(1'h0)] reg633 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg632 = (1'h0);
  reg [(3'h7):(1'h0)] reg631 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg630 = (1'h0);
  reg [(4'hf):(1'h0)] reg629 = (1'h0);
  reg [(3'h4):(1'h0)] reg628 = (1'h0);
  reg [(4'h9):(1'h0)] forvar627 = (1'h0);
  reg [(4'hd):(1'h0)] reg626 = (1'h0);
  reg [(4'hc):(1'h0)] reg625 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg624 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg623 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg622 = (1'h0);
  reg [(4'h9):(1'h0)] reg621 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg620 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg619 = (1'h0);
  reg [(4'ha):(1'h0)] forvar618 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar617 = (1'h0);
  reg [(4'hd):(1'h0)] reg616 = (1'h0);
  reg [(3'h5):(1'h0)] reg615 = (1'h0);
  reg [(4'hc):(1'h0)] reg614 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar613 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar612 = (1'h0);
  reg [(4'hd):(1'h0)] forvar611 = (1'h0);
  reg [(3'h7):(1'h0)] reg597 = (1'h0);
  reg [(5'h10):(1'h0)] reg598 = (1'h0);
  reg [(4'he):(1'h0)] reg610 = (1'h0);
  reg [(4'hd):(1'h0)] reg609 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg608 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg607 = (1'h0);
  reg [(4'h8):(1'h0)] forvar606 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg605 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg604 = (1'h0);
  reg [(4'h8):(1'h0)] forvar603 = (1'h0);
  reg [(4'hc):(1'h0)] reg602 = (1'h0);
  reg [(3'h7):(1'h0)] reg601 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg599 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar598 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar597 = (1'h0);
  reg [(3'h4):(1'h0)] reg596 = (1'h0);
  reg [(3'h7):(1'h0)] reg595 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg594 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg593 = (1'h0);
  reg [(4'ha):(1'h0)] reg592 = (1'h0);
  reg [(4'h8):(1'h0)] reg591 = (1'h0);
  reg [(5'h10):(1'h0)] reg590 = (1'h0);
  reg [(4'hb):(1'h0)] forvar589 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar588 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg587 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg586 = (1'h0);
  reg [(3'h7):(1'h0)] forvar585 = (1'h0);
  reg [(4'ha):(1'h0)] reg584 = (1'h0);
  reg [(4'hc):(1'h0)] reg583 = (1'h0);
  reg [(4'hd):(1'h0)] reg582 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar581 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg580 = (1'h0);
  reg [(3'h7):(1'h0)] reg579 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg578 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg577 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg576 = (1'h0);
  reg [(4'hb):(1'h0)] forvar575 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar574 = (1'h0);
  reg [(4'h8):(1'h0)] forvar573 = (1'h0);
  reg [(2'h2):(1'h0)] reg572 = (1'h0);
  reg [(4'hd):(1'h0)] forvar571 = (1'h0);
  reg [(4'h8):(1'h0)] forvar570 = (1'h0);
  reg [(2'h2):(1'h0)] reg569 = (1'h0);
  reg [(4'h8):(1'h0)] forvar549 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar539 = (1'h0);
  reg [(4'hf):(1'h0)] reg568 = (1'h0);
  reg [(4'hb):(1'h0)] reg567 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg566 = (1'h0);
  reg signed [(4'he):(1'h0)] reg565 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg564 = (1'h0);
  reg [(3'h7):(1'h0)] forvar563 = (1'h0);
  reg [(4'h8):(1'h0)] reg562 = (1'h0);
  reg [(4'hd):(1'h0)] reg561 = (1'h0);
  reg [(4'hd):(1'h0)] reg560 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg556 = (1'h0);
  reg [(4'hf):(1'h0)] reg552 = (1'h0);
  reg [(4'hd):(1'h0)] reg559 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg558 = (1'h0);
  reg [(3'h7):(1'h0)] reg557 = (1'h0);
  reg [(5'h10):(1'h0)] forvar556 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg555 = (1'h0);
  reg [(4'h9):(1'h0)] reg554 = (1'h0);
  reg signed [(4'he):(1'h0)] reg553 = (1'h0);
  reg [(4'hf):(1'h0)] forvar552 = (1'h0);
  reg [(4'hd):(1'h0)] reg551 = (1'h0);
  reg [(4'hd):(1'h0)] reg550 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg549 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar548 = (1'h0);
  reg [(4'hc):(1'h0)] reg540 = (1'h0);
  reg [(3'h6):(1'h0)] forvar538 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg534 = (1'h0);
  reg [(4'hf):(1'h0)] reg547 = (1'h0);
  reg [(4'h8):(1'h0)] reg546 = (1'h0);
  reg [(5'h10):(1'h0)] reg545 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg544 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg543 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg542 = (1'h0);
  reg [(2'h2):(1'h0)] reg541 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar540 = (1'h0);
  reg signed [(4'he):(1'h0)] reg539 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg538 = (1'h0);
  reg [(4'ha):(1'h0)] reg537 = (1'h0);
  reg [(3'h5):(1'h0)] reg536 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg535 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar534 = (1'h0);
  reg [(2'h2):(1'h0)] forvar533 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire532;
  wire signed [(4'he):(1'h0)] wire531;
  wire signed [(4'hb):(1'h0)] wire530;
  reg signed [(4'h8):(1'h0)] reg529 = (1'h0);
  reg [(4'h8):(1'h0)] reg528 = (1'h0);
  reg [(4'h8):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg526 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar525 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg524 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg523 = (1'h0);
  reg [(2'h3):(1'h0)] forvar522 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar521 = (1'h0);
  reg signed [(4'he):(1'h0)] reg520 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg519 = (1'h0);
  reg [(4'h8):(1'h0)] reg518 = (1'h0);
  reg signed [(4'he):(1'h0)] reg517 = (1'h0);
  reg [(2'h3):(1'h0)] reg516 = (1'h0);
  reg [(4'hc):(1'h0)] reg515 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar514 = (1'h0);
  reg [(4'he):(1'h0)] reg513 = (1'h0);
  reg [(4'hd):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg511 = (1'h0);
  reg [(3'h6):(1'h0)] reg510 = (1'h0);
  reg [(3'h7):(1'h0)] forvar509 = (1'h0);
  reg [(4'h8):(1'h0)] forvar508 = (1'h0);
  reg [(3'h7):(1'h0)] forvar507 = (1'h0);
  reg [(2'h2):(1'h0)] reg493 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar489 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg504 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar500 = (1'h0);
  reg [(4'hc):(1'h0)] reg496 = (1'h0);
  reg [(4'ha):(1'h0)] reg491 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg490 = (1'h0);
  reg [(3'h4):(1'h0)] reg506 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg505 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar504 = (1'h0);
  reg [(3'h4):(1'h0)] reg503 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg502 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar499 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg501 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg500 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg498 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg497 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar496 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg495 = (1'h0);
  reg [(3'h5):(1'h0)] reg494 = (1'h0);
  reg [(4'he):(1'h0)] forvar493 = (1'h0);
  reg [(3'h6):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar491 = (1'h0);
  reg [(2'h3):(1'h0)] forvar490 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg489 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg488 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg487 = (1'h0);
  reg [(4'hc):(1'h0)] reg486 = (1'h0);
  reg [(4'hf):(1'h0)] forvar485 = (1'h0);
  reg [(4'ha):(1'h0)] forvar484 = (1'h0);
  reg [(4'h9):(1'h0)] forvar483 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg482 = (1'h0);
  reg [(2'h3):(1'h0)] reg481 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg480 = (1'h0);
  reg [(4'h9):(1'h0)] forvar479 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg478 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg477 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg476 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg475 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar474 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg473 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg472 = (1'h0);
  reg [(4'hb):(1'h0)] reg471 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar469 = (1'h0);
  reg [(3'h5):(1'h0)] reg460 = (1'h0);
  reg [(4'hb):(1'h0)] forvar456 = (1'h0);
  reg [(3'h6):(1'h0)] forvar455 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar450 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar446 = (1'h0);
  reg [(4'h9):(1'h0)] reg443 = (1'h0);
  reg [(3'h7):(1'h0)] forvar442 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar440 = (1'h0);
  reg [(4'hc):(1'h0)] reg439 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg466 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg470 = (1'h0);
  reg signed [(4'he):(1'h0)] reg469 = (1'h0);
  reg [(4'hb):(1'h0)] reg468 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg467 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar466 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar465 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg464 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg453 = (1'h0);
  reg [(4'hc):(1'h0)] forvar451 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg448 = (1'h0);
  reg [(4'hd):(1'h0)] reg463 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg462 = (1'h0);
  reg signed [(4'he):(1'h0)] reg461 = (1'h0);
  reg [(3'h7):(1'h0)] forvar460 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg458 = (1'h0);
  reg [(2'h2):(1'h0)] reg457 = (1'h0);
  reg signed [(4'he):(1'h0)] reg456 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg454 = (1'h0);
  reg [(3'h4):(1'h0)] forvar453 = (1'h0);
  reg [(4'he):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg451 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg450 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg449 = (1'h0);
  reg [(2'h2):(1'h0)] forvar448 = (1'h0);
  reg [(4'hd):(1'h0)] reg447 = (1'h0);
  reg [(4'hc):(1'h0)] reg446 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg445 = (1'h0);
  reg [(5'h10):(1'h0)] forvar444 = (1'h0);
  reg [(3'h5):(1'h0)] forvar443 = (1'h0);
  reg [(4'he):(1'h0)] reg442 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg441 = (1'h0);
  reg [(3'h7):(1'h0)] reg440 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar439 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg438 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar437 = (1'h0);
  reg signed [(4'he):(1'h0)] reg436 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg435 = (1'h0);
  reg [(4'hf):(1'h0)] forvar434 = (1'h0);
  reg [(4'ha):(1'h0)] forvar433 = (1'h0);
  reg [(3'h6):(1'h0)] forvar432 = (1'h0);
  reg [(4'hf):(1'h0)] reg431 = (1'h0);
  wire [(4'hf):(1'h0)] wire430;
  wire signed [(3'h5):(1'h0)] wire429;
  wire signed [(2'h2):(1'h0)] wire186;
  wire [(3'h5):(1'h0)] wire22;
  wire [(4'hb):(1'h0)] wire21;
  wire [(4'he):(1'h0)] wire188;
  wire [(4'hc):(1'h0)] wire189;
  wire signed [(4'he):(1'h0)] wire427;
  assign y = {reg699,
                 reg698,
                 reg697,
                 reg696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 reg689,
                 forvar688,
                 reg687,
                 forvar686,
                 forvar685,
                 reg684,
                 reg683,
                 reg682,
                 reg681,
                 forvar680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 reg675,
                 reg674,
                 reg673,
                 reg672,
                 forvar671,
                 reg670,
                 forvar669,
                 reg662,
                 forvar659,
                 reg658,
                 forvar657,
                 forvar647,
                 forvar642,
                 forvar650,
                 forvar649,
                 forvar645,
                 reg637,
                 reg646,
                 reg651,
                 forvar643,
                 forvar638,
                 reg668,
                 reg667,
                 reg666,
                 forvar665,
                 reg664,
                 reg663,
                 forvar662,
                 reg661,
                 reg660,
                 reg659,
                 forvar658,
                 reg657,
                 forvar656,
                 reg655,
                 reg654,
                 reg653,
                 reg652,
                 forvar651,
                 reg650,
                 reg649,
                 reg648,
                 reg647,
                 forvar646,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg640,
                 reg639,
                 reg638,
                 forvar637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 forvar627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 reg619,
                 forvar618,
                 forvar617,
                 reg616,
                 reg615,
                 reg614,
                 forvar613,
                 forvar612,
                 forvar611,
                 reg597,
                 reg598,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 forvar606,
                 reg605,
                 reg604,
                 forvar603,
                 reg602,
                 reg601,
                 reg600,
                 reg599,
                 forvar598,
                 forvar597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 forvar589,
                 forvar588,
                 reg587,
                 reg586,
                 forvar585,
                 reg584,
                 reg583,
                 reg582,
                 forvar581,
                 reg580,
                 reg579,
                 reg578,
                 reg577,
                 reg576,
                 forvar575,
                 forvar574,
                 forvar573,
                 reg572,
                 forvar571,
                 forvar570,
                 reg569,
                 forvar549,
                 forvar539,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 reg564,
                 forvar563,
                 reg562,
                 reg561,
                 reg560,
                 reg556,
                 reg552,
                 reg559,
                 reg558,
                 reg557,
                 forvar556,
                 reg555,
                 reg554,
                 reg553,
                 forvar552,
                 reg551,
                 reg550,
                 reg549,
                 forvar548,
                 reg540,
                 forvar538,
                 reg534,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 reg543,
                 reg542,
                 reg541,
                 forvar540,
                 reg539,
                 reg538,
                 reg537,
                 reg536,
                 reg535,
                 forvar534,
                 forvar533,
                 wire532,
                 wire531,
                 wire530,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 forvar525,
                 reg524,
                 reg523,
                 forvar522,
                 forvar521,
                 reg520,
                 reg519,
                 reg518,
                 reg517,
                 reg516,
                 reg515,
                 forvar514,
                 reg513,
                 reg512,
                 reg511,
                 reg510,
                 forvar509,
                 forvar508,
                 forvar507,
                 reg493,
                 forvar489,
                 reg504,
                 forvar500,
                 reg496,
                 reg491,
                 reg490,
                 reg506,
                 reg505,
                 forvar504,
                 reg503,
                 reg502,
                 forvar499,
                 reg501,
                 reg500,
                 reg499,
                 reg498,
                 reg497,
                 forvar496,
                 reg495,
                 reg494,
                 forvar493,
                 reg492,
                 forvar491,
                 forvar490,
                 reg489,
                 reg488,
                 reg487,
                 reg486,
                 forvar485,
                 forvar484,
                 forvar483,
                 reg482,
                 reg481,
                 reg480,
                 forvar479,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 forvar474,
                 reg473,
                 reg472,
                 reg471,
                 forvar469,
                 reg460,
                 forvar456,
                 forvar455,
                 forvar450,
                 forvar446,
                 reg443,
                 forvar442,
                 forvar440,
                 reg439,
                 reg434,
                 reg466,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 forvar466,
                 forvar465,
                 reg464,
                 reg453,
                 forvar451,
                 reg448,
                 reg463,
                 reg462,
                 reg461,
                 forvar460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 forvar453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 forvar448,
                 reg447,
                 reg446,
                 reg445,
                 forvar444,
                 forvar443,
                 reg442,
                 reg441,
                 reg440,
                 forvar439,
                 reg438,
                 forvar437,
                 reg436,
                 reg435,
                 forvar434,
                 forvar433,
                 forvar432,
                 reg431,
                 wire430,
                 wire429,
                 wire186,
                 wire22,
                 wire21,
                 wire188,
                 wire189,
                 wire427,
                 (1'h0)};
  assign wire21 = ((!wire18) ?
                      {$unsigned(wire19)} : $signed($unsigned((wire16 ?
                          wire16 : wire16))));
  assign wire22 = (wire19 >> wire21[(4'hb):(4'h8)]);
  module23 modinst187 (wire186, clk, wire22, wire20, wire19, wire16, wire21);
  assign wire188 = ({wire21} ?
                       (|(wire20 ?
                           $signed(wire19) : (wire18 ?
                               wire19 : wire21))) : wire16);
  assign wire189 = ({{(wire16 * (8'hb5))}} & wire17);
  module190 modinst428 (wire427, clk, wire18, wire22, wire19, wire188, wire189);
  assign wire429 = ({{wire19}} ?
                       wire16 : (wire19[(2'h3):(2'h3)] ?
                           ($signed(wire18) >>> ((8'hb6) != wire19)) : {(wire20 ?
                                   wire188 : wire22)}));
  assign wire430 = $unsigned((((~^(8'ha9)) & (wire186 ?
                       wire20 : (8'hac))) || {$unsigned(wire21)}));
  always
    @(posedge clk) begin
      reg431 <= wire20;
      if (($signed(wire188) ?
          ((|wire189[(1'h0):(1'h0)]) ?
              $unsigned((~|wire188)) : $unsigned((^reg431))) : ($signed({wire430}) ?
              wire18[(3'h4):(1'h0)] : (+wire22[(2'h3):(2'h2)]))))
        begin
          for (forvar432 = (1'h0); (forvar432 < (1'h1)); forvar432 = (forvar432 + (1'h1)))
            begin
              for (forvar433 = (1'h0); (forvar433 < (2'h2)); forvar433 = (forvar433 + (1'h1)))
                begin
                  for (forvar434 = (1'h0); (forvar434 < (1'h1)); forvar434 = (forvar434 + (1'h1)))
                    begin
                      reg435 <= {(&$signed($unsigned(wire188)))};
                      reg436 <= wire16[(4'h8):(3'h4)];
                    end
                  for (forvar437 = (1'h0); (forvar437 < (1'h0)); forvar437 = (forvar437 + (1'h1)))
                    begin
                      reg438 <= (~|({reg431[(4'h8):(2'h2)]} + ((wire19 ?
                          forvar437 : (8'had)) >> forvar437[(4'h9):(3'h7)])));
                    end
                  for (forvar439 = (1'h0); (forvar439 < (2'h3)); forvar439 = (forvar439 + (1'h1)))
                    begin
                      reg440 <= {$unsigned({reg438})};
                      reg441 <= $signed({((wire189 | wire19) ?
                              $signed(forvar437) : (wire20 ?
                                  reg431 : (8'ha2)))});
                    end
                  reg442 <= $signed(((reg441[(4'h8):(4'h8)] ?
                      $unsigned((8'hab)) : wire16[(3'h6):(1'h0)]) - ((~|wire188) >> (forvar432 | wire16))));
                end
              for (forvar443 = (1'h0); (forvar443 < (1'h0)); forvar443 = (forvar443 + (1'h1)))
                begin
                  for (forvar444 = (1'h0); (forvar444 < (1'h0)); forvar444 = (forvar444 + (1'h1)))
                    begin
                      reg445 <= $signed((^~((wire188 ? forvar439 : wire20) ?
                          (wire430 <= wire427) : $signed(wire22))));
                      reg446 <= ($unsigned(((reg440 == forvar443) | (wire16 ?
                          wire19 : forvar433))) + wire20);
                      reg447 <= wire22;
                    end
                end
              if ((wire22[(2'h2):(2'h2)] == wire20))
                begin
                  for (forvar448 = (1'h0); (forvar448 < (2'h3)); forvar448 = (forvar448 + (1'h1)))
                    begin
                      reg449 <= ((wire430 + (forvar433[(3'h5):(1'h0)] ?
                              {reg435} : (reg445 ? forvar433 : wire427))) ?
                          (8'ha9) : reg436);
                      reg450 <= $unsigned(forvar437[(3'h4):(2'h3)]);
                      reg451 <= (reg431[(1'h1):(1'h1)] - (-reg440[(3'h5):(1'h1)]));
                      reg452 <= wire189[(2'h3):(2'h2)];
                    end
                  for (forvar453 = (1'h0); (forvar453 < (2'h2)); forvar453 = (forvar453 + (1'h1)))
                    begin
                      reg454 <= $unsigned(reg438[(3'h7):(1'h0)]);
                      reg455 <= (-{$unsigned(wire427)});
                    end
                  if ((^reg435[(1'h0):(1'h0)]))
                    begin
                      reg456 <= ($unsigned($unsigned($signed(forvar432))) ^~ $unsigned(((wire429 << reg440) ?
                          $signed(wire189) : (reg451 && reg435))));
                      reg457 <= (^~wire188);
                      reg458 <= (~|wire188);
                      reg459 <= $signed(reg452[(3'h7):(2'h3)]);
                    end
                  else
                    begin
                      reg456 <= $unsigned($unsigned($signed(((8'h9f) ~^ wire20))));
                      reg457 <= $signed((-$signed(wire189[(3'h6):(3'h5)])));
                    end
                  for (forvar460 = (1'h0); (forvar460 < (1'h0)); forvar460 = (forvar460 + (1'h1)))
                    begin
                      reg461 <= $signed($signed(($signed(forvar448) >= reg454[(3'h4):(2'h3)])));
                      reg462 <= reg452;
                      reg463 <= (8'ha9);
                    end
                end
              else
                begin
                  if ((((^wire427) ?
                          ($signed(reg452) ?
                              $signed(reg454) : $signed((8'hab))) : $unsigned($unsigned((8'ha0)))) ?
                      (wire18 ?
                          ($signed(reg436) ?
                              reg445[(2'h2):(1'h1)] : reg445[(3'h4):(3'h4)]) : (~^((8'hba) > reg442))) : $signed(($unsigned(reg440) ?
                          $signed(reg446) : $signed((8'hb0))))))
                    begin
                      reg448 <= ($signed($signed($unsigned(reg462))) ~^ (+(+(~|reg454))));
                      reg449 <= reg449[(3'h5):(1'h1)];
                    end
                  else
                    begin
                      reg448 <= $unsigned((|reg448[(4'ha):(3'h7)]));
                    end
                  reg450 <= (8'hac);
                  for (forvar451 = (1'h0); (forvar451 < (1'h0)); forvar451 = (forvar451 + (1'h1)))
                    begin
                      reg452 <= forvar453[(3'h4):(2'h2)];
                      reg453 <= wire189[(4'ha):(4'h9)];
                      reg454 <= {($unsigned(forvar443[(3'h5):(3'h4)]) ?
                              (~&reg451) : $signed((~|wire17)))};
                      reg455 <= (^(^{(~&reg442)}));
                    end
                  reg456 <= (^~($unsigned($signed(wire21)) ?
                      $signed((reg438 ? (8'ha9) : wire189)) : (|reg431)));
                end
            end
          reg464 <= (!$signed(wire20));
          for (forvar465 = (1'h0); (forvar465 < (2'h3)); forvar465 = (forvar465 + (1'h1)))
            begin
              if ((((reg449[(1'h0):(1'h0)] ?
                          reg436[(3'h6):(1'h1)] : (forvar439 ?
                              reg462 : reg454)) ?
                      $signed(reg438[(4'h8):(3'h4)]) : $signed($signed(reg453))) ?
                  $unsigned(({forvar448} ?
                      forvar437 : $unsigned(wire19))) : reg452))
                begin
                  for (forvar466 = (1'h0); (forvar466 < (1'h1)); forvar466 = (forvar466 + (1'h1)))
                    begin
                      reg467 <= (^wire189);
                      reg468 <= (|(&(^~((8'ha8) ? reg435 : reg449))));
                      reg469 <= reg447;
                      reg470 <= $unsigned($unsigned(reg464[(1'h1):(1'h1)]));
                    end
                end
              else
                begin
                  if ({$unsigned(((reg446 ^ (8'hae)) ?
                          (reg467 != reg431) : {reg470}))})
                    begin
                      reg466 <= $signed(((^wire20) >= (&(8'hb7))));
                      reg467 <= reg464[(1'h0):(1'h0)];
                      reg468 <= $signed((~&(reg453 ?
                          $unsigned(reg461) : $signed(reg456))));
                    end
                  else
                    begin
                      reg466 <= (wire186[(2'h2):(1'h0)] ?
                          reg431 : (~{(~^forvar451)}));
                      reg467 <= {$unsigned({$signed(wire19)})};
                    end
                end
            end
        end
      else
        begin
          for (forvar432 = (1'h0); (forvar432 < (2'h3)); forvar432 = (forvar432 + (1'h1)))
            begin
              for (forvar433 = (1'h0); (forvar433 < (2'h2)); forvar433 = (forvar433 + (1'h1)))
                begin
                  if ($signed((wire16[(2'h2):(1'h0)] ?
                      (reg442[(2'h2):(2'h2)] ?
                          (-(8'ha1)) : (~^forvar460)) : (-$signed(forvar448)))))
                    begin
                      reg434 <= $unsigned({(wire17[(3'h5):(2'h3)] ?
                              wire17 : {(8'hb9)})});
                      reg435 <= ($signed($unsigned(reg453)) ?
                          ($unsigned((-wire17)) ^ reg458) : (+$unsigned(reg468[(3'h7):(3'h6)])));
                      reg436 <= $unsigned(((((8'hba) ^ forvar466) | (forvar453 ?
                          wire188 : reg457)) ^ $unsigned($unsigned(wire17))));
                    end
                  else
                    begin
                      reg434 <= reg435[(3'h6):(2'h2)];
                      reg435 <= $unsigned(((^~$signed(wire21)) | (&((8'ha4) ^ wire189))));
                    end
                end
              for (forvar437 = (1'h0); (forvar437 < (2'h3)); forvar437 = (forvar437 + (1'h1)))
                begin
                  reg438 <= (reg440 ?
                      wire188 : ($unsigned((reg440 ?
                          forvar434 : forvar437)) >= (((8'h9c) == reg469) >> (forvar439 ?
                          wire18 : (8'hae)))));
                  reg439 <= reg470;
                  for (forvar440 = (1'h0); (forvar440 < (1'h1)); forvar440 = (forvar440 + (1'h1)))
                    begin
                      reg441 <= {wire427};
                    end
                  for (forvar442 = (1'h0); (forvar442 < (2'h2)); forvar442 = (forvar442 + (1'h1)))
                    begin
                      reg443 <= ($signed(($unsigned(forvar442) ?
                          (reg438 ?
                              reg462 : reg453) : (~|forvar448))) >>> reg453);
                    end
                end
              for (forvar444 = (1'h0); (forvar444 < (1'h1)); forvar444 = (forvar444 + (1'h1)))
                begin
                  if ($signed(forvar432[(1'h1):(1'h0)]))
                    begin
                      reg445 <= (-((8'hb0) <<< ((!reg443) ?
                          (reg450 != reg457) : reg451)));
                    end
                  else
                    begin
                      reg445 <= {$unsigned(($unsigned(wire430) ?
                              $unsigned(forvar465) : $signed(reg458)))};
                    end
                  for (forvar446 = (1'h0); (forvar446 < (1'h0)); forvar446 = (forvar446 + (1'h1)))
                    begin
                      reg447 <= (^~($unsigned(((8'hb4) == (8'hae))) ?
                          reg457 : reg462[(1'h1):(1'h1)]));
                    end
                  if (reg464)
                    begin
                      reg448 <= $unsigned((($signed(forvar437) ?
                              $signed(reg455) : forvar446) ?
                          reg451[(2'h3):(1'h1)] : reg453));
                    end
                  else
                    begin
                      reg448 <= (^~reg435[(2'h2):(2'h2)]);
                      reg449 <= (reg462[(2'h3):(1'h0)] ?
                          $signed(reg434[(3'h5):(2'h3)]) : {reg461});
                    end
                  for (forvar450 = (1'h0); (forvar450 < (1'h0)); forvar450 = (forvar450 + (1'h1)))
                    begin
                      reg451 <= $signed($unsigned($unsigned((reg464 >= forvar440))));
                      reg452 <= $unsigned($signed((8'ha4)));
                      reg453 <= reg451[(3'h5):(3'h4)];
                    end
                end
              reg454 <= forvar448;
            end
          for (forvar455 = (1'h0); (forvar455 < (1'h1)); forvar455 = (forvar455 + (1'h1)))
            begin
              for (forvar456 = (1'h0); (forvar456 < (1'h1)); forvar456 = (forvar456 + (1'h1)))
                begin
                  if ($unsigned((((forvar444 ? forvar450 : forvar433) ?
                      $unsigned(forvar439) : $unsigned(forvar437)) <<< $signed(forvar437[(3'h4):(3'h4)]))))
                    begin
                      reg457 <= {((&(wire186 ? reg434 : reg469)) || wire429)};
                    end
                  else
                    begin
                      reg457 <= ($signed($unsigned(wire186[(1'h0):(1'h0)])) ?
                          $signed(forvar466[(2'h2):(1'h1)]) : forvar432);
                      reg458 <= ((($signed((8'h9c)) * reg466) ?
                          ((forvar450 > reg449) ?
                              wire22 : {reg431}) : (+(8'h9c))) >>> ($unsigned(reg453[(3'h4):(2'h2)]) ?
                          ((&wire17) ^~ (forvar443 && reg434)) : reg466[(3'h6):(1'h0)]));
                      reg459 <= ((forvar456[(4'h8):(3'h7)] ?
                              $signed(reg436[(1'h0):(1'h0)]) : {$unsigned(forvar460)}) ?
                          (-(((8'h9f) ?
                              reg469 : reg440) > (reg456 > reg438))) : (reg464[(4'hb):(2'h3)] <<< {reg466[(4'hb):(2'h2)]}));
                      reg460 <= ($unsigned(reg468) >>> reg454[(3'h4):(2'h3)]);
                    end
                  if ((wire16 >> (^~$unsigned($signed(forvar446)))))
                    begin
                      reg461 <= forvar444;
                    end
                  else
                    begin
                      reg461 <= (reg457 != (({wire427} ?
                          $signed(reg454) : {forvar455}) || {$unsigned(reg448)}));
                    end
                  if (($signed($unsigned(reg442)) + $unsigned($signed((forvar466 ?
                      reg435 : reg453)))))
                    begin
                      reg462 <= ($signed((wire16 ?
                          forvar439 : (&reg457))) | ((reg450[(3'h5):(2'h3)] >>> (forvar448 & wire188)) + wire20));
                      reg463 <= ($signed((reg466 ?
                              (~|reg458) : ((8'h9d) ? forvar450 : reg464))) ?
                          (~$unsigned((~(8'h9c)))) : (~&(forvar437 ^~ (reg431 & forvar456))));
                      reg464 <= ($signed(((reg458 ?
                              forvar451 : forvar460) + forvar437[(4'hc):(4'h8)])) ?
                          ((!wire430[(3'h7):(3'h6)]) < ((!reg463) ?
                              $unsigned(wire16) : forvar434)) : {reg461});
                    end
                  else
                    begin
                      reg462 <= (~&{{wire429[(1'h0):(1'h0)]}});
                      reg463 <= $unsigned({$signed((wire188 <= forvar437))});
                      reg464 <= reg462;
                    end
                  for (forvar465 = (1'h0); (forvar465 < (1'h0)); forvar465 = (forvar465 + (1'h1)))
                    begin
                      reg466 <= reg448[(3'h4):(2'h2)];
                      reg467 <= $signed(reg455[(4'h9):(3'h5)]);
                      reg468 <= reg442[(4'hc):(4'ha)];
                    end
                end
              for (forvar469 = (1'h0); (forvar469 < (1'h0)); forvar469 = (forvar469 + (1'h1)))
                begin
                  if (reg462[(1'h0):(1'h0)])
                    begin
                      reg470 <= ((~|reg443) ?
                          (reg455 ?
                              reg463 : ((~&forvar451) | $unsigned(wire17))) : (~^$signed($signed(reg438))));
                      reg471 <= {{{(-wire188)}}};
                      reg472 <= (reg431[(4'hd):(3'h5)] >> reg451[(3'h5):(1'h0)]);
                    end
                  else
                    begin
                      reg470 <= $signed({$signed((reg470 ?
                              forvar437 : forvar442))});
                      reg471 <= wire429[(3'h4):(2'h3)];
                      reg472 <= (forvar439 ?
                          (^$signed((wire429 - reg463))) : forvar433[(3'h6):(1'h0)]);
                      reg473 <= wire21[(4'h8):(1'h0)];
                    end
                  for (forvar474 = (1'h0); (forvar474 < (2'h2)); forvar474 = (forvar474 + (1'h1)))
                    begin
                      reg475 <= (reg450 | forvar453);
                      reg476 <= ({(-$unsigned(forvar439))} ?
                          wire16 : (!((&reg445) ?
                              (reg468 < forvar469) : $unsigned(reg450))));
                    end
                  if ((^~((reg447 >= (reg459 ?
                      forvar474 : forvar456)) > reg453)))
                    begin
                      reg477 <= $unsigned($unsigned($signed({(8'ha6)})));
                      reg478 <= ({$signed(reg439)} ?
                          (^(8'hac)) : $signed((~|$signed(reg461))));
                    end
                  else
                    begin
                      reg477 <= reg467;
                    end
                  for (forvar479 = (1'h0); (forvar479 < (1'h0)); forvar479 = (forvar479 + (1'h1)))
                    begin
                      reg480 <= forvar469[(1'h1):(1'h0)];
                      reg481 <= $unsigned((forvar432[(1'h0):(1'h0)] <= reg436));
                      reg482 <= forvar443;
                    end
                end
            end
        end
      for (forvar483 = (1'h0); (forvar483 < (1'h0)); forvar483 = (forvar483 + (1'h1)))
        begin
          for (forvar484 = (1'h0); (forvar484 < (2'h3)); forvar484 = (forvar484 + (1'h1)))
            begin
              for (forvar485 = (1'h0); (forvar485 < (2'h3)); forvar485 = (forvar485 + (1'h1)))
                begin
                  if ((forvar460 ? reg454 : reg455[(3'h4):(1'h0)]))
                    begin
                      reg486 <= reg462;
                      reg487 <= (!(~(^{forvar432})));
                      reg488 <= $unsigned($unsigned(($signed(forvar443) ?
                          $signed(forvar466) : $unsigned(reg457))));
                    end
                  else
                    begin
                      reg486 <= (reg457[(1'h1):(1'h1)] ?
                          $unsigned($signed(wire18)) : $signed($unsigned((^forvar442))));
                    end
                end
            end
          if ({$signed((~^(reg460 - reg472)))})
            begin
              reg489 <= reg464;
              for (forvar490 = (1'h0); (forvar490 < (1'h1)); forvar490 = (forvar490 + (1'h1)))
                begin
                  for (forvar491 = (1'h0); (forvar491 < (2'h3)); forvar491 = (forvar491 + (1'h1)))
                    begin
                      reg492 <= reg478[(2'h2):(1'h1)];
                    end
                end
              for (forvar493 = (1'h0); (forvar493 < (2'h3)); forvar493 = (forvar493 + (1'h1)))
                begin
                  reg494 <= {forvar453[(1'h0):(1'h0)]};
                  reg495 <= reg453[(4'hb):(3'h7)];
                  for (forvar496 = (1'h0); (forvar496 < (1'h1)); forvar496 = (forvar496 + (1'h1)))
                    begin
                      reg497 <= ((8'ha7) ^ forvar450);
                      reg498 <= reg462;
                    end
                end
              if ({forvar446[(3'h4):(2'h3)]})
                begin
                  if ((wire427[(3'h5):(1'h0)] ?
                      $unsigned(((~|forvar456) ?
                          forvar442[(1'h0):(1'h0)] : reg461[(2'h2):(2'h2)])) : (~|reg461)))
                    begin
                      reg499 <= $unsigned(($unsigned(((8'haa) ?
                          reg460 : wire189)) > ((forvar465 * wire21) < reg438[(4'hb):(1'h1)])));
                      reg500 <= reg451[(2'h2):(1'h1)];
                      reg501 <= forvar446;
                    end
                  else
                    begin
                      reg499 <= reg497;
                      reg500 <= ((forvar453[(1'h1):(1'h0)] ?
                              forvar455 : {$unsigned(forvar493)}) ?
                          reg492[(2'h2):(2'h2)] : forvar432);
                      reg501 <= (8'haf);
                    end
                end
              else
                begin
                  for (forvar499 = (1'h0); (forvar499 < (2'h2)); forvar499 = (forvar499 + (1'h1)))
                    begin
                      reg500 <= reg469[(3'h7):(3'h4)];
                      reg501 <= ($signed($unsigned((reg436 ?
                              reg463 : wire16))) ?
                          ($signed($unsigned(wire16)) ?
                              reg455 : $unsigned($unsigned(reg462))) : (|((8'ha7) ?
                              (forvar490 ^ reg456) : forvar450)));
                      reg502 <= ($unsigned($signed({reg473})) || ((reg463[(3'h5):(1'h1)] ?
                          reg458 : $unsigned(wire430)) >>> $unsigned(forvar460[(1'h1):(1'h1)])));
                      reg503 <= $unsigned(((reg435 ?
                              (wire430 ?
                                  forvar484 : reg473) : reg478[(4'h8):(3'h4)]) ?
                          $unsigned(reg488) : (8'ha8)));
                    end
                  for (forvar504 = (1'h0); (forvar504 < (1'h1)); forvar504 = (forvar504 + (1'h1)))
                    begin
                      reg505 <= reg454[(3'h6):(2'h2)];
                      reg506 <= $signed({$unsigned({reg448})});
                    end
                end
            end
          else
            begin
              if ((forvar450[(2'h2):(2'h2)] ?
                  wire21 : ($unsigned($signed(wire16)) ?
                      $signed((8'hb5)) : ($signed(reg439) & $signed(reg471)))))
                begin
                  if ((forvar451[(4'h9):(2'h3)] < {((&(8'hb5)) & $unsigned(reg505))}))
                    begin
                      reg489 <= (($unsigned((~|wire186)) ?
                              ((|reg497) ?
                                  $unsigned(reg431) : wire189[(2'h2):(1'h1)]) : reg502) ?
                          reg489[(2'h3):(1'h0)] : (-$signed($signed(reg431))));
                      reg490 <= ({$unsigned((wire19 + reg499))} < (reg489 > reg452));
                      reg491 <= {$signed(reg443[(4'h9):(3'h4)])};
                      reg492 <= (wire427[(4'ha):(4'h9)] ?
                          $unsigned($unsigned(forvar474[(2'h3):(2'h3)])) : {forvar483});
                    end
                  else
                    begin
                      reg489 <= ({forvar450} ?
                          reg451[(4'ha):(2'h2)] : (~^(8'ha4)));
                      reg490 <= reg469[(2'h2):(1'h0)];
                      reg491 <= ((!forvar453) >= wire19[(3'h7):(3'h7)]);
                      reg492 <= reg446[(4'h9):(3'h5)];
                    end
                  for (forvar493 = (1'h0); (forvar493 < (2'h2)); forvar493 = (forvar493 + (1'h1)))
                    begin
                      reg494 <= (forvar484[(3'h4):(1'h1)] << ((((8'h9c) ?
                              forvar451 : (8'hb9)) ~^ (8'ha9)) ?
                          $signed((forvar493 ?
                              forvar451 : reg438)) : $signed({(8'hb7)})));
                      reg495 <= (reg435 != $unsigned($unsigned((forvar443 ?
                          reg438 : forvar446))));
                    end
                  if ($signed(wire20))
                    begin
                      reg496 <= {$signed(((~^reg489) ?
                              (+(8'hba)) : reg498[(4'h8):(3'h4)]))};
                      reg497 <= reg502;
                      reg498 <= reg503[(2'h2):(1'h1)];
                      reg499 <= $signed(reg466);
                    end
                  else
                    begin
                      reg496 <= $unsigned(reg468);
                      reg497 <= reg457[(1'h0):(1'h0)];
                      reg498 <= (8'h9f);
                      reg499 <= {reg446[(3'h4):(1'h0)]};
                    end
                  for (forvar500 = (1'h0); (forvar500 < (2'h2)); forvar500 = (forvar500 + (1'h1)))
                    begin
                      reg501 <= $unsigned((8'ha5));
                      reg502 <= (&{$unsigned((~&reg502))});
                      reg503 <= $signed({(8'hba)});
                      reg504 <= ($signed({(forvar434 <= forvar450)}) | wire429);
                    end
                end
              else
                begin
                  for (forvar489 = (1'h0); (forvar489 < (2'h2)); forvar489 = (forvar489 + (1'h1)))
                    begin
                      reg490 <= forvar434[(4'h9):(3'h6)];
                      reg491 <= reg441;
                      reg492 <= ((~|(reg454[(2'h2):(1'h1)] ?
                          reg481[(1'h1):(1'h0)] : $signed(reg488))) == forvar448[(1'h0):(1'h0)]);
                    end
                  if (reg431[(1'h0):(1'h0)])
                    begin
                      reg493 <= (($signed((~reg463)) >> ((wire16 ?
                              forvar456 : reg489) || (8'hb0))) ?
                          (8'hae) : reg453);
                      reg494 <= $unsigned((~$signed($unsigned(reg495))));
                    end
                  else
                    begin
                      reg493 <= reg431[(3'h5):(3'h5)];
                      reg494 <= {$unsigned(($unsigned(reg442) >>> forvar499))};
                      reg495 <= $signed($unsigned($signed((reg489 >= wire17))));
                    end
                end
            end
          for (forvar507 = (1'h0); (forvar507 < (1'h0)); forvar507 = (forvar507 + (1'h1)))
            begin
              for (forvar508 = (1'h0); (forvar508 < (1'h1)); forvar508 = (forvar508 + (1'h1)))
                begin
                  for (forvar509 = (1'h0); (forvar509 < (1'h1)); forvar509 = (forvar509 + (1'h1)))
                    begin
                      reg510 <= ((~^{$unsigned((8'haf))}) ?
                          (((reg454 || reg457) * forvar443) - reg470) : ((^(reg461 ?
                                  reg472 : reg494)) ?
                              $signed((reg434 ?
                                  reg463 : reg454)) : forvar455[(1'h0):(1'h0)]));
                      reg511 <= (^~reg497);
                      reg512 <= wire22;
                      reg513 <= forvar456[(3'h4):(1'h1)];
                    end
                  for (forvar514 = (1'h0); (forvar514 < (1'h1)); forvar514 = (forvar514 + (1'h1)))
                    begin
                      reg515 <= reg503[(3'h4):(1'h0)];
                      reg516 <= {reg494};
                    end
                  reg517 <= (~&($unsigned($signed(forvar448)) ?
                      ($unsigned(reg477) < (reg472 || forvar448)) : reg480));
                  if (((wire18 <<< {(reg434 >>> forvar489)}) <= wire189[(4'ha):(1'h0)]))
                    begin
                      reg518 <= $signed((8'hb4));
                    end
                  else
                    begin
                      reg518 <= (&reg489[(2'h3):(1'h0)]);
                      reg519 <= forvar500;
                      reg520 <= {$signed(($unsigned(reg494) | (~forvar443)))};
                    end
                end
              for (forvar521 = (1'h0); (forvar521 < (1'h0)); forvar521 = (forvar521 + (1'h1)))
                begin
                  for (forvar522 = (1'h0); (forvar522 < (1'h0)); forvar522 = (forvar522 + (1'h1)))
                    begin
                      reg523 <= (+$signed((reg459[(1'h1):(1'h1)] ?
                          reg515[(3'h6):(3'h5)] : reg466)));
                    end
                  if ({((forvar437 ? $unsigned(wire186) : {forvar521}) ?
                          ({forvar466} == $signed(wire189)) : $signed($signed(reg517)))})
                    begin
                      reg524 <= (reg513[(4'h8):(3'h5)] < $signed(forvar514));
                    end
                  else
                    begin
                      reg524 <= (({(reg494 < (8'ha3))} ?
                          $signed($signed(forvar437)) : ((reg480 ?
                              reg495 : (8'hb5)) ^~ (&(8'hb4)))) || reg500[(4'hf):(3'h7)]);
                    end
                  for (forvar525 = (1'h0); (forvar525 < (2'h2)); forvar525 = (forvar525 + (1'h1)))
                    begin
                      reg526 <= (^(+$unsigned($unsigned(reg505))));
                      reg527 <= $signed($signed(reg467[(3'h5):(2'h3)]));
                      reg528 <= ((|reg515) ~^ forvar493);
                      reg529 <= $signed((!reg528));
                    end
                end
            end
        end
    end
  assign wire530 = ($unsigned(((forvar446 ?
                       reg520 : forvar444) >>> reg477[(4'ha):(1'h1)])) > $unsigned(reg439[(4'h9):(1'h1)]));
  assign wire531 = (^~forvar525[(1'h1):(1'h1)]);
  assign wire532 = (~^(^($signed(reg524) && {(8'h9f)})));
  always
    @(posedge clk) begin
      for (forvar533 = (1'h0); (forvar533 < (1'h1)); forvar533 = (forvar533 + (1'h1)))
        begin
          if ($unsigned(reg460))
            begin
              if (reg487[(3'h5):(3'h5)])
                begin
                  for (forvar534 = (1'h0); (forvar534 < (1'h0)); forvar534 = (forvar534 + (1'h1)))
                    begin
                      reg535 <= (reg448 ?
                          reg526[(2'h2):(2'h2)] : $signed($unsigned((^reg527))));
                      reg536 <= (8'ha7);
                      reg537 <= forvar439;
                      reg538 <= {forvar433};
                    end
                  reg539 <= reg535;
                  for (forvar540 = (1'h0); (forvar540 < (1'h0)); forvar540 = (forvar540 + (1'h1)))
                    begin
                      reg541 <= (((8'ha7) ?
                          $signed($unsigned(forvar484)) : $signed((~wire19))) && ((^(reg526 ?
                              reg538 : reg487)) ?
                          (~(reg468 ?
                              reg449 : forvar437)) : reg537[(4'ha):(1'h0)]));
                      reg542 <= $unsigned((+(reg478 >>> $unsigned(reg438))));
                      reg543 <= {$unsigned(((forvar443 - reg454) > ((8'haf) * reg486)))};
                      reg544 <= ($signed(((reg516 ? reg520 : reg462) ?
                              $unsigned((8'hb4)) : forvar499)) ?
                          (({forvar451} ? (&reg449) : wire17[(2'h2):(2'h2)]) ?
                              {$unsigned(wire17)} : (reg515 * reg436)) : $signed(forvar455[(2'h3):(2'h2)]));
                    end
                  if (((8'h9c) ?
                      wire17 : (forvar493[(2'h3):(2'h3)] ?
                          (~$signed(wire22)) : (~|(+forvar490)))))
                    begin
                      reg545 <= ({{(reg538 ? forvar440 : reg475)}} ?
                          ((~|(reg535 && reg476)) ?
                              (((8'had) ~^ reg495) ?
                                  wire429 : $signed(forvar469)) : $signed($unsigned((8'ha0)))) : reg441[(4'h9):(1'h1)]);
                    end
                  else
                    begin
                      reg545 <= (reg502 & (((~&(8'h9c)) ?
                          {reg487} : {forvar446}) << reg523));
                      reg546 <= forvar446;
                      reg547 <= (((-$signed((8'ha1))) << $signed((&reg546))) ?
                          (forvar491[(3'h4):(1'h1)] ?
                              $signed((reg493 ?
                                  wire530 : forvar460)) : reg498) : ((reg524 ?
                                  reg515[(3'h4):(2'h2)] : forvar490[(2'h2):(1'h1)]) ?
                              $unsigned((reg518 ?
                                  forvar465 : reg443)) : ((reg452 ?
                                  forvar451 : reg468) < (^~reg517))));
                    end
                end
              else
                begin
                  if ((!(({wire21} ? reg492 : {wire21}) ?
                      reg455[(4'ha):(3'h5)] : reg440)))
                    begin
                      reg534 <= $signed($signed({$unsigned(reg448)}));
                      reg535 <= (^~(8'hae));
                    end
                  else
                    begin
                      reg534 <= {((wire532 ?
                              reg528 : {reg453}) >= $signed(forvar499[(3'h5):(1'h1)]))};
                      reg535 <= ((8'h9d) >>> $signed({$signed(reg524)}));
                      reg536 <= forvar493[(4'hd):(4'ha)];
                      reg537 <= ((|reg471) ^ (((forvar540 != reg547) <<< forvar432) && reg441));
                    end
                  for (forvar538 = (1'h0); (forvar538 < (2'h3)); forvar538 = (forvar538 + (1'h1)))
                    begin
                      reg539 <= (((reg489[(3'h5):(1'h1)] ?
                          (~^forvar460) : (reg500 ?
                              wire430 : reg495)) == forvar455[(1'h0):(1'h0)]) ^ $signed(wire427));
                      reg540 <= forvar474[(3'h7):(3'h6)];
                      reg541 <= reg506;
                      reg542 <= $unsigned(((~&(reg510 << reg463)) << {forvar479}));
                    end
                end
              if (((8'haa) <<< forvar444[(3'h4):(2'h2)]))
                begin
                  for (forvar548 = (1'h0); (forvar548 < (2'h3)); forvar548 = (forvar548 + (1'h1)))
                    begin
                      reg549 <= $signed(reg445);
                      reg550 <= reg431[(4'hf):(3'h7)];
                      reg551 <= ((reg482 < $signed((~reg500))) ?
                          ((reg494[(2'h2):(1'h1)] ?
                              reg491 : (-forvar507)) >> wire21[(2'h3):(1'h1)]) : ($signed(forvar440) ?
                              reg510[(2'h3):(1'h0)] : forvar439));
                    end
                  for (forvar552 = (1'h0); (forvar552 < (2'h2)); forvar552 = (forvar552 + (1'h1)))
                    begin
                      reg553 <= ($unsigned((~^(8'h9d))) ?
                          (|$unsigned($unsigned(reg523))) : $unsigned(((-wire19) < reg517[(4'he):(1'h1)])));
                      reg554 <= ($unsigned(($signed(forvar439) != (reg480 <<< reg448))) + (forvar509 ?
                          reg480[(3'h4):(2'h3)] : {(8'hb0)}));
                      reg555 <= reg528[(3'h7):(3'h4)];
                    end
                  for (forvar556 = (1'h0); (forvar556 < (2'h2)); forvar556 = (forvar556 + (1'h1)))
                    begin
                      reg557 <= $unsigned((~&reg501[(2'h2):(2'h2)]));
                    end
                  if ((8'hb3))
                    begin
                      reg558 <= reg490[(2'h2):(2'h2)];
                      reg559 <= ($signed((reg450 != (reg497 << (8'ha3)))) ?
                          {(~^(~forvar453))} : ($signed(reg517[(4'hb):(3'h7)]) ?
                              $unsigned((forvar451 < forvar444)) : reg446));
                    end
                  else
                    begin
                      reg558 <= $unsigned(reg505);
                    end
                end
              else
                begin
                  for (forvar548 = (1'h0); (forvar548 < (1'h1)); forvar548 = (forvar548 + (1'h1)))
                    begin
                      reg549 <= (^(8'hb7));
                    end
                  reg550 <= (&(^~$signed($unsigned(reg471))));
                  if (((~$signed($unsigned((8'hb9)))) & $signed(reg469)))
                    begin
                      reg551 <= $unsigned($signed(((reg466 >= forvar522) ?
                          $signed((8'h9d)) : {forvar465})));
                      reg552 <= reg528[(3'h4):(1'h1)];
                    end
                  else
                    begin
                      reg551 <= reg463[(3'h6):(3'h4)];
                      reg552 <= (~wire16);
                      reg553 <= ($signed(((~|(8'ha2)) & (^~reg453))) ?
                          $unsigned($signed($unsigned(reg558))) : {$signed(wire430)});
                    end
                  if (({((+(8'hb6)) ? {forvar440} : (forvar474 || (8'hb9)))} ?
                      ($signed(reg453) ~^ (|(8'hba))) : $signed(forvar552)))
                    begin
                      reg554 <= (($signed(reg526) <<< reg540) ?
                          wire20[(4'hb):(3'h4)] : (~$signed(wire530)));
                      reg555 <= $signed((+(^(|reg466))));
                      reg556 <= (~|$signed(wire188));
                      reg557 <= ($unsigned(((reg482 ? forvar548 : wire189) ?
                              $signed(reg440) : (!wire19))) ?
                          ((8'ha2) <= $unsigned((~reg462))) : $signed($unsigned((8'hab))));
                    end
                  else
                    begin
                      reg554 <= (~|$unsigned(((&reg488) <= $unsigned(reg456))));
                      reg555 <= $signed($signed($signed((wire17 ?
                          forvar552 : (8'hae)))));
                      reg556 <= reg536[(3'h4):(2'h3)];
                      reg557 <= $unsigned({{reg506}});
                    end
                end
              if (((((reg459 ? wire532 : reg478) ~^ (+forvar432)) ?
                  $unsigned((reg438 ?
                      wire531 : reg534)) : $signed((+forvar509))) == reg490))
                begin
                  reg560 <= (((+(~^forvar493)) > (~forvar433)) != (((8'ha7) >> {reg536}) ?
                      $unsigned(forvar469[(1'h1):(1'h0)]) : {$unsigned(reg477)}));
                end
              else
                begin
                  if ({reg440})
                    begin
                      reg560 <= $signed((-(|forvar456)));
                      reg561 <= $signed($signed(((^~reg487) ?
                          forvar442 : (!reg466))));
                      reg562 <= {reg442[(1'h1):(1'h0)]};
                    end
                  else
                    begin
                      reg560 <= $signed(((((8'haa) > reg472) > (8'hb0)) < forvar552[(4'hd):(4'ha)]));
                      reg561 <= $unsigned((~|{wire531}));
                      reg562 <= (($unsigned(reg497[(2'h2):(1'h0)]) != (forvar504[(1'h0):(1'h0)] ?
                              $unsigned(forvar434) : (wire188 ?
                                  reg467 : reg528))) ?
                          $signed(reg446) : (forvar556[(4'he):(4'h9)] == (^reg436[(4'hc):(3'h5)])));
                    end
                  for (forvar563 = (1'h0); (forvar563 < (1'h1)); forvar563 = (forvar563 + (1'h1)))
                    begin
                      reg564 <= forvar521;
                      reg565 <= (reg494[(2'h2):(2'h2)] >> reg543[(2'h2):(2'h2)]);
                      reg566 <= {reg565[(4'ha):(2'h2)]};
                      reg567 <= $signed(($unsigned((reg511 <= (8'hb6))) ^~ ((reg454 - reg490) ?
                          (reg513 == reg554) : $signed(wire531))));
                    end
                end
              reg568 <= {(((reg480 ? forvar548 : forvar491) ?
                      reg544 : (reg551 ?
                          (8'hb2) : forvar489)) != {(|(8'h9e))})};
            end
          else
            begin
              if (forvar525[(1'h1):(1'h0)])
                begin
                  for (forvar534 = (1'h0); (forvar534 < (1'h0)); forvar534 = (forvar534 + (1'h1)))
                    begin
                      reg535 <= $signed($signed(reg540[(1'h1):(1'h1)]));
                      reg536 <= (^reg567[(2'h2):(2'h2)]);
                      reg537 <= $signed(reg545[(3'h5):(3'h5)]);
                      reg538 <= (|$unsigned($unsigned((-(8'hb0)))));
                    end
                  for (forvar539 = (1'h0); (forvar539 < (2'h2)); forvar539 = (forvar539 + (1'h1)))
                    begin
                      reg540 <= $signed(forvar522);
                      reg541 <= forvar499;
                      reg542 <= (reg492 ?
                          reg450[(1'h1):(1'h1)] : {reg565[(4'hc):(3'h5)]});
                      reg543 <= ($signed((~&reg512[(4'ha):(3'h7)])) - ($signed(reg539[(2'h3):(1'h0)]) == (reg454 ?
                          reg516 : $signed((8'hb2)))));
                    end
                  if ({$signed(forvar443)})
                    begin
                      reg544 <= $signed(reg566[(3'h4):(2'h2)]);
                      reg545 <= $signed(reg440);
                      reg546 <= (8'haa);
                      reg547 <= (reg438[(2'h3):(2'h2)] ?
                          $signed(reg472) : forvar522[(2'h2):(2'h2)]);
                    end
                  else
                    begin
                      reg544 <= (forvar443[(1'h1):(1'h0)] ?
                          {({reg446} ?
                                  reg447 : (reg471 ?
                                      reg431 : reg517))} : (($signed(reg496) ^~ reg519[(3'h5):(3'h4)]) - ((wire18 > reg503) && reg469)));
                      reg545 <= {(~|(^(8'haf)))};
                      reg546 <= forvar490;
                      reg547 <= reg489;
                    end
                end
              else
                begin
                  for (forvar534 = (1'h0); (forvar534 < (2'h2)); forvar534 = (forvar534 + (1'h1)))
                    begin
                      reg535 <= wire22[(2'h3):(2'h3)];
                      reg536 <= ((({(8'h9c)} ?
                              $signed(forvar493) : $unsigned(reg445)) ?
                          $signed({reg436}) : (!(~&forvar496))) >> {{((8'ha1) ?
                                  forvar432 : wire429)}});
                    end
                end
              for (forvar548 = (1'h0); (forvar548 < (1'h1)); forvar548 = (forvar548 + (1'h1)))
                begin
                  for (forvar549 = (1'h0); (forvar549 < (1'h0)); forvar549 = (forvar549 + (1'h1)))
                    begin
                      reg550 <= reg535[(3'h4):(1'h1)];
                    end
                  reg551 <= {$unsigned($signed(reg436[(3'h4):(3'h4)]))};
                  for (forvar552 = (1'h0); (forvar552 < (1'h0)); forvar552 = (forvar552 + (1'h1)))
                    begin
                      reg553 <= (forvar507[(3'h4):(2'h3)] ^ forvar538);
                      reg554 <= ($signed(($signed(wire21) ?
                              forvar440[(3'h5):(2'h3)] : (~forvar533))) ?
                          $unsigned((8'hb8)) : (8'haa));
                      reg555 <= (^((~|(reg543 ?
                          (8'hae) : forvar443)) > reg560));
                    end
                end
            end
          reg569 <= $unsigned((((~wire18) ?
                  $unsigned(reg566) : $unsigned(reg489)) ?
              ($unsigned(reg524) ?
                  forvar465 : (reg493 >= (8'hac))) : reg475[(3'h4):(1'h1)]));
        end
      for (forvar570 = (1'h0); (forvar570 < (1'h1)); forvar570 = (forvar570 + (1'h1)))
        begin
          for (forvar571 = (1'h0); (forvar571 < (1'h0)); forvar571 = (forvar571 + (1'h1)))
            begin
              reg572 <= $unsigned({$signed(reg469[(4'hd):(3'h4)])});
            end
          for (forvar573 = (1'h0); (forvar573 < (2'h3)); forvar573 = (forvar573 + (1'h1)))
            begin
              for (forvar574 = (1'h0); (forvar574 < (1'h1)); forvar574 = (forvar574 + (1'h1)))
                begin
                  for (forvar575 = (1'h0); (forvar575 < (2'h3)); forvar575 = (forvar575 + (1'h1)))
                    begin
                      reg576 <= $signed($signed($unsigned($signed(reg455))));
                      reg577 <= (^($unsigned((&reg435)) >= reg481));
                      reg578 <= wire18;
                      reg579 <= $signed(reg578);
                    end
                  reg580 <= $signed(((~|$signed((8'hb9))) ?
                      ({forvar434} == ((8'ha7) <= reg497)) : {reg454[(3'h4):(1'h1)]}));
                  for (forvar581 = (1'h0); (forvar581 < (2'h3)); forvar581 = (forvar581 + (1'h1)))
                    begin
                      reg582 <= {$unsigned($signed($unsigned(reg495)))};
                      reg583 <= $signed($signed(forvar507));
                      reg584 <= $unsigned({reg440[(2'h3):(2'h3)]});
                    end
                  for (forvar585 = (1'h0); (forvar585 < (1'h0)); forvar585 = (forvar585 + (1'h1)))
                    begin
                      reg586 <= (({(reg463 ? wire531 : reg490)} ?
                              $signed((forvar474 ?
                                  forvar440 : forvar432)) : ($unsigned(reg535) >> {wire427})) ?
                          (^forvar514) : (~^reg494));
                      reg587 <= ((~((reg457 ?
                              forvar508 : reg467) > (wire531 <= reg562))) ?
                          (({reg447} || (forvar509 << forvar460)) ?
                              $signed(reg541) : ((^~forvar508) ?
                                  reg455[(1'h0):(1'h0)] : {reg434})) : $signed(reg482[(1'h1):(1'h0)]));
                    end
                end
              for (forvar588 = (1'h0); (forvar588 < (1'h1)); forvar588 = (forvar588 + (1'h1)))
                begin
                  for (forvar589 = (1'h0); (forvar589 < (1'h0)); forvar589 = (forvar589 + (1'h1)))
                    begin
                      reg590 <= {$signed((8'h9f))};
                      reg591 <= ((8'h9c) ? reg580 : (+$signed((~|reg586))));
                    end
                  if (reg496)
                    begin
                      reg592 <= (8'ha8);
                      reg593 <= forvar489[(1'h0):(1'h0)];
                      reg594 <= (reg495 ?
                          (!forvar514[(4'ha):(3'h5)]) : wire530[(4'h8):(4'h8)]);
                      reg595 <= $signed((8'hb6));
                    end
                  else
                    begin
                      reg592 <= (((&(~forvar448)) ?
                              ((reg538 ? forvar509 : reg440) ?
                                  $unsigned(reg446) : ((8'hb0) != reg592)) : {forvar581}) ?
                          reg513[(1'h1):(1'h1)] : $signed((^reg582[(4'hc):(4'h9)])));
                      reg593 <= {$unsigned(reg577[(2'h2):(1'h1)])};
                      reg594 <= forvar575[(3'h7):(3'h6)];
                      reg595 <= {$signed(reg480[(2'h2):(1'h1)])};
                    end
                end
            end
          if ($signed(reg546[(3'h5):(1'h0)]))
            begin
              reg596 <= reg516[(1'h0):(1'h0)];
              for (forvar597 = (1'h0); (forvar597 < (2'h3)); forvar597 = (forvar597 + (1'h1)))
                begin
                  for (forvar598 = (1'h0); (forvar598 < (1'h1)); forvar598 = (forvar598 + (1'h1)))
                    begin
                      reg599 <= {$unsigned((!(~&reg579)))};
                      reg600 <= reg590[(2'h3):(1'h0)];
                      reg601 <= (~|(~&$signed((forvar451 ? reg540 : reg431))));
                      reg602 <= $unsigned(($unsigned($signed(forvar442)) <= reg587));
                    end
                  for (forvar603 = (1'h0); (forvar603 < (2'h3)); forvar603 = (forvar603 + (1'h1)))
                    begin
                      reg604 <= $unsigned(($unsigned($unsigned(reg580)) & reg451[(4'h9):(1'h0)]));
                      reg605 <= (!(((+(8'had)) <<< reg449) ?
                          forvar444 : (~^$unsigned(reg540))));
                    end
                  for (forvar606 = (1'h0); (forvar606 < (1'h0)); forvar606 = (forvar606 + (1'h1)))
                    begin
                      reg607 <= ($unsigned(reg566[(2'h3):(1'h1)]) ?
                          (&$signed((reg565 ?
                              reg487 : reg550))) : ($unsigned($signed(reg517)) * forvar521));
                      reg608 <= (((forvar490 ?
                          $signed(reg524) : reg488[(2'h2):(1'h0)]) ^ (+(^~reg503))) || reg564);
                      reg609 <= $signed(forvar522);
                      reg610 <= (forvar439[(4'ha):(1'h1)] ?
                          ((8'ha5) * reg454) : (wire427 ?
                              reg445 : $signed((!(8'ha2)))));
                    end
                end
            end
          else
            begin
              reg596 <= ((8'had) ?
                  ((((8'hb1) ? wire189 : (8'hb2)) ?
                      (!wire530) : $signed((8'hb2))) | ((forvar585 ?
                          reg438 : forvar588) ?
                      reg448[(4'h8):(3'h4)] : $signed(reg527))) : (((reg590 ?
                          forvar585 : reg593) ?
                      (reg605 ?
                          reg552 : wire16) : reg516[(2'h2):(1'h1)]) || (+{reg439})));
              if ($signed(reg524[(3'h5):(2'h2)]))
                begin
                  for (forvar597 = (1'h0); (forvar597 < (1'h0)); forvar597 = (forvar597 + (1'h1)))
                    begin
                      reg598 <= ($unsigned(((~|(8'hb0)) ?
                              {reg557} : {reg511})) ?
                          $signed(((wire21 ~^ reg538) <= $unsigned(reg517))) : ((reg491[(3'h7):(2'h2)] ?
                                  (^~(8'ha6)) : forvar597) ?
                              (|(~^(8'ha0))) : reg579));
                      reg599 <= ((~$signed((reg535 && forvar446))) ?
                          $unsigned(reg541[(2'h2):(2'h2)]) : (reg435 > ((^~reg466) ?
                              (~^forvar508) : (reg557 ? (8'hb5) : reg591))));
                      reg600 <= ($unsigned($unsigned((-forvar465))) <= $unsigned($unsigned($signed(forvar508))));
                    end
                end
              else
                begin
                  if ($unsigned(($signed($signed(reg487)) ?
                      reg535[(4'hb):(3'h4)] : $unsigned((reg584 ?
                          reg551 : (8'hb7))))))
                    begin
                      reg597 <= (~^(-((forvar521 * reg431) ~^ (forvar474 >= reg523))));
                      reg598 <= $unsigned((reg461 + (reg473 ?
                          $unsigned(forvar437) : forvar585[(3'h7):(2'h2)])));
                    end
                  else
                    begin
                      reg597 <= reg469[(1'h0):(1'h0)];
                      reg598 <= (forvar460[(3'h6):(3'h5)] ?
                          {reg595[(3'h4):(2'h3)]} : $unsigned(($signed(reg534) ?
                              (^reg555) : forvar606)));
                      reg599 <= (^~$signed({$unsigned(reg467)}));
                    end
                end
            end
          for (forvar611 = (1'h0); (forvar611 < (1'h1)); forvar611 = (forvar611 + (1'h1)))
            begin
              for (forvar612 = (1'h0); (forvar612 < (1'h0)); forvar612 = (forvar612 + (1'h1)))
                begin
                  for (forvar613 = (1'h0); (forvar613 < (2'h2)); forvar613 = (forvar613 + (1'h1)))
                    begin
                      reg614 <= (~^forvar437[(2'h2):(1'h0)]);
                      reg615 <= reg567;
                      reg616 <= ((forvar611 >> (8'hb9)) ?
                          (|reg607[(3'h6):(2'h3)]) : reg584[(2'h2):(2'h2)]);
                    end
                end
              for (forvar617 = (1'h0); (forvar617 < (2'h3)); forvar617 = (forvar617 + (1'h1)))
                begin
                  for (forvar618 = (1'h0); (forvar618 < (2'h3)); forvar618 = (forvar618 + (1'h1)))
                    begin
                      reg619 <= reg584[(4'h9):(3'h5)];
                      reg620 <= $unsigned(reg542[(1'h1):(1'h1)]);
                      reg621 <= ($unsigned(reg550) ?
                          reg552 : $unsigned($signed((forvar549 ?
                              reg519 : reg452))));
                    end
                  if ($signed($unsigned((&reg561))))
                    begin
                      reg622 <= ($signed((~$unsigned((8'ha8)))) != (($signed(reg457) ?
                              (wire427 - reg604) : $unsigned((8'ha5))) ?
                          ((reg599 << wire532) ?
                              reg457[(1'h0):(1'h0)] : {reg490}) : reg597));
                      reg623 <= ({(8'hb4)} ?
                          ($signed((forvar606 >= reg499)) ?
                              reg596[(1'h0):(1'h0)] : $signed($unsigned(reg461))) : $unsigned($unsigned(reg610[(2'h3):(1'h1)])));
                      reg624 <= reg562;
                      reg625 <= forvar453;
                    end
                  else
                    begin
                      reg622 <= ((reg578 ?
                          $unsigned((^reg500)) : $unsigned((!wire189))) >>> $signed(forvar573));
                      reg623 <= reg557[(2'h2):(2'h2)];
                      reg624 <= {(reg490 ?
                              (&(reg461 + reg503)) : ((reg556 ?
                                      reg576 : reg482) ?
                                  $signed(forvar489) : wire21[(1'h0):(1'h0)]))};
                      reg625 <= (({(reg553 || forvar570)} <= (^~(reg535 ?
                              forvar589 : reg609))) ?
                          reg602 : (wire186[(2'h2):(2'h2)] * {(reg554 << reg496)}));
                    end
                  reg626 <= $unsigned($signed($unsigned(wire429)));
                end
              for (forvar627 = (1'h0); (forvar627 < (1'h1)); forvar627 = (forvar627 + (1'h1)))
                begin
                  if ((reg501 - $signed(reg528)))
                    begin
                      reg628 <= (reg569 & forvar456[(3'h6):(2'h2)]);
                    end
                  else
                    begin
                      reg628 <= $unsigned($unsigned(((wire188 <<< forvar612) + (~&reg477))));
                      reg629 <= ({reg468[(3'h5):(3'h5)]} < forvar440[(3'h7):(3'h6)]);
                      reg630 <= ((^(~&$signed(reg481))) > reg516);
                      reg631 <= {((-forvar499[(4'ha):(3'h6)]) != {forvar466})};
                    end
                  if ((reg610 & (($signed(reg559) ?
                      (~^reg596) : (reg454 ? reg608 : reg557)) >>> ({(8'ha4)} ?
                      reg501[(3'h5):(2'h3)] : forvar485[(3'h7):(1'h1)]))))
                    begin
                      reg632 <= reg454[(4'h8):(3'h6)];
                      reg633 <= $signed({forvar598[(3'h4):(2'h3)]});
                      reg634 <= reg549[(2'h2):(2'h2)];
                      reg635 <= {reg451[(4'hb):(3'h6)]};
                    end
                  else
                    begin
                      reg632 <= {(-$signed(reg486))};
                      reg633 <= {(~&reg536)};
                      reg634 <= forvar433[(3'h5):(2'h3)];
                    end
                  reg636 <= forvar627;
                end
            end
        end
      if (($unsigned(($unsigned((8'h9e)) ?
              (forvar489 ? wire22 : forvar443) : forvar466)) ?
          reg492[(2'h3):(1'h0)] : (((&reg619) ?
                  $signed(reg555) : (forvar442 ~^ (8'h9e))) ?
              {(reg569 ? (8'ha3) : reg456)} : $unsigned($signed((8'ha6))))))
        begin
          if (forvar589)
            begin
              for (forvar637 = (1'h0); (forvar637 < (1'h0)); forvar637 = (forvar637 + (1'h1)))
                begin
                  reg638 <= ($unsigned((reg534 << reg549[(2'h3):(2'h3)])) >> (reg513[(2'h2):(2'h2)] <= {$signed(reg569)}));
                  if (reg616)
                    begin
                      reg639 <= ((({reg506} ^ (^~reg599)) ?
                              reg566 : forvar453[(3'h4):(2'h3)]) ?
                          ((~$unsigned(reg555)) - reg456[(2'h3):(1'h0)]) : ($unsigned((~|reg469)) ^~ reg471[(4'hb):(3'h7)]));
                    end
                  else
                    begin
                      reg639 <= $unsigned({((~|reg604) * (!forvar479))});
                      reg640 <= ($unsigned(forvar606[(4'h8):(1'h0)]) < forvar581);
                      reg641 <= $signed(reg538[(2'h3):(1'h0)]);
                    end
                  if ((8'hb3))
                    begin
                      reg642 <= (!((((8'ha3) ? forvar485 : reg471) ?
                              (8'hab) : $signed((8'hb1))) ?
                          (8'hb4) : (8'hb4)));
                      reg643 <= $signed((+reg553));
                    end
                  else
                    begin
                      reg642 <= $unsigned($signed(reg538));
                      reg643 <= forvar493[(3'h7):(3'h7)];
                      reg644 <= {($signed(reg539[(4'hb):(4'hb)]) ?
                              ($unsigned(reg519) ?
                                  {reg635} : (forvar563 ?
                                      forvar499 : reg481)) : $signed($unsigned(reg551)))};
                      reg645 <= (!$unsigned($signed($signed(forvar479))));
                    end
                  for (forvar646 = (1'h0); (forvar646 < (2'h2)); forvar646 = (forvar646 + (1'h1)))
                    begin
                      reg647 <= ((((8'ha7) ~^ $unsigned(reg536)) ?
                          forvar522[(1'h1):(1'h1)] : ((wire17 ?
                                  reg493 : reg607) ?
                              (forvar443 ?
                                  reg626 : reg469) : $unsigned(forvar573))) - $unsigned(((forvar618 ^~ reg475) ?
                          (reg599 ? reg602 : reg481) : (forvar646 ?
                              (8'hab) : reg620))));
                      reg648 <= $unsigned($unsigned(reg439));
                      reg649 <= $signed(reg545[(4'hc):(4'h9)]);
                      reg650 <= (~|$unsigned(reg599));
                    end
                end
              for (forvar651 = (1'h0); (forvar651 < (1'h0)); forvar651 = (forvar651 + (1'h1)))
                begin
                  if (wire188[(4'h8):(3'h5)])
                    begin
                      reg652 <= $signed(forvar484[(1'h1):(1'h1)]);
                      reg653 <= (reg504[(4'hd):(4'ha)] - {forvar490});
                    end
                  else
                    begin
                      reg652 <= ($unsigned(($signed(forvar651) ?
                          (^~wire429) : reg462)) + $signed({(~^reg462)}));
                      reg653 <= $unsigned($unsigned((8'hb6)));
                      reg654 <= ((+(forvar613[(4'h9):(4'h9)] ?
                          (^reg551) : $unsigned(reg524))) * $unsigned(((forvar507 ?
                              forvar465 : reg601) ?
                          reg576 : (^forvar563))));
                      reg655 <= $signed(($unsigned($unsigned(forvar646)) & forvar627[(3'h7):(3'h6)]));
                    end
                end
              for (forvar656 = (1'h0); (forvar656 < (2'h2)); forvar656 = (forvar656 + (1'h1)))
                begin
                  reg657 <= (~^$signed(reg494));
                  for (forvar658 = (1'h0); (forvar658 < (1'h0)); forvar658 = (forvar658 + (1'h1)))
                    begin
                      reg659 <= reg644[(4'h8):(3'h4)];
                      reg660 <= {$signed(forvar606[(3'h5):(2'h3)])};
                      reg661 <= wire429;
                    end
                  for (forvar662 = (1'h0); (forvar662 < (2'h3)); forvar662 = (forvar662 + (1'h1)))
                    begin
                      reg663 <= {((~|(reg536 > (8'ha6))) ?
                              (reg537[(1'h0):(1'h0)] ?
                                  {reg501} : ((8'h9f) ?
                                      reg463 : reg545)) : forvar611)};
                      reg664 <= ((8'hb7) < $unsigned(reg614[(4'hc):(4'hc)]));
                    end
                  for (forvar665 = (1'h0); (forvar665 < (1'h0)); forvar665 = (forvar665 + (1'h1)))
                    begin
                      reg666 <= $signed((8'hb8));
                      reg667 <= reg564[(2'h2):(1'h0)];
                      reg668 <= ((~(~|reg622[(1'h1):(1'h1)])) ?
                          (~forvar603) : ($unsigned({reg605}) + {forvar499[(4'hc):(4'hb)]}));
                    end
                end
            end
          else
            begin
              for (forvar637 = (1'h0); (forvar637 < (1'h1)); forvar637 = (forvar637 + (1'h1)))
                begin
                  for (forvar638 = (1'h0); (forvar638 < (2'h2)); forvar638 = (forvar638 + (1'h1)))
                    begin
                      reg639 <= $unsigned((({reg560} >>> $unsigned((8'hb9))) ?
                          (wire430 ?
                              reg562[(3'h5):(3'h4)] : reg590[(1'h0):(1'h0)]) : {(reg495 > (8'hba))}));
                      reg640 <= forvar455;
                      reg641 <= wire20;
                      reg642 <= forvar439[(1'h1):(1'h1)];
                    end
                end
              if (($unsigned((reg664 ?
                  (reg550 ? (8'hb8) : forvar440) : (^~forvar575))) - reg602))
                begin
                  for (forvar643 = (1'h0); (forvar643 < (2'h2)); forvar643 = (forvar643 + (1'h1)))
                    begin
                      reg644 <= reg538;
                      reg645 <= ($unsigned({(reg488 ?
                              forvar556 : reg619)}) ^ $signed($signed((forvar432 ?
                          reg668 : wire18))));
                    end
                  for (forvar646 = (1'h0); (forvar646 < (2'h2)); forvar646 = (forvar646 + (1'h1)))
                    begin
                      reg647 <= $unsigned(reg621);
                      reg648 <= $unsigned($unsigned(((forvar585 <= reg448) ?
                          $unsigned((8'haa)) : $signed((8'hb2)))));
                    end
                  if ($unsigned($signed((reg431[(4'h9):(3'h5)] ?
                      $unsigned(wire188) : $signed(forvar574)))))
                    begin
                      reg649 <= $unsigned({$signed(reg626[(3'h4):(2'h3)])});
                      reg650 <= ((reg636 ?
                          (reg504 & (reg493 + reg577)) : reg564) - reg517);
                    end
                  else
                    begin
                      reg649 <= (((((8'ha5) == forvar465) >> reg478[(4'h8):(3'h4)]) | {((8'hb1) >>> (8'ha6))}) ?
                          ({forvar440} ^~ $signed(forvar479)) : reg482);
                      reg650 <= reg480;
                      reg651 <= $unsigned((+(reg517[(2'h3):(1'h1)] ?
                          reg511 : reg583)));
                    end
                end
              else
                begin
                  if (forvar466[(2'h2):(1'h0)])
                    begin
                      reg643 <= $unsigned(reg555);
                      reg644 <= (^$unsigned(reg449[(3'h6):(3'h5)]));
                    end
                  else
                    begin
                      reg643 <= {reg489};
                      reg644 <= (~($unsigned((reg553 ?
                          forvar521 : (8'hab))) << ($unsigned((8'hb4)) ?
                          (forvar442 ? forvar549 : reg449) : reg544)));
                      reg645 <= reg510[(2'h3):(1'h0)];
                    end
                  reg646 <= reg500[(4'hd):(4'hd)];
                end
            end
        end
      else
        begin
          if ($signed(((~&(reg567 != reg641)) - {{reg478}})))
            begin
              if (forvar443)
                begin
                  if (({($signed((8'hb3)) ?
                          (|reg561) : $unsigned(reg648))} <<< forvar442))
                    begin
                      reg637 <= (reg624 ?
                          reg451 : {((reg499 && reg464) - (reg519 == reg567))});
                      reg638 <= $signed($unsigned((reg503[(2'h2):(2'h2)] <<< forvar491[(1'h0):(1'h0)])));
                      reg639 <= $unsigned(($unsigned($unsigned(forvar575)) + reg526));
                    end
                  else
                    begin
                      reg637 <= reg547[(1'h1):(1'h1)];
                    end
                  if (forvar469)
                    begin
                      reg640 <= (+reg668);
                      reg641 <= $signed((wire17[(1'h1):(1'h0)] ?
                          ($signed(reg653) ?
                              (~&reg576) : $signed(reg470)) : $signed(reg604)));
                      reg642 <= ({(((8'haf) ? reg647 : (8'hae)) ?
                              reg504[(4'ha):(2'h2)] : (reg577 ?
                                  forvar455 : reg601))} - (reg640[(3'h5):(3'h4)] ?
                          reg436[(3'h5):(3'h4)] : ((reg541 * reg654) ?
                              {reg583} : forvar643)));
                    end
                  else
                    begin
                      reg640 <= (8'hb7);
                      reg641 <= (((^$unsigned(reg623)) ?
                          reg605 : (^$unsigned(reg601))) == forvar651[(2'h2):(1'h1)]);
                      reg642 <= $signed(reg539[(4'he):(4'h9)]);
                    end
                end
              else
                begin
                  if ($unsigned(($unsigned((forvar479 ? wire21 : reg620)) ?
                      ((8'ha2) ^ reg556[(2'h2):(2'h2)]) : (8'hb1))))
                    begin
                      reg637 <= reg448;
                      reg638 <= (reg492[(2'h3):(1'h0)] ?
                          reg558[(2'h2):(1'h0)] : (~|reg583));
                      reg639 <= $signed((~|reg604));
                      reg640 <= $signed(reg460);
                    end
                  else
                    begin
                      reg637 <= forvar490[(2'h3):(1'h1)];
                    end
                end
              if ($unsigned($signed(forvar508[(2'h2):(1'h1)])))
                begin
                  for (forvar643 = (1'h0); (forvar643 < (1'h1)); forvar643 = (forvar643 + (1'h1)))
                    begin
                      reg644 <= (forvar646 || {((reg434 ? wire430 : reg464) ?
                              {wire18} : $unsigned(reg547))});
                    end
                  for (forvar645 = (1'h0); (forvar645 < (1'h1)); forvar645 = (forvar645 + (1'h1)))
                    begin
                      reg646 <= ($signed({(reg557 ^~ reg470)}) ?
                          reg523 : (((~^reg655) ?
                                  {forvar606} : $signed(forvar440)) ?
                              ($unsigned(reg524) * $unsigned(reg595)) : ($signed(reg486) ?
                                  $unsigned(reg625) : $signed(forvar485))));
                    end
                end
              else
                begin
                  if ($signed((-reg632)))
                    begin
                      reg643 <= $signed({$signed((forvar570 + reg451))});
                      reg644 <= forvar508;
                      reg645 <= (~|$signed(($unsigned((8'hb7)) ?
                          reg599 : $signed((8'hb6)))));
                    end
                  else
                    begin
                      reg643 <= (forvar451[(4'h8):(4'h8)] < $unsigned(reg506));
                      reg644 <= (~&reg654);
                      reg645 <= $unsigned(($signed((^reg566)) == forvar540));
                    end
                  if ((reg469[(3'h5):(2'h2)] >>> (((-forvar483) ?
                      reg553 : (forvar637 ?
                          reg595 : reg492)) & ((+reg595) == (reg491 ~^ reg640)))))
                    begin
                      reg646 <= ((~&(reg446 ?
                          $signed(reg636) : $unsigned(reg496))) < (~|{(forvar588 ^ (8'hac))}));
                      reg647 <= forvar538[(3'h5):(3'h5)];
                    end
                  else
                    begin
                      reg646 <= forvar522[(1'h0):(1'h0)];
                      reg647 <= ($unsigned({(8'ha8)}) ?
                          $unsigned($signed($signed(reg645))) : (8'ha7));
                    end
                end
              reg648 <= reg651[(2'h2):(1'h0)];
              for (forvar649 = (1'h0); (forvar649 < (1'h0)); forvar649 = (forvar649 + (1'h1)))
                begin
                  for (forvar650 = (1'h0); (forvar650 < (2'h2)); forvar650 = (forvar650 + (1'h1)))
                    begin
                      reg651 <= ($signed((reg595 ?
                          forvar533 : $unsigned((8'ha1)))) << reg458);
                      reg652 <= $signed((reg562 ? wire16 : forvar456));
                    end
                  if ($unsigned(reg529[(3'h7):(1'h0)]))
                    begin
                      reg653 <= $unsigned(forvar645);
                      reg654 <= $unsigned((reg537[(1'h1):(1'h1)] ?
                          {forvar598} : (|reg462)));
                    end
                  else
                    begin
                      reg653 <= (~|$unsigned({$signed(reg649)}));
                      reg654 <= (&((~&$unsigned(forvar549)) ?
                          $signed($signed(reg440)) : $signed((reg527 ?
                              forvar662 : forvar509))));
                    end
                end
            end
          else
            begin
              for (forvar637 = (1'h0); (forvar637 < (1'h0)); forvar637 = (forvar637 + (1'h1)))
                begin
                  if ($unsigned({reg590}))
                    begin
                      reg638 <= reg511[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg638 <= $signed(reg661);
                      reg639 <= ($unsigned($unsigned((wire532 || reg580))) >= $unsigned((forvar556[(4'h9):(4'h9)] ?
                          (reg451 > (8'ha7)) : (8'ha3))));
                      reg640 <= reg586[(2'h2):(1'h0)];
                      reg641 <= (reg547[(4'hc):(3'h4)] ?
                          reg583[(4'h8):(1'h0)] : (~^reg529[(3'h4):(1'h0)]));
                    end
                  for (forvar642 = (1'h0); (forvar642 < (2'h2)); forvar642 = (forvar642 + (1'h1)))
                    begin
                      reg643 <= ((~|(|{reg529})) ?
                          (8'hb8) : (($signed(reg565) ?
                              reg621[(2'h2):(1'h0)] : $unsigned(reg619)) > forvar617));
                      reg644 <= reg594[(2'h2):(2'h2)];
                      reg645 <= (reg459[(4'h9):(1'h0)] & ((((8'ha6) ?
                                  (8'had) : reg593) ?
                              reg623[(2'h2):(1'h1)] : $unsigned(reg519)) ?
                          ({reg527} > forvar651[(3'h7):(3'h4)]) : ((reg597 & forvar451) ^ (reg544 ?
                              reg549 : forvar571))));
                      reg646 <= ((8'hb9) ?
                          (^~$unsigned(((8'ha5) - reg620))) : forvar585);
                    end
                end
              if ((8'ha4))
                begin
                  for (forvar647 = (1'h0); (forvar647 < (1'h0)); forvar647 = (forvar647 + (1'h1)))
                    begin
                      reg648 <= $signed(reg590[(4'hd):(1'h1)]);
                      reg649 <= $unsigned((((forvar439 | reg644) ?
                          ((8'h9d) + reg512) : (&(8'h9d))) & reg543[(3'h4):(3'h4)]));
                    end
                end
              else
                begin
                  if (reg555)
                    begin
                      reg647 <= (~{$signed($unsigned(forvar649))});
                      reg648 <= {$signed($unsigned(forvar504))};
                    end
                  else
                    begin
                      reg647 <= (~|{reg657});
                      reg648 <= forvar474[(3'h5):(3'h4)];
                    end
                end
            end
          reg655 <= forvar643[(2'h3):(2'h2)];
          for (forvar656 = (1'h0); (forvar656 < (2'h2)); forvar656 = (forvar656 + (1'h1)))
            begin
              if (reg497[(1'h0):(1'h0)])
                begin
                  for (forvar657 = (1'h0); (forvar657 < (1'h1)); forvar657 = (forvar657 + (1'h1)))
                    begin
                      reg658 <= ($unsigned((^~$signed(forvar490))) ^~ $signed($signed((~reg559))));
                      reg659 <= (!$unsigned((reg591[(1'h1):(1'h1)] ?
                          (reg463 | (8'hb2)) : reg642[(3'h6):(1'h0)])));
                      reg660 <= {reg636[(3'h7):(2'h2)]};
                    end
                  reg661 <= {(8'hb1)};
                end
              else
                begin
                  for (forvar657 = (1'h0); (forvar657 < (2'h3)); forvar657 = (forvar657 + (1'h1)))
                    begin
                      reg658 <= (^~$signed((~&{forvar446})));
                    end
                  for (forvar659 = (1'h0); (forvar659 < (1'h1)); forvar659 = (forvar659 + (1'h1)))
                    begin
                      reg660 <= forvar549[(3'h7):(3'h5)];
                      reg661 <= (^reg535[(4'he):(4'he)]);
                      reg662 <= (|$unsigned($signed({(8'h9d)})));
                      reg663 <= {reg644[(1'h1):(1'h0)]};
                    end
                  reg664 <= {(~^(!forvar617))};
                  for (forvar665 = (1'h0); (forvar665 < (2'h2)); forvar665 = (forvar665 + (1'h1)))
                    begin
                      reg666 <= reg447[(4'ha):(3'h6)];
                      reg667 <= reg599[(2'h3):(2'h2)];
                      reg668 <= ($signed($signed($signed(reg619))) ?
                          $signed((~&(wire18 << reg538))) : ({wire18[(3'h6):(2'h3)]} > ((reg526 ^ reg491) ^ (8'hb9))));
                    end
                end
            end
          for (forvar669 = (1'h0); (forvar669 < (2'h2)); forvar669 = (forvar669 + (1'h1)))
            begin
              reg670 <= (($unsigned((!reg520)) ?
                  (forvar496[(1'h1):(1'h0)] | reg615) : (~reg529)) >= ((forvar538[(2'h2):(1'h1)] ?
                  reg546[(2'h2):(1'h1)] : {reg487}) == (-(reg600 <<< forvar450))));
              for (forvar671 = (1'h0); (forvar671 < (1'h1)); forvar671 = (forvar671 + (1'h1)))
                begin
                  if ((8'ha7))
                    begin
                      reg672 <= $signed($signed(($signed(reg599) ?
                          (^reg650) : $unsigned(reg436))));
                      reg673 <= forvar575[(3'h7):(1'h0)];
                      reg674 <= reg467;
                      reg675 <= (^$signed($unsigned((reg523 ?
                          reg439 : (8'hb0)))));
                    end
                  else
                    begin
                      reg672 <= $unsigned(reg565);
                      reg673 <= ({(reg499[(3'h4):(3'h4)] || forvar647[(3'h4):(2'h3)])} ?
                          {$signed((~&(8'ha0)))} : $unsigned((reg478 ?
                              (forvar552 ?
                                  wire189 : reg453) : $unsigned(reg494))));
                      reg674 <= $signed((((forvar485 ? reg549 : forvar549) ?
                              ((8'h9d) ? reg516 : reg610) : (&reg478)) ?
                          reg503 : $unsigned(wire530)));
                    end
                  if (reg482[(4'h8):(3'h5)])
                    begin
                      reg676 <= (forvar671 ? {$unsigned({(8'ha0)})} : reg626);
                      reg677 <= $signed($unsigned(reg580[(3'h6):(3'h6)]));
                      reg678 <= (8'ha0);
                      reg679 <= forvar651[(1'h0):(1'h0)];
                    end
                  else
                    begin
                      reg676 <= reg535[(4'hb):(3'h5)];
                      reg677 <= (forvar491[(3'h4):(1'h0)] ?
                          (reg451 | forvar611[(1'h1):(1'h0)]) : (^~reg655[(3'h5):(3'h4)]));
                      reg678 <= $unsigned(({(reg482 >> reg652)} ?
                          reg470 : reg674[(4'hd):(4'h9)]));
                      reg679 <= {(+($signed(reg675) >= (^~(8'ha2))))};
                    end
                  for (forvar680 = (1'h0); (forvar680 < (2'h3)); forvar680 = (forvar680 + (1'h1)))
                    begin
                      reg681 <= $signed($signed({$unsigned(forvar646)}));
                      reg682 <= reg453[(4'h9):(3'h4)];
                      reg683 <= $unsigned((+{forvar499[(4'h8):(1'h0)]}));
                      reg684 <= ((((8'ha4) && forvar525) < (forvar617[(3'h4):(2'h2)] ?
                          (8'ha6) : reg516)) >> $unsigned((!$signed(forvar442))));
                    end
                end
              for (forvar685 = (1'h0); (forvar685 < (1'h1)); forvar685 = (forvar685 + (1'h1)))
                begin
                  for (forvar686 = (1'h0); (forvar686 < (1'h1)); forvar686 = (forvar686 + (1'h1)))
                    begin
                      reg687 <= $signed((^(&(~reg587))));
                    end
                  for (forvar688 = (1'h0); (forvar688 < (2'h2)); forvar688 = (forvar688 + (1'h1)))
                    begin
                      reg689 <= $signed(forvar522[(1'h0):(1'h0)]);
                      reg690 <= $signed((forvar549[(3'h6):(2'h3)] ?
                          (+(-reg659)) : ({reg489} ?
                              (forvar539 << forvar606) : (reg520 ?
                                  forvar450 : reg463))));
                      reg691 <= (-(($signed(forvar647) ^ ((8'h9c) | forvar680)) ?
                          (forvar484 ?
                              $signed(reg517) : (reg670 && forvar451)) : (reg436 ?
                              forvar484[(3'h6):(3'h5)] : (~^reg569))));
                    end
                  if ({reg473})
                    begin
                      reg692 <= $unsigned($unsigned($signed(forvar496[(1'h0):(1'h0)])));
                      reg693 <= $unsigned($signed(({wire532} ~^ $signed(forvar585))));
                      reg694 <= (^~$unsigned(((forvar538 ?
                          wire17 : (8'h9d)) + (forvar514 ? reg443 : wire531))));
                    end
                  else
                    begin
                      reg692 <= reg435[(3'h6):(3'h4)];
                      reg693 <= (({$signed(reg584)} ?
                          (8'ha1) : wire429[(1'h0):(1'h0)]) != $unsigned({$unsigned((8'hb1))}));
                    end
                  if ($signed(reg564))
                    begin
                      reg695 <= ((((reg567 ? reg549 : reg594) ?
                          $unsigned(wire186) : $signed(reg499)) > (^reg564[(4'ha):(1'h1)])) <<< (reg681[(1'h1):(1'h0)] ?
                          forvar456 : forvar603[(3'h6):(3'h4)]));
                      reg696 <= ((($unsigned(reg442) ?
                              $unsigned((8'ha5)) : $unsigned(forvar574)) > ($signed(reg455) ?
                              (-(8'h9e)) : wire17)) ?
                          ({(~(8'haf))} ?
                              (~|forvar656) : wire186) : $signed($signed(forvar548)));
                      reg697 <= ($unsigned((wire189[(3'h7):(3'h6)] ?
                          (reg535 + reg675) : (forvar442 > forvar485))) | forvar443);
                      reg698 <= (-({$unsigned(reg619)} * $signed($unsigned(reg564))));
                    end
                  else
                    begin
                      reg695 <= $signed((8'ha3));
                      reg696 <= reg450;
                      reg697 <= $signed((+reg491));
                      reg698 <= ($signed((8'hae)) ^~ {(forvar509[(3'h6):(2'h2)] ~^ reg486)});
                    end
                end
            end
        end
      reg699 <= {forvar453};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module190  (y, clk, wire195, wire194, wire193, wire192, wire191);
  output wire [(32'h99d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire195;
  input wire signed [(3'h5):(1'h0)] wire194;
  input wire [(4'ha):(1'h0)] wire193;
  input wire [(3'h7):(1'h0)] wire192;
  input wire [(3'h5):(1'h0)] wire191;
  reg signed [(4'ha):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg425 = (1'h0);
  reg [(3'h7):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg423 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg422 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar421 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg420 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg419 = (1'h0);
  reg [(4'hf):(1'h0)] reg418 = (1'h0);
  reg [(4'he):(1'h0)] reg417 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar416 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg415 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar414 = (1'h0);
  reg signed [(4'he):(1'h0)] reg413 = (1'h0);
  reg [(4'ha):(1'h0)] forvar412 = (1'h0);
  reg [(3'h7):(1'h0)] forvar411 = (1'h0);
  reg [(2'h3):(1'h0)] reg410 = (1'h0);
  reg [(4'hd):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg408 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg406 = (1'h0);
  reg [(3'h4):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg404 = (1'h0);
  reg [(4'hc):(1'h0)] forvar403 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg402 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg401 = (1'h0);
  reg [(3'h7):(1'h0)] forvar400 = (1'h0);
  reg [(3'h7):(1'h0)] forvar399 = (1'h0);
  reg [(2'h3):(1'h0)] reg398 = (1'h0);
  reg [(5'h10):(1'h0)] forvar397 = (1'h0);
  reg [(3'h7):(1'h0)] forvar396 = (1'h0);
  reg [(4'hc):(1'h0)] reg395 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar394 = (1'h0);
  reg [(4'ha):(1'h0)] reg393 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg392 = (1'h0);
  reg [(5'h10):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg390 = (1'h0);
  reg [(2'h3):(1'h0)] forvar389 = (1'h0);
  reg [(4'hd):(1'h0)] reg388 = (1'h0);
  reg [(4'hc):(1'h0)] reg387 = (1'h0);
  reg [(3'h5):(1'h0)] forvar386 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg385 = (1'h0);
  reg [(3'h6):(1'h0)] reg384 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg383 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar382 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar381 = (1'h0);
  reg [(4'hf):(1'h0)] forvar380 = (1'h0);
  reg [(4'hd):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg378 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar377 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg376 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg375 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar374 = (1'h0);
  reg [(2'h2):(1'h0)] reg373 = (1'h0);
  reg signed [(4'he):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg371 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg370 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar369 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar368 = (1'h0);
  reg [(4'hf):(1'h0)] forvar364 = (1'h0);
  reg [(4'ha):(1'h0)] reg358 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar355 = (1'h0);
  reg signed [(4'he):(1'h0)] reg353 = (1'h0);
  reg [(5'h10):(1'h0)] reg348 = (1'h0);
  reg [(4'he):(1'h0)] reg342 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg369 = (1'h0);
  reg [(3'h4):(1'h0)] reg368 = (1'h0);
  reg [(3'h5):(1'h0)] reg367 = (1'h0);
  reg [(4'h8):(1'h0)] reg366 = (1'h0);
  reg [(4'hb):(1'h0)] reg365 = (1'h0);
  reg [(3'h5):(1'h0)] reg364 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg362 = (1'h0);
  reg [(4'hb):(1'h0)] reg361 = (1'h0);
  reg [(4'he):(1'h0)] reg360 = (1'h0);
  reg [(4'he):(1'h0)] reg359 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg357 = (1'h0);
  reg [(3'h5):(1'h0)] reg356 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg355 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg354 = (1'h0);
  reg [(5'h10):(1'h0)] forvar353 = (1'h0);
  reg [(3'h6):(1'h0)] forvar352 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg347 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar344 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg343 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar341 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg352 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg351 = (1'h0);
  reg [(4'h9):(1'h0)] reg350 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar348 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar347 = (1'h0);
  reg [(2'h2):(1'h0)] reg346 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg345 = (1'h0);
  reg signed [(4'he):(1'h0)] reg344 = (1'h0);
  reg [(4'hb):(1'h0)] forvar343 = (1'h0);
  reg [(4'hf):(1'h0)] forvar342 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg341 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg340 = (1'h0);
  reg [(5'h10):(1'h0)] reg339 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg338 = (1'h0);
  reg [(4'he):(1'h0)] reg337 = (1'h0);
  reg [(4'ha):(1'h0)] reg336 = (1'h0);
  reg [(4'he):(1'h0)] reg335 = (1'h0);
  reg [(3'h4):(1'h0)] reg334 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg331 = (1'h0);
  reg [(4'hf):(1'h0)] reg333 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg332 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar331 = (1'h0);
  reg [(4'hb):(1'h0)] forvar330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg329 = (1'h0);
  reg [(4'hc):(1'h0)] forvar328 = (1'h0);
  reg [(2'h2):(1'h0)] reg327 = (1'h0);
  reg [(4'he):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg325 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg324 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg323 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg322 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg321 = (1'h0);
  reg [(3'h6):(1'h0)] forvar320 = (1'h0);
  reg signed [(4'he):(1'h0)] reg319 = (1'h0);
  reg [(4'hc):(1'h0)] reg318 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg317 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg316 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar315 = (1'h0);
  reg [(3'h4):(1'h0)] reg314 = (1'h0);
  reg [(4'hc):(1'h0)] forvar313 = (1'h0);
  reg [(3'h4):(1'h0)] reg312 = (1'h0);
  reg [(3'h7):(1'h0)] reg311 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg310 = (1'h0);
  reg [(4'h8):(1'h0)] reg309 = (1'h0);
  reg [(3'h4):(1'h0)] forvar308 = (1'h0);
  reg [(4'hd):(1'h0)] forvar299 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg298 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar295 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg293 = (1'h0);
  reg [(4'h9):(1'h0)] forvar290 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg307 = (1'h0);
  reg [(5'h10):(1'h0)] reg306 = (1'h0);
  reg [(3'h5):(1'h0)] reg305 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg304 = (1'h0);
  reg [(4'h9):(1'h0)] forvar303 = (1'h0);
  reg [(4'hf):(1'h0)] reg302 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg301 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg300 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg299 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar298 = (1'h0);
  reg [(3'h7):(1'h0)] reg297 = (1'h0);
  reg [(3'h7):(1'h0)] reg296 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg295 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg294 = (1'h0);
  reg [(3'h4):(1'h0)] forvar293 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg292 = (1'h0);
  reg [(3'h4):(1'h0)] reg291 = (1'h0);
  reg [(3'h6):(1'h0)] reg290 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg289 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg288 = (1'h0);
  reg [(4'hb):(1'h0)] forvar287 = (1'h0);
  reg [(2'h2):(1'h0)] reg285 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg283 = (1'h0);
  reg [(2'h2):(1'h0)] reg286 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar285 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg284 = (1'h0);
  reg [(4'hd):(1'h0)] forvar283 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar282 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg245 = (1'h0);
  reg [(4'hc):(1'h0)] reg281 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg280 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar279 = (1'h0);
  reg [(4'hd):(1'h0)] reg278 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg277 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg276 = (1'h0);
  reg [(4'hd):(1'h0)] reg275 = (1'h0);
  reg [(3'h5):(1'h0)] reg274 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg273 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg272 = (1'h0);
  reg [(3'h4):(1'h0)] reg271 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg270 = (1'h0);
  reg [(3'h4):(1'h0)] reg269 = (1'h0);
  reg [(4'ha):(1'h0)] reg268 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar267 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar266 = (1'h0);
  reg [(4'h9):(1'h0)] forvar261 = (1'h0);
  reg [(4'ha):(1'h0)] reg259 = (1'h0);
  reg signed [(4'he):(1'h0)] reg265 = (1'h0);
  reg [(4'hd):(1'h0)] reg264 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg263 = (1'h0);
  reg [(4'hc):(1'h0)] reg262 = (1'h0);
  reg [(4'hb):(1'h0)] reg261 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg260 = (1'h0);
  reg [(4'ha):(1'h0)] forvar259 = (1'h0);
  reg [(3'h5):(1'h0)] reg258 = (1'h0);
  reg [(3'h7):(1'h0)] reg257 = (1'h0);
  reg [(5'h10):(1'h0)] reg256 = (1'h0);
  reg [(3'h7):(1'h0)] reg255 = (1'h0);
  reg [(3'h4):(1'h0)] forvar254 = (1'h0);
  reg signed [(4'he):(1'h0)] reg253 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg252 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg250 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar249 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg248 = (1'h0);
  reg [(4'h8):(1'h0)] reg247 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg246 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar245 = (1'h0);
  reg [(4'he):(1'h0)] forvar244 = (1'h0);
  reg [(3'h6):(1'h0)] reg238 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg243 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg242 = (1'h0);
  reg [(4'h9):(1'h0)] forvar241 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg240 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg239 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar238 = (1'h0);
  reg [(3'h4):(1'h0)] reg237 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg236 = (1'h0);
  reg [(4'he):(1'h0)] reg235 = (1'h0);
  reg [(4'h8):(1'h0)] forvar234 = (1'h0);
  reg [(4'h8):(1'h0)] reg233 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg232 = (1'h0);
  reg [(3'h5):(1'h0)] reg231 = (1'h0);
  reg signed [(4'he):(1'h0)] reg230 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar228 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar227 = (1'h0);
  reg [(3'h6):(1'h0)] reg228 = (1'h0);
  reg [(4'h8):(1'h0)] reg227 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg226 = (1'h0);
  reg [(3'h7):(1'h0)] reg225 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg224 = (1'h0);
  reg [(4'ha):(1'h0)] reg223 = (1'h0);
  reg [(4'hd):(1'h0)] reg222 = (1'h0);
  reg [(4'h9):(1'h0)] reg221 = (1'h0);
  reg [(2'h2):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg219 = (1'h0);
  reg [(3'h5):(1'h0)] reg218 = (1'h0);
  reg [(3'h5):(1'h0)] forvar217 = (1'h0);
  reg [(4'h9):(1'h0)] forvar216 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg214 = (1'h0);
  reg signed [(4'he):(1'h0)] reg213 = (1'h0);
  reg [(4'hd):(1'h0)] reg212 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar211 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg210 = (1'h0);
  reg [(4'hf):(1'h0)] forvar209 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg208 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg207 = (1'h0);
  reg [(4'hb):(1'h0)] reg206 = (1'h0);
  reg [(3'h4):(1'h0)] reg205 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg204 = (1'h0);
  reg [(4'he):(1'h0)] forvar203 = (1'h0);
  reg [(3'h6):(1'h0)] forvar202 = (1'h0);
  reg [(4'h8):(1'h0)] reg202 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire201;
  wire [(4'he):(1'h0)] wire200;
  wire signed [(3'h7):(1'h0)] wire199;
  wire signed [(2'h3):(1'h0)] wire198;
  wire signed [(4'h9):(1'h0)] wire197;
  wire [(4'hb):(1'h0)] wire196;
  assign y = {reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 forvar421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 forvar416,
                 reg415,
                 forvar414,
                 reg413,
                 forvar412,
                 forvar411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 reg406,
                 reg405,
                 reg404,
                 forvar403,
                 reg402,
                 reg401,
                 forvar400,
                 forvar399,
                 reg398,
                 forvar397,
                 forvar396,
                 reg395,
                 forvar394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 forvar389,
                 reg388,
                 reg387,
                 forvar386,
                 reg385,
                 reg384,
                 reg383,
                 forvar382,
                 forvar381,
                 forvar380,
                 reg379,
                 reg378,
                 forvar377,
                 reg376,
                 reg375,
                 forvar374,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 forvar369,
                 forvar368,
                 forvar364,
                 reg358,
                 forvar355,
                 reg353,
                 reg348,
                 reg342,
                 reg369,
                 reg368,
                 reg367,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg359,
                 forvar358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 forvar353,
                 forvar352,
                 reg347,
                 forvar344,
                 reg343,
                 forvar341,
                 reg352,
                 reg351,
                 reg350,
                 reg349,
                 forvar348,
                 forvar347,
                 reg346,
                 reg345,
                 reg344,
                 forvar343,
                 forvar342,
                 reg341,
                 reg340,
                 reg339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg331,
                 reg333,
                 reg332,
                 forvar331,
                 forvar330,
                 reg329,
                 forvar328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 forvar320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 forvar315,
                 reg314,
                 forvar313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 forvar308,
                 forvar299,
                 reg298,
                 forvar295,
                 reg293,
                 forvar290,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 forvar303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 forvar298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 forvar293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 forvar287,
                 reg285,
                 reg283,
                 reg286,
                 forvar285,
                 reg284,
                 forvar283,
                 forvar282,
                 reg249,
                 reg245,
                 reg281,
                 reg280,
                 forvar279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg270,
                 reg269,
                 reg268,
                 forvar267,
                 forvar266,
                 forvar261,
                 reg259,
                 reg265,
                 reg264,
                 reg263,
                 reg262,
                 reg261,
                 reg260,
                 forvar259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 forvar254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 forvar249,
                 reg248,
                 reg247,
                 reg246,
                 forvar245,
                 forvar244,
                 reg238,
                 reg243,
                 reg242,
                 forvar241,
                 reg240,
                 reg239,
                 forvar238,
                 reg237,
                 reg236,
                 reg235,
                 forvar234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 forvar228,
                 forvar227,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 forvar217,
                 forvar216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 forvar211,
                 reg210,
                 forvar209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 forvar203,
                 forvar202,
                 reg202,
                 wire201,
                 wire200,
                 wire199,
                 wire198,
                 wire197,
                 wire196,
                 (1'h0)};
  assign wire196 = wire194[(2'h2):(1'h0)];
  assign wire197 = ((~|$unsigned((8'hb0))) ?
                       (~$unsigned((8'hb7))) : wire193[(1'h0):(1'h0)]);
  assign wire198 = $unsigned(wire191);
  assign wire199 = (wire193[(4'h9):(4'h8)] ?
                       {{wire191}} : $signed(wire195[(3'h5):(2'h3)]));
  assign wire200 = ($unsigned(wire198) ?
                       wire197[(3'h6):(3'h5)] : (((wire197 != wire196) <= ((8'ha8) ?
                           wire196 : wire199)) >> {{wire191}}));
  assign wire201 = ($signed((wire191 ?
                       $unsigned(wire196) : (wire200 ?
                           wire196 : wire194))) | $unsigned({wire196[(4'ha):(1'h1)]}));
  always
    @(posedge clk) begin
      if (($unsigned((~|wire194[(3'h5):(3'h5)])) || {(((8'hac) ^ wire191) == (wire193 & wire195))}))
        begin
          reg202 <= ($unsigned($unsigned($unsigned(wire198))) ?
              $signed({(wire196 ? wire194 : wire198)}) : wire193);
        end
      else
        begin
          for (forvar202 = (1'h0); (forvar202 < (2'h2)); forvar202 = (forvar202 + (1'h1)))
            begin
              if ($unsigned(($unsigned($unsigned(wire192)) | wire199)))
                begin
                  for (forvar203 = (1'h0); (forvar203 < (2'h2)); forvar203 = (forvar203 + (1'h1)))
                    begin
                      reg204 <= {$signed(wire193[(4'h8):(3'h6)])};
                      reg205 <= ((wire194 - $unsigned($signed(forvar202))) ?
                          ($signed($signed(wire200)) + $unsigned((wire195 >= (8'hab)))) : $unsigned({wire193}));
                      reg206 <= (!{($unsigned((8'hba)) == reg205)});
                      reg207 <= (($unsigned((reg205 ?
                              wire198 : wire199)) ^ $signed(wire197)) ?
                          $unsigned(reg204[(3'h6):(3'h4)]) : ($unsigned({reg205}) ?
                              $unsigned({forvar203}) : wire194));
                    end
                  if ((~|wire196))
                    begin
                      reg208 <= (|(|wire199));
                    end
                  else
                    begin
                      reg208 <= (($unsigned((wire192 ? reg204 : wire194)) ?
                          forvar203[(4'h9):(1'h0)] : {reg205[(1'h1):(1'h1)]}) | $signed((((8'hb7) ?
                              reg205 : (8'hac)) ?
                          $signed(wire192) : $signed((8'ha3)))));
                    end
                  for (forvar209 = (1'h0); (forvar209 < (1'h0)); forvar209 = (forvar209 + (1'h1)))
                    begin
                      reg210 <= wire196;
                    end
                  for (forvar211 = (1'h0); (forvar211 < (1'h1)); forvar211 = (forvar211 + (1'h1)))
                    begin
                      reg212 <= reg202;
                      reg213 <= ((~&(~(wire200 ? reg208 : reg212))) ?
                          (($unsigned(reg208) >>> reg208) ?
                              $unsigned($unsigned(reg207)) : $signed($signed((8'hb9)))) : (wire199 | wire198));
                      reg214 <= $unsigned(wire197);
                      reg215 <= (^~(reg207 ?
                          {$signed((8'hb0))} : $unsigned($unsigned(wire197))));
                    end
                end
              else
                begin
                  for (forvar203 = (1'h0); (forvar203 < (2'h2)); forvar203 = (forvar203 + (1'h1)))
                    begin
                      reg204 <= wire193;
                      reg205 <= $unsigned(forvar202[(3'h5):(3'h5)]);
                    end
                  reg206 <= (!{(+$signed(reg215))});
                end
            end
          for (forvar216 = (1'h0); (forvar216 < (1'h0)); forvar216 = (forvar216 + (1'h1)))
            begin
              for (forvar217 = (1'h0); (forvar217 < (2'h2)); forvar217 = (forvar217 + (1'h1)))
                begin
                  if ($unsigned({reg205[(1'h0):(1'h0)]}))
                    begin
                      reg218 <= {forvar203};
                      reg219 <= $signed((!$unsigned(reg214)));
                    end
                  else
                    begin
                      reg218 <= $signed(((wire199 ?
                          (!reg212) : $signed(reg212)) && (&$unsigned((8'hb7)))));
                    end
                  if ($unsigned(wire193))
                    begin
                      reg220 <= $unsigned((^$signed($unsigned((8'hb0)))));
                      reg221 <= $unsigned($unsigned(reg214));
                    end
                  else
                    begin
                      reg220 <= reg220[(2'h2):(1'h0)];
                    end
                  if ($signed($unsigned(($signed(reg212) + (~^reg219)))))
                    begin
                      reg222 <= reg204;
                      reg223 <= $signed(($unsigned(wire201[(3'h6):(3'h6)]) ?
                          (~(forvar211 ?
                              wire196 : forvar203)) : (((8'ha4) <= forvar202) ?
                              $signed(wire191) : forvar217)));
                    end
                  else
                    begin
                      reg222 <= (wire199 << ($unsigned((+(8'hb1))) ?
                          (8'hb1) : ({(8'hb3)} <<< {wire200})));
                    end
                  if (($unsigned($unsigned((~&reg218))) ?
                      (($signed(reg218) > reg222) ?
                          ((wire199 ? (8'ha4) : (8'ha3)) ?
                              wire193[(3'h6):(3'h6)] : {reg206}) : wire201) : (^$unsigned(wire199))))
                    begin
                      reg224 <= (reg215 ?
                          {(~|(reg202 ^ reg212))} : $unsigned($unsigned($unsigned(wire193))));
                      reg225 <= (((reg223 ?
                                  reg202[(2'h2):(1'h1)] : $unsigned(forvar209)) ?
                              wire198[(2'h3):(2'h2)] : (~|wire197[(3'h6):(1'h1)])) ?
                          {((forvar217 ? reg214 : reg213) ?
                                  reg212 : $signed(wire201))} : wire191);
                      reg226 <= ($unsigned({(~|wire196)}) ?
                          forvar217 : (reg222 | forvar203[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg224 <= reg206;
                      reg225 <= (wire201 ?
                          {$signed($unsigned(wire196))} : forvar203[(4'h9):(4'h9)]);
                    end
                end
            end
          if ((reg215[(3'h5):(1'h1)] ^ wire196[(3'h5):(3'h5)]))
            begin
              reg227 <= ($signed($unsigned(((8'ha5) >= wire201))) | (reg207 != $signed({reg219})));
              reg228 <= (wire200[(3'h7):(3'h6)] | ({$unsigned(reg220)} ?
                  forvar217[(2'h2):(1'h0)] : forvar217[(3'h5):(2'h3)]));
            end
          else
            begin
              for (forvar227 = (1'h0); (forvar227 < (2'h2)); forvar227 = (forvar227 + (1'h1)))
                begin
                  for (forvar228 = (1'h0); (forvar228 < (2'h3)); forvar228 = (forvar228 + (1'h1)))
                    begin
                      reg229 <= (wire191[(2'h2):(2'h2)] ?
                          $unsigned(reg224) : reg205);
                      reg230 <= ($signed(($unsigned(reg221) <= $unsigned((8'hb1)))) ?
                          ($unsigned((forvar211 && wire196)) ?
                              $signed(reg208) : $signed((wire201 * reg210))) : (^~$unsigned((reg205 ?
                              (8'haa) : (8'haa)))));
                      reg231 <= forvar228;
                      reg232 <= $signed((8'hb0));
                    end
                end
              reg233 <= ((8'hae) ?
                  (!(wire197[(3'h7):(1'h0)] && $unsigned((8'ha6)))) : (($signed(reg214) == $unsigned(reg219)) != wire200[(2'h2):(1'h0)]));
              for (forvar234 = (1'h0); (forvar234 < (2'h2)); forvar234 = (forvar234 + (1'h1)))
                begin
                  if ((8'hb2))
                    begin
                      reg235 <= forvar228;
                      reg236 <= {reg219};
                      reg237 <= (reg214 <= ((8'hb7) ~^ wire197[(4'h8):(3'h7)]));
                    end
                  else
                    begin
                      reg235 <= (&($signed(wire196[(4'hb):(3'h4)]) << $unsigned($unsigned((8'hae)))));
                      reg236 <= $unsigned($unsigned((reg225[(1'h1):(1'h0)] << (^~wire201))));
                    end
                end
              if (reg222)
                begin
                  for (forvar238 = (1'h0); (forvar238 < (2'h2)); forvar238 = (forvar238 + (1'h1)))
                    begin
                      reg239 <= (~&($unsigned(wire196[(3'h6):(2'h3)]) ?
                          reg219[(4'h8):(4'h8)] : $unsigned((reg208 ^ reg233))));
                      reg240 <= (-reg228);
                    end
                  for (forvar241 = (1'h0); (forvar241 < (2'h2)); forvar241 = (forvar241 + (1'h1)))
                    begin
                      reg242 <= $unsigned(reg212);
                      reg243 <= $unsigned(($unsigned(reg223[(1'h0):(1'h0)]) != ($signed((8'hb5)) <= (|reg237))));
                    end
                end
              else
                begin
                  reg238 <= {$unsigned(($unsigned(reg219) + ((8'ha2) ?
                          reg233 : wire191)))};
                end
            end
          if ($signed(reg227[(3'h6):(3'h5)]))
            begin
              for (forvar244 = (1'h0); (forvar244 < (1'h1)); forvar244 = (forvar244 + (1'h1)))
                begin
                  for (forvar245 = (1'h0); (forvar245 < (1'h0)); forvar245 = (forvar245 + (1'h1)))
                    begin
                      reg246 <= $unsigned($signed(((reg229 < (8'hb6)) & reg229)));
                      reg247 <= forvar227[(2'h3):(2'h2)];
                      reg248 <= (8'ha6);
                    end
                  for (forvar249 = (1'h0); (forvar249 < (2'h2)); forvar249 = (forvar249 + (1'h1)))
                    begin
                      reg250 <= (!reg242);
                      reg251 <= $signed($unsigned((reg224[(1'h1):(1'h0)] ^~ reg238[(2'h3):(1'h1)])));
                      reg252 <= {(reg222 || $unsigned(reg237[(2'h3):(1'h1)]))};
                      reg253 <= reg247;
                    end
                  for (forvar254 = (1'h0); (forvar254 < (2'h2)); forvar254 = (forvar254 + (1'h1)))
                    begin
                      reg255 <= (($signed({forvar249}) ^~ (^(wire198 ?
                              (8'haa) : forvar217))) ?
                          ((8'ha4) ?
                              reg246 : $signed((reg235 ?
                                  reg207 : reg236))) : (reg223 ?
                              ({forvar203} << (reg214 ?
                                  (8'ha1) : reg250)) : $unsigned((reg252 << wire201))));
                      reg256 <= (((8'ha9) ~^ (~(reg230 ?
                          reg237 : reg229))) | $signed(({forvar217} ?
                          (reg219 ? (8'ha9) : reg227) : reg253)));
                      reg257 <= $signed($unsigned(((~^forvar254) ^~ $signed(reg230))));
                      reg258 <= $signed($unsigned(forvar228));
                    end
                end
              if ($unsigned($signed({(-wire191)})))
                begin
                  for (forvar259 = (1'h0); (forvar259 < (1'h1)); forvar259 = (forvar259 + (1'h1)))
                    begin
                      reg260 <= $signed((!((forvar249 ?
                          reg250 : reg252) + $signed((8'hb8)))));
                      reg261 <= (((&forvar234) + wire193) != ($signed(forvar228[(3'h4):(1'h1)]) ?
                          $unsigned($unsigned(reg214)) : {$unsigned(reg256)}));
                      reg262 <= (-reg219[(4'h9):(3'h7)]);
                      reg263 <= reg238;
                    end
                  reg264 <= ($signed(({reg246} ?
                      reg253 : $signed(forvar203))) ^ (8'hb6));
                  reg265 <= forvar254[(3'h4):(2'h3)];
                end
              else
                begin
                  if (($unsigned(reg261) ?
                      forvar245 : $signed($signed((~|(8'hb0))))))
                    begin
                      reg259 <= $unsigned(reg264);
                      reg260 <= ((&(reg258 ?
                              (~(8'ha3)) : wire195[(4'ha):(3'h4)])) ?
                          ($unsigned(reg265) ?
                              ((^~reg236) << forvar217[(3'h5):(3'h5)]) : {(reg206 >= reg255)}) : ((-$unsigned(reg261)) && $signed(reg246[(4'h8):(1'h1)])));
                    end
                  else
                    begin
                      reg259 <= (8'haa);
                      reg260 <= reg204[(3'h6):(1'h1)];
                    end
                  for (forvar261 = (1'h0); (forvar261 < (1'h1)); forvar261 = (forvar261 + (1'h1)))
                    begin
                      reg262 <= $unsigned($signed(wire199[(2'h3):(2'h3)]));
                      reg263 <= ((forvar203 >= reg258[(2'h3):(2'h2)]) & (((reg224 ?
                                  wire191 : (8'h9f)) ?
                              $unsigned(reg260) : (forvar254 | reg219)) ?
                          $signed(forvar259) : $signed((reg235 ?
                              wire197 : reg253))));
                    end
                end
              for (forvar266 = (1'h0); (forvar266 < (1'h0)); forvar266 = (forvar266 + (1'h1)))
                begin
                  for (forvar267 = (1'h0); (forvar267 < (2'h3)); forvar267 = (forvar267 + (1'h1)))
                    begin
                      reg268 <= (!(|(~$signed(reg220))));
                      reg269 <= forvar202[(3'h4):(3'h4)];
                      reg270 <= (($unsigned(forvar216) ?
                          ((-(8'hb1)) ?
                              (forvar266 ?
                                  reg264 : reg246) : $signed(reg262)) : wire193) & $unsigned(wire201));
                      reg271 <= $signed(((^~$signed(reg253)) ?
                          $unsigned($signed((8'ha2))) : {(-wire199)}));
                    end
                  if (forvar234[(2'h3):(1'h0)])
                    begin
                      reg272 <= $signed($unsigned(reg255[(2'h3):(2'h2)]));
                    end
                  else
                    begin
                      reg272 <= (((8'hab) ?
                          ((-reg271) ?
                              $unsigned(reg261) : ((8'hb6) ?
                                  (8'hb4) : forvar254)) : $unsigned((reg222 && forvar202))) ~^ $signed($unsigned((reg218 - forvar228))));
                      reg273 <= $signed(reg233);
                      reg274 <= reg270;
                    end
                  if ($signed($signed($signed((forvar259 > (8'ha1))))))
                    begin
                      reg275 <= $unsigned((+reg260[(2'h3):(2'h3)]));
                      reg276 <= (($signed((forvar234 ? reg205 : wire201)) ?
                          (reg240 & wire193[(1'h0):(1'h0)]) : $unsigned((^~reg226))) <<< (&$signed(reg204[(2'h2):(2'h2)])));
                      reg277 <= $unsigned($unsigned(reg204));
                      reg278 <= forvar228;
                    end
                  else
                    begin
                      reg275 <= (reg231 ?
                          (wire193 ?
                              (8'hb7) : (!$signed((8'ha7)))) : reg229[(1'h1):(1'h1)]);
                      reg276 <= (reg213[(3'h4):(3'h4)] ^ forvar216);
                      reg277 <= (wire199[(1'h1):(1'h0)] * $unsigned($signed(forvar202)));
                    end
                  for (forvar279 = (1'h0); (forvar279 < (2'h2)); forvar279 = (forvar279 + (1'h1)))
                    begin
                      reg280 <= reg261;
                      reg281 <= $signed((reg205 + (~&(forvar209 & (8'ha7)))));
                    end
                end
            end
          else
            begin
              for (forvar244 = (1'h0); (forvar244 < (2'h3)); forvar244 = (forvar244 + (1'h1)))
                begin
                  if ($signed((!{(^wire199)})))
                    begin
                      reg245 <= (^~reg215[(3'h7):(3'h4)]);
                      reg246 <= ({reg236[(1'h0):(1'h0)]} ?
                          reg261 : reg274[(2'h3):(2'h2)]);
                    end
                  else
                    begin
                      reg245 <= ((($signed(reg247) ?
                          {wire199} : (wire201 >>> forvar227)) > $signed((reg235 >>> reg236))) <= $unsigned(reg264[(4'hb):(2'h3)]));
                      reg246 <= (forvar209 ?
                          wire197[(2'h2):(1'h0)] : {((~|reg261) ?
                                  (!reg218) : $signed(reg213))});
                    end
                  if ($unsigned((reg274[(3'h4):(2'h2)] & reg246)))
                    begin
                      reg247 <= $signed({($signed(forvar227) ?
                              (forvar202 ?
                                  reg271 : reg265) : forvar202[(2'h2):(2'h2)])});
                      reg248 <= $unsigned((|(reg230 ^~ (-(8'hb3)))));
                      reg249 <= ({reg237[(2'h2):(1'h1)]} ?
                          $unsigned($unsigned(reg222)) : ({{wire193}} == $signed(forvar228[(4'h8):(2'h2)])));
                    end
                  else
                    begin
                      reg247 <= wire197;
                      reg248 <= (-forvar259);
                    end
                end
            end
        end
      for (forvar282 = (1'h0); (forvar282 < (2'h3)); forvar282 = (forvar282 + (1'h1)))
        begin
          if ((^~forvar279))
            begin
              for (forvar283 = (1'h0); (forvar283 < (2'h2)); forvar283 = (forvar283 + (1'h1)))
                begin
                  reg284 <= reg232;
                end
            end
          else
            begin
              if ($signed($unsigned($unsigned((8'ha3)))))
                begin
                  for (forvar283 = (1'h0); (forvar283 < (1'h0)); forvar283 = (forvar283 + (1'h1)))
                    begin
                      reg284 <= $signed((((reg257 ?
                          reg207 : reg219) >>> reg275[(3'h7):(1'h0)]) < $unsigned(reg208[(4'h9):(3'h6)])));
                    end
                  for (forvar285 = (1'h0); (forvar285 < (1'h0)); forvar285 = (forvar285 + (1'h1)))
                    begin
                      reg286 <= $unsigned((~^(~&(!forvar209))));
                    end
                end
              else
                begin
                  if (($unsigned(((reg273 + (8'ha8)) ?
                          (reg207 + forvar217) : (reg286 ?
                              wire192 : forvar261))) ?
                      $unsigned({reg261}) : ({{reg222}} ?
                          $unsigned((reg258 * reg277)) : $signed(forvar203[(4'hd):(3'h6)]))))
                    begin
                      reg283 <= reg229;
                      reg284 <= ((^~{((8'hb7) <<< (8'ha4))}) ?
                          (reg235 == $signed(forvar238[(2'h3):(1'h0)])) : ((8'h9d) - $unsigned(reg238[(1'h0):(1'h0)])));
                      reg285 <= ($signed((+reg233[(3'h6):(2'h2)])) ?
                          $unsigned(((^~reg230) <<< (~wire195))) : reg284[(3'h5):(2'h2)]);
                      reg286 <= $signed($unsigned($signed((~|reg242))));
                    end
                  else
                    begin
                      reg283 <= (forvar209[(4'hd):(4'h8)] << $signed(wire197));
                    end
                  for (forvar287 = (1'h0); (forvar287 < (2'h2)); forvar287 = (forvar287 + (1'h1)))
                    begin
                      reg288 <= (^~($unsigned(forvar209) >= {$unsigned(reg271)}));
                      reg289 <= (-((|$unsigned(reg229)) ?
                          forvar209 : $signed((+(8'hb1)))));
                    end
                end
              if (reg206[(3'h4):(2'h2)])
                begin
                  if ({$unsigned((~(wire200 ^ (8'h9e))))})
                    begin
                      reg290 <= {($unsigned(forvar245) ?
                              ({reg210} ?
                                  $unsigned(reg231) : ((8'hb6) <= (8'hb7))) : (^$unsigned(reg229)))};
                      reg291 <= forvar279;
                    end
                  else
                    begin
                      reg290 <= reg250[(3'h7):(3'h4)];
                      reg291 <= (^~$signed($unsigned(forvar259)));
                      reg292 <= reg208;
                    end
                  for (forvar293 = (1'h0); (forvar293 < (2'h3)); forvar293 = (forvar293 + (1'h1)))
                    begin
                      reg294 <= ($signed(reg240) >>> reg226[(3'h4):(1'h0)]);
                      reg295 <= reg262[(2'h3):(1'h1)];
                      reg296 <= ((($signed((8'h9f)) ?
                          (reg252 ?
                              reg240 : reg230) : reg219[(4'h8):(3'h5)]) || reg264) ^ ((reg272[(4'hd):(3'h6)] ?
                              reg283[(3'h5):(1'h1)] : (reg213 ?
                                  reg242 : reg260)) ?
                          ((~^reg237) ?
                              $signed(reg247) : $unsigned((8'hb1))) : $unsigned(reg247[(3'h7):(3'h5)])));
                      reg297 <= {(~reg239)};
                    end
                  for (forvar298 = (1'h0); (forvar298 < (1'h0)); forvar298 = (forvar298 + (1'h1)))
                    begin
                      reg299 <= reg281[(3'h5):(2'h3)];
                      reg300 <= $unsigned($signed(reg268[(4'ha):(1'h0)]));
                      reg301 <= {$signed($unsigned({forvar282}))};
                      reg302 <= (forvar266 ?
                          ((~$signed(reg251)) ?
                              (+(~reg233)) : (+forvar259)) : $signed(((reg260 ?
                              (8'h9d) : reg258) > reg214)));
                    end
                  for (forvar303 = (1'h0); (forvar303 < (2'h3)); forvar303 = (forvar303 + (1'h1)))
                    begin
                      reg304 <= ($signed($unsigned((forvar202 ?
                          reg242 : forvar227))) << $unsigned(((forvar211 >= reg212) & (reg278 && reg301))));
                      reg305 <= ((|($unsigned(wire197) ?
                              reg281[(4'h8):(2'h2)] : (|(8'ha5)))) ?
                          $unsigned(reg295) : (^((reg272 >> reg269) ^~ $signed(forvar285))));
                      reg306 <= (reg246[(4'h9):(1'h1)] ?
                          {reg257[(3'h5):(3'h5)]} : $signed($signed(((8'ha5) ?
                              reg275 : reg260))));
                      reg307 <= forvar234;
                    end
                end
              else
                begin
                  for (forvar290 = (1'h0); (forvar290 < (2'h3)); forvar290 = (forvar290 + (1'h1)))
                    begin
                      reg291 <= (forvar267 ?
                          ($signed(reg307[(2'h3):(2'h2)]) ?
                              (~^(reg257 ~^ reg307)) : $signed({reg297})) : reg264);
                    end
                  if ($signed(reg208))
                    begin
                      reg292 <= {reg257[(2'h3):(2'h3)]};
                      reg293 <= reg302;
                      reg294 <= $unsigned((|reg238));
                    end
                  else
                    begin
                      reg292 <= reg233[(2'h2):(1'h0)];
                    end
                  for (forvar295 = (1'h0); (forvar295 < (2'h2)); forvar295 = (forvar295 + (1'h1)))
                    begin
                      reg296 <= ($signed($unsigned($signed(forvar279))) << reg293);
                      reg297 <= reg299[(2'h2):(2'h2)];
                      reg298 <= reg249;
                    end
                  for (forvar299 = (1'h0); (forvar299 < (1'h0)); forvar299 = (forvar299 + (1'h1)))
                    begin
                      reg300 <= (~forvar228);
                      reg301 <= reg256;
                    end
                end
              for (forvar308 = (1'h0); (forvar308 < (2'h3)); forvar308 = (forvar308 + (1'h1)))
                begin
                  if ((reg204[(3'h6):(3'h5)] & $signed(reg263)))
                    begin
                      reg309 <= (8'hb6);
                      reg310 <= ($unsigned(reg264[(3'h5):(2'h2)]) > {$unsigned({reg212})});
                      reg311 <= $unsigned(reg227[(2'h2):(1'h1)]);
                      reg312 <= ((forvar261[(3'h4):(2'h3)] ?
                          wire200 : (reg207 ? wire193 : reg309)) << reg245);
                    end
                  else
                    begin
                      reg309 <= ({{(~forvar308)}} ?
                          $signed(((reg250 ? reg257 : reg301) ?
                              reg296[(1'h0):(1'h0)] : ((8'ha0) ?
                                  reg206 : forvar279))) : ((!(forvar228 ?
                              (8'haf) : (8'ha9))) | wire200[(3'h5):(1'h1)]));
                      reg310 <= forvar287[(3'h4):(1'h1)];
                      reg311 <= {reg205};
                    end
                  for (forvar313 = (1'h0); (forvar313 < (1'h0)); forvar313 = (forvar313 + (1'h1)))
                    begin
                      reg314 <= reg272;
                    end
                  for (forvar315 = (1'h0); (forvar315 < (2'h3)); forvar315 = (forvar315 + (1'h1)))
                    begin
                      reg316 <= ((~^(reg206[(3'h5):(1'h0)] | (reg204 ?
                          reg306 : reg298))) & ($signed((8'ha0)) == reg290[(1'h1):(1'h0)]));
                      reg317 <= reg300[(3'h4):(1'h1)];
                      reg318 <= forvar295[(3'h7):(3'h6)];
                      reg319 <= $signed(reg311[(3'h6):(1'h1)]);
                    end
                end
              if ((~&{reg310}))
                begin
                  for (forvar320 = (1'h0); (forvar320 < (2'h2)); forvar320 = (forvar320 + (1'h1)))
                    begin
                      reg321 <= $unsigned(wire197);
                    end
                end
              else
                begin
                  for (forvar320 = (1'h0); (forvar320 < (2'h3)); forvar320 = (forvar320 + (1'h1)))
                    begin
                      reg321 <= $unsigned(forvar267);
                      reg322 <= ((&(reg280 ?
                          (forvar283 ? reg258 : reg236) : (&reg206))) - reg250);
                      reg323 <= reg286;
                    end
                  if ($unsigned((reg318 ?
                      ((8'ha7) ?
                          (reg210 ? reg277 : reg205) : (|reg249)) : (8'hb7))))
                    begin
                      reg324 <= {reg252[(3'h7):(1'h1)]};
                      reg325 <= reg276[(3'h5):(1'h1)];
                      reg326 <= (reg306[(1'h1):(1'h0)] && forvar267);
                    end
                  else
                    begin
                      reg324 <= $signed($signed((^forvar308[(2'h3):(2'h2)])));
                      reg325 <= (+(8'ha0));
                      reg326 <= $unsigned($unsigned($signed(reg250)));
                      reg327 <= ($unsigned(forvar238) + ((8'hb2) ?
                          reg276[(2'h3):(2'h3)] : (8'h9e)));
                    end
                  for (forvar328 = (1'h0); (forvar328 < (2'h3)); forvar328 = (forvar328 + (1'h1)))
                    begin
                      reg329 <= ($signed($unsigned((forvar315 ?
                          reg233 : reg291))) == {(reg314 * $signed(reg310))});
                    end
                end
            end
          if ($signed(($signed($signed(forvar303)) ?
              reg207 : $unsigned((reg219 ? forvar245 : reg205)))))
            begin
              for (forvar330 = (1'h0); (forvar330 < (2'h3)); forvar330 = (forvar330 + (1'h1)))
                begin
                  for (forvar331 = (1'h0); (forvar331 < (1'h0)); forvar331 = (forvar331 + (1'h1)))
                    begin
                      reg332 <= ((~reg286) * {(~&(!reg329))});
                      reg333 <= ({reg242[(2'h2):(1'h1)]} ?
                          ((reg284 >> (~^wire198)) <<< (reg311 * $unsigned(reg212))) : ({$signed(reg237)} ^~ (reg295 ^ {reg307})));
                    end
                end
            end
          else
            begin
              for (forvar330 = (1'h0); (forvar330 < (2'h2)); forvar330 = (forvar330 + (1'h1)))
                begin
                  if ($signed($signed(reg280)))
                    begin
                      reg331 <= wire200[(4'h9):(3'h4)];
                      reg332 <= {($unsigned((forvar285 && reg312)) ?
                              reg271[(1'h1):(1'h1)] : (~(~wire199)))};
                    end
                  else
                    begin
                      reg331 <= $unsigned((reg214[(3'h5):(1'h1)] >>> forvar320));
                      reg332 <= ($unsigned(reg295[(1'h0):(1'h0)]) ?
                          (reg228 <= ((-reg290) + (reg292 ^~ reg333))) : forvar254);
                      reg333 <= $unsigned(reg283[(4'h9):(1'h0)]);
                    end
                  if ({(~&(reg301[(4'hd):(3'h6)] ?
                          $signed(reg305) : forvar266))})
                    begin
                      reg334 <= {((((8'hb1) >> reg238) ^ forvar287[(3'h4):(2'h3)]) ?
                              (~&$signed(reg257)) : (+$unsigned(reg227)))};
                      reg335 <= ({$unsigned((reg207 ?
                              reg298 : reg292))} ^~ $unsigned((reg280[(3'h5):(1'h1)] ?
                          forvar238 : (forvar313 ^~ reg281))));
                      reg336 <= reg236;
                    end
                  else
                    begin
                      reg334 <= (^~($signed((!reg206)) ?
                          ($unsigned(wire198) >= (reg206 ?
                              reg312 : reg289)) : $unsigned(reg269[(1'h1):(1'h1)])));
                    end
                  if ($unsigned(($unsigned((reg242 * reg309)) != {$signed(reg276)})))
                    begin
                      reg337 <= $unsigned((reg294 < ((!wire191) < reg220[(1'h1):(1'h1)])));
                      reg338 <= reg245[(2'h2):(1'h0)];
                      reg339 <= ((~^reg295) ?
                          $signed((+reg236[(4'h8):(3'h5)])) : reg232);
                    end
                  else
                    begin
                      reg337 <= reg277[(1'h0):(1'h0)];
                      reg338 <= $unsigned(reg331);
                    end
                end
              reg340 <= (&{(reg213[(3'h5):(1'h0)] ?
                      (reg229 ? forvar249 : (8'hac)) : reg238)});
            end
        end
      if ((&((reg248 << $signed((8'ha2))) >>> (~&reg263))))
        begin
          reg341 <= $unsigned(($signed($signed(reg289)) ?
              ((reg296 || reg264) <<< reg213) : $signed((&reg259))));
          for (forvar342 = (1'h0); (forvar342 < (2'h2)); forvar342 = (forvar342 + (1'h1)))
            begin
              for (forvar343 = (1'h0); (forvar343 < (2'h3)); forvar343 = (forvar343 + (1'h1)))
                begin
                  if ((reg215 >>> $signed($signed((reg340 || forvar308)))))
                    begin
                      reg344 <= ((((reg240 <<< reg307) ?
                              (~reg205) : (reg301 ? forvar303 : reg226)) ?
                          (wire196 * $signed(forvar295)) : $signed((^~(8'ha6)))) ~^ $signed((reg213[(1'h1):(1'h1)] ?
                          $unsigned(reg273) : reg275[(3'h7):(3'h4)])));
                    end
                  else
                    begin
                      reg344 <= forvar238;
                      reg345 <= $signed(($unsigned((-reg302)) + forvar211[(2'h3):(1'h1)]));
                      reg346 <= reg205[(3'h4):(1'h0)];
                    end
                end
              for (forvar347 = (1'h0); (forvar347 < (2'h3)); forvar347 = (forvar347 + (1'h1)))
                begin
                  for (forvar348 = (1'h0); (forvar348 < (2'h2)); forvar348 = (forvar348 + (1'h1)))
                    begin
                      reg349 <= $unsigned(reg261);
                      reg350 <= $unsigned($signed((~reg349)));
                    end
                  reg351 <= ({forvar259[(1'h0):(1'h0)]} ?
                      (reg274[(1'h0):(1'h0)] ?
                          $signed($unsigned(reg208)) : $signed((reg206 < (8'ha3)))) : (~^($unsigned(reg317) ?
                          reg326[(3'h5):(3'h5)] : {(8'h9e)})));
                  reg352 <= (reg288[(4'hb):(4'hb)] ?
                      reg327[(1'h0):(1'h0)] : wire195);
                end
            end
        end
      else
        begin
          if ($unsigned($unsigned($signed((forvar315 * (8'had))))))
            begin
              for (forvar341 = (1'h0); (forvar341 < (2'h3)); forvar341 = (forvar341 + (1'h1)))
                begin
                  for (forvar342 = (1'h0); (forvar342 < (2'h2)); forvar342 = (forvar342 + (1'h1)))
                    begin
                      reg343 <= ((+reg298[(4'h9):(3'h4)]) ?
                          reg220[(2'h2):(1'h1)] : (^reg250));
                    end
                  for (forvar344 = (1'h0); (forvar344 < (1'h0)); forvar344 = (forvar344 + (1'h1)))
                    begin
                      reg345 <= $unsigned($signed($signed((8'hb1))));
                      reg346 <= (($signed((reg333 ? reg273 : reg350)) ?
                          {forvar298} : $unsigned($signed(reg212))) << $unsigned((^~(^reg296))));
                      reg347 <= $signed($unsigned((reg307[(3'h6):(3'h6)] ?
                          reg302 : reg341[(3'h5):(3'h5)])));
                    end
                  for (forvar348 = (1'h0); (forvar348 < (2'h2)); forvar348 = (forvar348 + (1'h1)))
                    begin
                      reg349 <= (~&forvar343[(3'h5):(2'h3)]);
                      reg350 <= $signed($unsigned((!$unsigned((8'haa)))));
                      reg351 <= reg272[(4'hc):(1'h0)];
                    end
                end
              for (forvar352 = (1'h0); (forvar352 < (1'h0)); forvar352 = (forvar352 + (1'h1)))
                begin
                  for (forvar353 = (1'h0); (forvar353 < (1'h0)); forvar353 = (forvar353 + (1'h1)))
                    begin
                      reg354 <= $unsigned($signed(({forvar211} ^ (reg297 == reg331))));
                      reg355 <= reg334;
                      reg356 <= $unsigned((&$unsigned((&forvar342))));
                      reg357 <= (wire192[(3'h5):(2'h2)] ?
                          {{(~reg251)}} : $signed($signed((|(8'had)))));
                    end
                end
              for (forvar358 = (1'h0); (forvar358 < (1'h0)); forvar358 = (forvar358 + (1'h1)))
                begin
                  if ((|($signed(reg331[(2'h2):(1'h0)]) << (reg305 ?
                      reg236 : reg247))))
                    begin
                      reg359 <= wire195[(3'h7):(3'h7)];
                      reg360 <= (((&{reg312}) ?
                              (reg293[(2'h2):(1'h0)] ?
                                  reg245[(1'h0):(1'h0)] : reg319[(3'h5):(2'h3)]) : reg222[(3'h7):(2'h2)]) ?
                          forvar299[(2'h2):(1'h1)] : ((^forvar249) ?
                              reg208 : (^forvar295)));
                      reg361 <= $signed((({reg355} * $signed((8'ha2))) + (8'hb2)));
                      reg362 <= forvar211;
                    end
                  else
                    begin
                      reg359 <= reg306;
                    end
                  if (((&((^reg273) * $unsigned(reg311))) ?
                      reg284 : reg210[(2'h3):(2'h2)]))
                    begin
                      reg363 <= $signed((~&$unsigned($unsigned(reg231))));
                      reg364 <= ((({reg265} >> forvar342[(4'h9):(1'h1)]) ?
                          reg249 : reg218[(2'h2):(1'h1)]) | reg339[(2'h3):(2'h3)]);
                      reg365 <= reg240;
                      reg366 <= $signed(($unsigned($unsigned(reg345)) ?
                          (reg240 ^ reg354) : $signed((reg212 ?
                              reg208 : forvar267))));
                    end
                  else
                    begin
                      reg363 <= (~$signed($unsigned(reg364[(1'h0):(1'h0)])));
                    end
                  if (({forvar299[(4'hc):(1'h1)]} ~^ $signed((~&(reg341 >>> reg300)))))
                    begin
                      reg367 <= ((reg326[(2'h2):(2'h2)] ?
                              wire200[(2'h2):(1'h0)] : (reg283[(3'h4):(2'h3)] ?
                                  (~&reg253) : (|reg236))) ?
                          reg260[(4'h8):(2'h3)] : reg259[(4'h8):(3'h7)]);
                    end
                  else
                    begin
                      reg367 <= ({reg347} ? (8'hb7) : (~|reg255));
                      reg368 <= (({{reg269}} ?
                              ((reg339 ? reg219 : (8'hb6)) ?
                                  forvar295 : {(8'had)}) : (~|(reg295 * (8'ha0)))) ?
                          reg240[(3'h4):(2'h3)] : $unsigned({forvar330[(4'h8):(3'h4)]}));
                      reg369 <= $unsigned(($signed((wire200 >> reg344)) ?
                          reg237[(2'h3):(1'h0)] : reg364[(2'h2):(2'h2)]));
                    end
                end
            end
          else
            begin
              if ({$signed($signed(((8'haf) ^ (8'ha6))))})
                begin
                  if (((~&$unsigned((reg298 ?
                      forvar344 : forvar227))) || forvar308[(2'h3):(1'h1)]))
                    begin
                      reg341 <= ((|forvar313) ?
                          reg237 : $unsigned((~|reg219[(3'h6):(2'h3)])));
                      reg342 <= $signed(({(forvar347 ? (8'hac) : reg355)} ?
                          ((reg343 ? (8'hb0) : forvar259) ?
                              forvar228[(4'hb):(2'h3)] : $signed(reg365)) : $signed((|reg253))));
                    end
                  else
                    begin
                      reg341 <= forvar211[(3'h6):(2'h3)];
                      reg342 <= $unsigned(reg207[(2'h2):(1'h0)]);
                    end
                  if ((|$signed((((8'h9e) ? (8'hb5) : reg232) ?
                      reg344 : $signed(reg338)))))
                    begin
                      reg343 <= (($unsigned(reg293[(1'h0):(1'h0)]) & $signed((reg236 != (8'haa)))) >= reg223);
                      reg344 <= ((|($unsigned(reg311) - (reg336 ?
                          forvar279 : forvar282))) > {reg300});
                      reg345 <= ((~^(^~$unsigned((8'hba)))) ?
                          {reg318} : $signed((8'h9f)));
                      reg346 <= reg299;
                    end
                  else
                    begin
                      reg343 <= {$unsigned(reg357[(4'hc):(4'h8)])};
                    end
                  if (((reg260[(4'h9):(1'h1)] < ($signed(forvar330) ?
                      forvar328 : reg296[(2'h3):(1'h0)])) != (reg368[(1'h0):(1'h0)] || {$signed(forvar287)})))
                    begin
                      reg347 <= (((!$signed(forvar244)) - (reg335 ?
                              {(8'ha4)} : (+(8'h9e)))) ?
                          forvar353 : reg268);
                      reg348 <= $signed($unsigned(((reg264 & reg318) << $unsigned(reg223))));
                    end
                  else
                    begin
                      reg347 <= $signed(reg236);
                    end
                  if (reg345[(3'h7):(3'h7)])
                    begin
                      reg349 <= reg226;
                      reg350 <= ((+$unsigned($unsigned(reg349))) ?
                          wire195 : (forvar245[(3'h4):(3'h4)] > {$signed(reg230)}));
                      reg351 <= (reg208 ^~ $signed(reg213));
                    end
                  else
                    begin
                      reg349 <= forvar330[(3'h7):(3'h5)];
                      reg350 <= reg312;
                    end
                end
              else
                begin
                  for (forvar341 = (1'h0); (forvar341 < (1'h0)); forvar341 = (forvar341 + (1'h1)))
                    begin
                      reg342 <= reg247;
                      reg343 <= (($signed((forvar341 ? reg242 : (8'hb0))) ?
                              reg208 : $unsigned(wire195)) ?
                          {reg250[(3'h4):(2'h3)]} : {$signed($signed(reg300))});
                      reg344 <= reg304;
                      reg345 <= {forvar287};
                    end
                end
              if (forvar202[(1'h1):(1'h1)])
                begin
                  if (($signed($signed(forvar282)) ^ ($unsigned(reg365[(4'h8):(3'h7)]) * $signed((8'hb2)))))
                    begin
                      reg352 <= ($unsigned(($signed(reg341) ^~ reg269)) ?
                          reg346[(1'h0):(1'h0)] : ((reg335 ?
                                  {reg270} : $unsigned(reg293)) ?
                              {$signed(wire196)} : (~|$signed(forvar348))));
                      reg353 <= $signed(reg230);
                    end
                  else
                    begin
                      reg352 <= {{(!(reg368 ? forvar238 : (8'had)))}};
                      reg353 <= forvar315;
                      reg354 <= reg323[(4'he):(4'hb)];
                    end
                  for (forvar355 = (1'h0); (forvar355 < (2'h2)); forvar355 = (forvar355 + (1'h1)))
                    begin
                      reg356 <= reg290[(3'h5):(3'h4)];
                      reg357 <= $unsigned($signed((~|(reg322 ^~ reg316))));
                      reg358 <= ($signed($unsigned($unsigned(reg356))) ?
                          {((forvar295 ? reg350 : reg233) ?
                                  (~|forvar331) : reg324[(3'h4):(2'h3)])} : {{(reg212 ?
                                      reg355 : reg291)}});
                      reg359 <= {forvar352};
                    end
                  if ((^~reg277))
                    begin
                      reg360 <= reg348;
                    end
                  else
                    begin
                      reg360 <= ((^~forvar254) ?
                          $unsigned($unsigned(forvar295[(3'h5):(3'h5)])) : $signed((~^(forvar290 ?
                              forvar287 : reg367))));
                      reg361 <= (8'ha0);
                      reg362 <= ((~&(~(forvar328 ? forvar254 : forvar330))) ?
                          ($unsigned((reg259 < forvar287)) == $unsigned((+forvar355))) : {wire191});
                      reg363 <= $unsigned((~reg272));
                    end
                  for (forvar364 = (1'h0); (forvar364 < (2'h2)); forvar364 = (forvar364 + (1'h1)))
                    begin
                      reg365 <= reg240[(3'h5):(1'h0)];
                      reg366 <= reg318;
                      reg367 <= ($unsigned((+((8'ha1) ?
                          forvar344 : wire201))) ^~ ({(~^reg360)} * reg255));
                    end
                end
              else
                begin
                  if (forvar227)
                    begin
                      reg352 <= (({reg361} ?
                          $signed($unsigned((8'h9f))) : reg298) | (^(reg301[(4'h8):(1'h0)] > {reg277})));
                      reg353 <= $unsigned($signed(((reg361 ? reg323 : reg205) ?
                          $signed(reg324) : {forvar344})));
                      reg354 <= ({wire201} <<< ((reg299[(4'h8):(3'h4)] ^ $signed((8'ha1))) ?
                          $unsigned(forvar279[(4'h8):(3'h4)]) : reg314[(2'h3):(1'h0)]));
                    end
                  else
                    begin
                      reg352 <= $unsigned((8'hb4));
                      reg353 <= reg301;
                      reg354 <= (({reg324} >>> $unsigned(wire201[(4'ha):(1'h1)])) | ((~&$signed(reg220)) - (forvar216[(1'h1):(1'h1)] ?
                          (forvar202 ? reg326 : reg229) : {reg337})));
                    end
                  for (forvar355 = (1'h0); (forvar355 < (1'h0)); forvar355 = (forvar355 + (1'h1)))
                    begin
                      reg356 <= $signed((!reg268[(3'h6):(2'h2)]));
                      reg357 <= (^~reg343);
                      reg358 <= reg290[(1'h1):(1'h0)];
                    end
                end
              for (forvar368 = (1'h0); (forvar368 < (1'h0)); forvar368 = (forvar368 + (1'h1)))
                begin
                  for (forvar369 = (1'h0); (forvar369 < (2'h2)); forvar369 = (forvar369 + (1'h1)))
                    begin
                      reg370 <= reg363;
                      reg371 <= $signed((^~$unsigned($unsigned(reg346))));
                      reg372 <= $signed(reg369);
                      reg373 <= forvar331[(1'h0):(1'h0)];
                    end
                  for (forvar374 = (1'h0); (forvar374 < (1'h0)); forvar374 = (forvar374 + (1'h1)))
                    begin
                      reg375 <= $unsigned((8'h9c));
                      reg376 <= (!(8'hb3));
                    end
                  for (forvar377 = (1'h0); (forvar377 < (2'h2)); forvar377 = (forvar377 + (1'h1)))
                    begin
                      reg378 <= forvar295[(3'h6):(3'h4)];
                    end
                end
              reg379 <= reg258[(1'h0):(1'h0)];
            end
          for (forvar380 = (1'h0); (forvar380 < (1'h1)); forvar380 = (forvar380 + (1'h1)))
            begin
              for (forvar381 = (1'h0); (forvar381 < (2'h3)); forvar381 = (forvar381 + (1'h1)))
                begin
                  for (forvar382 = (1'h0); (forvar382 < (1'h1)); forvar382 = (forvar382 + (1'h1)))
                    begin
                      reg383 <= ((~&$unsigned((reg331 ?
                          (8'hb8) : reg253))) + {$signed({reg376})});
                      reg384 <= ($signed((~&(reg317 << forvar217))) ?
                          (8'ha2) : reg327);
                    end
                  reg385 <= $signed($unsigned(reg273));
                  for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
                    begin
                      reg387 <= $unsigned((reg314[(1'h1):(1'h1)] ?
                          (reg253 | (reg229 | reg256)) : (forvar295 << forvar261[(2'h3):(1'h1)])));
                      reg388 <= $signed($signed($signed((^~forvar279))));
                    end
                  for (forvar389 = (1'h0); (forvar389 < (2'h2)); forvar389 = (forvar389 + (1'h1)))
                    begin
                      reg390 <= $signed(forvar267);
                    end
                end
              if (($unsigned((~|(reg252 ?
                  reg302 : (8'hac)))) << {$signed($signed(reg278))}))
                begin
                  if ($signed((~|reg348)))
                    begin
                      reg391 <= ((-($signed(forvar266) ?
                              forvar358[(1'h0):(1'h0)] : $unsigned((8'hb3)))) ?
                          $unsigned(reg265) : (~|(^{reg318})));
                      reg392 <= reg202;
                      reg393 <= reg305;
                    end
                  else
                    begin
                      reg391 <= reg379[(1'h1):(1'h0)];
                      reg392 <= ($unsigned($signed($signed((8'h9c)))) ?
                          wire196 : ((-reg242) ?
                              $unsigned($unsigned((8'ha8))) : reg261[(4'ha):(1'h0)]));
                      reg393 <= (($unsigned(((8'hb1) <= forvar261)) + (reg239[(2'h2):(2'h2)] ?
                              $unsigned((8'hb8)) : (&reg272))) ?
                          (reg344[(3'h6):(1'h1)] <= (~&$signed(forvar238))) : ((~((8'hb4) ?
                                  reg240 : (8'h9e))) ?
                              $unsigned((reg288 >>> reg296)) : forvar342[(4'hc):(3'h7)]));
                    end
                  for (forvar394 = (1'h0); (forvar394 < (1'h0)); forvar394 = (forvar394 + (1'h1)))
                    begin
                      reg395 <= $unsigned({(+$signed(reg235))});
                    end
                end
              else
                begin
                  if (((($unsigned(reg363) ?
                          reg295[(4'ha):(3'h4)] : (8'h9e)) - (reg307[(3'h6):(2'h2)] ?
                          {reg226} : $signed((8'ha3)))) ?
                      {(~|(reg318 * reg309))} : $signed(reg391)))
                    begin
                      reg391 <= {(reg219 == $signed(forvar244))};
                      reg392 <= reg252[(4'h8):(3'h5)];
                    end
                  else
                    begin
                      reg391 <= reg384[(3'h4):(1'h0)];
                      reg392 <= forvar282;
                      reg393 <= (8'haa);
                    end
                end
              for (forvar396 = (1'h0); (forvar396 < (1'h0)); forvar396 = (forvar396 + (1'h1)))
                begin
                  for (forvar397 = (1'h0); (forvar397 < (1'h1)); forvar397 = (forvar397 + (1'h1)))
                    begin
                      reg398 <= $unsigned($signed((!reg368[(1'h1):(1'h0)])));
                    end
                end
            end
          for (forvar399 = (1'h0); (forvar399 < (2'h2)); forvar399 = (forvar399 + (1'h1)))
            begin
              for (forvar400 = (1'h0); (forvar400 < (1'h0)); forvar400 = (forvar400 + (1'h1)))
                begin
                  reg401 <= reg356[(3'h5):(1'h1)];
                  reg402 <= $signed((forvar266[(4'hc):(2'h2)] ?
                      reg356[(2'h3):(1'h0)] : (reg316 ?
                          (+reg289) : $unsigned(reg319))));
                  for (forvar403 = (1'h0); (forvar403 < (1'h1)); forvar403 = (forvar403 + (1'h1)))
                    begin
                      reg404 <= (&(reg272[(3'h7):(2'h2)] + ((8'hae) ?
                          reg343 : (reg373 ? forvar234 : forvar369))));
                      reg405 <= $signed($unsigned((+(reg252 ?
                          reg225 : forvar293))));
                      reg406 <= $signed(forvar396[(3'h4):(1'h0)]);
                      reg407 <= (!$unsigned($signed((reg237 < reg213))));
                    end
                  if ($signed($signed({((8'hb8) ? reg227 : forvar241)})))
                    begin
                      reg408 <= $signed((!(~^$signed(forvar315))));
                      reg409 <= ((8'hb4) && (&forvar358));
                      reg410 <= $unsigned(reg352);
                    end
                  else
                    begin
                      reg408 <= $signed($signed($signed($unsigned(reg264))));
                    end
                end
            end
        end
      for (forvar411 = (1'h0); (forvar411 < (2'h3)); forvar411 = (forvar411 + (1'h1)))
        begin
          for (forvar412 = (1'h0); (forvar412 < (1'h1)); forvar412 = (forvar412 + (1'h1)))
            begin
              reg413 <= reg214[(3'h5):(1'h1)];
              for (forvar414 = (1'h0); (forvar414 < (2'h3)); forvar414 = (forvar414 + (1'h1)))
                begin
                  reg415 <= reg358[(2'h3):(2'h3)];
                end
              for (forvar416 = (1'h0); (forvar416 < (2'h3)); forvar416 = (forvar416 + (1'h1)))
                begin
                  if (reg259[(2'h3):(1'h1)])
                    begin
                      reg417 <= $signed($signed(reg208));
                      reg418 <= (~&reg243);
                      reg419 <= (8'had);
                      reg420 <= (forvar227[(4'hb):(1'h1)] < forvar287);
                    end
                  else
                    begin
                      reg417 <= forvar244[(4'hb):(4'h8)];
                      reg418 <= (!reg334[(2'h2):(1'h0)]);
                      reg419 <= (reg352[(4'hb):(4'h9)] >> (((forvar244 ?
                                  reg213 : reg358) ?
                              (reg208 == reg372) : (8'ha1)) ?
                          $unsigned(reg375[(1'h1):(1'h0)]) : reg350));
                    end
                  for (forvar421 = (1'h0); (forvar421 < (2'h2)); forvar421 = (forvar421 + (1'h1)))
                    begin
                      reg422 <= {($signed((!reg291)) | reg343[(1'h0):(1'h0)])};
                      reg423 <= (($unsigned((!reg310)) ?
                          reg314[(1'h1):(1'h1)] : (&$signed(forvar331))) == reg307[(3'h5):(3'h5)]);
                      reg424 <= $signed(({$unsigned(reg336)} - $unsigned(reg226[(1'h1):(1'h1)])));
                      reg425 <= reg262[(4'ha):(4'ha)];
                    end
                end
            end
          reg426 <= forvar352;
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module23
#(parameter param185 = {(8'hb4)})
(y, clk, wire28, wire27, wire26, wire25, wire24);
  output wire [(32'h63f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire28;
  input wire [(4'hb):(1'h0)] wire27;
  input wire [(4'ha):(1'h0)] wire26;
  input wire signed [(4'hf):(1'h0)] wire25;
  input wire signed [(4'h9):(1'h0)] wire24;
  wire signed [(3'h4):(1'h0)] wire184;
  wire signed [(4'hf):(1'h0)] wire183;
  wire signed [(4'hd):(1'h0)] wire182;
  reg [(4'hc):(1'h0)] reg181 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg180 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg179 = (1'h0);
  reg [(4'he):(1'h0)] reg178 = (1'h0);
  reg [(4'ha):(1'h0)] reg177 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar176 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg175 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg174 = (1'h0);
  reg [(3'h5):(1'h0)] forvar173 = (1'h0);
  reg [(4'hb):(1'h0)] reg172 = (1'h0);
  reg [(4'he):(1'h0)] reg171 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg170 = (1'h0);
  reg [(4'hc):(1'h0)] reg169 = (1'h0);
  reg [(4'h9):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg [(3'h4):(1'h0)] reg165 = (1'h0);
  reg [(4'h8):(1'h0)] forvar164 = (1'h0);
  reg [(4'hc):(1'h0)] reg163 = (1'h0);
  reg [(4'ha):(1'h0)] reg162 = (1'h0);
  reg [(4'h8):(1'h0)] reg161 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg160 = (1'h0);
  reg [(3'h6):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar158 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg157 = (1'h0);
  reg signed [(4'he):(1'h0)] reg156 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg155 = (1'h0);
  reg signed [(4'he):(1'h0)] reg154 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar152 = (1'h0);
  reg [(3'h5):(1'h0)] reg150 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg153 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg152 = (1'h0);
  reg [(5'h10):(1'h0)] reg151 = (1'h0);
  reg [(4'hb):(1'h0)] forvar150 = (1'h0);
  reg [(4'hb):(1'h0)] forvar149 = (1'h0);
  reg [(2'h2):(1'h0)] reg148 = (1'h0);
  reg [(3'h5):(1'h0)] forvar147 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg146 = (1'h0);
  reg [(4'hd):(1'h0)] reg145 = (1'h0);
  reg [(4'h8):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg143 = (1'h0);
  reg [(3'h5):(1'h0)] reg142 = (1'h0);
  reg [(3'h6):(1'h0)] forvar141 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg140 = (1'h0);
  reg [(3'h5):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg138 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg137 = (1'h0);
  reg [(4'he):(1'h0)] reg132 = (1'h0);
  reg [(4'hb):(1'h0)] reg136 = (1'h0);
  reg [(3'h6):(1'h0)] reg135 = (1'h0);
  reg signed [(4'he):(1'h0)] reg134 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar132 = (1'h0);
  reg [(3'h7):(1'h0)] reg131 = (1'h0);
  reg [(5'h10):(1'h0)] forvar130 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg129 = (1'h0);
  reg [(3'h7):(1'h0)] reg128 = (1'h0);
  reg [(4'hd):(1'h0)] reg127 = (1'h0);
  reg [(4'hd):(1'h0)] reg126 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg125 = (1'h0);
  reg [(4'ha):(1'h0)] reg124 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg123 = (1'h0);
  reg signed [(4'he):(1'h0)] reg122 = (1'h0);
  reg [(5'h10):(1'h0)] forvar121 = (1'h0);
  reg [(2'h2):(1'h0)] reg120 = (1'h0);
  reg [(3'h5):(1'h0)] reg119 = (1'h0);
  reg [(3'h7):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg117 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg116 = (1'h0);
  reg [(4'ha):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg114 = (1'h0);
  reg [(5'h10):(1'h0)] reg113 = (1'h0);
  reg [(3'h7):(1'h0)] reg112 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar109 = (1'h0);
  reg [(4'h9):(1'h0)] reg111 = (1'h0);
  reg [(4'hf):(1'h0)] reg110 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg108 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg107 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar106 = (1'h0);
  reg [(4'he):(1'h0)] forvar105 = (1'h0);
  reg signed [(4'he):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg103 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar100 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg100 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar99 = (1'h0);
  wire signed [(4'he):(1'h0)] wire98;
  wire signed [(2'h2):(1'h0)] wire97;
  reg [(2'h3):(1'h0)] reg96 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg95 = (1'h0);
  reg [(4'he):(1'h0)] forvar94 = (1'h0);
  reg [(4'hd):(1'h0)] forvar93 = (1'h0);
  reg [(4'h8):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg91 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg90 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar89 = (1'h0);
  reg [(4'ha):(1'h0)] reg88 = (1'h0);
  reg [(4'h9):(1'h0)] reg87 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg86 = (1'h0);
  reg [(4'h8):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg84 = (1'h0);
  reg [(3'h7):(1'h0)] reg83 = (1'h0);
  reg [(4'he):(1'h0)] reg82 = (1'h0);
  reg [(3'h5):(1'h0)] reg81 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar80 = (1'h0);
  reg [(4'he):(1'h0)] reg79 = (1'h0);
  reg [(3'h4):(1'h0)] reg78 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg77 = (1'h0);
  reg [(3'h6):(1'h0)] reg76 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar75 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar74 = (1'h0);
  reg [(2'h3):(1'h0)] reg73 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar72 = (1'h0);
  reg [(4'hd):(1'h0)] reg71 = (1'h0);
  reg [(3'h7):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg69 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg68 = (1'h0);
  reg [(3'h7):(1'h0)] forvar67 = (1'h0);
  reg [(4'hb):(1'h0)] forvar63 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg67 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg66 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg65 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg64 = (1'h0);
  reg [(4'ha):(1'h0)] reg63 = (1'h0);
  reg [(4'hd):(1'h0)] reg62 = (1'h0);
  reg [(4'he):(1'h0)] reg61 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg60 = (1'h0);
  reg [(5'h10):(1'h0)] forvar59 = (1'h0);
  reg [(3'h7):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg57 = (1'h0);
  reg [(4'hd):(1'h0)] reg56 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg55 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar54 = (1'h0);
  reg [(4'hc):(1'h0)] reg53 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg52 = (1'h0);
  reg [(4'hf):(1'h0)] reg51 = (1'h0);
  reg [(2'h2):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar47 = (1'h0);
  reg [(4'h9):(1'h0)] reg49 = (1'h0);
  reg [(4'hb):(1'h0)] reg48 = (1'h0);
  reg [(2'h3):(1'h0)] reg47 = (1'h0);
  reg [(3'h5):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg45 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg44 = (1'h0);
  reg [(4'hc):(1'h0)] reg43 = (1'h0);
  reg signed [(4'he):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg41 = (1'h0);
  reg [(4'h8):(1'h0)] reg40 = (1'h0);
  reg [(4'he):(1'h0)] forvar39 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar38 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar37 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar36 = (1'h0);
  wire [(4'he):(1'h0)] wire35;
  wire [(2'h2):(1'h0)] wire34;
  wire signed [(4'h9):(1'h0)] wire33;
  wire signed [(4'hd):(1'h0)] wire32;
  wire [(4'hc):(1'h0)] wire31;
  wire signed [(3'h5):(1'h0)] wire30;
  wire [(4'hc):(1'h0)] wire29;
  assign y = {wire184,
                 wire183,
                 wire182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 forvar176,
                 reg175,
                 reg174,
                 forvar173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 forvar164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 forvar158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 forvar152,
                 reg150,
                 reg153,
                 reg152,
                 reg151,
                 forvar150,
                 forvar149,
                 reg148,
                 forvar147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 forvar141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg132,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 forvar132,
                 reg131,
                 forvar130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 forvar121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 forvar109,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 forvar106,
                 forvar105,
                 reg104,
                 reg103,
                 reg102,
                 forvar100,
                 reg101,
                 reg100,
                 forvar99,
                 wire98,
                 wire97,
                 reg96,
                 reg95,
                 forvar94,
                 forvar93,
                 reg92,
                 reg91,
                 reg90,
                 forvar89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 forvar80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 forvar75,
                 forvar74,
                 reg73,
                 forvar72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 forvar67,
                 forvar63,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 forvar59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 forvar54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 forvar47,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 forvar39,
                 forvar38,
                 forvar37,
                 forvar36,
                 wire35,
                 wire34,
                 wire33,
                 wire32,
                 wire31,
                 wire30,
                 wire29,
                 (1'h0)};
  assign wire29 = ($unsigned(wire27[(2'h3):(2'h2)]) > (8'ha7));
  assign wire30 = ($signed(wire29[(2'h3):(1'h0)]) ?
                      $signed((wire27 == (~|wire29))) : (wire27[(3'h6):(3'h4)] ?
                          (wire24 ?
                              wire24[(1'h1):(1'h1)] : wire27[(4'h9):(4'h9)]) : ((wire27 ?
                                  wire25 : wire26) ?
                              wire29[(4'ha):(4'h8)] : $unsigned(wire28))));
  assign wire31 = (((wire30[(3'h4):(2'h2)] == (8'h9c)) ?
                      $unsigned($signed(wire29)) : $signed(wire25[(4'hf):(4'ha)])) ^ wire29[(4'h9):(4'h8)]);
  assign wire32 = wire31;
  assign wire33 = wire30[(2'h2):(1'h1)];
  assign wire34 = (-wire33);
  assign wire35 = ({wire34} < wire25);
  always
    @(posedge clk) begin
      for (forvar36 = (1'h0); (forvar36 < (2'h3)); forvar36 = (forvar36 + (1'h1)))
        begin
          for (forvar37 = (1'h0); (forvar37 < (2'h2)); forvar37 = (forvar37 + (1'h1)))
            begin
              for (forvar38 = (1'h0); (forvar38 < (2'h3)); forvar38 = (forvar38 + (1'h1)))
                begin
                  for (forvar39 = (1'h0); (forvar39 < (2'h3)); forvar39 = (forvar39 + (1'h1)))
                    begin
                      reg40 <= (~^wire33);
                    end
                  if (wire24)
                    begin
                      reg41 <= (^(~&$signed(((8'h9d) > (8'ha9)))));
                      reg42 <= (^wire35[(4'he):(4'ha)]);
                    end
                  else
                    begin
                      reg41 <= (+(~&({forvar36} ?
                          (wire32 && forvar36) : (8'h9c))));
                      reg42 <= wire29;
                      reg43 <= $signed((($unsigned(wire35) ?
                          $signed(reg40) : (wire27 ?
                              (8'ha4) : (8'hb5))) <= (forvar37[(2'h3):(2'h2)] > (wire26 + wire30))));
                      reg44 <= ($signed((reg43 ? (~&wire32) : {wire28})) ?
                          forvar37[(4'ha):(4'h8)] : (~^forvar39[(3'h4):(1'h0)]));
                    end
                  if (($signed(($unsigned((8'hb4)) ?
                          $signed(forvar39) : forvar37[(3'h5):(3'h4)])) ?
                      ($unsigned($signed(reg42)) ?
                          wire28[(2'h3):(2'h2)] : wire24) : ((&(forvar36 ?
                          wire31 : (8'h9f))) <= ((~&wire26) ~^ reg44))))
                    begin
                      reg45 <= $signed($unsigned((^~(|wire32))));
                      reg46 <= wire25;
                    end
                  else
                    begin
                      reg45 <= $unsigned($unsigned(((&forvar39) ?
                          $unsigned(wire26) : (^reg42))));
                      reg46 <= $signed($signed((forvar39 ~^ (reg45 ?
                          reg40 : wire33))));
                    end
                end
              if (({wire27} ^ wire24[(3'h5):(1'h1)]))
                begin
                  if ($signed(forvar39[(2'h2):(2'h2)]))
                    begin
                      reg47 <= (&((reg41[(4'hb):(4'ha)] ?
                          {reg44} : reg44[(3'h7):(3'h6)]) < {(&wire28)}));
                      reg48 <= $signed(wire25);
                      reg49 <= (wire26 > $signed({(^reg46)}));
                    end
                  else
                    begin
                      reg47 <= $signed((~|forvar39[(4'h9):(3'h4)]));
                      reg48 <= forvar37[(1'h1):(1'h0)];
                    end
                end
              else
                begin
                  for (forvar47 = (1'h0); (forvar47 < (2'h3)); forvar47 = (forvar47 + (1'h1)))
                    begin
                      reg48 <= ($unsigned($signed(wire26)) ?
                          (~&(^((8'ha6) ? wire35 : wire33))) : wire26);
                      reg49 <= wire24;
                      reg50 <= $signed(($unsigned((wire29 >= (8'hb4))) + forvar39[(1'h1):(1'h0)]));
                      reg51 <= (^~(^$unsigned($unsigned((8'ha2)))));
                    end
                  if (wire33[(3'h7):(2'h2)])
                    begin
                      reg52 <= $signed(wire26[(2'h2):(1'h0)]);
                    end
                  else
                    begin
                      reg52 <= $unsigned((~({wire24} <<< reg45[(2'h2):(1'h0)])));
                      reg53 <= reg46;
                    end
                end
              for (forvar54 = (1'h0); (forvar54 < (1'h1)); forvar54 = (forvar54 + (1'h1)))
                begin
                  reg55 <= {reg52[(4'h9):(1'h0)]};
                  if ((&(reg42[(3'h4):(2'h3)] <= $unsigned(((8'hb7) ^ reg53)))))
                    begin
                      reg56 <= $signed({((!reg46) << $unsigned(wire33))});
                      reg57 <= ($signed($unsigned((wire35 ?
                          reg48 : reg48))) || ($unsigned((wire34 - reg41)) ?
                          reg46[(3'h5):(2'h2)] : ((&reg53) ?
                              (^reg55) : (reg45 ? (8'ha4) : wire34))));
                      reg58 <= (~|{reg53[(1'h1):(1'h1)]});
                    end
                  else
                    begin
                      reg56 <= (((^~{wire31}) * $signed($signed(reg42))) ?
                          reg42[(3'h5):(1'h0)] : reg53);
                      reg57 <= $unsigned($signed(((~^wire25) ?
                          {(8'ha4)} : $signed(forvar37))));
                      reg58 <= {(reg41 ?
                              ((8'ha9) ? reg45 : {(8'ha4)}) : {reg44})};
                    end
                  for (forvar59 = (1'h0); (forvar59 < (2'h3)); forvar59 = (forvar59 + (1'h1)))
                    begin
                      reg60 <= (((~|$signed(wire25)) ?
                          {$signed(reg50)} : wire25[(3'h5):(3'h5)]) | (~&reg56));
                      reg61 <= ($signed((~|(+(8'had)))) * (((forvar39 != reg49) ?
                              (forvar47 ? wire24 : reg60) : reg50) ?
                          reg48 : forvar39[(4'hb):(2'h3)]));
                      reg62 <= reg53[(3'h4):(2'h3)];
                    end
                end
              if ($unsigned(reg41[(3'h6):(1'h1)]))
                begin
                  reg63 <= (&$unsigned(($signed(wire35) ?
                      (|reg55) : $signed(reg61))));
                  if (reg55[(1'h1):(1'h0)])
                    begin
                      reg64 <= $unsigned(reg43[(4'ha):(4'ha)]);
                      reg65 <= (~^(reg63 <<< ($unsigned((8'hb8)) ?
                          $signed(reg42) : (wire33 ? reg45 : wire24))));
                    end
                  else
                    begin
                      reg64 <= wire31[(2'h2):(1'h1)];
                      reg65 <= ($unsigned(reg48[(3'h6):(2'h3)]) ?
                          reg48 : wire30);
                      reg66 <= $signed($signed((&$signed(wire28))));
                    end
                  reg67 <= $unsigned({$unsigned((!forvar37))});
                end
              else
                begin
                  for (forvar63 = (1'h0); (forvar63 < (2'h2)); forvar63 = (forvar63 + (1'h1)))
                    begin
                      reg64 <= reg49[(2'h2):(1'h0)];
                      reg65 <= reg46[(1'h1):(1'h0)];
                      reg66 <= forvar39[(4'hc):(1'h0)];
                    end
                  for (forvar67 = (1'h0); (forvar67 < (1'h1)); forvar67 = (forvar67 + (1'h1)))
                    begin
                      reg68 <= $unsigned((reg57[(2'h3):(1'h1)] ?
                          $unsigned(reg58) : reg46));
                      reg69 <= (8'ha1);
                      reg70 <= wire24;
                    end
                end
            end
          reg71 <= $unsigned(((~reg45) << $signed((!reg42))));
          for (forvar72 = (1'h0); (forvar72 < (1'h0)); forvar72 = (forvar72 + (1'h1)))
            begin
              reg73 <= (wire31 && reg70[(2'h3):(1'h0)]);
              for (forvar74 = (1'h0); (forvar74 < (1'h0)); forvar74 = (forvar74 + (1'h1)))
                begin
                  for (forvar75 = (1'h0); (forvar75 < (2'h2)); forvar75 = (forvar75 + (1'h1)))
                    begin
                      reg76 <= reg56;
                      reg77 <= $signed({(reg68[(2'h3):(2'h3)] ?
                              $unsigned(wire32) : wire25)});
                      reg78 <= ((&$unsigned((|forvar38))) ?
                          wire31[(4'h9):(3'h5)] : $unsigned(((8'ha7) ?
                              {wire25} : $unsigned((8'hba)))));
                      reg79 <= (reg51 && reg69);
                    end
                  for (forvar80 = (1'h0); (forvar80 < (2'h3)); forvar80 = (forvar80 + (1'h1)))
                    begin
                      reg81 <= $signed({forvar39});
                      reg82 <= ((|reg50) ?
                          (-reg77) : (($signed(reg55) ?
                                  wire35 : (forvar59 - (8'ha6))) ?
                              (+((8'h9e) && reg50)) : (forvar37 ?
                                  reg47[(2'h3):(1'h0)] : $signed(reg44))));
                      reg83 <= reg40;
                      reg84 <= {(&$unsigned((~^reg73)))};
                    end
                  if ((reg66[(2'h2):(1'h1)] << wire24[(3'h4):(2'h2)]))
                    begin
                      reg85 <= ($signed((+(reg67 ?
                          reg51 : reg65))) && (~^wire27));
                      reg86 <= $signed((~|reg43));
                      reg87 <= reg50;
                      reg88 <= $signed($signed(wire24));
                    end
                  else
                    begin
                      reg85 <= reg71[(3'h4):(2'h2)];
                      reg86 <= ((^~$unsigned($signed((8'ha2)))) ?
                          reg86[(2'h2):(1'h1)] : (($unsigned(reg88) ?
                              (forvar39 ~^ (8'ha0)) : $unsigned((8'hac))) > $unsigned($signed(reg73))));
                    end
                  for (forvar89 = (1'h0); (forvar89 < (2'h2)); forvar89 = (forvar89 + (1'h1)))
                    begin
                      reg90 <= $signed($unsigned(reg77));
                      reg91 <= ((|$signed(wire29[(4'h8):(1'h0)])) ?
                          $unsigned(reg57) : ({(forvar75 ?
                                  reg70 : forvar39)} || ((|wire27) ?
                              (forvar72 || forvar74) : (forvar38 ^~ reg45))));
                    end
                end
              reg92 <= (8'h9d);
              for (forvar93 = (1'h0); (forvar93 < (2'h2)); forvar93 = (forvar93 + (1'h1)))
                begin
                  for (forvar94 = (1'h0); (forvar94 < (1'h0)); forvar94 = (forvar94 + (1'h1)))
                    begin
                      reg95 <= reg91;
                      reg96 <= ({(((8'ha9) ? reg81 : reg67) ?
                              (~reg76) : (^(8'haf)))} == reg61[(3'h7):(1'h0)]);
                    end
                end
            end
        end
    end
  assign wire97 = $signed(forvar72[(3'h7):(1'h0)]);
  assign wire98 = {reg40[(3'h4):(2'h3)]};
  always
    @(posedge clk) begin
      for (forvar99 = (1'h0); (forvar99 < (2'h2)); forvar99 = (forvar99 + (1'h1)))
        begin
          if (((~|{wire34[(1'h1):(1'h0)]}) != $unsigned($unsigned((+reg57)))))
            begin
              reg100 <= (+reg90[(3'h5):(1'h1)]);
            end
          else
            begin
              if ((~^forvar93[(3'h7):(3'h4)]))
                begin
                  reg100 <= $unsigned(((-$unsigned(reg47)) ^~ (^(wire26 > reg84))));
                  reg101 <= (wire34[(1'h0):(1'h0)] ^ (($signed(wire34) ?
                          $signed(reg53) : {forvar89}) ?
                      wire98 : reg44[(2'h3):(1'h1)]));
                end
              else
                begin
                  for (forvar100 = (1'h0); (forvar100 < (2'h2)); forvar100 = (forvar100 + (1'h1)))
                    begin
                      reg101 <= (reg68 + $signed(({(8'ha4)} ?
                          (forvar38 >>> reg68) : $signed(reg81))));
                      reg102 <= reg73;
                      reg103 <= {(((^reg85) ?
                                  {forvar54} : reg55[(3'h6):(1'h0)]) ?
                              {{reg70}} : (~&reg47[(1'h0):(1'h0)]))};
                      reg104 <= $unsigned(reg70);
                    end
                end
              for (forvar105 = (1'h0); (forvar105 < (1'h1)); forvar105 = (forvar105 + (1'h1)))
                begin
                  for (forvar106 = (1'h0); (forvar106 < (2'h2)); forvar106 = (forvar106 + (1'h1)))
                    begin
                      reg107 <= ($signed(wire24[(4'h9):(2'h3)]) == forvar39[(4'hb):(4'h9)]);
                      reg108 <= ({{(reg58 ? reg61 : forvar63)}} ?
                          $signed($unsigned($unsigned(reg53))) : $unsigned(reg83[(3'h6):(2'h2)]));
                    end
                end
              if (reg90)
                begin
                  if (reg67[(3'h4):(1'h1)])
                    begin
                      reg109 <= wire24[(4'h8):(2'h2)];
                      reg110 <= $unsigned((reg103[(2'h3):(2'h2)] && ((&forvar80) <= $unsigned(forvar93))));
                      reg111 <= ($signed($signed((+reg79))) ?
                          ($signed((reg100 ?
                              wire25 : wire29)) ^~ {((8'hb6) << reg90)}) : $signed(({forvar74} <<< ((8'hae) ?
                              reg103 : forvar80))));
                    end
                  else
                    begin
                      reg109 <= $signed(reg79[(1'h0):(1'h0)]);
                      reg110 <= $signed(($unsigned(reg56[(4'h9):(3'h6)]) ?
                          ($unsigned(wire35) << (forvar80 ?
                              reg104 : forvar74)) : {$unsigned(reg49)}));
                      reg111 <= $unsigned(forvar105[(3'h7):(1'h1)]);
                    end
                end
              else
                begin
                  for (forvar109 = (1'h0); (forvar109 < (2'h3)); forvar109 = (forvar109 + (1'h1)))
                    begin
                      reg110 <= $signed(wire31);
                      reg111 <= (^~(~|$signed($unsigned(reg40))));
                      reg112 <= {$unsigned(reg57[(1'h1):(1'h0)])};
                      reg113 <= forvar94;
                    end
                  if (reg58[(3'h5):(2'h3)])
                    begin
                      reg114 <= $signed((~(~^{(8'hb2)})));
                      reg115 <= (8'hba);
                    end
                  else
                    begin
                      reg114 <= $signed({$signed(reg69[(3'h5):(2'h3)])});
                      reg115 <= wire29;
                      reg116 <= (!reg100);
                      reg117 <= {$signed((reg71[(2'h2):(2'h2)] ?
                              {forvar47} : reg88[(1'h1):(1'h0)]))};
                    end
                end
            end
          reg118 <= $signed({(~{(8'hb8)})});
          if ({reg91})
            begin
              reg119 <= reg50;
            end
          else
            begin
              if (wire33[(1'h1):(1'h1)])
                begin
                  if (((^~reg117[(3'h7):(2'h3)]) & {((wire34 * wire31) <= $signed(forvar109))}))
                    begin
                      reg119 <= ($unsigned((reg77 ?
                          (reg114 > reg83) : $signed(reg65))) <= $signed((wire26 ?
                          reg79[(4'h9):(3'h7)] : reg51[(4'hc):(3'h7)])));
                    end
                  else
                    begin
                      reg119 <= (~|{{forvar37[(2'h2):(1'h1)]}});
                    end
                end
              else
                begin
                  reg119 <= wire35[(3'h5):(1'h1)];
                  reg120 <= ($unsigned({(reg90 ? forvar105 : forvar80)}) ?
                      reg73[(1'h0):(1'h0)] : $signed((+reg116)));
                  for (forvar121 = (1'h0); (forvar121 < (1'h0)); forvar121 = (forvar121 + (1'h1)))
                    begin
                      reg122 <= (((8'hb7) ?
                              $unsigned($unsigned(wire25)) : (reg76 * reg117[(3'h4):(1'h1)])) ?
                          {((reg42 ? reg115 : reg77) ?
                                  (reg120 ?
                                      reg112 : reg60) : $unsigned(reg79))} : ($signed((~^reg91)) != $signed($signed(forvar89))));
                      reg123 <= reg103;
                      reg124 <= {(reg90 ?
                              {(reg115 <<< forvar93)} : ({reg119} + reg48))};
                      reg125 <= forvar39;
                    end
                  if (reg91)
                    begin
                      reg126 <= (($signed($unsigned(reg52)) - reg60[(1'h0):(1'h0)]) ?
                          (($signed(reg44) ?
                                  (wire25 ? reg90 : reg65) : forvar36) ?
                              (^reg44) : (!forvar75[(3'h6):(2'h2)])) : (~|reg87));
                      reg127 <= $signed($unsigned(reg120[(1'h0):(1'h0)]));
                    end
                  else
                    begin
                      reg126 <= (wire98[(1'h0):(1'h0)] ^~ ((~^(reg78 - wire97)) ?
                          $unsigned($signed(reg104)) : ((forvar100 ^ reg84) ?
                              reg68 : (forvar99 ? reg56 : reg83))));
                      reg127 <= (+(((forvar93 ? wire29 : (8'ha7)) != (reg63 ?
                          (8'hb8) : reg63)) <= $unsigned(((8'ha4) ?
                          reg56 : forvar39))));
                      reg128 <= (~&$signed(((reg87 ?
                          forvar121 : reg42) * (reg107 ? wire31 : wire25))));
                      reg129 <= ($signed($unsigned($unsigned(forvar99))) - wire32[(3'h5):(2'h3)]);
                    end
                end
              if (reg115)
                begin
                  for (forvar130 = (1'h0); (forvar130 < (2'h2)); forvar130 = (forvar130 + (1'h1)))
                    begin
                      reg131 <= {$unsigned(((^~reg122) != {wire34}))};
                    end
                  for (forvar132 = (1'h0); (forvar132 < (2'h3)); forvar132 = (forvar132 + (1'h1)))
                    begin
                      reg133 <= (reg71 ?
                          $signed(reg61[(4'hc):(2'h2)]) : $signed(wire34));
                      reg134 <= $unsigned(reg50[(2'h2):(1'h0)]);
                      reg135 <= (~|reg50);
                      reg136 <= forvar132;
                    end
                end
              else
                begin
                  for (forvar130 = (1'h0); (forvar130 < (2'h2)); forvar130 = (forvar130 + (1'h1)))
                    begin
                      reg131 <= (^reg111);
                      reg132 <= ({$signed(reg83)} > ((-$unsigned(reg116)) ?
                          $signed(reg113[(4'ha):(1'h1)]) : (8'ha0)));
                      reg133 <= $unsigned(($signed(((8'had) >> reg111)) ?
                          {(reg129 == reg112)} : (!(reg131 >>> forvar36))));
                      reg134 <= $signed({{$unsigned(reg136)}});
                    end
                  if ($signed((8'h9c)))
                    begin
                      reg135 <= ($unsigned(reg95) ? reg110 : (8'hb2));
                      reg136 <= (-($unsigned((~(8'ha4))) ?
                          ({(8'had)} >> {wire98}) : ((forvar39 ^ wire27) << (|(8'hb3)))));
                    end
                  else
                    begin
                      reg135 <= $signed(($unsigned((reg53 <<< wire24)) | (reg101[(4'ha):(3'h7)] == (!forvar105))));
                      reg136 <= $unsigned(($unsigned(reg48) ?
                          (reg95[(1'h1):(1'h0)] ?
                              (reg52 ?
                                  (8'ha7) : reg57) : forvar89) : forvar67));
                      reg137 <= $unsigned($signed(reg77[(1'h0):(1'h0)]));
                    end
                  if (wire33)
                    begin
                      reg138 <= (~&($signed((~reg129)) ?
                          ($signed((8'hb2)) ?
                              (reg132 ?
                                  (8'hb5) : reg133) : $unsigned(reg132)) : (~^reg42[(3'h6):(3'h4)])));
                    end
                  else
                    begin
                      reg138 <= wire97;
                      reg139 <= ((8'h9e) + (($signed(reg101) >= $signed(forvar130)) || (reg67 & $unsigned(reg135))));
                      reg140 <= (reg111 ?
                          reg125[(1'h0):(1'h0)] : (forvar63[(3'h4):(2'h3)] > ($signed(reg112) - (-reg65))));
                    end
                  for (forvar141 = (1'h0); (forvar141 < (2'h2)); forvar141 = (forvar141 + (1'h1)))
                    begin
                      reg142 <= ($signed((reg107 - wire28[(1'h0):(1'h0)])) || {$signed((~(8'ha9)))});
                      reg143 <= $signed((!(!((8'hb1) + (8'hab)))));
                      reg144 <= ($signed(reg137) + $signed(($unsigned((8'hb0)) << reg126[(4'h8):(3'h7)])));
                    end
                end
            end
        end
      reg145 <= $signed(forvar67);
      reg146 <= $signed((($signed(reg64) ? reg140 : (!(8'ha7))) ?
          reg129 : ({wire27} ?
              ((8'ha4) ? reg96 : (8'ha2)) : $unsigned(reg107))));
      for (forvar147 = (1'h0); (forvar147 < (2'h2)); forvar147 = (forvar147 + (1'h1)))
        begin
          reg148 <= {(~|$signed(forvar74))};
          for (forvar149 = (1'h0); (forvar149 < (1'h1)); forvar149 = (forvar149 + (1'h1)))
            begin
              if ($unsigned({(~^$signed((8'ha9)))}))
                begin
                  for (forvar150 = (1'h0); (forvar150 < (2'h2)); forvar150 = (forvar150 + (1'h1)))
                    begin
                      reg151 <= (8'ha5);
                      reg152 <= reg107[(4'h8):(3'h4)];
                      reg153 <= {(!$unsigned(reg146))};
                    end
                end
              else
                begin
                  reg150 <= forvar100[(4'h8):(3'h4)];
                  reg151 <= (|($signed(reg62[(3'h7):(3'h6)]) ?
                      forvar94[(4'he):(3'h7)] : $unsigned({reg70})));
                  for (forvar152 = (1'h0); (forvar152 < (1'h1)); forvar152 = (forvar152 + (1'h1)))
                    begin
                      reg153 <= (({(forvar130 << forvar93)} != (forvar121 && wire29)) ?
                          ((^~$unsigned(forvar80)) ?
                              $signed(wire34[(1'h1):(1'h1)]) : wire32[(3'h5):(2'h2)]) : forvar37);
                      reg154 <= reg134;
                      reg155 <= $unsigned(({reg43} ?
                          ((reg78 <<< reg113) & $unsigned(wire30)) : reg56));
                      reg156 <= $signed((reg42[(4'h8):(4'h8)] ?
                          $unsigned((^wire24)) : {wire97}));
                    end
                  reg157 <= (reg129 - (8'hba));
                end
              for (forvar158 = (1'h0); (forvar158 < (2'h3)); forvar158 = (forvar158 + (1'h1)))
                begin
                  if ({(((reg51 ? reg145 : reg125) ?
                              $signed(forvar141) : reg115) ?
                          ($unsigned(reg81) && ((8'ha7) ?
                              (8'h9f) : reg91)) : ((forvar141 ~^ forvar67) ?
                              $unsigned(reg101) : $signed(reg58)))})
                    begin
                      reg159 <= (8'haa);
                    end
                  else
                    begin
                      reg159 <= $signed($signed(reg108[(1'h0):(1'h0)]));
                    end
                  if ((($signed((|reg63)) <<< $unsigned($signed(reg96))) != (reg41[(2'h3):(2'h2)] * reg104)))
                    begin
                      reg160 <= forvar63;
                      reg161 <= $unsigned({wire98[(1'h1):(1'h1)]});
                      reg162 <= $unsigned($unsigned((!forvar152[(3'h5):(2'h3)])));
                      reg163 <= reg42;
                    end
                  else
                    begin
                      reg160 <= ((&reg103[(2'h3):(2'h2)]) >= reg151);
                      reg161 <= ($signed((~wire30)) ?
                          reg66[(1'h1):(1'h0)] : (~&(~$signed(reg114))));
                      reg162 <= ($signed(((reg82 ?
                              forvar150 : forvar100) * (forvar94 ^~ reg148))) ?
                          ($signed((8'ha5)) > (^$signed(forvar47))) : (^~wire32));
                    end
                  for (forvar164 = (1'h0); (forvar164 < (1'h1)); forvar164 = (forvar164 + (1'h1)))
                    begin
                      reg165 <= {$unsigned(forvar72[(3'h7):(2'h3)])};
                      reg166 <= (($unsigned($signed(reg115)) >> (~^$unsigned(reg88))) ?
                          {{reg51[(3'h5):(2'h3)]}} : ((reg117[(1'h1):(1'h0)] ?
                                  (reg41 && reg57) : (forvar93 << reg155)) ?
                              {$signed(reg142)} : $signed((~|(8'h9d)))));
                      reg167 <= $signed({$unsigned(reg155[(3'h4):(1'h1)])});
                      reg168 <= wire97;
                    end
                  if ((~|$unsigned(((~^reg144) ? (reg41 * wire28) : reg104))))
                    begin
                      reg169 <= reg133;
                    end
                  else
                    begin
                      reg169 <= reg133[(1'h0):(1'h0)];
                      reg170 <= reg102[(4'h9):(4'h9)];
                      reg171 <= reg150[(3'h4):(2'h3)];
                    end
                end
              reg172 <= (forvar152[(3'h5):(1'h1)] > reg165[(1'h1):(1'h1)]);
            end
          for (forvar173 = (1'h0); (forvar173 < (2'h2)); forvar173 = (forvar173 + (1'h1)))
            begin
              reg174 <= (((reg103 <= ((8'hb0) >> (8'ha7))) ?
                  reg165 : ((wire34 ? forvar93 : reg62) ~^ (reg77 ?
                      reg169 : reg115))) ^~ ($unsigned(reg69[(4'hc):(4'ha)]) | (~(~&forvar54))));
              reg175 <= (|reg45[(3'h5):(2'h3)]);
              for (forvar176 = (1'h0); (forvar176 < (1'h1)); forvar176 = (forvar176 + (1'h1)))
                begin
                  if (forvar121[(4'he):(4'hb)])
                    begin
                      reg177 <= ((^~(((8'haa) && reg101) > (|reg126))) && wire28[(3'h4):(2'h2)]);
                      reg178 <= ($signed((~|reg88)) ?
                          reg91[(4'h8):(2'h2)] : reg53);
                      reg179 <= (reg45[(3'h5):(3'h5)] ?
                          {($signed(reg157) ?
                                  {reg116} : reg171[(1'h1):(1'h1)])} : ($signed(forvar59[(4'h8):(2'h3)]) ?
                              reg122 : reg161[(2'h3):(1'h1)]));
                    end
                  else
                    begin
                      reg177 <= ((8'h9f) ?
                          ((+reg162[(3'h6):(2'h3)]) <<< (reg85[(3'h6):(3'h4)] ?
                              $signed(forvar74) : reg116)) : reg78);
                      reg178 <= ((~|(!reg47)) ? ({{reg67}} + reg143) : (8'ha6));
                      reg179 <= (&($signed((reg172 ?
                          (8'hac) : (8'hb4))) - ($signed((8'hb5)) ?
                          (reg122 ? forvar36 : reg48) : $signed((8'hb8)))));
                      reg180 <= (reg103 <= (reg52 && (reg118[(2'h3):(2'h3)] == forvar47)));
                    end
                end
              reg181 <= {$signed(($unsigned(reg122) ?
                      reg46[(3'h5):(1'h0)] : (wire27 ? forvar150 : wire98)))};
            end
        end
    end
  assign wire182 = reg122;
  assign wire183 = (reg175 >= (^((reg108 ?
                       forvar158 : wire30) == $unsigned(forvar106))));
  assign wire184 = (|reg126[(3'h6):(1'h0)]);
endmodule