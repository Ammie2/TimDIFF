module top
#( parameter param451 = (({((8'hac) ? (-(8'hbf)) : {(8'ha7)}), ((!(8'had)) ? ((7'h42) || (8'hbb)) : {(8'ha8)})} >>> (8'hb5)) > ((+(((7'h44) || (8'hab)) ? ((8'ha3) ^~ (8'ha6)) : (-(8'ha3)))) ^ ((((8'ha5) * (8'ha0)) ? ((7'h44) + (8'hb0)) : ((8'ha6) ? (8'ha0) : (8'haa))) ^ (((8'hb6) ^ (8'ha8)) ? {(8'ha2)} : ((8'ha5) ? (8'hbc) : (8'ha1)))))) )
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h39b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire3;
  input wire signed [(5'h11):(1'h0)] wire2;
  input wire signed [(2'h2):(1'h0)] wire1;
  input wire signed [(4'h9):(1'h0)] wire0;
  wire [(3'h7):(1'h0)] wire450;
  wire [(4'he):(1'h0)] wire441;
  wire signed [(3'h5):(1'h0)] wire191;
  reg signed [(4'he):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg189 = (1'h0);
  reg [(3'h5):(1'h0)] reg188 = (1'h0);
  reg [(4'he):(1'h0)] reg187 = (1'h0);
  reg [(2'h2):(1'h0)] reg186 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg185 = (1'h0);
  reg [(4'hd):(1'h0)] reg184 = (1'h0);
  reg [(4'hc):(1'h0)] reg183 = (1'h0);
  reg [(3'h6):(1'h0)] reg182 = (1'h0);
  reg [(4'hb):(1'h0)] reg181 = (1'h0);
  reg [(3'h5):(1'h0)] reg180 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg179 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg178 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg176 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg174 = (1'h0);
  reg [(5'h13):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg171 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg170 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg167 = (1'h0);
  reg [(4'hc):(1'h0)] reg166 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg165 = (1'h0);
  reg [(3'h4):(1'h0)] reg164 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg163 = (1'h0);
  reg [(5'h13):(1'h0)] reg162 = (1'h0);
  reg [(3'h5):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg160 = (1'h0);
  reg [(4'h8):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg158 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg157 = (1'h0);
  reg [(4'hb):(1'h0)] reg156 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg154 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg152 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg151 = (1'h0);
  reg [(5'h13):(1'h0)] reg150 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg149 = (1'h0);
  reg [(5'h11):(1'h0)] reg148 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire146;
  wire [(4'hb):(1'h0)] wire26;
  reg [(4'hc):(1'h0)] reg25 = (1'h0);
  reg [(5'h14):(1'h0)] reg24 = (1'h0);
  reg [(3'h6):(1'h0)] reg23 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg22 = (1'h0);
  reg [(4'he):(1'h0)] reg21 = (1'h0);
  wire signed [(5'h13):(1'h0)] wire20;
  wire signed [(5'h14):(1'h0)] wire19;
  reg signed [(5'h12):(1'h0)] reg18 = (1'h0);
  reg [(4'hd):(1'h0)] reg17 = (1'h0);
  reg [(5'h13):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg14 = (1'h0);
  reg [(5'h10):(1'h0)] reg13 = (1'h0);
  reg [(5'h13):(1'h0)] reg12 = (1'h0);
  reg signed [(4'he):(1'h0)] reg11 = (1'h0);
  reg [(3'h7):(1'h0)] reg10 = (1'h0);
  reg [(4'hf):(1'h0)] reg9 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire8;
  wire [(4'he):(1'h0)] wire7;
  wire [(5'h12):(1'h0)] wire6;
  wire signed [(2'h2):(1'h0)] wire5;
  wire signed [(2'h3):(1'h0)] wire4;
  reg signed [(5'h10):(1'h0)] reg443 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire444;
  wire [(3'h5):(1'h0)] wire445;
  wire signed [(4'hc):(1'h0)] wire446;
  wire [(5'h11):(1'h0)] wire447;
  wire signed [(4'hc):(1'h0)] wire448;
  assign y = {wire450,
                 wire441,
                 wire191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 wire146,
                 wire26,
                 reg25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 wire20,
                 wire19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg9,
                 wire8,
                 wire7,
                 wire6,
                 wire5,
                 wire4,
                 reg443,
                 wire444,
                 wire445,
                 wire446,
                 wire447,
                 wire448,
                 (1'h0)};
  assign wire4 = (((wire3[(4'hd):(3'h4)] || $signed(wire3)) ?
                     (^~(wire2 && $unsigned(wire0))) : (+wire1)) * (wire1[(1'h1):(1'h0)] >> ($signed((^~wire1)) ?
                     (wire0 ? wire2 : (!wire3)) : wire0[(3'h4):(1'h1)])));
  assign wire5 = ($unsigned($signed(((wire1 ? wire0 : wire0) - (wire0 ?
                         wire4 : wire1)))) ?
                     {{(wire2 ~^ wire1[(1'h1):(1'h0)]),
                             {(^~wire2), ((8'hb6) != wire3)}},
                         $unsigned((~|wire0[(3'h7):(2'h3)]))} : $signed(wire1));
  assign wire6 = $unsigned(wire1[(2'h2):(2'h2)]);
  assign wire7 = wire5[(1'h0):(1'h0)];
  assign wire8 = wire5;
  always
    @(posedge clk) begin
      reg9 <= $unsigned(wire3);
      if (wire5)
        begin
          reg10 <= ($unsigned($unsigned(((wire7 >> wire8) <= $unsigned(reg9)))) ?
              (wire3[(1'h0):(1'h0)] ?
                  {$unsigned($signed(wire3))} : wire1) : (wire0 ?
                  $unsigned($signed(wire3)) : {$unsigned($signed(wire6)),
                      wire1[(2'h2):(2'h2)]}));
          reg11 <= $unsigned(($signed((((8'ha7) ?
              wire7 : wire2) <= $unsigned(wire3))) & $unsigned((^$signed(wire5)))));
          if ({wire6, wire3})
            begin
              reg12 <= $unsigned($unsigned((8'hb7)));
              reg13 <= $signed((($signed($unsigned(wire2)) >= wire1) ?
                  ({(~reg11)} ? wire0[(4'h8):(3'h5)] : reg9) : {((~|wire8) ?
                          (wire4 ^~ reg12) : (!(8'ha9)))}));
              reg14 = reg9;
              reg15 = wire1;
            end
          else
            begin
              reg12 <= reg12[(3'h7):(3'h6)];
              reg13 <= (-$signed((reg14 - ((wire6 ? reg9 : (8'ha6)) ?
                  reg12 : (reg13 ? wire1 : reg9)))));
              reg14 <= (~^($unsigned(($signed((8'hb6)) ?
                  $signed(wire8) : (8'h9f))) * ($signed($signed(wire5)) & wire4)));
              reg15 = $unsigned(wire4[(1'h0):(1'h0)]);
            end
        end
      else
        begin
          reg10 <= $signed($signed((wire1 ?
              (reg13 >= reg13[(4'hd):(1'h1)]) : (^~(wire7 ? wire2 : wire0)))));
          if ({($signed($unsigned(wire6[(4'hf):(4'hc)])) ?
                  (~$signed($signed(reg11))) : $signed(wire1[(2'h2):(1'h1)]))})
            begin
              reg11 = wire0[(4'h8):(1'h1)];
              reg12 = reg13[(3'h6):(1'h0)];
            end
          else
            begin
              reg11 <= $unsigned(reg9);
              reg12 <= (reg9 <= $signed(($signed((reg14 >> (8'had))) ?
                  {$signed((8'hbb)),
                      (wire3 != (8'ha4))} : wire6[(5'h10):(1'h0)])));
              reg13 = reg11[(3'h6):(3'h6)];
              reg14 <= wire0[(3'h7):(3'h5)];
            end
          reg15 <= (^~($unsigned(reg15[(4'hd):(4'hd)]) ?
              $unsigned(wire7[(4'he):(4'he)]) : {($signed(wire1) <<< reg14[(2'h2):(2'h2)]),
                  {reg11[(4'hb):(2'h2)], (wire4 ? (8'hb0) : reg14)}}));
          reg16 = wire7;
        end
      reg17 <= $signed(reg16);
      reg18 <= ($unsigned($unsigned($signed($unsigned(reg14)))) ?
          wire8 : (reg17 ^~ $signed(wire3[(5'h10):(4'ha)])));
    end
  assign wire19 = $unsigned($unsigned(wire4));
  assign wire20 = reg14;
  always
    @(posedge clk) begin
      reg21 <= (($signed($signed(((8'h9f) >= wire1))) ?
          $signed(((reg12 ? reg9 : reg18) ?
              $unsigned(reg12) : reg10)) : (($signed((8'hac)) ?
                  $unsigned(reg14) : wire20) ?
              (&$unsigned(wire2)) : ((&wire0) >>> $signed(wire6)))) <= ((8'haa) ?
          (-wire19[(3'h6):(1'h1)]) : (reg12[(4'he):(4'h8)] <<< (wire0[(3'h4):(3'h4)] ?
              ((8'ha4) && wire6) : (8'hb7)))));
      reg22 <= wire0;
      reg23 <= (wire19[(4'h9):(1'h0)] ?
          $unsigned((reg13 == $signed($signed((7'h43))))) : (wire5[(1'h1):(1'h0)] & $unsigned(wire0)));
      reg24 = reg23[(2'h3):(1'h1)];
      reg25 <= $unsigned((wire2[(2'h3):(1'h0)] ?
          {$unsigned($unsigned(reg15)),
              (reg17 != $signed(reg22))} : (&(~|(|(8'hbd))))));
    end
  assign wire26 = ((~&$unsigned((-(reg10 ^ reg17)))) ?
                      reg12 : (!{$unsigned(wire8),
                          (wire8[(3'h7):(3'h7)] ?
                              reg25[(4'hb):(1'h0)] : wire5)}));
  module27 modinst147 (.wire29(reg11), .wire28(reg10), .clk(clk), .wire30(wire20), .y(wire146), .wire31(wire3));
  always
    @(posedge clk) begin
      if ({(^((wire5 & (wire26 < reg12)) + (!{reg21, wire5}))), reg11})
        begin
          if ((((-reg11) ?
              reg24 : (|(reg24[(3'h5):(1'h0)] != {wire6}))) ^ ({($unsigned(reg15) ?
                      $unsigned(reg22) : $unsigned(wire0))} ?
              $signed((8'hb4)) : ({(reg10 ? wire3 : reg17),
                  {(7'h42)}} > $signed({(7'h44)})))))
            begin
              reg148 = reg14[(2'h2):(1'h1)];
              reg149 = $unsigned($signed(wire5));
              reg150 <= {(!({wire5} ?
                      (+(reg11 | reg10)) : reg13[(2'h2):(2'h2)])),
                  $signed((($unsigned((8'ha5)) & reg25[(3'h6):(3'h4)]) ?
                      $signed($signed(wire8)) : wire3))};
            end
          else
            begin
              reg148 <= wire146;
              reg149 <= $unsigned((($unsigned(reg10[(1'h0):(1'h0)]) ?
                      (!(!reg13)) : reg148) ?
                  {($unsigned(reg24) != (8'hb1)),
                      (wire146 ~^ {reg21})} : reg23));
            end
          reg151 <= ($unsigned($unsigned($signed($unsigned(wire0)))) ?
              reg149[(1'h0):(1'h0)] : ({$unsigned((^~reg22)),
                  ((reg18 + reg9) >> wire20)} <= (reg22[(2'h3):(1'h1)] ?
                  reg16 : $signed(reg10[(2'h2):(1'h1)]))));
          if ((!$unsigned(reg15)))
            begin
              reg152 = wire2[(5'h11):(4'ha)];
              reg153 = wire20[(4'ha):(2'h2)];
              reg154 = $signed(({(!$signed(reg25))} ? reg21 : wire5));
            end
          else
            begin
              reg152 = wire1[(2'h2):(2'h2)];
            end
          if ($signed((~&$unsigned((^$signed(reg18))))))
            begin
              reg155 = $unsigned((~|(reg148[(4'h8):(1'h0)] <= $unsigned($unsigned(reg25)))));
            end
          else
            begin
              reg155 <= $signed($unsigned({reg12}));
              reg156 <= ($signed({reg22[(2'h3):(1'h1)]}) ?
                  reg155[(3'h6):(3'h4)] : ((~|reg13) ?
                      (8'hb3) : ($signed((7'h42)) == (~$signed(reg22)))));
              reg157 <= ((7'h44) ?
                  $unsigned(reg23[(1'h1):(1'h1)]) : $signed(((~&wire7) ?
                      ($signed(wire26) >>> $signed(reg17)) : (+(~|(8'h9f))))));
              reg158 <= $unsigned(((7'h43) ?
                  $signed({wire4[(1'h0):(1'h0)],
                      $unsigned(reg149)}) : (8'haf)));
            end
          if ($signed($signed(({reg24, (~&wire1)} ?
              wire0 : $unsigned((wire3 ? reg12 : (8'ha9)))))))
            begin
              reg159 = (8'hb7);
              reg160 <= (((wire6[(3'h7):(3'h4)] & $signed({reg10})) - (~^(~^(wire26 ?
                  wire20 : wire5)))) < $unsigned($unsigned((-reg157[(2'h3):(1'h0)]))));
              reg161 <= reg18[(2'h2):(2'h2)];
              reg162 <= ($unsigned((((~reg150) ?
                          wire0[(1'h0):(1'h0)] : (reg23 + reg14)) ?
                      wire2[(5'h10):(4'h9)] : (^~{reg14}))) ?
                  wire8[(2'h2):(2'h2)] : $unsigned(reg161[(2'h2):(1'h1)]));
            end
          else
            begin
              reg159 = reg162;
              reg160 <= $signed(($unsigned(((~^reg149) ?
                      $signed(reg153) : $signed((8'hab)))) ?
                  ($signed({reg154,
                      reg25}) | reg148[(4'hd):(3'h7)]) : ($signed(((8'hb2) ?
                          reg162 : reg160)) ?
                      $unsigned((wire19 >= reg18)) : wire3)));
              reg161 <= (|(($unsigned((8'h9c)) > (~&((8'h9f) ?
                  reg18 : reg153))) * ($unsigned((~^reg15)) ^ $unsigned($signed(reg153)))));
              reg162 <= reg24[(4'ha):(3'h5)];
            end
        end
      else
        begin
          reg148 = (reg155[(4'h9):(1'h0)] || reg11);
          reg149 <= ((^reg158) == ({$signed({wire26})} ?
              (+$signed((reg162 && reg161))) : wire0));
          if ($signed($signed(reg10[(3'h5):(1'h0)])))
            begin
              reg150 <= {{$signed(((~^wire6) || {reg157})),
                      wire7[(3'h5):(1'h1)]},
                  reg14};
              reg151 <= {(^((reg23[(3'h5):(2'h3)] ?
                      wire20[(3'h4):(2'h2)] : reg154[(4'ha):(3'h6)]) >> $signed(wire20))),
                  ($signed(wire5) ? wire8 : $unsigned(wire0[(4'h9):(4'h9)]))};
              reg152 = wire8[(4'h8):(3'h7)];
              reg153 = reg162;
              reg154 <= $signed($unsigned((~|(!$unsigned(reg158)))));
            end
          else
            begin
              reg150 <= ($unsigned(wire5) ?
                  $unsigned({(+(wire26 ~^ reg18))}) : reg153[(3'h7):(3'h5)]);
              reg151 = reg162[(5'h10):(2'h3)];
              reg152 = $signed(reg21);
              reg153 <= $unsigned(reg24[(3'h7):(2'h3)]);
              reg154 = $unsigned(reg15[(4'h9):(1'h0)]);
            end
          if ((($unsigned((~$unsigned(reg21))) << wire7[(4'hc):(3'h4)]) ?
              $signed(((wire7[(4'he):(4'he)] ?
                      (reg10 == (8'haa)) : $signed(reg162)) ?
                  wire4 : ((reg10 || (8'hb6)) <<< $signed(reg159)))) : (reg10 >> $signed($unsigned($signed(reg13))))))
            begin
              reg155 = wire5[(1'h0):(1'h0)];
            end
          else
            begin
              reg155 <= $unsigned(($signed(((~|wire8) ?
                      {reg11} : $unsigned(reg149))) ?
                  ({reg9, $signed(wire5)} ?
                      $signed({reg12, reg159}) : ($unsigned(reg154) ?
                          $unsigned(reg150) : $unsigned((8'haf)))) : ((wire26 ?
                      (wire2 ? wire8 : reg151) : reg21) >>> ((~reg23) ?
                      (~^reg149) : (7'h40)))));
              reg156 = (~($unsigned($unsigned($unsigned(reg16))) && wire5));
            end
          if ((reg16[(4'h8):(2'h3)] ?
              ((reg12[(3'h6):(1'h1)] ?
                  (|wire5[(1'h0):(1'h0)]) : ((reg18 ? reg162 : reg15) ?
                      $unsigned(wire3) : $unsigned((8'h9d)))) < (($signed(reg22) ?
                      {wire146, reg159} : (wire6 ? reg156 : reg10)) ?
                  (|$signed((7'h44))) : (reg18[(5'h11):(1'h0)] ?
                      wire20 : (reg150 ?
                          reg161 : reg16)))) : $signed(((reg14[(2'h2):(1'h1)] | $signed(wire3)) ?
                  ((reg22 ? wire20 : reg9) > reg149) : ($signed(wire3) ?
                      (wire8 > (8'haf)) : {reg11, reg13})))))
            begin
              reg157 <= $signed($signed((wire0 && $unsigned((wire0 ?
                  wire20 : wire1)))));
              reg158 = reg157;
              reg159 <= $signed((((~^wire20[(5'h10):(4'hf)]) ?
                  reg149[(1'h0):(1'h0)] : {$signed(reg155),
                      reg14[(1'h0):(1'h0)]}) && (~(wire146[(5'h13):(4'hf)] + (reg22 ?
                  reg23 : reg11)))));
              reg160 <= $signed((reg24 ?
                  $unsigned(reg12[(3'h7):(2'h2)]) : {reg157}));
            end
          else
            begin
              reg157 <= (wire1[(1'h1):(1'h0)] ?
                  (wire19[(5'h11):(2'h3)] != $signed((wire26 + ((8'haa) || reg155)))) : {$unsigned((8'hb0))});
              reg158 = ($unsigned((~$signed(reg160[(4'he):(1'h0)]))) >= {$unsigned(reg9[(4'hb):(4'h9)])});
              reg159 = reg18;
              reg160 <= (^~reg157);
              reg161 <= (wire2[(3'h5):(1'h1)] != ((reg21 ?
                      reg149 : $unsigned((wire7 ? reg13 : reg18))) ?
                  $unsigned($signed(wire2[(3'h4):(3'h4)])) : wire8[(3'h7):(1'h1)]));
            end
        end
      reg163 = (^~{(^$unsigned((8'had)))});
      if ((-$signed((8'hbb))))
        begin
          reg164 = ($unsigned((~|(8'ha6))) - (~^{$unsigned((~^reg159))}));
          reg165 <= ((|({reg11, (~|reg15)} ?
                  reg9 : $unsigned((reg157 ? (8'hb1) : reg160)))) ?
              ($signed(reg18) & $unsigned(wire6)) : reg154[(5'h10):(1'h0)]);
          reg166 <= {{(($signed(reg162) ?
                          $signed(reg10) : (wire3 ? (7'h41) : wire146)) ?
                      wire1 : ((reg150 && reg21) ? (^~(8'ha6)) : reg14))}};
          reg167 = wire0[(3'h5):(2'h3)];
        end
      else
        begin
          reg164 <= $unsigned(((+$signed($unsigned(reg17))) ?
              $unsigned($signed({reg158})) : ((~^$unsigned(reg159)) ^ reg167)));
          if ($unsigned({(~&$unsigned($unsigned(reg165)))}))
            begin
              reg165 = wire3;
            end
          else
            begin
              reg165 <= $unsigned($unsigned((({(8'h9c)} ?
                  (&reg10) : $unsigned(reg9)) == $signed((&wire1)))));
              reg166 <= $unsigned(((($unsigned(reg159) - wire2) ?
                  {(reg166 ?
                          (8'hb7) : wire6)} : (reg21[(2'h2):(2'h2)] || $unsigned(wire3))) > reg149));
              reg167 = reg15;
            end
          reg168 <= {((((~^reg159) ?
                          (wire26 && reg11) : (wire2 ? (8'ha6) : reg164)) ?
                      ((^wire8) >= (+reg156)) : (&(reg153 ? reg167 : wire6))) ?
                  reg153 : (+(wire8[(3'h6):(1'h1)] < reg150[(5'h11):(1'h1)])))};
          if (($signed(reg155[(1'h0):(1'h0)]) + ($unsigned(reg17) ?
              $signed($signed($signed(reg162))) : $signed(reg18))))
            begin
              reg169 = reg165;
              reg170 = (8'ha5);
              reg171 <= $unsigned((reg14[(2'h3):(2'h2)] ?
                  $unsigned((~&$signed(reg18))) : {$signed((reg18 <<< wire1)),
                      ((-(8'ha7)) ? $signed(reg167) : $signed(wire26))}));
              reg172 = $signed($signed(reg153[(3'h4):(2'h2)]));
            end
          else
            begin
              reg169 <= {$signed((|{$signed(wire26)})),
                  (reg164 ?
                      reg160 : ((^(~&reg156)) ?
                          (wire0[(2'h3):(1'h0)] ?
                              (wire5 ?
                                  wire146 : reg10) : (~&wire5)) : (^~wire6[(4'he):(4'hc)])))};
              reg170 = reg24;
              reg171 = (~^reg161);
              reg172 = (wire3[(3'h4):(1'h1)] ? $unsigned((8'ha7)) : reg15);
              reg173 <= ((reg159 <= {$unsigned({wire20}), (!(&wire5))}) ?
                  reg153 : (|$unsigned((-wire5))));
            end
        end
      if ((8'haf))
        begin
          reg174 = reg159[(2'h3):(2'h3)];
          reg175 <= (($unsigned((^~(reg160 ? reg171 : reg24))) ?
                  reg14[(1'h1):(1'h1)] : reg159) ?
              reg13[(4'h9):(2'h3)] : reg16[(5'h11):(2'h2)]);
          reg176 = $signed((reg158 * {{(reg173 >>> (8'hbc))}}));
          reg177 <= $signed(($signed(($unsigned(reg150) ?
                  reg152 : $signed((8'h9d)))) ?
              ((wire5[(2'h2):(1'h0)] ? reg9[(4'hb):(4'h8)] : wire7) ?
                  (^reg164[(2'h3):(2'h2)]) : $unsigned(reg170)) : reg25[(2'h3):(2'h2)]));
        end
      else
        begin
          reg174 = reg154[(4'he):(4'hc)];
          reg175 <= ((($signed((^~(8'hac))) ?
                  $signed({(7'h43)}) : $signed((reg156 ?
                      (8'ha7) : wire5))) * $unsigned(((8'h9e) < {reg173}))) ?
              wire1 : {{({reg175} ? (reg167 != reg165) : (reg153 == (8'hbf))),
                      (8'hae)}});
          reg176 = wire8[(3'h4):(1'h1)];
          reg177 = wire146[(5'h12):(3'h7)];
        end
    end
  always
    @(posedge clk) begin
      reg178 <= $signed($signed({(|reg151), {$unsigned((8'hb6))}}));
      reg179 <= reg158[(2'h2):(1'h1)];
      if ($unsigned(((~($unsigned(reg15) >= (!reg177))) | (((reg172 ^~ reg170) ?
          reg162 : $unsigned(reg13)) <= reg164[(2'h2):(1'h0)]))))
        begin
          reg180 <= reg149[(1'h0):(1'h0)];
          if (($signed((~^((reg14 ? (8'ha3) : reg165) ^ $signed((8'ha2))))) ?
              reg162[(5'h11):(4'ha)] : $signed($signed(((+reg180) * (wire2 < reg177))))))
            begin
              reg181 = reg176[(1'h0):(1'h0)];
              reg182 = (!(^~reg17));
            end
          else
            begin
              reg181 <= $signed((reg151[(1'h1):(1'h0)] ?
                  (reg178[(3'h4):(1'h1)] ?
                      {((8'h9d) ?
                              reg14 : (8'ha3))} : {$signed(reg152)}) : reg18[(4'h8):(3'h5)]));
              reg182 = (+(|reg157[(3'h4):(1'h1)]));
            end
          reg183 = (8'hae);
          reg184 = reg17[(3'h6):(3'h5)];
        end
      else
        begin
          reg180 = $signed(reg18[(3'h4):(2'h3)]);
          reg181 = reg10;
          reg182 <= (~|reg161);
          if (wire146[(4'hb):(2'h2)])
            begin
              reg183 <= ((+($unsigned($signed((8'haa))) <<< (~^$signed(wire19)))) ?
                  {wire20} : $unsigned($unsigned(({reg21} & (+reg182)))));
              reg184 = (~&(+reg179));
              reg185 = $unsigned(reg21[(2'h3):(1'h1)]);
            end
          else
            begin
              reg183 = reg9;
            end
        end
      if ($unsigned($signed((($signed(reg9) > $signed(reg24)) == $signed(wire26[(4'ha):(4'h8)])))))
        begin
          reg186 <= $unsigned((reg153 != $unsigned(((8'haa) ?
              $unsigned(reg17) : $unsigned(wire2)))));
          reg187 = reg150[(4'h9):(3'h4)];
          reg188 = reg165[(3'h4):(1'h1)];
        end
      else
        begin
          reg186 = reg172[(5'h14):(5'h10)];
          if ($unsigned(reg9))
            begin
              reg187 <= ({({((8'ha6) & reg148),
                      $unsigned(wire7)} == {reg24[(4'ha):(1'h1)]})} >> $unsigned($unsigned($signed($unsigned(reg18)))));
            end
          else
            begin
              reg187 = $signed(reg165[(1'h1):(1'h0)]);
              reg188 = reg13;
              reg189 <= (({(^(8'ha0)), reg13} ?
                      reg169[(4'h8):(3'h6)] : reg150[(5'h12):(4'h9)]) ?
                  ({(|(reg12 < (8'h9f)))} << $signed((!$unsigned((8'ha1))))) : $signed(reg24[(4'ha):(1'h0)]));
            end
          reg190 <= $unsigned(({(reg22[(1'h1):(1'h0)] ?
                  {wire8} : {reg148,
                      (8'hb9)})} * $signed($unsigned((~|reg17)))));
        end
    end
  assign wire191 = $signed(reg151);
  module192 modinst442 (wire441, clk, reg184, reg14, reg150, reg158, reg16);
  always
    @(posedge clk) begin
      reg443 = reg11;
    end
  assign wire444 = $unsigned({($unsigned(reg183[(3'h5):(1'h0)]) ?
                           $signed((wire191 || reg179)) : reg180[(1'h1):(1'h0)]),
                       reg23[(1'h0):(1'h0)]});
  assign wire445 = reg175[(2'h2):(2'h2)];
  assign wire446 = reg17[(4'h9):(3'h5)];
  assign wire447 = reg182[(3'h5):(1'h1)];
  module192 modinst449 (wire448, clk, reg190, reg12, reg152, reg154, reg176);
  assign wire450 = $unsigned(wire4[(2'h3):(1'h0)]);
endmodule

module module192  (y, clk, wire197, wire196, wire195, wire194, wire193);
  output wire [(32'h26d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire197;
  input wire signed [(5'h13):(1'h0)] wire196;
  input wire [(4'hb):(1'h0)] wire195;
  input wire [(3'h7):(1'h0)] wire194;
  input wire signed [(5'h13):(1'h0)] wire193;
  wire signed [(4'hf):(1'h0)] wire439;
  reg [(4'he):(1'h0)] reg438 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg436 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire403;
  wire [(5'h15):(1'h0)] wire375;
  wire [(4'h8):(1'h0)] wire354;
  wire signed [(3'h7):(1'h0)] wire352;
  wire [(4'h9):(1'h0)] wire295;
  reg [(4'hc):(1'h0)] reg294 = (1'h0);
  reg signed [(4'he):(1'h0)] reg293 = (1'h0);
  reg [(2'h3):(1'h0)] reg292 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg291 = (1'h0);
  reg [(3'h5):(1'h0)] reg290 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg289 = (1'h0);
  reg [(3'h5):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg286 = (1'h0);
  wire [(5'h13):(1'h0)] wire285;
  reg [(5'h15):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg283 = (1'h0);
  reg [(4'hf):(1'h0)] reg282 = (1'h0);
  reg [(4'hc):(1'h0)] reg281 = (1'h0);
  reg [(5'h15):(1'h0)] reg280 = (1'h0);
  reg [(5'h15):(1'h0)] reg279 = (1'h0);
  reg [(5'h15):(1'h0)] reg278 = (1'h0);
  reg [(3'h7):(1'h0)] reg277 = (1'h0);
  reg [(2'h2):(1'h0)] reg276 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg275 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg274 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg273 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg272 = (1'h0);
  reg [(5'h10):(1'h0)] reg271 = (1'h0);
  wire [(3'h6):(1'h0)] wire270;
  wire [(5'h12):(1'h0)] wire269;
  wire [(4'he):(1'h0)] wire268;
  wire signed [(5'h15):(1'h0)] wire267;
  wire [(5'h14):(1'h0)] wire266;
  wire [(4'ha):(1'h0)] wire265;
  wire [(5'h13):(1'h0)] wire263;
  reg [(5'h15):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg406 = (1'h0);
  reg [(2'h3):(1'h0)] reg407 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg408 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg409 = (1'h0);
  wire [(5'h13):(1'h0)] wire410;
  wire [(3'h6):(1'h0)] wire411;
  wire [(4'hf):(1'h0)] wire434;
  assign y = {wire439,
                 reg438,
                 reg437,
                 reg436,
                 wire403,
                 wire375,
                 wire354,
                 wire352,
                 wire295,
                 reg294,
                 reg293,
                 reg292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 wire285,
                 reg284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 wire270,
                 wire269,
                 wire268,
                 wire267,
                 wire266,
                 wire265,
                 wire263,
                 reg405,
                 reg406,
                 reg407,
                 reg408,
                 reg409,
                 wire410,
                 wire411,
                 wire434,
                 (1'h0)};
  module198 modinst264 (.wire200(wire193), .wire199(wire195), .wire202(wire197), .y(wire263), .wire201(wire196), .clk(clk));
  assign wire265 = ((|wire195) ?
                       {$signed(wire197[(4'h9):(3'h4)]),
                           ($signed((|wire197)) ?
                               wire194[(2'h2):(2'h2)] : wire193)} : wire196[(4'hd):(3'h4)]);
  assign wire266 = (~&(($signed((wire193 ^ wire193)) >>> wire196[(3'h7):(2'h3)]) != {{wire265[(1'h1):(1'h1)],
                           $signed(wire196)}}));
  assign wire267 = wire266[(2'h3):(1'h0)];
  assign wire268 = (~&(7'h42));
  assign wire269 = (({{$signed(wire268)}} ?
                       wire267[(3'h7):(2'h3)] : {((|wire267) <<< {wire194,
                               (8'hb9)}),
                           $signed(wire194)}) & $signed((8'hbb)));
  assign wire270 = $unsigned(wire267[(5'h12):(4'hf)]);
  always
    @(posedge clk) begin
      if (wire263)
        begin
          reg271 <= (-wire269[(1'h1):(1'h0)]);
          if ({{(+(^~$unsigned(wire270)))},
              ({($signed(wire263) ? (8'hbd) : (wire197 ? (8'haa) : wire269)),
                      (~|$unsigned(wire193))} ?
                  (((wire268 || wire194) * (reg271 ? wire266 : wire196)) ?
                      (~&(wire195 ? wire268 : wire194)) : {(&wire265),
                          (!wire269)}) : (((wire268 ^ wire268) ?
                          (~&wire269) : wire195[(3'h6):(2'h3)]) ?
                      ($signed(wire193) ~^ (!wire193)) : $unsigned((~^(8'h9f)))))})
            begin
              reg272 <= $signed(({(!(wire270 > wire265))} < reg271[(4'hd):(1'h0)]));
              reg273 = reg271[(4'hc):(1'h1)];
              reg274 = $unsigned((reg272 == $signed(wire265)));
              reg275 = (8'hb4);
            end
          else
            begin
              reg272 <= reg272[(3'h5):(1'h0)];
              reg273 <= (reg272[(3'h5):(3'h5)] >> reg274[(1'h0):(1'h0)]);
              reg274 <= ((-(((wire270 >> wire195) <= ((8'hb2) ?
                      reg271 : reg271)) != $unsigned($unsigned(reg275)))) ?
                  (($unsigned(wire263) | wire197) ?
                      (($signed(wire197) ? (~^reg274) : $unsigned(reg272)) ?
                          {$unsigned(wire197),
                              wire265[(2'h3):(1'h0)]} : (wire268 >> {(8'hbd)})) : ($unsigned((^~wire267)) + $signed({wire269}))) : (!((wire266 ?
                      wire194[(2'h2):(2'h2)] : $unsigned(wire194)) | $signed((wire194 ^ wire270)))));
              reg275 <= $unsigned((((((8'hbd) ?
                  wire195 : reg273) >> wire269[(2'h2):(1'h0)]) ~^ $unsigned($unsigned(wire270))) != wire193));
              reg276 = reg272[(2'h2):(1'h1)];
            end
          reg277 <= (^~{$signed($unsigned($signed(reg272))),
              wire267[(3'h5):(1'h0)]});
          reg278 = (7'h40);
        end
      else
        begin
          reg271 <= (wire269[(3'h5):(1'h0)] ?
              {$unsigned({(wire267 >= wire197), (~reg275)}),
                  $unsigned(reg277[(3'h7):(3'h7)])} : (wire196 ?
                  reg274[(3'h5):(2'h2)] : $signed($unsigned({wire193}))));
          reg272 <= {$unsigned(wire196),
              $signed($signed($unsigned({wire263})))};
          reg273 = $unsigned(($signed(reg276[(2'h2):(2'h2)]) <<< (8'hbe)));
          reg274 <= wire266;
          reg275 <= ($unsigned(wire267[(4'hc):(4'h8)]) >> (~^$signed((~^$signed(wire267)))));
        end
      reg279 <= reg278;
      reg280 <= (((((wire196 * wire196) > $unsigned(reg277)) ?
              wire263 : reg274[(3'h7):(2'h3)]) ?
          wire267 : ((^~((8'hae) + wire193)) ?
              ((reg276 ? wire195 : reg279) ?
                  wire195 : (wire269 >> wire266)) : wire267)) & reg279[(4'h9):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg281 <= ((+($unsigned((reg277 ^ reg280)) ?
              (reg279[(4'h8):(3'h7)] < {wire266}) : $signed(wire269))) ?
          reg280[(3'h7):(3'h7)] : ((wire194[(1'h1):(1'h0)] ?
                  $signed({wire263}) : {$unsigned((7'h41))}) ?
              $unsigned({wire270[(1'h0):(1'h0)]}) : wire195));
      reg282 = reg276;
      reg283 <= $signed(($signed((!(|reg278))) >>> $signed(((8'had) ?
          (reg272 && reg277) : wire269))));
      reg284 = (^~$unsigned(reg278));
    end
  assign wire285 = $unsigned($signed((!$signed((reg272 ? reg278 : (8'hb3))))));
  always
    @(posedge clk) begin
      reg286 <= $signed({(~&($unsigned((8'ha5)) >> ((8'ha4) ?
              wire195 : wire196)))});
      reg287 <= reg281;
      if (wire269)
        begin
          if ((((~^$signed((wire266 && reg280))) ^ (wire195[(4'h8):(3'h5)] ^ wire196[(4'h8):(4'h8)])) ?
              reg283[(3'h4):(2'h3)] : (wire263[(4'hd):(1'h1)] ?
                  (&(wire270 ?
                      $signed(wire193) : wire270)) : ($signed((wire266 ?
                      reg276 : reg274)) << (^(reg281 ^ reg278))))))
            begin
              reg288 = $signed((-$unsigned((^wire195))));
            end
          else
            begin
              reg288 = reg284[(5'h15):(5'h10)];
              reg289 = reg287;
              reg290 <= (((reg280 ?
                  (wire195 ?
                      reg280 : $signed(wire266)) : $signed($signed(reg278))) | wire266[(4'hf):(4'h8)]) != reg271[(1'h1):(1'h1)]);
              reg291 <= ($signed(reg277[(1'h0):(1'h0)]) ?
                  reg272[(1'h1):(1'h1)] : (~|reg283));
            end
          reg292 = ((-(($unsigned(reg282) || wire268) ^~ reg281)) || reg281[(1'h1):(1'h0)]);
          reg293 = (^wire269);
          reg294 = (!reg272[(3'h5):(3'h5)]);
        end
      else
        begin
          reg288 = wire194[(2'h3):(2'h3)];
        end
    end
  assign wire295 = (((^~((reg273 ? reg283 : wire193) <<< (wire263 ?
                           wire195 : wire195))) ?
                       {{(reg283 ? reg281 : reg286)},
                           wire263} : $signed((!reg283[(3'h4):(1'h0)]))) || (~^reg274));
  module296 modinst353 (.wire299(reg283), .y(wire352), .wire298(reg282), .wire300(wire194), .clk(clk), .wire297(wire268));
  assign wire354 = {$signed(((^(wire270 ? reg274 : (8'hb3))) <<< wire193))};
  module355 modinst376 (.wire359(wire285), .y(wire375), .wire358(wire268), .clk(clk), .wire356(reg293), .wire357(reg291));
  module377 modinst404 (.y(wire403), .wire381(reg271), .wire380(wire375), .wire378(reg280), .clk(clk), .wire379(reg289), .wire382(reg281));
  always
    @(posedge clk) begin
      reg405 = $signed((~|(|($unsigned(wire197) >>> $unsigned(wire197)))));
      reg406 = $unsigned($signed($unsigned(wire354[(2'h3):(2'h2)])));
      reg407 <= ($signed($unsigned($signed((wire196 ~^ (8'hbf))))) != ((($signed(wire267) ?
                  (reg279 ? wire194 : wire263) : $unsigned((8'hb7))) ?
              (~^(wire197 && reg271)) : ($signed(reg287) ?
                  ((8'haa) & reg277) : (wire196 ? wire193 : reg286))) ?
          $signed((~^(reg277 ?
              wire285 : reg279))) : ($unsigned($signed(reg294)) ?
              (~^wire268) : $signed((|wire265)))));
      reg408 = $unsigned(wire270);
      reg409 = wire354[(3'h6):(3'h5)];
    end
  assign wire410 = {wire195};
  assign wire411 = reg278[(1'h1):(1'h1)];
  module412 modinst435 (.y(wire434), .wire413(reg409), .wire416(reg405), .wire417(wire269), .wire414(reg273), .wire415(reg408), .clk(clk));
  always
    @(posedge clk) begin
      reg436 = wire194[(3'h7):(3'h4)];
      reg437 = (~&reg294);
      reg438 <= ((wire269 < (reg271 ?
          wire196 : (^{(8'hbd), (8'ha0)}))) && wire267[(5'h12):(3'h6)]);
    end
  module355 modinst440 (.wire359(wire263), .wire356(wire375), .y(wire439), .wire357(wire295), .wire358(reg291), .clk(clk));
endmodule

module module27
#( parameter param145 = ((((+((8'hb8) >> (8'hb8))) ? {(~(8'hb5))} : (((8'hac) ? (7'h41) : (8'hb8)) > ((8'hbc) ? (7'h40) : (8'h9d)))) ? (((~|(8'h9c)) ? ((8'hbc) ? (8'ha8) : (8'h9f)) : ((8'had) ? (8'haf) : (8'ha4))) ? (((8'h9c) - (8'hb0)) ^~ ((8'ha5) < (8'hb0))) : (!((8'hb3) ? (8'ha8) : (8'hbd)))) : {(8'hbc)}) ? (((-(~&(8'hbc))) ? (&((8'hba) ? (8'hbd) : (8'hb3))) : (+(~^(8'hb0)))) ? (({(8'hb2)} - {(8'hbd), (8'hba)}) <= (((7'h42) > (8'hba)) && ((8'haf) < (8'hb3)))) : (^(((8'ha5) <<< (8'hbe)) ? {(8'hba)} : {(8'ha2), (8'ha9)}))) : {((((8'hbf) <<< (8'hb2)) && ((8'hac) | (7'h43))) << ({(8'haf), (8'hae)} ? ((8'hbd) & (8'hae)) : ((8'ha9) ~^ (8'ha5))))}) )
(y, clk, wire28, wire29, wire30, wire31);
  output wire [(32'h15b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire28;
  input wire [(4'ha):(1'h0)] wire29;
  input wire signed [(5'h13):(1'h0)] wire30;
  input wire [(3'h6):(1'h0)] wire31;
  wire signed [(4'h9):(1'h0)] wire144;
  wire signed [(4'hb):(1'h0)] wire143;
  wire [(4'hb):(1'h0)] wire142;
  wire signed [(2'h2):(1'h0)] wire141;
  wire signed [(4'he):(1'h0)] wire140;
  wire [(5'h13):(1'h0)] wire139;
  wire signed [(4'h8):(1'h0)] wire138;
  wire [(5'h15):(1'h0)] wire137;
  wire [(4'hb):(1'h0)] wire136;
  wire [(5'h12):(1'h0)] wire135;
  wire [(3'h4):(1'h0)] wire134;
  wire signed [(3'h7):(1'h0)] wire133;
  wire signed [(3'h4):(1'h0)] wire132;
  wire signed [(5'h13):(1'h0)] wire32;
  wire signed [(5'h13):(1'h0)] wire33;
  reg [(5'h12):(1'h0)] reg34 = (1'h0);
  reg signed [(4'he):(1'h0)] reg35 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg37 = (1'h0);
  reg [(4'h8):(1'h0)] reg38 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg39 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg41 = (1'h0);
  reg [(4'hf):(1'h0)] reg42 = (1'h0);
  reg [(4'hf):(1'h0)] reg43 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire60;
  wire signed [(5'h15):(1'h0)] wire130;
  assign y = {wire144,
                 wire143,
                 wire142,
                 wire141,
                 wire140,
                 wire139,
                 wire138,
                 wire137,
                 wire136,
                 wire135,
                 wire134,
                 wire133,
                 wire132,
                 wire32,
                 wire33,
                 reg34,
                 reg35,
                 reg36,
                 reg37,
                 reg38,
                 reg39,
                 reg40,
                 reg41,
                 reg42,
                 reg43,
                 wire60,
                 wire130,
                 (1'h0)};
  assign wire32 = wire31;
  assign wire33 = (((&wire31[(1'h0):(1'h0)]) ?
                          $unsigned(wire32[(1'h1):(1'h1)]) : (8'h9c)) ?
                      wire30 : $signed((!{{wire30}})));
  always
    @(posedge clk) begin
      if ({($unsigned($unsigned((8'hbf))) >> ({{wire29}, (~|wire29)} ?
              (^wire28[(1'h0):(1'h0)]) : $unsigned(((7'h44) <= wire28))))})
        begin
          reg34 <= (($signed((+wire29[(4'h8):(3'h7)])) & (&wire29[(4'h8):(2'h3)])) ?
              wire28 : $signed($signed((~(wire29 ^~ (8'ha0))))));
          reg35 = reg34[(4'h8):(1'h0)];
          reg36 <= ($unsigned(((wire33[(4'h8):(3'h5)] ?
                  wire32 : ((8'hbc) ? (8'hb8) : reg34)) ?
              $unsigned(wire29[(1'h1):(1'h1)]) : $unsigned((wire29 ?
                  wire33 : wire29)))) && wire28);
        end
      else
        begin
          reg34 <= reg34;
          reg35 <= ($unsigned((~^$signed($signed(wire32)))) ?
              wire29 : ($signed(wire31) << (wire29[(4'h8):(3'h7)] ?
                  wire31 : (~&((7'h42) ^~ reg35)))));
          reg36 <= (($signed((~wire28)) ?
                  ($unsigned({wire29}) ?
                      ($unsigned(wire31) ?
                          (8'h9f) : reg36[(4'ha):(1'h1)]) : {(wire32 - reg36),
                          reg36[(3'h5):(1'h0)]}) : (~&$signed((wire30 >>> reg34)))) ?
              (($unsigned((wire31 ? wire28 : reg36)) ?
                  ((&wire32) ? reg34 : (wire29 >> reg36)) : {$signed(reg35),
                      $unsigned(wire31)}) > ((~|wire33) <<< wire29)) : $signed(wire32[(4'h8):(1'h0)]));
        end
      reg37 <= (({(wire28 >= $signed(reg34))} + (8'hac)) ?
          $signed((wire33[(4'h8):(1'h0)] ?
              $unsigned(wire29[(1'h1):(1'h0)]) : ((wire33 ? reg34 : reg35) ?
                  $signed(reg34) : ((7'h40) || reg35)))) : reg35[(1'h1):(1'h1)]);
      if (reg37[(4'h9):(3'h5)])
        begin
          reg38 <= $signed($signed($signed((((8'ha0) ?
              wire31 : wire31) + (reg34 ? wire28 : reg34)))));
          if (reg34[(3'h5):(1'h0)])
            begin
              reg39 <= {$signed({($signed(wire28) ?
                          (wire30 ^~ wire28) : (~|wire28))}),
                  ((|(wire30 ?
                      $signed((8'hb1)) : wire30[(3'h4):(1'h0)])) && ((wire29[(3'h7):(3'h5)] ?
                      (!wire30) : ((8'ha3) ?
                          reg37 : reg34)) >= {$unsigned(reg36), (|reg35)}))};
              reg40 <= wire31;
              reg41 <= $signed((reg37[(4'h8):(1'h0)] >> (!($signed((8'hac)) ?
                  (reg39 * wire31) : $unsigned((8'hab))))));
              reg42 <= (~&reg37);
              reg43 <= ((~^(~&$signed($unsigned(reg38)))) ?
                  (~&(~|((reg37 ? reg40 : reg36) ?
                      (^reg36) : {(8'hb8)}))) : {((+$unsigned(reg41)) ?
                          ((wire32 ?
                              reg42 : wire32) ^ $signed(wire29)) : (^~(reg40 | reg41)))});
            end
          else
            begin
              reg39 = (8'h9c);
            end
        end
      else
        begin
          reg38 = {(&reg39)};
        end
    end
  module44 modinst61 (.wire48(reg39), .wire45(reg35), .clk(clk), .wire47(wire32), .y(wire60), .wire46(reg42));
  module62 modinst131 (.clk(clk), .wire63(reg40), .y(wire130), .wire66(reg38), .wire65(wire32), .wire67(wire30), .wire64(reg41));
  assign wire132 = ((+wire28[(3'h5):(2'h2)]) >= (~^reg41[(1'h0):(1'h0)]));
  assign wire133 = {$unsigned(wire30)};
  assign wire134 = (~reg38);
  assign wire135 = wire31;
  assign wire136 = reg39;
  assign wire137 = ($unsigned((7'h43)) + {wire135, $unsigned(reg40)});
  assign wire138 = reg43[(3'h4):(1'h1)];
  assign wire139 = $unsigned(wire28);
  assign wire140 = (!wire135[(4'h9):(1'h1)]);
  assign wire141 = {(&$signed($signed(wire30[(4'ha):(1'h1)])))};
  assign wire142 = {(^$signed(wire138)), {$unsigned(reg40[(3'h5):(1'h0)])}};
  assign wire143 = wire141[(2'h2):(1'h1)];
  assign wire144 = reg42;
endmodule

module module62  (y, clk, wire67, wire66, wire65, wire64, wire63);
  output wire [(32'h313):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire67;
  input wire signed [(4'h8):(1'h0)] wire66;
  input wire [(5'h10):(1'h0)] wire65;
  input wire signed [(5'h14):(1'h0)] wire64;
  input wire [(3'h7):(1'h0)] wire63;
  wire [(4'h8):(1'h0)] wire129;
  wire [(3'h5):(1'h0)] wire128;
  wire signed [(3'h7):(1'h0)] wire127;
  wire signed [(5'h15):(1'h0)] wire126;
  wire signed [(5'h12):(1'h0)] wire125;
  wire [(2'h3):(1'h0)] wire124;
  reg [(5'h13):(1'h0)] reg123 = (1'h0);
  reg [(5'h12):(1'h0)] reg122 = (1'h0);
  reg [(5'h12):(1'h0)] reg121 = (1'h0);
  reg [(2'h3):(1'h0)] reg120 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg117 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg116 = (1'h0);
  reg [(4'h8):(1'h0)] reg115 = (1'h0);
  reg [(4'hd):(1'h0)] reg114 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg113 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire112;
  reg signed [(4'he):(1'h0)] reg111 = (1'h0);
  reg [(5'h11):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg109 = (1'h0);
  reg [(2'h2):(1'h0)] reg108 = (1'h0);
  wire [(3'h5):(1'h0)] wire107;
  wire signed [(3'h6):(1'h0)] wire106;
  wire [(4'hc):(1'h0)] wire105;
  reg signed [(4'he):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg103 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg102 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg101 = (1'h0);
  reg [(3'h4):(1'h0)] reg100 = (1'h0);
  reg [(5'h14):(1'h0)] reg99 = (1'h0);
  reg [(3'h7):(1'h0)] reg98 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg97 = (1'h0);
  reg [(2'h2):(1'h0)] reg96 = (1'h0);
  reg [(2'h3):(1'h0)] reg95 = (1'h0);
  reg signed [(4'he):(1'h0)] reg94 = (1'h0);
  wire [(4'hf):(1'h0)] wire93;
  wire signed [(4'h9):(1'h0)] wire92;
  wire [(4'he):(1'h0)] wire91;
  wire [(5'h10):(1'h0)] wire90;
  wire signed [(5'h11):(1'h0)] wire89;
  reg signed [(5'h12):(1'h0)] reg88 = (1'h0);
  reg [(5'h14):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg86 = (1'h0);
  reg [(4'hd):(1'h0)] reg85 = (1'h0);
  reg [(5'h12):(1'h0)] reg84 = (1'h0);
  reg [(5'h13):(1'h0)] reg83 = (1'h0);
  reg [(3'h4):(1'h0)] reg82 = (1'h0);
  reg [(3'h5):(1'h0)] reg81 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg79 = (1'h0);
  reg [(4'ha):(1'h0)] reg78 = (1'h0);
  reg [(4'h8):(1'h0)] reg77 = (1'h0);
  reg [(4'ha):(1'h0)] reg76 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg75 = (1'h0);
  reg [(5'h11):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg72 = (1'h0);
  reg [(2'h3):(1'h0)] reg71 = (1'h0);
  reg [(5'h11):(1'h0)] reg70 = (1'h0);
  reg [(4'hb):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg68 = (1'h0);
  assign y = {wire129,
                 wire128,
                 wire127,
                 wire126,
                 wire125,
                 wire124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 wire112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 wire107,
                 wire106,
                 wire105,
                 reg104,
                 reg103,
                 reg102,
                 reg101,
                 reg100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 wire93,
                 wire92,
                 wire91,
                 wire90,
                 wire89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((($signed({(7'h43)}) ~^ (+{wire66})) > $unsigned((^$unsigned(wire67[(3'h6):(3'h4)])))))
        begin
          reg68 <= $signed((8'h9e));
          if ({($signed($unsigned($signed(reg68))) ?
                  wire65[(3'h5):(1'h0)] : wire65[(4'hb):(3'h7)])})
            begin
              reg69 = wire64;
              reg70 <= {($signed(($unsigned((8'ha0)) ? {wire63} : wire67)) ?
                      (&(|reg68)) : $signed(((wire65 >>> wire67) < (~&wire65))))};
              reg71 <= (($signed((-(reg70 ? (8'ha9) : wire66))) ?
                      (8'h9f) : ((((8'ha7) == wire63) ?
                          $signed(wire66) : $signed(reg70)) < wire63[(2'h2):(1'h0)])) ?
                  $signed(((&$signed(wire67)) >> ($unsigned(reg68) <<< (reg68 | wire66)))) : (wire66 ~^ {(wire63[(3'h6):(1'h0)] != reg70)}));
            end
          else
            begin
              reg69 <= reg69[(2'h2):(1'h0)];
              reg70 <= reg70;
              reg71 <= $unsigned($signed((-{wire63[(3'h4):(1'h0)],
                  (^~reg69)})));
              reg72 = wire66[(2'h2):(1'h1)];
              reg73 <= {(+(wire65 - wire65[(5'h10):(3'h6)])),
                  (-((reg70[(1'h0):(1'h0)] ^ wire67) >>> (reg69[(1'h0):(1'h0)] + (reg69 ?
                      reg69 : (7'h44)))))};
            end
          reg74 = (reg69 >= reg69[(3'h4):(3'h4)]);
        end
      else
        begin
          if (wire63[(3'h4):(2'h3)])
            begin
              reg68 = wire65[(1'h0):(1'h0)];
            end
          else
            begin
              reg68 <= (^~reg68);
              reg69 <= (((+reg71[(1'h0):(1'h0)]) ?
                  (reg68 > $signed({wire67,
                      wire66})) : (~$unsigned((8'ha5)))) || reg72[(5'h12):(4'hf)]);
              reg70 <= ($unsigned((~{wire66,
                  wire65[(4'h8):(3'h5)]})) != {{($unsigned(wire64) ?
                          ((8'h9d) ^ reg73) : reg72)}});
            end
          reg71 <= $signed(($signed(((wire65 ? wire67 : reg72) ?
              {reg73, reg74} : $signed(wire64))) && {$signed((reg73 ?
                  wire64 : wire67)),
              wire64[(3'h6):(1'h1)]}));
        end
      reg75 <= reg74;
      reg76 <= (((-(~|reg71[(2'h3):(2'h3)])) | $unsigned((^~reg70[(4'hd):(4'hc)]))) ?
          (($signed(wire66) ? wire63 : $signed((reg74 ? reg68 : reg75))) ?
              (&(~|wire66)) : $unsigned((&reg69[(3'h6):(1'h1)]))) : reg69);
      if (({reg71} ^ ({(reg72[(1'h1):(1'h1)] ^ $unsigned(wire64)),
              (~^(wire65 * reg73))} ?
          $unsigned($unsigned((wire63 == wire63))) : {$signed(reg72[(5'h13):(5'h10)]),
              $unsigned((reg74 ? wire65 : wire64))})))
        begin
          if ((~|reg68[(1'h1):(1'h1)]))
            begin
              reg77 = (~|(&reg74[(2'h2):(2'h2)]));
              reg78 = wire64;
              reg79 = $unsigned(((reg71[(1'h1):(1'h0)] ^~ ($unsigned(reg74) < (-wire63))) <<< $signed(reg74)));
            end
          else
            begin
              reg77 <= ($unsigned(reg72[(5'h14):(3'h4)]) >> (&$unsigned((wire67[(3'h5):(2'h3)] ?
                  (~^reg78) : $unsigned((8'hae))))));
              reg78 <= reg71[(1'h0):(1'h0)];
              reg79 <= reg69;
              reg80 <= ($unsigned((!(8'hbb))) ?
                  {{{(reg75 ? (8'hb9) : reg79)}, (!reg79[(4'ha):(4'h9)])},
                      reg74[(5'h11):(4'hf)]} : wire64);
            end
          if ((~|$unsigned($unsigned((8'ha1)))))
            begin
              reg81 <= ({{reg73}} ? reg78[(3'h4):(2'h2)] : $signed(reg78));
              reg82 = wire66;
              reg83 = $signed($unsigned(($signed(wire67) <= {reg71})));
              reg84 <= $signed(({reg79[(4'he):(4'hd)],
                      ($unsigned((8'had)) ? $signed(reg80) : reg77)} ?
                  (((reg71 ~^ reg69) > (~|wire66)) ?
                      $signed(reg81[(2'h3):(1'h0)]) : reg73) : $unsigned(($unsigned(reg79) <= wire65))));
              reg85 = wire65;
            end
          else
            begin
              reg81 <= $signed({(((+(8'h9e)) ? $signed((7'h44)) : (+reg84)) ?
                      $signed($signed(reg70)) : (~^{reg80, reg68}))});
              reg82 <= $signed((((&(wire66 ? wire64 : reg80)) ?
                      $unsigned((~^reg69)) : {(reg71 | reg68), (~^reg83)}) ?
                  {reg69[(2'h3):(1'h0)],
                      reg85[(3'h5):(3'h4)]} : (~&{(wire67 != reg75)})));
            end
          reg86 <= (((reg75 + (reg83 + (reg75 < (7'h40)))) >>> $unsigned(((reg77 ?
                  reg74 : reg80) >>> (~reg70)))) ?
              reg69[(1'h0):(1'h0)] : $unsigned((($signed(reg83) >> (~wire67)) - reg82[(3'h4):(1'h1)])));
          reg87 <= $signed({(({reg77, (8'h9c)} ?
                  (reg69 ^~ (8'hb2)) : (8'hb2)) <= (8'hac))});
          reg88 = (8'hb2);
        end
      else
        begin
          if ((wire64 <= $unsigned($signed(reg83[(3'h5):(1'h1)]))))
            begin
              reg77 = reg76;
            end
          else
            begin
              reg77 <= {reg77[(3'h5):(2'h2)]};
              reg78 <= {(reg81[(3'h4):(2'h2)] ?
                      (wire63[(1'h0):(1'h0)] ?
                          $unsigned(((8'ha8) ? reg69 : reg69)) : ((reg81 ?
                                  reg82 : reg75) ?
                              reg68 : (reg73 >= (8'hbb)))) : reg71[(1'h0):(1'h0)])};
              reg79 = (^wire63);
              reg80 <= $unsigned((((8'h9f) ^~ (8'hbd)) ?
                  $unsigned(((reg82 <= (8'hb3)) ?
                      $unsigned((8'hbe)) : reg86[(2'h2):(1'h0)])) : ({reg73} <= ((|reg69) >= (reg77 ?
                      reg68 : reg83)))));
            end
        end
    end
  assign wire89 = (~reg69);
  assign wire90 = (-({wire63[(3'h4):(3'h4)],
                      $unsigned(reg77)} >= $unsigned({reg85[(4'hb):(2'h2)]})));
  assign wire91 = $signed(reg70[(4'h9):(1'h0)]);
  assign wire92 = {(+reg86)};
  assign wire93 = ((((((8'hb5) <<< reg70) ?
                          wire66[(1'h0):(1'h0)] : (reg82 ?
                              (8'ha0) : reg71)) ^ reg71) < ((^~$unsigned(wire92)) ?
                          reg87 : (^(&wire63)))) ?
                      wire90 : (8'hb6));
  always
    @(posedge clk) begin
      reg94 <= {$unsigned(wire89)};
      reg95 <= (~|((~^(!(reg81 ?
          wire93 : reg77))) <= $unsigned(($signed(wire65) >= ((8'hb6) ?
          (7'h42) : reg79)))));
      if (reg71[(2'h3):(2'h3)])
        begin
          if ({$unsigned(reg81[(2'h2):(1'h1)])})
            begin
              reg96 = reg84;
            end
          else
            begin
              reg96 = reg86;
              reg97 <= (+(($signed($unsigned((8'hb3))) > $unsigned({reg83})) ?
                  $unsigned($unsigned($unsigned(reg87))) : ((~^$unsigned(reg78)) ^~ reg79[(4'he):(3'h7)])));
              reg98 = $signed((8'h9f));
              reg99 = (^reg82);
            end
          reg100 <= ($unsigned((reg75[(1'h1):(1'h0)] > {(^reg95),
                  $signed(wire93)})) ?
              (wire66[(1'h1):(1'h1)] == (7'h44)) : (~|{reg95[(1'h0):(1'h0)],
                  {$signed(reg95)}}));
          if ($unsigned(reg96))
            begin
              reg101 <= (($signed(reg99[(4'h8):(3'h4)]) & {$unsigned((&wire89))}) - ((+$signed((reg76 ?
                  wire89 : (8'hbc)))) ~^ {$signed({reg73})}));
              reg102 <= (-($signed(((^wire90) ~^ $signed(wire67))) ?
                  reg81[(1'h0):(1'h0)] : reg84[(3'h6):(1'h0)]));
              reg103 = reg81[(1'h1):(1'h0)];
              reg104 = $signed(reg88);
            end
          else
            begin
              reg101 <= (({{(reg104 > reg69)}, $unsigned((wire91 ~^ reg80))} ?
                  $unsigned(reg100[(2'h3):(1'h0)]) : ((~^((8'ha5) - reg96)) >> ((~&wire65) ?
                      (reg78 ^~ wire64) : (reg104 ?
                          reg78 : reg75)))) ^~ ($unsigned(((wire91 ?
                          reg94 : reg95) ?
                      $signed(reg69) : ((8'hab) ^~ reg72))) ?
                  ($unsigned((!wire67)) >>> reg84) : $unsigned($signed((reg84 ?
                      reg75 : wire93)))));
            end
        end
      else
        begin
          reg96 <= (+{$signed(($signed(reg81) ? (^~reg87) : {wire89})),
              $unsigned(((reg102 ? reg95 : reg70) >>> reg80[(2'h3):(2'h2)]))});
          reg97 = $unsigned($signed($unsigned($unsigned($signed(reg99)))));
          reg98 <= (+$signed({{(~reg74), (reg103 ? reg95 : reg88)},
              $signed(reg80[(4'hc):(3'h4)])}));
        end
    end
  assign wire105 = ($signed(reg71) ?
                       {{(|$unsigned(reg100)),
                               {reg85[(4'hd):(4'h8)],
                                   ((8'hbc) ? wire92 : reg79)}}} : {reg70,
                           reg97[(4'hd):(2'h2)]});
  assign wire106 = (^(8'ha7));
  assign wire107 = $unsigned(reg102);
  always
    @(posedge clk) begin
      reg108 = reg94[(4'ha):(3'h4)];
      if (($signed(reg74[(4'ha):(1'h0)]) ?
          $unsigned({reg81,
              wire63}) : (($signed((~|wire89)) + (~&reg103[(3'h7):(2'h3)])) ?
              reg102[(2'h3):(1'h0)] : (reg80 == (reg69 ?
                  reg73[(1'h1):(1'h1)] : (reg104 ? reg96 : reg79))))))
        begin
          reg109 <= (~^{($signed({(7'h44)}) ?
                  ((reg79 >= reg85) != $signed((8'ha5))) : reg83[(4'hc):(4'h9)]),
              reg98[(3'h5):(3'h4)]});
          reg110 = reg72;
        end
      else
        begin
          reg109 = $signed($signed($signed((~$signed(reg74)))));
          reg110 <= $unsigned($signed(($signed((reg88 >= reg80)) ?
              reg103[(5'h10):(5'h10)] : wire91)));
          reg111 <= $signed({((reg77[(3'h6):(1'h1)] > {reg103}) ?
                  reg77[(1'h1):(1'h1)] : (+$unsigned((8'hbf)))),
              reg84});
        end
    end
  assign wire112 = (^$signed(reg100));
  always
    @(posedge clk) begin
      reg113 <= reg84;
      reg114 <= $signed(reg81);
      reg115 = reg108;
      if ((wire92 ?
          (((wire63[(2'h3):(1'h0)] ? reg85 : reg75) >> {(reg81 ? reg98 : reg82),
                  (reg71 ^~ reg111)}) ?
              $signed($unsigned((^reg84))) : $signed((&{reg87}))) : reg85[(4'hb):(3'h5)]))
        begin
          if (reg70)
            begin
              reg116 = reg69[(3'h7):(2'h3)];
              reg117 = (-($unsigned($signed((-(8'ha8)))) > {$signed(reg70[(4'ha):(2'h2)])}));
            end
          else
            begin
              reg116 <= $unsigned({{{reg103[(4'hb):(3'h4)],
                          (reg104 ? (8'hb1) : reg71)}}});
              reg117 = (!((&wire67) ? (^$signed((^wire107))) : (8'hb9)));
              reg118 = {(~|reg68), reg74};
            end
          reg119 = reg86;
          reg120 <= $unsigned($unsigned($signed({$signed(reg73),
              $signed(wire91)})));
          reg121 = reg94;
        end
      else
        begin
          if ($unsigned(wire89))
            begin
              reg116 = $signed((~|reg96));
              reg117 <= (($signed(((reg85 + (8'hae)) >= reg96[(1'h0):(1'h0)])) ?
                      $unsigned((~|reg73)) : ($unsigned((reg109 ^~ reg85)) ?
                          reg85[(3'h5):(2'h3)] : (wire64 ?
                              reg111[(2'h2):(2'h2)] : {reg69, reg79}))) ?
                  reg76 : (reg99[(5'h13):(4'h9)] + ((reg78 & reg98[(2'h2):(1'h0)]) ?
                      ((reg95 >= (7'h41)) ?
                          (reg96 ? wire112 : reg111) : {wire64}) : reg86)));
              reg118 = $unsigned(reg82);
            end
          else
            begin
              reg116 = $unsigned(reg99[(5'h12):(4'h9)]);
              reg117 <= $signed($signed((reg84[(4'he):(3'h5)] * {(reg98 ?
                      reg77 : reg73),
                  (reg117 + reg78)})));
            end
          if (($unsigned((reg109[(3'h4):(2'h2)] <= {reg74[(4'h9):(3'h7)]})) ?
              wire112 : $unsigned(reg114[(1'h0):(1'h0)])))
            begin
              reg119 <= (^(((!reg75) && $unsigned({reg71})) <= (reg121 ?
                  (8'hb0) : $unsigned(reg113))));
              reg120 <= (reg95 ?
                  (reg77 ?
                      (~&wire105) : $unsigned((~|$signed(reg103)))) : {reg113,
                      {(8'hbc),
                          ($signed(reg98) ? (reg108 && reg100) : reg99)}});
            end
          else
            begin
              reg119 <= reg109[(3'h6):(3'h6)];
              reg120 <= (|(($signed($signed(reg84)) ?
                      wire90 : $signed($signed(reg87))) ?
                  (~^({wire63, reg85} ?
                      (reg73 ?
                          reg85 : reg103) : $unsigned(reg94))) : $unsigned(($unsigned(reg87) ?
                      reg119 : $signed(wire65)))));
            end
          reg121 <= (reg116[(1'h0):(1'h0)] ?
              ({$signed($signed((8'ha2))),
                  (|((8'hb0) ? reg98 : reg104))} <= {$unsigned((wire105 ?
                      reg114 : reg80))}) : (!{($signed(wire64) > reg101)}));
          reg122 = (-$unsigned($signed(reg83)));
          reg123 = (~&$signed(reg121[(4'ha):(2'h2)]));
        end
    end
  assign wire124 = ((8'hb2) | {((reg110 ?
                           $signed(reg79) : $unsigned((8'hab))) && $unsigned($unsigned(reg74))),
                       (reg120[(1'h0):(1'h0)] && $signed(reg98[(3'h7):(3'h5)]))});
  assign wire125 = (|reg71[(1'h0):(1'h0)]);
  assign wire126 = (((reg81[(2'h2):(1'h0)] && (!(^wire66))) == ($unsigned({reg96}) ?
                           $unsigned(reg83[(2'h2):(1'h1)]) : (|reg72))) ?
                       (~wire67) : {{(((8'hbe) > wire63) != $unsigned(reg119))}});
  assign wire127 = $signed(reg117);
  assign wire128 = ($unsigned({(reg99 ?
                               (reg111 ? reg118 : wire64) : $signed(reg119)),
                           (((8'hb7) ? wire92 : (8'hb5)) + wire64)}) ?
                       $unsigned({$signed($signed(wire112))}) : reg98[(3'h4):(1'h0)]);
  assign wire129 = {(8'h9d)};
endmodule

module module44
#(parameter param58 = (8'hb7), parameter param59 = param58)
(y, clk, wire48, wire47, wire46, wire45);
  output wire [(32'h7d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'ha):(1'h0)] wire48;
  input wire [(5'h13):(1'h0)] wire47;
  input wire [(2'h3):(1'h0)] wire46;
  input wire signed [(4'he):(1'h0)] wire45;
  wire signed [(4'he):(1'h0)] wire57;
  wire [(5'h14):(1'h0)] wire56;
  wire signed [(5'h12):(1'h0)] wire55;
  wire [(5'h14):(1'h0)] wire54;
  wire signed [(3'h5):(1'h0)] wire53;
  wire [(3'h4):(1'h0)] wire52;
  wire signed [(4'hc):(1'h0)] wire51;
  wire signed [(4'hd):(1'h0)] wire50;
  wire [(5'h12):(1'h0)] wire49;
  assign y = {wire57,
                 wire56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire49,
                 (1'h0)};
  assign wire49 = $signed(wire48);
  assign wire50 = wire49;
  assign wire51 = wire47;
  assign wire52 = (8'hb7);
  assign wire53 = ((+($unsigned(wire46[(2'h2):(1'h0)]) ?
                      wire52 : {$unsigned(wire47), wire51})) + (+wire46));
  assign wire54 = ((&wire52) ?
                      {((^(wire49 ? wire49 : wire48)) ?
                              $unsigned(((8'hae) ?
                                  wire51 : wire47)) : ((^wire47) || wire47[(4'h8):(3'h5)]))} : ({(&$signed(wire52))} ?
                          wire51 : (-$signed($signed(wire47)))));
  assign wire55 = $signed((~$signed($signed((~(8'hb4))))));
  assign wire56 = wire53;
  assign wire57 = {wire53[(3'h5):(1'h0)]};
endmodule

module module412  (y, clk, wire417, wire416, wire415, wire414, wire413);
  output wire [(32'h9f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire417;
  input wire signed [(5'h15):(1'h0)] wire416;
  input wire signed [(4'h9):(1'h0)] wire415;
  input wire [(3'h4):(1'h0)] wire414;
  input wire [(4'h9):(1'h0)] wire413;
  wire [(3'h7):(1'h0)] wire433;
  wire signed [(5'h15):(1'h0)] wire432;
  reg [(3'h4):(1'h0)] reg431 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg430 = (1'h0);
  reg [(3'h7):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg428 = (1'h0);
  reg [(4'he):(1'h0)] reg427 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg426 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg425 = (1'h0);
  reg [(4'ha):(1'h0)] reg424 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg423 = (1'h0);
  reg [(3'h4):(1'h0)] reg422 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg420 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg419 = (1'h0);
  wire signed [(4'he):(1'h0)] wire418;
  assign y = {wire433,
                 wire432,
                 reg431,
                 reg430,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 wire418,
                 (1'h0)};
  assign wire418 = $unsigned($unsigned(wire415));
  always
    @(posedge clk) begin
      reg419 <= $unsigned((($signed((wire415 >= wire413)) ? (8'hba) : wire416) ?
          (~&$unsigned(wire415[(4'h8):(3'h6)])) : wire418[(4'h8):(3'h5)]));
      reg420 <= (&wire416);
      if ((wire416 << {(reg419 != (~^wire417[(5'h12):(3'h5)])),
          (($unsigned(wire413) & (|wire417)) ?
              ($unsigned(wire416) >>> $unsigned(wire413)) : wire416)}))
        begin
          if (wire414)
            begin
              reg421 <= wire414[(1'h0):(1'h0)];
              reg422 = wire417[(4'he):(1'h1)];
              reg423 <= $unsigned(reg421[(2'h2):(1'h1)]);
              reg424 <= ($signed({$signed((wire417 >>> wire415))}) << {((!$unsigned(reg423)) ?
                      $signed(wire413[(3'h4):(1'h1)]) : $signed(wire416[(5'h15):(3'h4)]))});
            end
          else
            begin
              reg421 <= (wire413 ?
                  $unsigned($unsigned((^~(reg423 ?
                      wire418 : reg423)))) : wire415);
              reg422 <= (((({(8'ha8), reg423} ?
                      (reg423 | (8'h9c)) : $unsigned(wire414)) ?
                  {$signed(reg419)} : $signed($signed(wire417))) <= $signed((reg420[(4'hf):(4'hc)] >>> $signed(wire417)))) <<< $signed($unsigned($signed(reg422))));
            end
          reg425 <= reg422[(1'h0):(1'h0)];
          reg426 = {{$unsigned($signed(reg420[(4'hd):(4'hb)]))}};
          reg427 = reg425[(1'h0):(1'h0)];
        end
      else
        begin
          reg421 <= $signed((wire414 <= ({$unsigned(wire417)} || ($unsigned(wire413) >> $signed(reg420)))));
          if (reg424)
            begin
              reg422 = reg425[(2'h3):(1'h1)];
              reg423 <= $unsigned(((~&(8'ha6)) ?
                  (~&((wire416 >>> reg426) ?
                      wire415 : {wire417,
                          reg424})) : $signed(reg427[(2'h2):(1'h0)])));
            end
          else
            begin
              reg422 = $signed(wire415);
              reg423 = {wire416, $signed(reg425)};
            end
          reg424 <= ((8'hb7) >>> (|$unsigned(((|(8'haa)) & $signed((8'ha5))))));
          reg425 <= (~reg421);
        end
      if ($unsigned($signed((reg419[(1'h0):(1'h0)] ?
          (^~$unsigned(wire418)) : $unsigned(wire414[(3'h4):(3'h4)])))))
        begin
          reg428 <= ($unsigned((reg423[(1'h1):(1'h0)] ?
              reg427[(2'h2):(1'h0)] : $signed((7'h41)))) >> (reg423[(3'h5):(3'h4)] ?
              $signed(({(7'h44)} ?
                  $signed(wire417) : (reg420 ^~ reg427))) : ((~$unsigned(wire417)) >= reg422[(2'h2):(1'h1)])));
          reg429 = (-(reg420 == reg422));
        end
      else
        begin
          if ((reg425 + $unsigned(wire415)))
            begin
              reg428 = {wire414[(2'h3):(2'h3)]};
            end
          else
            begin
              reg428 <= $unsigned((^(wire418 ^~ $unsigned((wire413 ?
                  reg423 : wire415)))));
            end
          reg429 <= $signed(({wire417, (8'hbb)} <<< ((((8'hae) ?
                      wire414 : reg429) ?
                  reg421[(1'h1):(1'h1)] : {reg423}) ?
              $signed(wire417[(2'h3):(1'h1)]) : ($unsigned(reg424) != (reg422 <= reg421)))));
          reg430 = $unsigned((&reg427));
        end
      reg431 = (reg427 || (^reg423));
    end
  assign wire432 = wire416;
  assign wire433 = wire417[(4'hd):(4'hd)];
endmodule

module module377
#( parameter param401 = (~&(!((((7'h42) ? (8'hae) : (8'hb3)) || {(8'ha4)}) ? ({(8'hac)} <<< (^~(8'hbe))) : (~&((8'haf) ~^ (8'ha8))))))
, parameter param402 = param401 )
(y, clk, wire382, wire381, wire380, wire379, wire378);
  output wire [(32'hb1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire382;
  input wire [(3'h7):(1'h0)] wire381;
  input wire [(3'h5):(1'h0)] wire380;
  input wire signed [(3'h4):(1'h0)] wire379;
  input wire signed [(4'hc):(1'h0)] wire378;
  wire signed [(5'h13):(1'h0)] wire400;
  wire signed [(4'h9):(1'h0)] wire399;
  wire signed [(4'h9):(1'h0)] wire398;
  wire [(5'h11):(1'h0)] wire397;
  wire signed [(2'h3):(1'h0)] wire396;
  reg [(4'ha):(1'h0)] reg395 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg394 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg393 = (1'h0);
  reg [(2'h3):(1'h0)] reg392 = (1'h0);
  reg [(3'h5):(1'h0)] reg391 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg390 = (1'h0);
  reg [(2'h2):(1'h0)] reg389 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg388 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg387 = (1'h0);
  reg [(3'h7):(1'h0)] reg386 = (1'h0);
  reg [(4'ha):(1'h0)] reg385 = (1'h0);
  reg [(5'h14):(1'h0)] reg384 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire383;
  assign y = {wire400,
                 wire399,
                 wire398,
                 wire397,
                 wire396,
                 reg395,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg390,
                 reg389,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg384,
                 wire383,
                 (1'h0)};
  assign wire383 = {{wire379[(2'h2):(1'h1)]},
                       ({((wire382 ? wire380 : wire379) ?
                               wire381[(3'h6):(3'h5)] : {wire378}),
                           {wire380, $unsigned((7'h40))}} != wire379)};
  always
    @(posedge clk) begin
      reg384 <= (8'ha4);
      if ($unsigned((wire382[(4'hc):(4'h9)] ?
          {(&(~wire378))} : $unsigned((~wire379[(2'h3):(1'h0)])))))
        begin
          reg385 <= (wire378[(4'h8):(4'h8)] == wire378[(3'h6):(2'h3)]);
          if ($signed($unsigned($unsigned(($unsigned(wire380) > {wire378,
              wire379})))))
            begin
              reg386 = {(~^{(^(^~(8'ha1)))})};
              reg387 <= {reg385[(3'h4):(3'h4)], (8'ha8)};
              reg388 <= reg387[(2'h3):(1'h0)];
              reg389 = (-reg388);
            end
          else
            begin
              reg386 = reg385[(2'h2):(2'h2)];
              reg387 <= (|(wire379[(2'h3):(1'h0)] ?
                  wire378[(4'h9):(1'h1)] : ((~wire380[(1'h0):(1'h0)]) ~^ ($signed(wire378) ?
                      (wire379 <= wire383) : {wire382}))));
              reg388 = (&$signed((((reg389 | (8'h9d)) & wire379[(3'h4):(1'h0)]) >>> wire381)));
              reg389 <= (-$signed($unsigned(reg387[(1'h1):(1'h1)])));
            end
          reg390 = (!($signed((8'h9c)) ~^ reg385));
          reg391 <= $unsigned((($signed((reg386 ?
                  wire380 : wire379)) || ($unsigned((8'haa)) != (|wire382))) ?
              $signed(reg387[(1'h0):(1'h0)]) : wire378));
        end
      else
        begin
          if ({reg389[(1'h1):(1'h1)]})
            begin
              reg385 <= reg385[(4'h8):(2'h2)];
              reg386 <= reg386;
              reg387 = ((~$signed($signed($unsigned(reg384)))) <<< $unsigned(reg390[(3'h5):(3'h4)]));
              reg388 <= $signed(($signed($unsigned(((7'h44) - reg389))) ?
                  $unsigned($signed((|reg384))) : reg385[(3'h4):(2'h3)]));
            end
          else
            begin
              reg385 <= $signed($signed(reg388));
              reg386 <= $signed((&(~|((wire379 <= reg389) + (reg386 <= reg385)))));
              reg387 <= {(|$unsigned($unsigned($unsigned(reg390)))),
                  {reg384,
                      ($unsigned($unsigned(reg391)) >>> ((!(8'hb6)) ?
                          (&reg384) : (~|(8'hb5))))}};
            end
          if ({wire380[(3'h5):(1'h1)]})
            begin
              reg389 = wire382[(2'h2):(1'h0)];
            end
          else
            begin
              reg389 = {$unsigned(wire379)};
              reg390 <= wire381[(3'h4):(1'h1)];
              reg391 <= ((~&wire381) ~^ ((+((-reg390) ?
                      (reg387 ? reg387 : wire382) : (8'ha5))) ?
                  $unsigned(wire383) : $unsigned(wire381)));
            end
          reg392 <= $unsigned((wire380 ?
              ((^~{reg387,
                  (8'hbe)}) ~^ ($signed((8'hb4)) ^~ (~^reg387))) : $signed($signed(reg386[(2'h3):(2'h2)]))));
          reg393 <= {reg388, reg388[(1'h1):(1'h0)]};
          reg394 = ($unsigned((!((wire382 <<< reg393) >= {reg392}))) & $signed(($unsigned($unsigned(reg392)) << reg389[(2'h2):(1'h0)])));
        end
      reg395 = $signed($signed($unsigned(($signed(reg390) ^~ $signed(reg386)))));
    end
  assign wire396 = $unsigned(reg385);
  assign wire397 = (!$signed(wire380[(3'h4):(3'h4)]));
  assign wire398 = (!$unsigned($unsigned((+reg386))));
  assign wire399 = $unsigned($unsigned((~wire396)));
  assign wire400 = wire396;
endmodule

module module355
#( parameter param374 = ((((&((7'h43) ? (8'hb3) : (8'h9c))) ? (~((8'hab) ? (8'hbd) : (8'hac))) : ((+(8'had)) ? ((8'hb0) ? (7'h42) : (8'h9e)) : ((8'hbf) ? (8'hac) : (8'hb6)))) ? ({((8'ha4) ? (8'had) : (8'ha6))} + ((^(7'h41)) + ((8'ha9) ? (8'ha4) : (8'hb8)))) : (~|(((8'ha2) == (8'ha4)) ? (~^(8'hb3)) : (8'ha6)))) ? ({(&((7'h43) ? (8'ha6) : (8'ha3))), ((^(8'ha0)) ? (~|(8'hbd)) : ((8'hb7) ? (8'hbc) : (8'hbd)))} ? ((((8'hbb) | (8'hb9)) | {(7'h41), (8'hac)}) + (|((8'ha6) >= (8'hbd)))) : (({(8'hb1)} ? {(8'ha6), (8'hab)} : ((8'hb6) ? (8'hb2) : (8'hb2))) << (|(-(8'hb3))))) : (^((|((8'hb6) > (8'hae))) ? (((8'ha7) != (8'ha7)) ~^ ((8'ha5) >>> (7'h44))) : {(^(8'ha4)), ((8'hae) >> (8'ha3))}))) )
(y, clk, wire359, wire358, wire357, wire356);
  output wire [(32'haf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire359;
  input wire [(3'h5):(1'h0)] wire358;
  input wire [(3'h7):(1'h0)] wire357;
  input wire [(4'he):(1'h0)] wire356;
  wire [(4'h8):(1'h0)] wire373;
  wire signed [(2'h2):(1'h0)] wire372;
  wire [(4'hc):(1'h0)] wire371;
  wire [(5'h10):(1'h0)] wire370;
  wire [(4'hc):(1'h0)] wire369;
  wire signed [(3'h7):(1'h0)] wire368;
  wire signed [(5'h15):(1'h0)] wire367;
  wire [(5'h11):(1'h0)] wire366;
  wire [(4'hd):(1'h0)] wire365;
  wire signed [(4'ha):(1'h0)] wire364;
  wire [(3'h7):(1'h0)] wire363;
  wire signed [(5'h14):(1'h0)] wire362;
  wire [(5'h15):(1'h0)] wire361;
  wire signed [(4'h8):(1'h0)] wire360;
  assign y = {wire373,
                 wire372,
                 wire371,
                 wire370,
                 wire369,
                 wire368,
                 wire367,
                 wire366,
                 wire365,
                 wire364,
                 wire363,
                 wire362,
                 wire361,
                 wire360,
                 (1'h0)};
  assign wire360 = wire357[(1'h1):(1'h1)];
  assign wire361 = ((wire356[(4'h8):(3'h6)] ?
                           ($unsigned((|wire359)) ?
                               ((~^wire357) ?
                                   (wire356 != wire357) : (wire356 + wire360)) : wire360[(3'h6):(2'h2)]) : wire356[(4'hb):(4'hb)]) ?
                       ((($unsigned(wire360) - (wire357 ? wire360 : wire360)) ?
                           $signed(wire357) : ({(8'hb2), wire357} ?
                               (+(7'h42)) : {wire358,
                                   wire359})) <= ($signed(wire359[(5'h11):(1'h1)]) != ((wire358 ?
                           wire360 : wire356) >= $signed(wire357)))) : wire356[(1'h0):(1'h0)]);
  assign wire362 = {(&$unsigned(((wire360 ?
                           wire356 : wire356) ^~ (~&wire359))))};
  assign wire363 = ((wire361[(4'hb):(3'h6)] ?
                       $unsigned((~&$unsigned(wire362))) : (wire359 ?
                           ((-wire362) ?
                               $signed((8'hae)) : (-wire358)) : wire356)) & {((~^{wire357,
                               wire356}) ?
                           wire358 : wire357),
                       wire359[(4'ha):(2'h3)]});
  assign wire364 = $signed(wire360[(2'h3):(2'h3)]);
  assign wire365 = $signed(wire361[(1'h1):(1'h0)]);
  assign wire366 = wire362;
  assign wire367 = $unsigned($signed(wire357));
  assign wire368 = {(~{$signed($signed(wire361))}),
                       $signed(($signed((-wire361)) * (8'ha1)))};
  assign wire369 = $unsigned(wire367);
  assign wire370 = ((($signed((~^wire366)) ?
                               wire360[(1'h1):(1'h1)] : $signed($signed(wire356))) ?
                           wire358[(2'h2):(1'h0)] : wire366[(2'h2):(1'h0)]) ?
                       (wire365[(4'h8):(3'h7)] != (wire367 >> $unsigned((wire357 ?
                           wire362 : (7'h43))))) : (wire364 ^ ({wire361[(4'hc):(3'h5)]} && $unsigned(((7'h41) ?
                           wire361 : wire363)))));
  assign wire371 = (8'haa);
  assign wire372 = {(({(wire361 >> wire365), $unsigned((8'hb8))} ?
                               ($unsigned(wire361) ?
                                   ((8'hb3) >>> wire371) : $signed((8'ha4))) : $unsigned((^wire371))) ?
                           $signed($unsigned(wire365)) : wire366[(3'h6):(3'h6)]),
                       (((((8'hb0) ? wire357 : wire365) ?
                                   $signed(wire359) : $unsigned(wire362)) ?
                               wire371 : wire356) ?
                           (($unsigned(wire368) ?
                               $signed(wire356) : (wire366 ?
                                   wire356 : wire365)) - $unsigned($signed(wire364))) : $signed((~wire358)))};
  assign wire373 = ((&(-$unsigned((+(8'ha8))))) ?
                       $unsigned($signed((~^wire367[(4'h8):(2'h2)]))) : wire365);
endmodule

module module296
#( parameter param350 = (~|(-{(((8'hb6) ? (8'had) : (7'h44)) ? ((8'ha6) >= (8'ha2)) : (~&(8'hb8))), (((8'haa) ? (8'h9e) : (8'hb2)) ? ((8'hb7) | (8'hab)) : (8'ha5))}))
, parameter param351 = ((^(((!param350) ^ {param350, param350}) ? param350 : (!{param350}))) >= (!(|((~param350) ? (param350 + (8'ha4)) : (-param350))))) )
(y, clk, wire300, wire299, wire298, wire297);
  output wire [(32'h241):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire300;
  input wire [(4'ha):(1'h0)] wire299;
  input wire signed [(2'h2):(1'h0)] wire298;
  input wire signed [(4'h8):(1'h0)] wire297;
  wire signed [(2'h3):(1'h0)] wire349;
  wire [(4'h9):(1'h0)] wire348;
  wire [(5'h14):(1'h0)] wire347;
  wire [(4'he):(1'h0)] wire346;
  wire signed [(2'h3):(1'h0)] wire345;
  wire [(4'ha):(1'h0)] wire344;
  reg signed [(5'h11):(1'h0)] reg343 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg341 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire340;
  wire [(5'h12):(1'h0)] wire339;
  reg signed [(4'h8):(1'h0)] reg338 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg337 = (1'h0);
  reg [(4'hd):(1'h0)] reg336 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire335;
  wire signed [(2'h2):(1'h0)] wire334;
  wire [(5'h15):(1'h0)] wire333;
  wire [(2'h3):(1'h0)] wire332;
  wire [(4'hc):(1'h0)] wire331;
  reg signed [(4'h9):(1'h0)] reg330 = (1'h0);
  reg [(3'h5):(1'h0)] reg329 = (1'h0);
  reg [(5'h13):(1'h0)] reg328 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg327 = (1'h0);
  reg [(4'hb):(1'h0)] reg326 = (1'h0);
  reg [(4'h8):(1'h0)] reg325 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg324 = (1'h0);
  reg [(5'h12):(1'h0)] reg323 = (1'h0);
  reg [(5'h11):(1'h0)] reg322 = (1'h0);
  reg [(3'h7):(1'h0)] reg321 = (1'h0);
  reg [(3'h5):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg319 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg318 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg317 = (1'h0);
  reg [(5'h11):(1'h0)] reg316 = (1'h0);
  reg [(4'h8):(1'h0)] reg315 = (1'h0);
  reg [(3'h6):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg313 = (1'h0);
  reg [(5'h14):(1'h0)] reg312 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg311 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg310 = (1'h0);
  reg [(4'h8):(1'h0)] reg309 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg308 = (1'h0);
  reg [(3'h5):(1'h0)] reg307 = (1'h0);
  wire signed [(4'hb):(1'h0)] wire306;
  wire [(2'h3):(1'h0)] wire305;
  wire [(3'h4):(1'h0)] wire304;
  wire [(5'h12):(1'h0)] wire303;
  wire [(5'h15):(1'h0)] wire302;
  wire signed [(5'h15):(1'h0)] wire301;
  assign y = {wire349,
                 wire348,
                 wire347,
                 wire346,
                 wire345,
                 wire344,
                 reg343,
                 reg342,
                 reg341,
                 wire340,
                 wire339,
                 reg338,
                 reg337,
                 reg336,
                 wire335,
                 wire334,
                 wire333,
                 wire332,
                 wire331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 wire306,
                 wire305,
                 wire304,
                 wire303,
                 wire302,
                 wire301,
                 (1'h0)};
  assign wire301 = $unsigned(wire300[(2'h2):(2'h2)]);
  assign wire302 = {($signed(wire298) ?
                           (~($signed(wire299) <<< $unsigned(wire297))) : (!(^wire299[(4'h8):(3'h6)]))),
                       wire298};
  assign wire303 = (8'hb9);
  assign wire304 = wire298[(1'h1):(1'h1)];
  assign wire305 = wire302[(5'h15):(4'h9)];
  assign wire306 = $signed($signed(wire305[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      reg307 <= $signed(wire300);
      reg308 <= $unsigned(wire305[(1'h0):(1'h0)]);
      reg309 <= wire301[(5'h13):(5'h11)];
      if (((wire306[(3'h6):(2'h2)] ?
              (~((~&wire302) ?
                  wire299[(3'h6):(2'h2)] : {wire305,
                      wire306})) : wire306[(3'h4):(1'h1)]) ?
          $signed($signed((reg307[(1'h0):(1'h0)] + (wire301 > wire305)))) : $signed(({reg308[(4'h9):(1'h1)]} ?
              $unsigned((wire305 ? reg307 : wire303)) : ((wire302 > wire305) ?
                  $signed(wire304) : (wire299 ? (7'h43) : wire298))))))
        begin
          reg310 <= (wire297 ^~ (!{wire305,
              ($unsigned(wire298) < (wire301 ? wire298 : (8'hbc)))}));
          reg311 = $unsigned(wire304);
        end
      else
        begin
          if ($signed(wire304))
            begin
              reg310 <= ((((^~$signed(reg309)) ?
                          ($unsigned(reg310) ?
                              (wire306 ?
                                  wire300 : reg309) : (wire303 - wire304)) : $unsigned((-reg309))) ?
                      ((^{reg309}) ?
                          wire300[(1'h0):(1'h0)] : wire305[(1'h0):(1'h0)]) : ((reg309 >> wire305[(2'h2):(1'h1)]) <<< {wire302[(4'he):(4'hd)],
                          (!wire297)})) ?
                  (&(((wire304 ?
                      wire299 : wire298) ^~ reg311) - wire298[(1'h0):(1'h0)])) : $signed((8'hbf)));
              reg311 <= $unsigned(($signed((wire299 ^~ (^reg309))) ?
                  wire297 : {($signed((8'ha6)) << (wire301 ?
                          wire306 : wire300)),
                      wire302}));
            end
          else
            begin
              reg310 <= (^(({(wire299 >= wire306)} <<< ((+reg310) | (&wire298))) >>> ((~&(~&wire299)) ?
                  $unsigned(reg307[(2'h2):(1'h1)]) : ($unsigned(reg309) ?
                      {wire306} : $unsigned(reg309)))));
              reg311 = $signed(wire297[(3'h7):(1'h0)]);
              reg312 = wire298[(2'h2):(1'h0)];
            end
          if ((~$unsigned($signed($unsigned((8'hb1))))))
            begin
              reg313 <= $unsigned((~reg310));
              reg314 <= $signed(wire299[(4'h8):(1'h0)]);
              reg315 <= {((^~($unsigned(reg312) | (reg307 ?
                      reg313 : (8'haf)))) & $signed((|$signed(reg314))))};
              reg316 = $unsigned({$signed($signed({(8'hbe), reg309}))});
            end
          else
            begin
              reg313 = reg314[(3'h5):(3'h4)];
              reg314 <= ({(((|wire300) - wire299) ?
                          {wire300, reg316} : $unsigned((~reg310))),
                      $unsigned(reg307)} ?
                  ($unsigned(reg314[(1'h0):(1'h0)]) ^~ ($unsigned((reg310 >> wire300)) * ($unsigned(wire303) ^~ wire297[(3'h7):(3'h4)]))) : $unsigned(({$signed(reg311)} ?
                      {(8'hb3)} : $unsigned((-(8'ha3))))));
              reg315 <= $signed((+({(+reg312)} ?
                  (reg315 ~^ (wire306 && reg316)) : (^~reg315[(3'h5):(1'h1)]))));
              reg316 <= $unsigned($signed(wire304[(1'h0):(1'h0)]));
            end
          reg317 <= reg309;
          reg318 <= (($signed(reg311) ?
                  (!{(reg312 << wire303),
                      $unsigned(wire304)}) : ((+$signed(wire303)) >= ({reg316,
                      reg310} ~^ (reg310 >>> reg312)))) ?
              ($unsigned(reg313[(3'h7):(3'h7)]) ?
                  $unsigned($unsigned(reg317)) : (|wire300[(1'h1):(1'h1)])) : $unsigned($signed((+reg310[(3'h6):(2'h3)]))));
          if ({(&(~reg312[(5'h13):(4'hf)])), wire300[(1'h1):(1'h0)]})
            begin
              reg319 = reg313;
              reg320 = (-$signed((~^wire300[(3'h6):(1'h1)])));
            end
          else
            begin
              reg319 = {wire305, wire304};
            end
        end
      if ({reg317})
        begin
          reg321 <= (8'ha4);
          reg322 <= wire297;
          if ((($unsigned($signed($signed(reg314))) ?
                  $unsigned(reg316) : (($signed((7'h42)) && (wire303 ?
                      reg317 : reg320)) <= ($signed(reg307) - {reg317}))) ?
              ((($unsigned((8'h9f)) ? {reg307} : $unsigned(reg317)) ?
                      (wire299 ? $signed(reg311) : wire303) : (|reg321)) ?
                  (($signed(wire305) <<< reg312[(1'h0):(1'h0)]) ?
                      ($unsigned(wire302) - reg312) : reg313) : $signed(reg318)) : {$signed(($signed(reg312) > (~|wire303)))}))
            begin
              reg323 <= ({{(reg318 ? $signed(wire304) : wire297),
                      (+(reg321 ?
                          (8'h9f) : (8'h9f)))}} || wire306[(3'h4):(1'h0)]);
            end
          else
            begin
              reg323 <= (reg323[(3'h4):(2'h3)] ?
                  (wire305[(2'h2):(2'h2)] ?
                      reg317[(1'h1):(1'h0)] : reg316) : $signed(reg309[(3'h4):(2'h2)]));
              reg324 = reg322;
              reg325 <= ($signed(((-(wire298 || reg317)) & reg309)) ?
                  {wire300,
                      reg310[(5'h10):(4'h8)]} : (wire299[(2'h3):(2'h2)] <<< ((wire297 ?
                      reg314[(1'h1):(1'h1)] : (wire302 ^ reg319)) ~^ reg313)));
            end
          if ((($unsigned(wire299[(1'h1):(1'h1)]) * $signed((!((8'hbf) ?
                  reg320 : wire301)))) ?
              wire303[(1'h1):(1'h0)] : ($unsigned({wire299}) ?
                  wire298 : (($signed(reg324) && reg316) ?
                      (!(!reg320)) : $signed({reg314})))))
            begin
              reg326 = ($signed(reg308) && $unsigned($signed((+$unsigned(reg312)))));
              reg327 = wire300[(3'h7):(3'h4)];
            end
          else
            begin
              reg326 = $signed((wire298 >> (8'ha3)));
              reg327 <= (wire300 ?
                  (8'hba) : $signed($unsigned((~^$unsigned(wire306)))));
              reg328 = ($signed($unsigned($unsigned(wire298[(1'h0):(1'h0)]))) <= $unsigned(wire300));
              reg329 = (!(^((wire301[(5'h14):(3'h4)] > $unsigned(reg317)) | (~$unsigned(reg319)))));
            end
          reg330 = $unsigned((~^reg316));
        end
      else
        begin
          reg321 = reg327[(4'hc):(2'h3)];
          reg322 = (^{reg307[(1'h1):(1'h1)]});
        end
    end
  assign wire331 = reg308[(3'h4):(1'h0)];
  assign wire332 = $signed((8'ha4));
  assign wire333 = ((^~reg314) ?
                       reg320[(3'h4):(2'h3)] : $signed($signed(reg327[(3'h7):(2'h3)])));
  assign wire334 = $unsigned((!{reg321[(1'h0):(1'h0)]}));
  assign wire335 = ((|$signed($signed($unsigned(reg320)))) ^ $unsigned(((reg310 <<< reg307[(1'h0):(1'h0)]) ?
                       ((reg310 ? reg318 : wire302) ?
                           $unsigned(wire306) : (reg330 & reg327)) : {reg315[(1'h0):(1'h0)]})));
  always
    @(posedge clk) begin
      reg336 = reg308[(1'h1):(1'h1)];
      reg337 <= (~|{(((wire331 * reg318) ^~ $unsigned(wire304)) <<< (8'h9d)),
          ({(wire302 < reg311), {(8'hbc), reg321}} - reg318)});
      reg338 = $signed((~|$signed($unsigned($signed(wire297)))));
    end
  assign wire339 = {((^~reg310) + (reg321 ?
                           wire298 : ((!wire297) > (~^wire302)))),
                       (($unsigned((reg337 ? reg320 : reg319)) ?
                               $signed((&wire301)) : reg324[(4'ha):(1'h1)]) ?
                           (8'hbc) : $signed((reg310 ?
                               $signed(reg328) : $unsigned(wire306))))};
  assign wire340 = $unsigned($signed((wire297[(3'h7):(3'h5)] ?
                       ($signed(reg329) ?
                           (wire306 ?
                               reg338 : reg324) : $signed(reg330)) : ($unsigned(reg317) + $signed(reg327)))));
  always
    @(posedge clk) begin
      if (reg323[(3'h7):(3'h6)])
        begin
          reg341 <= $signed($unsigned($unsigned(((reg313 ?
              reg311 : reg312) || (^~reg325)))));
          reg342 = wire305;
        end
      else
        begin
          reg341 = (8'hbb);
          reg342 <= $unsigned({{(wire333 ? wire334 : (8'hbe)), reg342}});
        end
      reg343 = wire299[(3'h6):(2'h3)];
    end
  assign wire344 = {$unsigned(reg311[(4'hd):(4'h8)])};
  assign wire345 = $unsigned($signed((!((wire340 ? wire298 : wire300) ?
                       reg314 : (reg322 ? reg311 : wire334)))));
  assign wire346 = reg316;
  assign wire347 = $unsigned(wire340[(2'h3):(1'h0)]);
  assign wire348 = (~^$signed((~reg313[(4'he):(3'h6)])));
  assign wire349 = $signed($signed($unsigned({reg309[(3'h7):(3'h5)],
                       ((8'ha7) & wire339)})));
endmodule

module module198  (y, clk, wire202, wire201, wire200, wire199);
  output wire [(32'h28e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire202;
  input wire [(5'h13):(1'h0)] wire201;
  input wire signed [(5'h13):(1'h0)] wire200;
  input wire signed [(2'h3):(1'h0)] wire199;
  wire [(3'h6):(1'h0)] wire262;
  reg [(4'h8):(1'h0)] reg261 = (1'h0);
  reg [(4'hb):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg259 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg258 = (1'h0);
  reg [(4'ha):(1'h0)] reg257 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg256 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg255 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg254 = (1'h0);
  reg [(2'h2):(1'h0)] reg253 = (1'h0);
  reg [(4'hc):(1'h0)] reg252 = (1'h0);
  wire [(5'h10):(1'h0)] wire251;
  wire [(4'hf):(1'h0)] wire250;
  wire signed [(5'h11):(1'h0)] wire249;
  reg signed [(3'h4):(1'h0)] reg248 = (1'h0);
  reg [(4'ha):(1'h0)] reg247 = (1'h0);
  reg [(4'he):(1'h0)] reg246 = (1'h0);
  reg [(3'h6):(1'h0)] reg245 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg244 = (1'h0);
  reg [(4'h8):(1'h0)] reg243 = (1'h0);
  reg [(5'h14):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg241 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg239 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg238 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg237 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg236 = (1'h0);
  reg [(2'h2):(1'h0)] reg235 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg234 = (1'h0);
  reg [(5'h15):(1'h0)] reg233 = (1'h0);
  reg [(5'h11):(1'h0)] reg232 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg231 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg229 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg228 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg227 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg226 = (1'h0);
  reg [(4'hc):(1'h0)] reg225 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg224 = (1'h0);
  wire [(4'h9):(1'h0)] wire223;
  wire [(5'h12):(1'h0)] wire222;
  wire signed [(5'h11):(1'h0)] wire221;
  wire signed [(3'h6):(1'h0)] wire220;
  wire [(4'h8):(1'h0)] wire219;
  wire signed [(5'h13):(1'h0)] wire218;
  wire [(4'h8):(1'h0)] wire217;
  reg signed [(4'he):(1'h0)] reg216 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg214 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg213 = (1'h0);
  reg [(5'h11):(1'h0)] reg212 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg211 = (1'h0);
  reg [(4'hd):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg209 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg208 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg207 = (1'h0);
  reg [(5'h11):(1'h0)] reg206 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire205;
  wire signed [(3'h7):(1'h0)] wire204;
  wire signed [(3'h6):(1'h0)] wire203;
  assign y = {wire262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 wire251,
                 wire250,
                 wire249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 reg228,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 wire223,
                 wire222,
                 wire221,
                 wire220,
                 wire219,
                 wire218,
                 wire217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 wire205,
                 wire204,
                 wire203,
                 (1'h0)};
  assign wire203 = {$unsigned((~({(8'hac)} ? (&(8'ha6)) : wire202))),
                       (wire200 ?
                           ($unsigned($signed(wire200)) << $signed(wire202)) : ($signed(wire202) ?
                               wire199[(2'h2):(1'h0)] : wire200[(5'h10):(1'h0)]))};
  assign wire204 = (~&wire199);
  assign wire205 = $signed(wire199[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      reg206 <= $unsigned(wire199[(2'h3):(2'h2)]);
      reg207 <= ($signed($signed($signed((~|reg206)))) ?
          wire205 : (wire203[(1'h0):(1'h0)] ?
              ({reg206, (~wire200)} ?
                  {wire204} : (!(^~reg206))) : ((~|$unsigned(wire200)) && wire202)));
      if (((((wire201[(5'h13):(3'h5)] ?
              (wire199 ? reg207 : wire203) : $unsigned(wire201)) ?
          wire201 : $signed($signed(wire204))) || wire199) ~^ wire203))
        begin
          reg208 = wire203[(2'h2):(2'h2)];
        end
      else
        begin
          reg208 <= (((~&{{wire204, wire203},
              wire204[(3'h6):(1'h1)]}) >>> (-reg208[(1'h1):(1'h0)])) || $signed((^wire203)));
        end
      if (($unsigned(($unsigned((wire199 ? wire200 : wire202)) ?
          ((~^wire204) ^~ $signed((8'hb6))) : (~|(reg206 <= (8'haf))))) >>> (({(-wire199),
              $signed(wire202)} ?
          wire203[(3'h5):(1'h0)] : $unsigned((+reg207))) & ((wire205 ?
          reg208[(4'h9):(3'h4)] : wire201[(4'h8):(3'h7)]) != $signed(wire204)))))
        begin
          reg209 = ($signed(wire205) ? (~&reg208) : $signed(reg206));
          reg210 <= $signed((($unsigned((7'h42)) & wire200[(3'h5):(3'h4)]) ?
              wire203[(3'h6):(2'h3)] : (~^reg207)));
          reg211 = $unsigned((-wire199[(2'h2):(1'h1)]));
          reg212 = (+$signed(reg207));
          reg213 = $unsigned(reg210);
        end
      else
        begin
          reg209 <= ($unsigned((8'ha6)) | (^~(|(+(wire202 ?
              wire205 : reg210)))));
          reg210 <= (^$signed(wire204[(2'h2):(1'h0)]));
          reg211 <= $signed(((reg213 ?
                  ((reg211 ? wire202 : reg211) ?
                      (^reg210) : (!reg211)) : {(8'haf)}) ?
              wire199[(1'h1):(1'h1)] : wire204[(2'h3):(2'h3)]));
          reg212 <= ((($unsigned((8'ha8)) ?
              $signed(wire204) : {$signed((8'ha2))}) && ($unsigned($unsigned(wire201)) ?
              (~$unsigned(reg206)) : wire200)) | reg209[(5'h11):(3'h5)]);
        end
      reg214 = $signed(($signed(wire205) - $signed((~|{reg206}))));
    end
  always
    @(posedge clk) begin
      reg215 = reg207;
      reg216 = $signed($unsigned((~&reg208[(1'h0):(1'h0)])));
    end
  assign wire217 = wire202;
  assign wire218 = (8'ha6);
  assign wire219 = $unsigned($signed((({reg213} ?
                           reg209 : reg214[(3'h7):(3'h7)]) ?
                       $signed((reg214 == reg210)) : ($unsigned(wire201) ?
                           ((7'h41) ^~ wire202) : $unsigned(wire199)))));
  assign wire220 = ($unsigned((-(~&(reg206 ? reg216 : reg208)))) ?
                       reg213[(4'h8):(2'h2)] : ($signed($signed(reg216)) ?
                           (&((wire204 * reg208) * (~^reg215))) : {wire205[(1'h1):(1'h1)]}));
  assign wire221 = {(7'h43),
                       ({reg207[(2'h2):(1'h1)],
                           $unsigned($signed(reg216))} >>> $signed($signed({reg207})))};
  assign wire222 = (~((wire201[(4'he):(4'hc)] || (-(&(8'hae)))) ?
                       wire219[(3'h6):(3'h5)] : ((((8'h9e) ? wire201 : reg210) ?
                               $unsigned(reg206) : ((8'hbf) ?
                                   reg216 : wire221)) ?
                           ((reg214 >= wire205) ?
                               reg210[(4'h9):(1'h0)] : reg210[(4'ha):(4'h9)]) : ($signed((8'hb9)) - reg211))));
  assign wire223 = (|{((|$signed(reg213)) || (~&wire201[(4'h9):(3'h4)]))});
  always
    @(posedge clk) begin
      if ((&$unsigned($unsigned((-((7'h44) & wire221))))))
        begin
          reg224 = reg216[(4'ha):(4'h9)];
          reg225 = wire219;
          if (wire200[(4'hc):(1'h0)])
            begin
              reg226 = reg214[(3'h4):(1'h1)];
              reg227 = $signed(((8'hbc) >= (~&{reg206[(1'h1):(1'h1)]})));
            end
          else
            begin
              reg226 = (8'hb4);
            end
          reg228 <= (($unsigned((^~$unsigned(reg210))) && reg206[(4'hf):(2'h3)]) << ((~^({reg211,
                      reg206} ?
                  $signed(wire218) : $unsigned(reg211))) ?
              (reg216 ?
                  ((wire222 ? wire203 : wire202) ?
                      $signed(wire204) : ((8'hba) > wire203)) : wire220) : ({{wire203,
                          (8'hb4)},
                      {wire201, wire204}} ?
                  (reg215[(3'h6):(1'h0)] ?
                      ((8'hb2) ?
                          reg209 : wire202) : $signed(wire219)) : ((reg211 ?
                      reg209 : reg207) + reg206))));
        end
      else
        begin
          reg224 <= {$signed(($signed((wire222 >>> reg225)) ?
                  ($signed((8'ha6)) < $signed((7'h43))) : reg225[(1'h0):(1'h0)])),
              (((|wire199[(1'h0):(1'h0)]) < (8'hbc)) ?
                  ($unsigned($signed(wire223)) & ((reg226 ? wire221 : reg227) ?
                      $unsigned(reg216) : (&(8'hb3)))) : {reg216[(3'h4):(1'h1)],
                      wire223[(3'h5):(2'h2)]})};
          if ($unsigned((((wire203 ? reg212 : reg206) ?
                  reg226 : {(wire221 & (8'hb7))}) ?
              $unsigned({$unsigned(wire200),
                  wire204[(3'h4):(3'h4)]}) : reg228[(3'h5):(1'h1)])))
            begin
              reg225 <= $signed((~(^wire221[(4'h9):(4'h9)])));
              reg226 <= $unsigned(($signed(wire218) ?
                  (wire222 ?
                      wire199[(2'h2):(1'h0)] : {(wire203 ?
                              reg225 : reg228)}) : (~^((reg206 ?
                      reg224 : reg207) || (8'hab)))));
              reg227 <= (((reg212 - ({(8'hbd)} ? reg212 : $signed(reg207))) ?
                  $signed((^reg227[(3'h6):(1'h0)])) : ($unsigned(reg208) + $unsigned((wire218 ~^ reg210)))) <<< {$unsigned($unsigned(wire219))});
            end
          else
            begin
              reg225 <= {{(((~&wire220) ?
                          $signed(reg213) : (~|(8'hbc))) * reg225)},
                  (^{(8'hb0), $signed(wire218)})};
              reg226 <= (wire199 ?
                  (((reg216[(4'ha):(4'h8)] <<< $signed(reg207)) ?
                      reg215[(3'h6):(3'h4)] : wire199) >= ({reg225} ?
                      wire217 : {$unsigned((8'ha8)),
                          $signed(reg216)})) : (($unsigned((7'h43)) != reg213) ?
                      (reg213[(4'he):(2'h3)] ?
                          $signed((wire220 ^~ wire222)) : {$signed(reg207)}) : ($signed((!reg209)) ?
                          $signed(((8'hac) - wire220)) : $unsigned({wire223}))));
              reg227 = (+wire199);
              reg228 <= $signed($signed(($signed($signed(reg215)) ?
                  ((wire202 ? reg208 : reg212) ?
                      ((8'hb3) ?
                          reg212 : reg210) : {wire221}) : (~&$signed((8'hab))))));
            end
          reg229 <= (($signed(wire220) ?
                  (~|(wire201 & (reg212 != wire217))) : $signed($unsigned((reg225 ^ (8'hbc))))) ?
              wire218[(5'h12):(2'h3)] : (($unsigned($signed((8'hb7))) ?
                      $signed((~wire200)) : $unsigned(reg213)) ?
                  ((reg210 ?
                      (reg211 > reg211) : (wire220 - reg224)) <= ($signed(wire220) ?
                      {(8'hbb)} : ((8'hbc) ?
                          wire199 : reg209))) : $signed(((&reg208) ?
                      (wire221 > reg209) : wire202[(4'h9):(2'h2)]))));
        end
      if ($signed(((wire219 ?
              ({(8'hb4)} ?
                  reg216[(1'h0):(1'h0)] : reg214[(4'h9):(3'h5)]) : $unsigned(reg225[(2'h2):(1'h1)])) ?
          reg225[(3'h5):(1'h1)] : wire220[(2'h2):(1'h1)])))
        begin
          reg230 = $signed(($unsigned(wire220) | $unsigned((((8'hb2) ^ reg224) != (~reg228)))));
          if (reg214)
            begin
              reg231 <= $signed((-wire202[(3'h4):(1'h1)]));
              reg232 <= {((!($unsigned(wire220) ?
                      (8'ha5) : reg212)) << (((wire221 ? reg224 : wire203) ?
                      reg211 : (^~reg206)) < wire204[(1'h0):(1'h0)]))};
              reg233 <= $unsigned((-$unsigned(($signed((8'hbb)) ?
                  reg231 : {reg216}))));
            end
          else
            begin
              reg231 = $signed(reg233);
            end
          reg234 = $signed($signed($signed({(8'hbe), $signed(reg229)})));
        end
      else
        begin
          reg230 <= reg228[(2'h3):(2'h2)];
          reg231 <= $unsigned($unsigned($unsigned(($signed(reg232) ?
              reg215[(3'h4):(2'h2)] : reg213[(2'h3):(2'h3)]))));
          reg232 <= (~(~^($unsigned((wire221 ?
              wire201 : (8'hb3))) > {(~|(7'h41)), $signed(reg232)})));
          if (reg207)
            begin
              reg233 = (~reg211[(4'h9):(4'h8)]);
              reg234 <= (({(reg211[(3'h7):(2'h3)] >>> reg210),
                      ((reg230 && reg212) ?
                          $signed(wire217) : reg211)} > ($signed((wire219 - reg231)) ?
                      wire220[(1'h0):(1'h0)] : wire200)) ?
                  $signed((8'ha5)) : {(reg211[(1'h0):(1'h0)] ?
                          reg208 : {reg213})});
              reg235 = wire204;
              reg236 = $signed($unsigned($signed(((8'hb2) ^~ $signed(reg216)))));
              reg237 = wire221[(4'he):(3'h5)];
            end
          else
            begin
              reg233 = $unsigned(wire220);
            end
          reg238 = $signed(wire201[(4'ha):(1'h1)]);
        end
      reg239 <= ((((~(+wire203)) ^ wire205) + reg208[(1'h0):(1'h0)]) >>> $unsigned(((+$unsigned(reg209)) ~^ {((8'had) ?
              (8'hb9) : reg229)})));
      reg240 <= $signed({$unsigned(wire202[(4'hd):(4'hd)])});
      if ($signed(reg216[(4'hd):(3'h7)]))
        begin
          reg241 = $signed(($unsigned(reg216) < $signed(reg240[(3'h7):(3'h5)])));
          reg242 = wire221;
          reg243 = wire200;
          reg244 <= $signed($signed({($signed(wire199) <<< wire204[(1'h0):(1'h0)]),
              {reg238[(1'h0):(1'h0)]}}));
          if (wire218)
            begin
              reg245 = (~^$unsigned($unsigned((reg225 ^~ (^reg210)))));
              reg246 <= (reg213[(4'hb):(4'ha)] ^~ ({(reg212 ?
                          ((8'hb9) || reg209) : wire201),
                      wire221} ?
                  (wire201[(3'h7):(3'h5)] ?
                      reg226 : $signed((wire200 ?
                          wire200 : (8'hb9)))) : $signed(reg225[(4'hb):(1'h0)])));
              reg247 = $signed(reg235);
              reg248 = $unsigned(reg214[(3'h7):(3'h6)]);
            end
          else
            begin
              reg245 = (reg213 * wire200[(3'h4):(1'h0)]);
            end
        end
      else
        begin
          reg241 = wire220;
        end
    end
  assign wire249 = (($unsigned($unsigned($signed((7'h41)))) ?
                           $signed((reg239[(3'h7):(3'h4)] != $signed(reg233))) : $unsigned(((^~reg243) ?
                               (reg215 ?
                                   reg242 : reg241) : $unsigned(wire219)))) ?
                       $unsigned($unsigned($unsigned((wire218 != reg238)))) : wire218[(4'h8):(1'h0)]);
  assign wire250 = wire200[(3'h6):(3'h4)];
  assign wire251 = reg226;
  always
    @(posedge clk) begin
      reg252 = {wire200, wire251};
    end
  always
    @(posedge clk) begin
      reg253 = reg240;
      reg254 = reg227[(1'h1):(1'h1)];
      reg255 = (7'h41);
    end
  always
    @(posedge clk) begin
      if (($unsigned((~^$unsigned((8'hba)))) + ($signed((reg243 ?
          reg243[(4'h8):(4'h8)] : (-reg234))) ^~ wire251)))
        begin
          reg256 <= ({((reg206 && (reg210 ? (8'hb1) : reg253)) ?
                  wire219[(4'h8):(2'h3)] : reg253[(1'h1):(1'h1)])} <<< ({((wire202 ?
                      (8'hb3) : (8'ha8)) ?
                  (|reg245) : reg235),
              reg212[(2'h3):(1'h1)]} || $unsigned(($signed(wire217) ^ (reg235 ?
              wire202 : wire222)))));
          reg257 <= (^~$signed((reg211 ?
              $unsigned((reg255 ?
                  (8'hb3) : (7'h44))) : wire217[(3'h4):(1'h0)])));
          reg258 <= ((reg243 >>> (^$signed((|wire219)))) ?
              $signed((wire218[(5'h12):(2'h2)] ?
                  (reg241 >> $unsigned(reg255)) : ((reg228 <= wire201) ?
                      (reg213 ? wire250 : reg212) : {reg248,
                          wire251}))) : (($unsigned($unsigned(reg232)) || $unsigned(reg228)) ?
                  (reg216[(3'h6):(2'h3)] ?
                      (reg234[(1'h0):(1'h0)] && (reg245 ?
                          reg239 : reg206)) : $unsigned({reg209,
                          wire202})) : (8'hb9)));
          reg259 = reg208;
          reg260 = (^$signed($signed(reg208[(2'h2):(1'h0)])));
        end
      else
        begin
          reg256 <= $unsigned(($signed(wire201) ?
              reg255[(1'h0):(1'h0)] : reg237));
          reg257 = (-$signed((^~{(wire249 ? reg244 : reg229)})));
        end
      reg261 = (wire201 ? (8'hb8) : reg207);
    end
  assign wire262 = $signed((8'hbf));
endmodule